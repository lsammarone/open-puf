magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< metal1 >>
rect 18580 27001 18626 27046
rect 4286 26662 4411 26737
rect 6437 17954 6539 18043
rect 23626 16080 23678 16086
rect 23626 16016 23678 16028
rect 23626 15958 23678 15964
tri 22957 15892 22965 15900 se
rect 22965 15892 23017 15957
rect 22957 15886 23017 15892
rect 23009 15885 23017 15886
tri 23009 15877 23017 15885 nw
rect 23045 15892 23097 15957
rect 23125 15932 23177 15957
tri 23177 15932 23186 15941 sw
rect 23125 15926 23186 15932
tri 23125 15917 23134 15926 ne
rect 23134 15925 23186 15926
tri 23097 15892 23105 15900 sw
rect 23045 15886 23105 15892
rect 23045 15885 23053 15886
tri 23045 15877 23053 15885 ne
rect 22957 15822 23009 15834
rect 22957 15764 23009 15770
rect 23053 15822 23105 15834
rect 23134 15861 23186 15873
rect 25592 15812 25711 15930
rect 23134 15803 23186 15809
rect 23053 15764 23105 15770
rect 2905 15235 2911 15243
rect 2904 15191 2911 15235
rect 2963 15191 2975 15243
rect 3027 15235 3033 15243
rect 23466 15235 23472 15243
rect 3027 15191 23472 15235
rect 23524 15191 23536 15243
rect 23588 15191 23594 15243
rect 23173 14930 23179 14938
rect 2996 14924 23179 14930
rect 3048 14886 23179 14924
rect 23231 14886 23243 14938
rect 23295 14886 23301 14938
rect 2996 14860 3048 14872
rect 2996 14802 3048 14808
rect 3088 14804 3094 14856
rect 3146 14804 3158 14856
rect 3210 14854 3216 14856
rect 23343 14854 23349 14862
rect 3210 14810 23349 14854
rect 23401 14810 23413 14862
rect 23465 14810 23471 14862
rect 3210 14804 3216 14810
rect 10043 14120 10107 14152
rect 8397 13471 8437 13503
rect 10741 11936 10936 12030
rect 2382 8577 2692 8746
rect 1982 7609 2123 7747
tri 2862 7142 2919 7199 ne
rect 2919 7117 3248 7199
tri 3248 7142 3305 7199 nw
rect 2919 7065 2925 7117
rect 2977 7065 2992 7117
rect 3044 7065 3058 7117
rect 3110 7065 3124 7117
rect 3176 7065 3190 7117
rect 3242 7065 3248 7117
rect 22371 1902 22619 2181
rect 24019 1796 24074 1802
rect 23083 1691 23154 1780
rect 24019 1744 24020 1796
rect 24072 1744 24074 1796
rect 24019 1732 24074 1744
rect 24019 1680 24020 1732
rect 24072 1680 24074 1732
tri 23988 1579 24019 1610 se
rect 24019 1579 24074 1680
rect 22649 1527 22655 1579
rect 22707 1527 22719 1579
rect 22771 1532 24074 1579
rect 22771 1527 22777 1532
rect 16454 912 16460 964
rect 16512 912 16524 964
rect 16576 957 16582 964
rect 16576 951 20950 957
rect 16576 912 20898 951
rect 11258 831 11264 883
rect 11316 831 11328 883
rect 11380 831 11386 883
rect 11544 856 11550 908
rect 11602 856 11614 908
rect 11666 856 11672 908
rect 20898 887 20950 899
rect 20898 829 20950 835
tri 12993 803 13013 823 se
rect 13013 803 13141 823
rect 12691 771 12752 803
rect 12964 771 13141 803
tri 12985 743 13013 771 ne
rect 13013 743 13141 771
rect 13100 50 13141 743
rect 21058 267 21779 268
rect 21058 215 21064 267
rect 21116 215 21130 267
rect 21182 215 21196 267
rect 21248 215 21262 267
rect 21314 215 21328 267
rect 21380 215 21394 267
rect 21446 215 21460 267
rect 21512 215 21526 267
rect 21578 215 21591 267
rect 21643 215 21656 267
rect 21708 215 21721 267
rect 21773 215 21779 267
rect 21058 197 21779 215
rect 21058 145 21064 197
rect 21116 145 21130 197
rect 21182 145 21196 197
rect 21248 145 21262 197
rect 21314 145 21328 197
rect 21380 145 21394 197
rect 21446 145 21460 197
rect 21512 145 21526 197
rect 21578 145 21591 197
rect 21643 145 21656 197
rect 21708 145 21721 197
rect 21773 145 21779 197
rect 21058 127 21779 145
rect 21058 75 21064 127
rect 21116 75 21130 127
rect 21182 75 21196 127
rect 21248 75 21262 127
rect 21314 75 21328 127
rect 21380 75 21394 127
rect 21446 75 21460 127
rect 21512 75 21526 127
rect 21578 75 21591 127
rect 21643 75 21656 127
rect 21708 75 21721 127
rect 21773 75 21779 127
rect 21058 74 21779 75
rect 13058 -2 13064 50
rect 13116 -2 13128 50
rect 13180 -2 13186 50
rect 24884 -321 24890 -269
rect 24942 -321 24954 -269
rect 25006 -321 25120 -269
rect 25172 -321 25184 -269
rect 25236 -321 25242 -269
rect 13024 -2255 13030 -2203
rect 13082 -2255 13094 -2203
rect 13146 -2255 19791 -2203
rect 19843 -2255 19855 -2203
rect 19907 -2255 20476 -2203
rect 20528 -2255 20540 -2203
rect 20592 -2255 20598 -2203
rect 20662 -2255 24936 -2203
<< via1 >>
rect 23626 16028 23678 16080
rect 23626 15964 23678 16016
rect 22957 15834 23009 15886
rect 22957 15770 23009 15822
rect 23053 15834 23105 15886
rect 23053 15770 23105 15822
rect 23134 15873 23186 15925
rect 23134 15809 23186 15861
rect 2911 15191 2963 15243
rect 2975 15191 3027 15243
rect 23472 15191 23524 15243
rect 23536 15191 23588 15243
rect 2996 14872 3048 14924
rect 23179 14886 23231 14938
rect 23243 14886 23295 14938
rect 2996 14808 3048 14860
rect 3094 14804 3146 14856
rect 3158 14804 3210 14856
rect 23349 14810 23401 14862
rect 23413 14810 23465 14862
rect 2925 7065 2977 7117
rect 2992 7065 3044 7117
rect 3058 7065 3110 7117
rect 3124 7065 3176 7117
rect 3190 7065 3242 7117
rect 24020 1744 24072 1796
rect 24020 1680 24072 1732
rect 22655 1527 22707 1579
rect 22719 1527 22771 1579
rect 16460 912 16512 964
rect 16524 912 16576 964
rect 11264 831 11316 883
rect 11328 831 11380 883
rect 11550 856 11602 908
rect 11614 856 11666 908
rect 20898 899 20950 951
rect 20898 835 20950 887
rect 21064 215 21116 267
rect 21130 215 21182 267
rect 21196 215 21248 267
rect 21262 215 21314 267
rect 21328 215 21380 267
rect 21394 215 21446 267
rect 21460 215 21512 267
rect 21526 215 21578 267
rect 21591 215 21643 267
rect 21656 215 21708 267
rect 21721 215 21773 267
rect 21064 145 21116 197
rect 21130 145 21182 197
rect 21196 145 21248 197
rect 21262 145 21314 197
rect 21328 145 21380 197
rect 21394 145 21446 197
rect 21460 145 21512 197
rect 21526 145 21578 197
rect 21591 145 21643 197
rect 21656 145 21708 197
rect 21721 145 21773 197
rect 21064 75 21116 127
rect 21130 75 21182 127
rect 21196 75 21248 127
rect 21262 75 21314 127
rect 21328 75 21380 127
rect 21394 75 21446 127
rect 21460 75 21512 127
rect 21526 75 21578 127
rect 21591 75 21643 127
rect 21656 75 21708 127
rect 21721 75 21773 127
rect 13064 -2 13116 50
rect 13128 -2 13180 50
rect 24890 -321 24942 -269
rect 24954 -321 25006 -269
rect 25120 -321 25172 -269
rect 25184 -321 25236 -269
rect 13030 -2255 13082 -2203
rect 13094 -2255 13146 -2203
rect 19791 -2255 19843 -2203
rect 19855 -2255 19907 -2203
rect 20476 -2255 20528 -2203
rect 20540 -2255 20592 -2203
<< metal2 >>
rect 2629 33702 3522 33703
rect 2629 33646 2638 33702
rect 2694 33646 2720 33702
rect 2776 33646 2802 33702
rect 2858 33646 2884 33702
rect 2940 33646 2966 33702
rect 3022 33646 3048 33702
rect 3104 33646 3130 33702
rect 3186 33646 3212 33702
rect 3268 33646 3294 33702
rect 3350 33646 3376 33702
rect 3432 33646 3457 33702
rect 3513 33646 3522 33702
rect 2629 33592 3522 33646
rect 2629 33536 2638 33592
rect 2694 33536 2720 33592
rect 2776 33536 2802 33592
rect 2858 33536 2884 33592
rect 2940 33536 2966 33592
rect 3022 33536 3048 33592
rect 3104 33536 3130 33592
rect 3186 33536 3212 33592
rect 3268 33536 3294 33592
rect 3350 33536 3376 33592
rect 3432 33536 3457 33592
rect 3513 33536 3522 33592
rect 2629 33482 3522 33536
rect 2629 33426 2638 33482
rect 2694 33426 2720 33482
rect 2776 33426 2802 33482
rect 2858 33426 2884 33482
rect 2940 33426 2966 33482
rect 3022 33426 3048 33482
rect 3104 33426 3130 33482
rect 3186 33426 3212 33482
rect 3268 33426 3294 33482
rect 3350 33426 3376 33482
rect 3432 33426 3457 33482
rect 3513 33426 3522 33482
rect 2629 33425 3522 33426
rect 4377 28824 4386 28880
rect 4442 28824 4471 28880
rect 4527 28824 4555 28880
rect 4611 28824 4639 28880
rect 4695 28824 4723 28880
rect 4779 28824 4807 28880
rect 4863 28824 4891 28880
rect 4947 28824 4956 28880
rect 4377 28768 4956 28824
rect 4377 28712 4386 28768
rect 4442 28712 4471 28768
rect 4527 28712 4555 28768
rect 4611 28712 4639 28768
rect 4695 28712 4723 28768
rect 4779 28712 4807 28768
rect 4863 28712 4891 28768
rect 4947 28712 4956 28768
rect 4377 28656 4956 28712
rect 4377 28600 4386 28656
rect 4442 28600 4471 28656
rect 4527 28600 4555 28656
rect 4611 28600 4639 28656
rect 4695 28600 4723 28656
rect 4779 28600 4807 28656
rect 4863 28600 4891 28656
rect 4947 28600 4956 28656
rect 6180 28824 6189 28880
rect 6245 28824 6274 28880
rect 6330 28824 6358 28880
rect 6414 28824 6442 28880
rect 6498 28824 6526 28880
rect 6582 28824 6610 28880
rect 6666 28824 6694 28880
rect 6750 28824 6759 28880
rect 6180 28768 6759 28824
rect 6180 28712 6189 28768
rect 6245 28712 6274 28768
rect 6330 28712 6358 28768
rect 6414 28712 6442 28768
rect 6498 28712 6526 28768
rect 6582 28712 6610 28768
rect 6666 28712 6694 28768
rect 6750 28712 6759 28768
rect 6180 28656 6759 28712
rect 6180 28600 6189 28656
rect 6245 28600 6274 28656
rect 6330 28600 6358 28656
rect 6414 28600 6442 28656
rect 6498 28600 6526 28656
rect 6582 28600 6610 28656
rect 6666 28600 6694 28656
rect 6750 28600 6759 28656
rect 7658 28824 7667 28880
rect 7723 28824 7752 28880
rect 7808 28824 7836 28880
rect 7892 28824 7920 28880
rect 7976 28824 8004 28880
rect 8060 28824 8088 28880
rect 8144 28824 8172 28880
rect 8228 28824 8237 28880
rect 7658 28768 8237 28824
rect 7658 28712 7667 28768
rect 7723 28712 7752 28768
rect 7808 28712 7836 28768
rect 7892 28712 7920 28768
rect 7976 28712 8004 28768
rect 8060 28712 8088 28768
rect 8144 28712 8172 28768
rect 8228 28712 8237 28768
rect 7658 28656 8237 28712
rect 7658 28600 7667 28656
rect 7723 28600 7752 28656
rect 7808 28600 7836 28656
rect 7892 28600 7920 28656
rect 7976 28600 8004 28656
rect 8060 28600 8088 28656
rect 8144 28600 8172 28656
rect 8228 28600 8237 28656
rect 9453 28824 9462 28880
rect 9518 28824 9547 28880
rect 9603 28824 9631 28880
rect 9687 28824 9715 28880
rect 9771 28824 9799 28880
rect 9855 28824 9883 28880
rect 9939 28824 9967 28880
rect 10023 28824 10032 28880
rect 9453 28768 10032 28824
rect 9453 28712 9462 28768
rect 9518 28712 9547 28768
rect 9603 28712 9631 28768
rect 9687 28712 9715 28768
rect 9771 28712 9799 28768
rect 9855 28712 9883 28768
rect 9939 28712 9967 28768
rect 10023 28712 10032 28768
rect 9453 28656 10032 28712
rect 9453 28600 9462 28656
rect 9518 28600 9547 28656
rect 9603 28600 9631 28656
rect 9687 28600 9715 28656
rect 9771 28600 9799 28656
rect 9855 28600 9883 28656
rect 9939 28600 9967 28656
rect 10023 28600 10032 28656
rect 11257 28824 11266 28880
rect 11322 28824 11351 28880
rect 11407 28824 11435 28880
rect 11491 28824 11519 28880
rect 11575 28824 11603 28880
rect 11659 28824 11687 28880
rect 11743 28824 11771 28880
rect 11827 28824 11836 28880
rect 11257 28768 11836 28824
rect 11257 28712 11266 28768
rect 11322 28712 11351 28768
rect 11407 28712 11435 28768
rect 11491 28712 11519 28768
rect 11575 28712 11603 28768
rect 11659 28712 11687 28768
rect 11743 28712 11771 28768
rect 11827 28712 11836 28768
rect 11257 28656 11836 28712
rect 11257 28600 11266 28656
rect 11322 28600 11351 28656
rect 11407 28600 11435 28656
rect 11491 28600 11519 28656
rect 11575 28600 11603 28656
rect 11659 28600 11687 28656
rect 11743 28600 11771 28656
rect 11827 28600 11836 28656
rect 23395 28134 24184 28143
rect 23395 28078 23397 28134
rect 23453 28078 23477 28134
rect 23533 28078 23557 28134
rect 23613 28078 23637 28134
rect 23693 28078 24184 28134
rect 23395 28052 24184 28078
rect 23395 27996 23397 28052
rect 23453 27996 23477 28052
rect 23533 27996 23557 28052
rect 23613 27996 23637 28052
rect 23693 27996 24184 28052
rect 23395 27970 24184 27996
rect 23395 27914 23397 27970
rect 23453 27914 23477 27970
rect 23533 27914 23557 27970
rect 23613 27914 23637 27970
rect 23693 27914 24184 27970
rect 23395 27888 24184 27914
rect 23395 27832 23397 27888
rect 23453 27832 23477 27888
rect 23533 27832 23557 27888
rect 23613 27832 23637 27888
rect 23693 27832 24184 27888
rect 23395 27805 24184 27832
rect 23395 27749 23397 27805
rect 23453 27749 23477 27805
rect 23533 27749 23557 27805
rect 23613 27749 23637 27805
rect 23693 27749 24184 27805
rect 23395 27722 24184 27749
rect 23395 27666 23397 27722
rect 23453 27666 23477 27722
rect 23533 27666 23557 27722
rect 23613 27666 23637 27722
rect 23693 27666 24184 27722
rect 23395 27657 24184 27666
rect 23395 26788 24184 26797
rect 23395 26732 23397 26788
rect 23453 26732 23477 26788
rect 23533 26732 23557 26788
rect 23613 26732 23637 26788
rect 23693 26732 24184 26788
rect 23395 26706 24184 26732
rect 23395 26650 23397 26706
rect 23453 26650 23477 26706
rect 23533 26650 23557 26706
rect 23613 26650 23637 26706
rect 23693 26650 24184 26706
rect 23395 26624 24184 26650
rect 23395 26568 23397 26624
rect 23453 26568 23477 26624
rect 23533 26568 23557 26624
rect 23613 26568 23637 26624
rect 23693 26568 24184 26624
rect 23395 26541 24184 26568
rect 23395 26485 23397 26541
rect 23453 26485 23477 26541
rect 23533 26485 23557 26541
rect 23613 26485 23637 26541
rect 23693 26485 24184 26541
rect 23395 26458 24184 26485
rect 23395 26402 23397 26458
rect 23453 26402 23477 26458
rect 23533 26402 23557 26458
rect 23613 26402 23637 26458
rect 23693 26402 24184 26458
rect 23395 26375 24184 26402
rect 23395 26319 23397 26375
rect 23453 26319 23477 26375
rect 23533 26319 23557 26375
rect 23613 26319 23637 26375
rect 23693 26319 24184 26375
rect 23395 26310 24184 26319
rect 2904 15243 2956 20589
rect 18742 17511 19020 17520
rect 18742 17455 18743 17511
rect 18799 17455 18853 17511
rect 18909 17455 18963 17511
rect 19019 17455 19020 17511
rect 18742 17424 19020 17455
rect 18742 17368 18743 17424
rect 18799 17368 18853 17424
rect 18909 17368 18963 17424
rect 19019 17368 19020 17424
rect 18742 17337 19020 17368
rect 18742 17281 18743 17337
rect 18799 17281 18853 17337
rect 18909 17281 18963 17337
rect 19019 17281 19020 17337
rect 18742 17250 19020 17281
rect 18742 17194 18743 17250
rect 18799 17194 18853 17250
rect 18909 17194 18963 17250
rect 19019 17194 19020 17250
rect 18742 17163 19020 17194
rect 18742 17107 18743 17163
rect 18799 17107 18853 17163
rect 18909 17107 18963 17163
rect 19019 17107 19020 17163
rect 18742 17076 19020 17107
rect 18742 17020 18743 17076
rect 18799 17020 18853 17076
rect 18909 17020 18963 17076
rect 19019 17020 19020 17076
rect 18742 16988 19020 17020
rect 18742 16932 18743 16988
rect 18799 16932 18853 16988
rect 18909 16932 18963 16988
rect 19019 16932 19020 16988
rect 18742 16900 19020 16932
rect 18742 16844 18743 16900
rect 18799 16844 18853 16900
rect 18909 16844 18963 16900
rect 19019 16844 19020 16900
rect 18742 16812 19020 16844
rect 18742 16756 18743 16812
rect 18799 16756 18853 16812
rect 18909 16756 18963 16812
rect 19019 16756 19020 16812
rect 18742 16724 19020 16756
rect 18742 16668 18743 16724
rect 18799 16668 18853 16724
rect 18909 16668 18963 16724
rect 19019 16668 19020 16724
rect 18742 16636 19020 16668
rect 18742 16580 18743 16636
rect 18799 16580 18853 16636
rect 18909 16580 18963 16636
rect 19019 16580 19020 16636
rect 18742 16571 19020 16580
rect 23624 16103 23680 16112
rect 23624 16028 23626 16047
rect 23678 16028 23680 16047
rect 23624 16023 23680 16028
rect 23624 15964 23626 15967
rect 23678 15964 23680 15967
rect 23624 15958 23680 15964
rect 23134 15925 23186 15931
rect 22957 15886 23009 15892
rect 22957 15822 23009 15834
rect 2904 15191 2911 15243
rect 2963 15191 2975 15243
rect 3027 15191 3033 15243
rect 2904 13789 2956 15191
rect 2996 14924 3048 14967
rect 2996 14860 3048 14872
tri 2913 13480 2996 13563 se
rect 2996 13532 3048 14808
rect 3088 14856 3140 14967
rect 22957 14886 23009 15770
rect 23053 15886 23105 15892
rect 23053 15822 23105 15834
rect 23053 14938 23105 15770
rect 23134 15861 23186 15873
rect 23134 15243 23186 15809
tri 23186 15243 23216 15273 sw
rect 23134 15239 23216 15243
tri 23216 15239 23220 15243 sw
tri 23462 15239 23466 15243 se
rect 23466 15239 23472 15243
rect 23134 15191 23472 15239
rect 23524 15191 23536 15243
rect 23588 15191 23594 15243
tri 23105 14938 23143 14976 sw
rect 23053 14916 23179 14938
tri 23053 14892 23077 14916 ne
rect 23077 14892 23179 14916
tri 23009 14886 23015 14892 sw
tri 23077 14886 23083 14892 ne
rect 23083 14886 23179 14892
rect 23231 14886 23243 14938
rect 23295 14886 23301 14938
rect 22957 14862 23015 14886
tri 23015 14862 23039 14886 sw
rect 22957 14858 23039 14862
tri 23039 14858 23043 14862 sw
tri 23339 14858 23343 14862 se
rect 23343 14858 23349 14862
rect 3088 14804 3094 14856
rect 3146 14804 3158 14856
rect 3210 14804 3216 14856
rect 22957 14810 23349 14858
rect 23401 14810 23413 14862
rect 23465 14810 23471 14862
rect 3088 14177 3140 14804
rect 3533 14228 3585 14268
rect 3077 14125 3140 14177
rect 3077 13852 3123 14125
rect 3077 13800 3140 13852
tri 2996 13480 3048 13532 nw
tri 2830 13397 2913 13480 se
tri 2913 13397 2996 13480 nw
tri 2812 13379 2830 13397 se
rect 2830 13379 2895 13397
tri 2895 13379 2913 13397 nw
rect 2812 13233 2864 13379
tri 2864 13348 2895 13379 nw
rect 3088 13175 3140 13800
rect 2536 12352 2588 12430
tri 2803 9407 2852 9456 se
rect 2852 9434 2904 9629
rect 2852 9407 2877 9434
tri 2877 9407 2904 9434 nw
rect 2803 9296 2859 9407
tri 2859 9389 2877 9407 nw
rect 2803 9216 2859 9240
rect 2803 9151 2859 9160
rect 2915 7063 2924 7119
rect 2980 7117 3012 7119
rect 3068 7117 3100 7119
rect 3156 7117 3187 7119
rect 2980 7065 2992 7117
rect 3176 7065 3187 7117
rect 2980 7063 3012 7065
rect 3068 7063 3100 7065
rect 3156 7063 3187 7065
rect 3243 7063 3252 7119
rect 21434 5601 23680 5610
rect 21434 5570 23624 5601
rect 21434 3067 21472 5570
rect 23624 5521 23680 5545
rect 23624 5456 23680 5465
rect 21195 3029 21472 3067
rect 21195 2099 21233 3029
rect 25158 2793 25214 2802
rect 25158 2713 25214 2737
rect 25158 2648 25214 2657
rect 20897 2090 21233 2099
rect 20953 2061 21233 2090
rect 20897 2010 20953 2034
rect 18818 1945 20819 1985
rect 20897 1945 20953 1954
rect 18818 1922 18858 1945
rect 16678 1882 18858 1922
rect 20779 1897 20819 1945
rect 20779 1889 21587 1897
rect 16678 1823 16718 1882
rect 20779 1857 22281 1889
rect 21547 1849 22281 1857
rect 16658 1783 16718 1823
tri 15723 912 15775 964 se
rect 15775 918 16460 964
rect 15775 912 15790 918
tri 15790 912 15796 918 nw
rect 16454 912 16460 918
rect 16512 912 16524 964
rect 16576 912 16582 964
tri 15721 910 15723 912 se
rect 15723 910 15780 912
rect 11544 908 12795 910
rect 11258 831 11264 883
rect 11316 831 11328 883
rect 11380 856 11386 883
tri 11386 856 11413 883 sw
rect 11544 856 11550 908
rect 11602 856 11614 908
rect 11666 902 12795 908
tri 12795 902 12803 910 sw
tri 15713 902 15721 910 se
rect 15721 902 15780 910
tri 15780 902 15790 912 nw
rect 11666 899 15777 902
tri 15777 899 15780 902 nw
rect 11666 887 15765 899
tri 15765 887 15777 899 nw
rect 11666 856 15734 887
tri 15734 856 15765 887 nw
tri 16653 856 16658 861 se
rect 16658 856 16717 1783
rect 22241 1659 22281 1849
rect 24020 1796 25210 1802
rect 24072 1750 25210 1796
rect 24020 1732 24072 1744
rect 25158 1732 25210 1750
rect 23062 1708 23118 1717
rect 22241 1652 23062 1659
rect 24020 1674 24072 1680
rect 22241 1628 23118 1652
rect 22241 1619 23062 1628
rect 22649 1527 22655 1579
rect 22707 1527 22719 1579
rect 22771 1527 22777 1579
rect 23062 1563 23118 1572
tri 22563 1441 22649 1527 se
rect 22649 1441 22667 1527
tri 22667 1441 22753 1527 nw
rect 11380 835 11413 856
tri 11413 835 11434 856 sw
tri 16632 835 16653 856 se
rect 16653 835 16717 856
rect 11380 831 11434 835
tri 11434 831 11438 835 sw
tri 16628 831 16632 835 se
rect 16632 831 16717 835
tri 11346 827 11350 831 ne
rect 11350 827 11438 831
tri 11438 827 11442 831 sw
tri 16624 827 16628 831 se
rect 16628 827 16717 831
tri 11350 791 11386 827 ne
rect 11386 791 16717 827
rect 20897 952 20953 961
rect 20897 887 20953 896
rect 20897 872 20898 887
rect 20950 872 20953 887
rect 20897 807 20953 816
tri 11386 773 11404 791 ne
rect 11404 773 16717 791
tri 14737 285 14775 323 se
rect 14775 285 20725 323
tri 20725 285 20763 323 sw
tri 14727 275 14737 285 se
rect 14737 282 20763 285
rect 14737 275 14795 282
tri 14795 275 14802 282 nw
tri 20686 275 20693 282 ne
rect 20693 275 20763 282
rect 14727 267 14787 275
tri 14787 267 14795 275 nw
tri 20693 267 20701 275 ne
rect 20701 268 20763 275
tri 20763 268 20780 285 sw
rect 20701 267 20780 268
tri 20780 267 20781 268 sw
rect 21058 267 21779 268
tri 14725 75 14727 77 se
rect 14727 75 14777 267
tri 14777 257 14787 267 nw
tri 20701 257 20711 267 ne
rect 20711 257 20781 267
tri 20711 215 20753 257 ne
rect 20753 215 20781 257
tri 20781 215 20833 267 sw
rect 21058 215 21064 267
rect 21116 265 21130 267
rect 21182 265 21196 267
rect 21248 265 21262 267
rect 21314 265 21328 267
rect 21380 265 21394 267
rect 21446 265 21460 267
rect 21512 265 21526 267
rect 21578 265 21591 267
rect 21643 265 21656 267
rect 21708 265 21721 267
rect 21126 215 21130 265
rect 21380 215 21391 265
rect 21447 215 21460 265
rect 21708 215 21711 265
rect 21773 215 21779 267
tri 20753 205 20763 215 ne
rect 20763 205 20833 215
tri 20833 205 20843 215 sw
rect 21058 209 21070 215
rect 21126 209 21151 215
rect 21207 209 21231 215
rect 21287 209 21311 215
rect 21367 209 21391 215
rect 21447 209 21471 215
rect 21527 209 21551 215
rect 21607 209 21631 215
rect 21687 209 21711 215
rect 21767 209 21779 215
tri 20763 197 20771 205 ne
rect 20771 197 20843 205
tri 20843 197 20851 205 sw
rect 21058 197 21779 209
tri 20771 145 20823 197 ne
rect 20823 145 20851 197
tri 20851 145 20903 197 sw
rect 21058 145 21064 197
rect 21116 145 21130 197
rect 21182 145 21196 197
rect 21248 145 21262 197
rect 21314 145 21328 197
rect 21380 145 21394 197
rect 21446 145 21460 197
rect 21512 145 21526 197
rect 21578 145 21591 197
rect 21643 145 21656 197
rect 21708 145 21721 197
rect 21773 145 21779 197
tri 20823 127 20841 145 ne
rect 20841 127 20903 145
tri 20903 127 20921 145 sw
rect 21058 133 21779 145
rect 21058 127 21070 133
rect 21126 127 21151 133
rect 21207 127 21231 133
rect 21287 127 21311 133
rect 21367 127 21391 133
rect 21447 127 21471 133
rect 21527 127 21551 133
rect 21607 127 21631 133
rect 21687 127 21711 133
rect 21767 127 21779 133
tri 20841 125 20843 127 ne
rect 20843 125 20921 127
tri 20921 125 20923 127 sw
tri 20843 77 20891 125 ne
rect 20891 77 20923 125
tri 20891 75 20893 77 ne
rect 20893 75 20923 77
tri 20923 75 20973 125 sw
rect 21058 75 21064 127
rect 21126 77 21130 127
rect 21380 77 21391 127
rect 21447 77 21460 127
rect 21708 77 21711 127
rect 21116 75 21130 77
rect 21182 75 21196 77
rect 21248 75 21262 77
rect 21314 75 21328 77
rect 21380 75 21394 77
rect 21446 75 21460 77
rect 21512 75 21526 77
rect 21578 75 21591 77
rect 21643 75 21656 77
rect 21708 75 21721 77
rect 21773 75 21779 127
tri 14700 50 14725 75 se
rect 14725 53 14777 75
tri 20893 53 20915 75 ne
rect 20915 74 20973 75
tri 20973 74 20974 75 sw
rect 21058 74 21779 75
tri 22561 74 22563 76 se
rect 22563 74 22607 1441
tri 22607 1381 22667 1441 nw
rect 20915 53 20974 74
rect 14725 50 14774 53
tri 14774 50 14777 53 nw
tri 20915 50 20918 53 ne
rect 20918 50 20974 53
tri 20974 50 20998 74 sw
tri 22537 50 22561 74 se
rect 22561 50 22607 74
rect 13058 -2 13064 50
rect 13116 -2 13128 50
rect 13180 45 14769 50
tri 14769 45 14774 50 nw
tri 20918 45 20923 50 ne
rect 20923 45 20998 50
tri 20998 45 21003 50 sw
tri 22532 45 22537 50 se
rect 22537 45 22607 50
rect 13180 -2 14722 45
tri 14722 -2 14769 45 nw
tri 20923 4 20964 45 ne
rect 20964 4 22607 45
rect 13100 -269 13141 -114
tri 13141 -269 13183 -227 sw
rect 13100 -277 13183 -269
tri 13183 -277 13191 -269 sw
rect 13100 -405 13189 -277
rect 24884 -321 24890 -269
rect 24942 -321 24954 -269
rect 25006 -321 25012 -269
rect 25114 -321 25120 -269
rect 25172 -321 25184 -269
rect 25236 -321 25242 -269
tri 13066 -2203 13100 -2169 se
rect 13100 -2203 13152 -405
tri 13152 -439 13186 -405 nw
tri 24850 -2043 24884 -2009 se
rect 24884 -2043 24936 -321
tri 24936 -355 24970 -321 nw
rect 20470 -2203 20598 -2095
rect 13024 -2255 13030 -2203
rect 13082 -2255 13094 -2203
rect 13146 -2255 13152 -2203
rect 19785 -2255 19791 -2203
rect 19843 -2255 19855 -2203
rect 19907 -2255 19913 -2203
rect 20470 -2255 20476 -2203
rect 20528 -2255 20540 -2203
rect 20592 -2255 20598 -2203
<< via2 >>
rect 2638 33646 2694 33702
rect 2720 33646 2776 33702
rect 2802 33646 2858 33702
rect 2884 33646 2940 33702
rect 2966 33646 3022 33702
rect 3048 33646 3104 33702
rect 3130 33646 3186 33702
rect 3212 33646 3268 33702
rect 3294 33646 3350 33702
rect 3376 33646 3432 33702
rect 3457 33646 3513 33702
rect 2638 33536 2694 33592
rect 2720 33536 2776 33592
rect 2802 33536 2858 33592
rect 2884 33536 2940 33592
rect 2966 33536 3022 33592
rect 3048 33536 3104 33592
rect 3130 33536 3186 33592
rect 3212 33536 3268 33592
rect 3294 33536 3350 33592
rect 3376 33536 3432 33592
rect 3457 33536 3513 33592
rect 2638 33426 2694 33482
rect 2720 33426 2776 33482
rect 2802 33426 2858 33482
rect 2884 33426 2940 33482
rect 2966 33426 3022 33482
rect 3048 33426 3104 33482
rect 3130 33426 3186 33482
rect 3212 33426 3268 33482
rect 3294 33426 3350 33482
rect 3376 33426 3432 33482
rect 3457 33426 3513 33482
rect 4386 28824 4442 28880
rect 4471 28824 4527 28880
rect 4555 28824 4611 28880
rect 4639 28824 4695 28880
rect 4723 28824 4779 28880
rect 4807 28824 4863 28880
rect 4891 28824 4947 28880
rect 4386 28712 4442 28768
rect 4471 28712 4527 28768
rect 4555 28712 4611 28768
rect 4639 28712 4695 28768
rect 4723 28712 4779 28768
rect 4807 28712 4863 28768
rect 4891 28712 4947 28768
rect 4386 28600 4442 28656
rect 4471 28600 4527 28656
rect 4555 28600 4611 28656
rect 4639 28600 4695 28656
rect 4723 28600 4779 28656
rect 4807 28600 4863 28656
rect 4891 28600 4947 28656
rect 6189 28824 6245 28880
rect 6274 28824 6330 28880
rect 6358 28824 6414 28880
rect 6442 28824 6498 28880
rect 6526 28824 6582 28880
rect 6610 28824 6666 28880
rect 6694 28824 6750 28880
rect 6189 28712 6245 28768
rect 6274 28712 6330 28768
rect 6358 28712 6414 28768
rect 6442 28712 6498 28768
rect 6526 28712 6582 28768
rect 6610 28712 6666 28768
rect 6694 28712 6750 28768
rect 6189 28600 6245 28656
rect 6274 28600 6330 28656
rect 6358 28600 6414 28656
rect 6442 28600 6498 28656
rect 6526 28600 6582 28656
rect 6610 28600 6666 28656
rect 6694 28600 6750 28656
rect 7667 28824 7723 28880
rect 7752 28824 7808 28880
rect 7836 28824 7892 28880
rect 7920 28824 7976 28880
rect 8004 28824 8060 28880
rect 8088 28824 8144 28880
rect 8172 28824 8228 28880
rect 7667 28712 7723 28768
rect 7752 28712 7808 28768
rect 7836 28712 7892 28768
rect 7920 28712 7976 28768
rect 8004 28712 8060 28768
rect 8088 28712 8144 28768
rect 8172 28712 8228 28768
rect 7667 28600 7723 28656
rect 7752 28600 7808 28656
rect 7836 28600 7892 28656
rect 7920 28600 7976 28656
rect 8004 28600 8060 28656
rect 8088 28600 8144 28656
rect 8172 28600 8228 28656
rect 9462 28824 9518 28880
rect 9547 28824 9603 28880
rect 9631 28824 9687 28880
rect 9715 28824 9771 28880
rect 9799 28824 9855 28880
rect 9883 28824 9939 28880
rect 9967 28824 10023 28880
rect 9462 28712 9518 28768
rect 9547 28712 9603 28768
rect 9631 28712 9687 28768
rect 9715 28712 9771 28768
rect 9799 28712 9855 28768
rect 9883 28712 9939 28768
rect 9967 28712 10023 28768
rect 9462 28600 9518 28656
rect 9547 28600 9603 28656
rect 9631 28600 9687 28656
rect 9715 28600 9771 28656
rect 9799 28600 9855 28656
rect 9883 28600 9939 28656
rect 9967 28600 10023 28656
rect 11266 28824 11322 28880
rect 11351 28824 11407 28880
rect 11435 28824 11491 28880
rect 11519 28824 11575 28880
rect 11603 28824 11659 28880
rect 11687 28824 11743 28880
rect 11771 28824 11827 28880
rect 11266 28712 11322 28768
rect 11351 28712 11407 28768
rect 11435 28712 11491 28768
rect 11519 28712 11575 28768
rect 11603 28712 11659 28768
rect 11687 28712 11743 28768
rect 11771 28712 11827 28768
rect 11266 28600 11322 28656
rect 11351 28600 11407 28656
rect 11435 28600 11491 28656
rect 11519 28600 11575 28656
rect 11603 28600 11659 28656
rect 11687 28600 11743 28656
rect 11771 28600 11827 28656
rect 23397 28078 23453 28134
rect 23477 28078 23533 28134
rect 23557 28078 23613 28134
rect 23637 28078 23693 28134
rect 23397 27996 23453 28052
rect 23477 27996 23533 28052
rect 23557 27996 23613 28052
rect 23637 27996 23693 28052
rect 23397 27914 23453 27970
rect 23477 27914 23533 27970
rect 23557 27914 23613 27970
rect 23637 27914 23693 27970
rect 23397 27832 23453 27888
rect 23477 27832 23533 27888
rect 23557 27832 23613 27888
rect 23637 27832 23693 27888
rect 23397 27749 23453 27805
rect 23477 27749 23533 27805
rect 23557 27749 23613 27805
rect 23637 27749 23693 27805
rect 23397 27666 23453 27722
rect 23477 27666 23533 27722
rect 23557 27666 23613 27722
rect 23637 27666 23693 27722
rect 23397 26732 23453 26788
rect 23477 26732 23533 26788
rect 23557 26732 23613 26788
rect 23637 26732 23693 26788
rect 23397 26650 23453 26706
rect 23477 26650 23533 26706
rect 23557 26650 23613 26706
rect 23637 26650 23693 26706
rect 23397 26568 23453 26624
rect 23477 26568 23533 26624
rect 23557 26568 23613 26624
rect 23637 26568 23693 26624
rect 23397 26485 23453 26541
rect 23477 26485 23533 26541
rect 23557 26485 23613 26541
rect 23637 26485 23693 26541
rect 23397 26402 23453 26458
rect 23477 26402 23533 26458
rect 23557 26402 23613 26458
rect 23637 26402 23693 26458
rect 23397 26319 23453 26375
rect 23477 26319 23533 26375
rect 23557 26319 23613 26375
rect 23637 26319 23693 26375
rect 18743 17455 18799 17511
rect 18853 17455 18909 17511
rect 18963 17455 19019 17511
rect 18743 17368 18799 17424
rect 18853 17368 18909 17424
rect 18963 17368 19019 17424
rect 18743 17281 18799 17337
rect 18853 17281 18909 17337
rect 18963 17281 19019 17337
rect 18743 17194 18799 17250
rect 18853 17194 18909 17250
rect 18963 17194 19019 17250
rect 18743 17107 18799 17163
rect 18853 17107 18909 17163
rect 18963 17107 19019 17163
rect 18743 17020 18799 17076
rect 18853 17020 18909 17076
rect 18963 17020 19019 17076
rect 18743 16932 18799 16988
rect 18853 16932 18909 16988
rect 18963 16932 19019 16988
rect 18743 16844 18799 16900
rect 18853 16844 18909 16900
rect 18963 16844 19019 16900
rect 18743 16756 18799 16812
rect 18853 16756 18909 16812
rect 18963 16756 19019 16812
rect 18743 16668 18799 16724
rect 18853 16668 18909 16724
rect 18963 16668 19019 16724
rect 18743 16580 18799 16636
rect 18853 16580 18909 16636
rect 18963 16580 19019 16636
rect 23624 16080 23680 16103
rect 23624 16047 23626 16080
rect 23626 16047 23678 16080
rect 23678 16047 23680 16080
rect 23624 16016 23680 16023
rect 23624 15967 23626 16016
rect 23626 15967 23678 16016
rect 23678 15967 23680 16016
rect 2803 9240 2859 9296
rect 2803 9160 2859 9216
rect 2924 7117 2980 7119
rect 3012 7117 3068 7119
rect 3100 7117 3156 7119
rect 3187 7117 3243 7119
rect 2924 7065 2925 7117
rect 2925 7065 2977 7117
rect 2977 7065 2980 7117
rect 3012 7065 3044 7117
rect 3044 7065 3058 7117
rect 3058 7065 3068 7117
rect 3100 7065 3110 7117
rect 3110 7065 3124 7117
rect 3124 7065 3156 7117
rect 3187 7065 3190 7117
rect 3190 7065 3242 7117
rect 3242 7065 3243 7117
rect 2924 7063 2980 7065
rect 3012 7063 3068 7065
rect 3100 7063 3156 7065
rect 3187 7063 3243 7065
rect 23624 5545 23680 5601
rect 23624 5465 23680 5521
rect 25158 2737 25214 2793
rect 25158 2657 25214 2713
rect 20897 2034 20953 2090
rect 20897 1954 20953 2010
rect 23062 1652 23118 1708
rect 23062 1572 23118 1628
rect 20897 951 20953 952
rect 20897 899 20898 951
rect 20898 899 20950 951
rect 20950 899 20953 951
rect 20897 896 20953 899
rect 20897 835 20898 872
rect 20898 835 20950 872
rect 20950 835 20953 872
rect 20897 816 20953 835
rect 21070 215 21116 265
rect 21116 215 21126 265
rect 21151 215 21182 265
rect 21182 215 21196 265
rect 21196 215 21207 265
rect 21231 215 21248 265
rect 21248 215 21262 265
rect 21262 215 21287 265
rect 21311 215 21314 265
rect 21314 215 21328 265
rect 21328 215 21367 265
rect 21391 215 21394 265
rect 21394 215 21446 265
rect 21446 215 21447 265
rect 21471 215 21512 265
rect 21512 215 21526 265
rect 21526 215 21527 265
rect 21551 215 21578 265
rect 21578 215 21591 265
rect 21591 215 21607 265
rect 21631 215 21643 265
rect 21643 215 21656 265
rect 21656 215 21687 265
rect 21711 215 21721 265
rect 21721 215 21767 265
rect 21070 209 21126 215
rect 21151 209 21207 215
rect 21231 209 21287 215
rect 21311 209 21367 215
rect 21391 209 21447 215
rect 21471 209 21527 215
rect 21551 209 21607 215
rect 21631 209 21687 215
rect 21711 209 21767 215
rect 21070 127 21126 133
rect 21151 127 21207 133
rect 21231 127 21287 133
rect 21311 127 21367 133
rect 21391 127 21447 133
rect 21471 127 21527 133
rect 21551 127 21607 133
rect 21631 127 21687 133
rect 21711 127 21767 133
rect 21070 77 21116 127
rect 21116 77 21126 127
rect 21151 77 21182 127
rect 21182 77 21196 127
rect 21196 77 21207 127
rect 21231 77 21248 127
rect 21248 77 21262 127
rect 21262 77 21287 127
rect 21311 77 21314 127
rect 21314 77 21328 127
rect 21328 77 21367 127
rect 21391 77 21394 127
rect 21394 77 21446 127
rect 21446 77 21447 127
rect 21471 77 21512 127
rect 21512 77 21526 127
rect 21526 77 21527 127
rect 21551 77 21578 127
rect 21578 77 21591 127
rect 21591 77 21607 127
rect 21631 77 21643 127
rect 21643 77 21656 127
rect 21656 77 21687 127
rect 21711 77 21721 127
rect 21721 77 21767 127
<< metal3 >>
rect 2627 33702 3523 33708
rect 2627 33646 2638 33702
rect 2694 33646 2720 33702
rect 2776 33646 2802 33702
rect 2858 33646 2884 33702
rect 2940 33646 2966 33702
rect 3022 33646 3048 33702
rect 3104 33646 3130 33702
rect 3186 33646 3212 33702
rect 3268 33646 3294 33702
rect 3350 33646 3376 33702
rect 3432 33646 3457 33702
rect 3513 33646 3523 33702
rect 2627 33592 3523 33646
rect 2627 33536 2638 33592
rect 2694 33536 2720 33592
rect 2776 33536 2802 33592
rect 2858 33536 2884 33592
rect 2940 33536 2966 33592
rect 3022 33536 3048 33592
rect 3104 33536 3130 33592
rect 3186 33536 3212 33592
rect 3268 33536 3294 33592
rect 3350 33536 3376 33592
rect 3432 33536 3457 33592
rect 3513 33536 3523 33592
rect 2627 33482 3523 33536
rect 2627 33426 2638 33482
rect 2694 33426 2720 33482
rect 2776 33426 2802 33482
rect 2858 33426 2884 33482
rect 2940 33426 2966 33482
rect 3022 33426 3048 33482
rect 3104 33426 3130 33482
rect 3186 33426 3212 33482
rect 3268 33426 3294 33482
rect 3350 33426 3376 33482
rect 3432 33426 3457 33482
rect 3513 33426 3523 33482
rect 1189 27807 1249 27867
rect 1309 27806 1369 27866
rect 1429 27806 1489 27866
rect 2174 27784 2228 27844
rect 2627 23589 3523 33426
rect 27651 32483 27999 32585
rect 23395 30012 23695 30018
rect 23459 29948 23513 30012
rect 23577 29948 23631 30012
rect 23395 29929 23695 29948
rect 23459 29865 23513 29929
rect 23577 29865 23631 29929
rect 23395 29846 23695 29865
rect 23459 29782 23513 29846
rect 23577 29782 23631 29846
rect 23395 29763 23695 29782
rect 23459 29699 23513 29763
rect 23577 29699 23631 29763
rect 23395 29680 23695 29699
rect 23459 29616 23513 29680
rect 23577 29616 23631 29680
rect 23395 29597 23695 29616
rect 23459 29533 23513 29597
rect 23577 29533 23631 29597
rect 23395 29514 23695 29533
rect 23459 29450 23513 29514
rect 23577 29450 23631 29514
rect 23395 29431 23695 29450
rect 23459 29367 23513 29431
rect 23577 29367 23631 29431
rect 23395 29348 23695 29367
rect 23459 29284 23513 29348
rect 23577 29284 23631 29348
rect 23395 29265 23695 29284
rect 23459 29201 23513 29265
rect 23577 29201 23631 29265
rect 23395 29182 23695 29201
rect 23459 29118 23513 29182
rect 23577 29118 23631 29182
rect 23395 29098 23695 29118
rect 23459 29034 23513 29098
rect 23577 29034 23631 29098
rect 23395 29014 23695 29034
rect 23459 28950 23513 29014
rect 23577 28950 23631 29014
rect 4381 28880 4952 28885
rect 4381 28824 4386 28880
rect 4442 28824 4471 28880
rect 4527 28824 4555 28880
rect 4611 28824 4639 28880
rect 4695 28824 4723 28880
rect 4779 28824 4807 28880
rect 4863 28824 4891 28880
rect 4947 28824 4952 28880
rect 4381 28768 4952 28824
rect 4381 28712 4386 28768
rect 4442 28712 4471 28768
rect 4527 28712 4555 28768
rect 4611 28712 4639 28768
rect 4695 28712 4723 28768
rect 4779 28712 4807 28768
rect 4863 28712 4891 28768
rect 4947 28712 4952 28768
rect 4381 28656 4952 28712
rect 4381 28600 4386 28656
rect 4442 28600 4471 28656
rect 4527 28600 4555 28656
rect 4611 28600 4639 28656
rect 4695 28600 4723 28656
rect 4779 28600 4807 28656
rect 4863 28600 4891 28656
rect 4947 28600 4952 28656
rect 4381 28595 4952 28600
rect 6184 28880 6755 28885
rect 6184 28824 6189 28880
rect 6245 28824 6274 28880
rect 6330 28824 6358 28880
rect 6414 28824 6442 28880
rect 6498 28824 6526 28880
rect 6582 28824 6610 28880
rect 6666 28824 6694 28880
rect 6750 28824 6755 28880
rect 6184 28768 6755 28824
rect 6184 28712 6189 28768
rect 6245 28712 6274 28768
rect 6330 28712 6358 28768
rect 6414 28712 6442 28768
rect 6498 28712 6526 28768
rect 6582 28712 6610 28768
rect 6666 28712 6694 28768
rect 6750 28712 6755 28768
rect 6184 28656 6755 28712
rect 6184 28600 6189 28656
rect 6245 28600 6274 28656
rect 6330 28600 6358 28656
rect 6414 28600 6442 28656
rect 6498 28600 6526 28656
rect 6582 28600 6610 28656
rect 6666 28600 6694 28656
rect 6750 28600 6755 28656
rect 6184 28595 6755 28600
rect 7662 28880 8233 28885
rect 7662 28824 7667 28880
rect 7723 28824 7752 28880
rect 7808 28824 7836 28880
rect 7892 28824 7920 28880
rect 7976 28824 8004 28880
rect 8060 28824 8088 28880
rect 8144 28824 8172 28880
rect 8228 28824 8233 28880
rect 7662 28768 8233 28824
rect 7662 28712 7667 28768
rect 7723 28712 7752 28768
rect 7808 28712 7836 28768
rect 7892 28712 7920 28768
rect 7976 28712 8004 28768
rect 8060 28712 8088 28768
rect 8144 28712 8172 28768
rect 8228 28712 8233 28768
rect 7662 28656 8233 28712
rect 7662 28600 7667 28656
rect 7723 28600 7752 28656
rect 7808 28600 7836 28656
rect 7892 28600 7920 28656
rect 7976 28600 8004 28656
rect 8060 28600 8088 28656
rect 8144 28600 8172 28656
rect 8228 28600 8233 28656
rect 7662 28595 8233 28600
rect 9457 28880 10028 28885
rect 9457 28824 9462 28880
rect 9518 28824 9547 28880
rect 9603 28824 9631 28880
rect 9687 28824 9715 28880
rect 9771 28824 9799 28880
rect 9855 28824 9883 28880
rect 9939 28824 9967 28880
rect 10023 28824 10028 28880
rect 9457 28768 10028 28824
rect 9457 28712 9462 28768
rect 9518 28712 9547 28768
rect 9603 28712 9631 28768
rect 9687 28712 9715 28768
rect 9771 28712 9799 28768
rect 9855 28712 9883 28768
rect 9939 28712 9967 28768
rect 10023 28712 10028 28768
rect 9457 28656 10028 28712
rect 9457 28600 9462 28656
rect 9518 28600 9547 28656
rect 9603 28600 9631 28656
rect 9687 28600 9715 28656
rect 9771 28600 9799 28656
rect 9855 28600 9883 28656
rect 9939 28600 9967 28656
rect 10023 28600 10028 28656
rect 9457 28595 10028 28600
rect 11261 28880 11832 28885
rect 11261 28824 11266 28880
rect 11322 28824 11351 28880
rect 11407 28824 11435 28880
rect 11491 28824 11519 28880
rect 11575 28824 11603 28880
rect 11659 28824 11687 28880
rect 11743 28824 11771 28880
rect 11827 28824 11832 28880
rect 11261 28768 11832 28824
rect 11261 28712 11266 28768
rect 11322 28712 11351 28768
rect 11407 28712 11435 28768
rect 11491 28712 11519 28768
rect 11575 28712 11603 28768
rect 11659 28712 11687 28768
rect 11743 28712 11771 28768
rect 11827 28712 11832 28768
rect 11261 28656 11832 28712
rect 11261 28600 11266 28656
rect 11322 28600 11351 28656
rect 11407 28600 11435 28656
rect 11491 28600 11519 28656
rect 11575 28600 11603 28656
rect 11659 28600 11687 28656
rect 11743 28600 11771 28656
rect 11827 28600 11832 28656
rect 11261 28595 11832 28600
rect 17953 28367 18013 28427
rect 18098 28362 18158 28422
rect 23395 28143 23695 28950
rect 23390 28134 23700 28143
rect 23390 28078 23397 28134
rect 23453 28078 23477 28134
rect 23533 28078 23557 28134
rect 23613 28078 23637 28134
rect 23693 28078 23700 28134
rect 23390 28052 23700 28078
rect 23390 27996 23397 28052
rect 23453 27996 23477 28052
rect 23533 27996 23557 28052
rect 23613 27996 23637 28052
rect 23693 27996 23700 28052
rect 23390 27970 23700 27996
rect 23390 27914 23397 27970
rect 23453 27914 23477 27970
rect 23533 27914 23557 27970
rect 23613 27914 23637 27970
rect 23693 27914 23700 27970
rect 23390 27888 23700 27914
rect 23390 27832 23397 27888
rect 23453 27832 23477 27888
rect 23533 27832 23557 27888
rect 23613 27832 23637 27888
rect 23693 27832 23700 27888
rect 23390 27805 23700 27832
rect 23390 27749 23397 27805
rect 23453 27749 23477 27805
rect 23533 27749 23557 27805
rect 23613 27749 23637 27805
rect 23693 27749 23700 27805
rect 23390 27722 23700 27749
rect 23390 27666 23397 27722
rect 23453 27666 23477 27722
rect 23533 27666 23557 27722
rect 23613 27666 23637 27722
rect 23693 27666 23700 27722
rect 23390 27657 23700 27666
rect 23395 26797 23695 27657
rect 23390 26788 23700 26797
rect 23390 26732 23397 26788
rect 23453 26732 23477 26788
rect 23533 26732 23557 26788
rect 23613 26732 23637 26788
rect 23693 26732 23700 26788
rect 23390 26706 23700 26732
rect 23390 26650 23397 26706
rect 23453 26650 23477 26706
rect 23533 26650 23557 26706
rect 23613 26650 23637 26706
rect 23693 26650 23700 26706
rect 23390 26624 23700 26650
rect 23390 26568 23397 26624
rect 23453 26568 23477 26624
rect 23533 26568 23557 26624
rect 23613 26568 23637 26624
rect 23693 26568 23700 26624
rect 23390 26541 23700 26568
rect 23390 26485 23397 26541
rect 23453 26485 23477 26541
rect 23533 26485 23557 26541
rect 23613 26485 23637 26541
rect 23693 26485 23700 26541
rect 23390 26458 23700 26485
rect 23390 26402 23397 26458
rect 23453 26402 23477 26458
rect 23533 26402 23557 26458
rect 23613 26402 23637 26458
rect 23693 26402 23700 26458
rect 23390 26375 23700 26402
rect 23390 26319 23397 26375
rect 23453 26319 23477 26375
rect 23533 26319 23557 26375
rect 23613 26319 23637 26375
rect 23693 26319 23700 26375
rect 23390 26310 23700 26319
tri 3523 23589 3840 23906 sw
rect 2627 23250 3840 23589
tri 2627 22933 2944 23250 ne
rect 2742 18488 2775 18511
tri 2775 18488 2798 18511 sw
rect 2742 18445 2798 18488
tri 2798 18445 2841 18488 sw
tri 2747 18394 2798 18445 ne
rect 2798 18422 2841 18445
tri 2841 18422 2864 18445 sw
rect 2798 9296 2864 18422
rect 2798 9240 2803 9296
rect 2859 9240 2864 9296
rect 2798 9216 2864 9240
rect 2798 9160 2803 9216
rect 2859 9160 2864 9216
rect 2798 9151 2864 9160
rect 2944 12745 3840 23250
rect 18737 17511 19055 17527
rect 18737 17455 18743 17511
rect 18799 17455 18853 17511
rect 18909 17455 18963 17511
rect 19019 17455 19055 17511
rect 18737 17424 19055 17455
rect 18737 17368 18743 17424
rect 18799 17368 18853 17424
rect 18909 17368 18963 17424
rect 19019 17368 19055 17424
rect 18737 17337 19055 17368
rect 18737 17281 18743 17337
rect 18799 17281 18853 17337
rect 18909 17281 18963 17337
rect 19019 17281 19055 17337
rect 18737 17250 19055 17281
rect 18737 17194 18743 17250
rect 18799 17194 18853 17250
rect 18909 17194 18963 17250
rect 19019 17194 19055 17250
rect 18737 17163 19055 17194
rect 18737 17107 18743 17163
rect 18799 17107 18853 17163
rect 18909 17107 18963 17163
rect 19019 17107 19055 17163
rect 18737 17076 19055 17107
rect 18737 17020 18743 17076
rect 18799 17020 18853 17076
rect 18909 17020 18963 17076
rect 19019 17020 19055 17076
rect 18737 16988 19055 17020
rect 18737 16932 18743 16988
rect 18799 16932 18853 16988
rect 18909 16932 18963 16988
rect 19019 16932 19055 16988
rect 18737 16900 19055 16932
rect 18737 16844 18743 16900
rect 18799 16844 18853 16900
rect 18909 16844 18963 16900
rect 19019 16844 19055 16900
rect 18737 16812 19055 16844
rect 18737 16756 18743 16812
rect 18799 16756 18853 16812
rect 18909 16756 18963 16812
rect 19019 16756 19055 16812
rect 18737 16724 19055 16756
rect 18737 16668 18743 16724
rect 18799 16668 18853 16724
rect 18909 16668 18963 16724
rect 19019 16668 19055 16724
rect 18737 16636 19055 16668
rect 18737 16580 18743 16636
rect 18799 16580 18853 16636
rect 18909 16580 18963 16636
rect 19019 16580 19055 16636
tri 18602 15656 18737 15791 se
rect 18737 15656 19055 16580
rect 23619 16103 23685 16108
tri 23052 16047 23067 16062 sw
rect 23619 16047 23624 16103
rect 23680 16047 23685 16103
rect 23052 16035 23067 16047
tri 23067 16035 23079 16047 sw
rect 22929 16023 23079 16035
tri 23079 16023 23091 16035 sw
rect 23619 16023 23685 16047
rect 22929 16001 23091 16023
tri 22929 15967 22963 16001 ne
rect 22963 15967 23091 16001
tri 23091 15967 23147 16023 sw
rect 23619 15967 23624 16023
rect 23680 15967 23685 16023
tri 22963 15937 22993 15967 ne
rect 22993 15937 23147 15967
tri 23147 15937 23177 15967 sw
tri 22993 15878 23052 15937 ne
rect 23052 15878 23177 15937
tri 23052 15873 23057 15878 ne
rect 2944 12681 2965 12745
rect 3029 12681 3053 12745
rect 3117 12681 3141 12745
rect 3205 12681 3229 12745
rect 3293 12681 3317 12745
rect 3381 12681 3405 12745
rect 3469 12681 3493 12745
rect 3557 12681 3581 12745
rect 3645 12681 3669 12745
rect 3733 12681 3757 12745
rect 3821 12681 3840 12745
rect 2944 12665 3840 12681
rect 2944 12601 2965 12665
rect 3029 12601 3053 12665
rect 3117 12601 3141 12665
rect 3205 12601 3229 12665
rect 3293 12601 3317 12665
rect 3381 12601 3405 12665
rect 3469 12601 3493 12665
rect 3557 12601 3581 12665
rect 3645 12601 3669 12665
rect 3733 12601 3757 12665
rect 3821 12601 3840 12665
rect 2944 12585 3840 12601
rect 2944 12521 2965 12585
rect 3029 12521 3053 12585
rect 3117 12521 3141 12585
rect 3205 12521 3229 12585
rect 3293 12521 3317 12585
rect 3381 12521 3405 12585
rect 3469 12521 3493 12585
rect 3557 12521 3581 12585
rect 3645 12521 3669 12585
rect 3733 12521 3757 12585
rect 3821 12521 3840 12585
rect 2944 12505 3840 12521
rect 2944 12441 2965 12505
rect 3029 12441 3053 12505
rect 3117 12441 3141 12505
rect 3205 12441 3229 12505
rect 3293 12441 3317 12505
rect 3381 12441 3405 12505
rect 3469 12441 3493 12505
rect 3557 12441 3581 12505
rect 3645 12441 3669 12505
rect 3733 12441 3757 12505
rect 3821 12441 3840 12505
rect 2944 12425 3840 12441
rect 2944 12361 2965 12425
rect 3029 12361 3053 12425
rect 3117 12361 3141 12425
rect 3205 12361 3229 12425
rect 3293 12361 3317 12425
rect 3381 12361 3405 12425
rect 3469 12361 3493 12425
rect 3557 12361 3581 12425
rect 3645 12361 3669 12425
rect 3733 12361 3757 12425
rect 3821 12361 3840 12425
rect 2944 12345 3840 12361
rect 2944 12281 2965 12345
rect 3029 12281 3053 12345
rect 3117 12281 3141 12345
rect 3205 12281 3229 12345
rect 3293 12281 3317 12345
rect 3381 12281 3405 12345
rect 3469 12281 3493 12345
rect 3557 12281 3581 12345
rect 3645 12281 3669 12345
rect 3733 12281 3757 12345
rect 3821 12281 3840 12345
rect 2944 12265 3840 12281
rect 2944 12201 2965 12265
rect 3029 12201 3053 12265
rect 3117 12201 3141 12265
rect 3205 12201 3229 12265
rect 3293 12201 3317 12265
rect 3381 12201 3405 12265
rect 3469 12201 3493 12265
rect 3557 12201 3581 12265
rect 3645 12201 3669 12265
rect 3733 12201 3757 12265
rect 3821 12201 3840 12265
rect 2944 12185 3840 12201
rect 2944 12121 2965 12185
rect 3029 12121 3053 12185
rect 3117 12121 3141 12185
rect 3205 12121 3229 12185
rect 3293 12121 3317 12185
rect 3381 12121 3405 12185
rect 3469 12121 3493 12185
rect 3557 12121 3581 12185
rect 3645 12121 3669 12185
rect 3733 12121 3757 12185
rect 3821 12121 3840 12185
rect 2944 12105 3840 12121
rect 2944 12041 2965 12105
rect 3029 12041 3053 12105
rect 3117 12041 3141 12105
rect 3205 12041 3229 12105
rect 3293 12041 3317 12105
rect 3381 12041 3405 12105
rect 3469 12041 3493 12105
rect 3557 12041 3581 12105
rect 3645 12041 3669 12105
rect 3733 12041 3757 12105
rect 3821 12041 3840 12105
rect 2944 12025 3840 12041
rect 2944 11961 2965 12025
rect 3029 11961 3053 12025
rect 3117 11961 3141 12025
rect 3205 11961 3229 12025
rect 3293 11961 3317 12025
rect 3381 11961 3405 12025
rect 3469 11961 3493 12025
rect 3557 11961 3581 12025
rect 3645 11961 3669 12025
rect 3733 11961 3757 12025
rect 3821 11961 3840 12025
rect 2944 11945 3840 11961
rect 2944 11881 2965 11945
rect 3029 11881 3053 11945
rect 3117 11881 3141 11945
rect 3205 11881 3229 11945
rect 3293 11881 3317 11945
rect 3381 11881 3405 11945
rect 3469 11881 3493 11945
rect 3557 11881 3581 11945
rect 3645 11881 3669 11945
rect 3733 11881 3757 11945
rect 3821 11881 3840 11945
rect 2944 11865 3840 11881
rect 2944 11801 2965 11865
rect 3029 11801 3053 11865
rect 3117 11801 3141 11865
rect 3205 11801 3229 11865
rect 3293 11801 3317 11865
rect 3381 11801 3405 11865
rect 3469 11801 3493 11865
rect 3557 11801 3581 11865
rect 3645 11801 3669 11865
rect 3733 11801 3757 11865
rect 3821 11801 3840 11865
rect 2944 11785 3840 11801
rect 2944 11721 2965 11785
rect 3029 11721 3053 11785
rect 3117 11721 3141 11785
rect 3205 11721 3229 11785
rect 3293 11721 3317 11785
rect 3381 11721 3405 11785
rect 3469 11721 3493 11785
rect 3557 11721 3581 11785
rect 3645 11721 3669 11785
rect 3733 11721 3757 11785
rect 3821 11721 3840 11785
rect 2944 11705 3840 11721
rect 2944 11641 2965 11705
rect 3029 11641 3053 11705
rect 3117 11641 3141 11705
rect 3205 11641 3229 11705
rect 3293 11641 3317 11705
rect 3381 11641 3405 11705
rect 3469 11641 3493 11705
rect 3557 11641 3581 11705
rect 3645 11641 3669 11705
rect 3733 11641 3757 11705
rect 3821 11641 3840 11705
rect 2944 11625 3840 11641
rect 2944 11561 2965 11625
rect 3029 11561 3053 11625
rect 3117 11561 3141 11625
rect 3205 11561 3229 11625
rect 3293 11561 3317 11625
rect 3381 11561 3405 11625
rect 3469 11561 3493 11625
rect 3557 11561 3581 11625
rect 3645 11561 3669 11625
rect 3733 11561 3757 11625
rect 3821 11561 3840 11625
rect 2944 11545 3840 11561
rect 2944 11481 2965 11545
rect 3029 11481 3053 11545
rect 3117 11481 3141 11545
rect 3205 11481 3229 11545
rect 3293 11481 3317 11545
rect 3381 11481 3405 11545
rect 3469 11481 3493 11545
rect 3557 11481 3581 11545
rect 3645 11481 3669 11545
rect 3733 11481 3757 11545
rect 3821 11481 3840 11545
rect 2944 11465 3840 11481
rect 2944 11401 2965 11465
rect 3029 11401 3053 11465
rect 3117 11401 3141 11465
rect 3205 11401 3229 11465
rect 3293 11401 3317 11465
rect 3381 11401 3405 11465
rect 3469 11401 3493 11465
rect 3557 11401 3581 11465
rect 3645 11401 3669 11465
rect 3733 11401 3757 11465
rect 3821 11401 3840 11465
rect 2944 11385 3840 11401
rect 2944 11321 2965 11385
rect 3029 11321 3053 11385
rect 3117 11321 3141 11385
rect 3205 11321 3229 11385
rect 3293 11321 3317 11385
rect 3381 11321 3405 11385
rect 3469 11321 3493 11385
rect 3557 11321 3581 11385
rect 3645 11321 3669 11385
rect 3733 11321 3757 11385
rect 3821 11321 3840 11385
rect 2944 11305 3840 11321
rect 2944 11241 2965 11305
rect 3029 11241 3053 11305
rect 3117 11241 3141 11305
rect 3205 11241 3229 11305
rect 3293 11241 3317 11305
rect 3381 11241 3405 11305
rect 3469 11241 3493 11305
rect 3557 11241 3581 11305
rect 3645 11241 3669 11305
rect 3733 11241 3757 11305
rect 3821 11241 3840 11305
rect 2944 11225 3840 11241
rect 2944 11161 2965 11225
rect 3029 11161 3053 11225
rect 3117 11161 3141 11225
rect 3205 11161 3229 11225
rect 3293 11161 3317 11225
rect 3381 11161 3405 11225
rect 3469 11161 3493 11225
rect 3557 11161 3581 11225
rect 3645 11161 3669 11225
rect 3733 11161 3757 11225
rect 3821 11161 3840 11225
rect 2944 11145 3840 11161
rect 2944 11081 2965 11145
rect 3029 11081 3053 11145
rect 3117 11081 3141 11145
rect 3205 11081 3229 11145
rect 3293 11081 3317 11145
rect 3381 11081 3405 11145
rect 3469 11081 3493 11145
rect 3557 11081 3581 11145
rect 3645 11081 3669 11145
rect 3733 11081 3757 11145
rect 3821 11081 3840 11145
rect 2944 11065 3840 11081
rect 2944 11001 2965 11065
rect 3029 11001 3053 11065
rect 3117 11001 3141 11065
rect 3205 11001 3229 11065
rect 3293 11001 3317 11065
rect 3381 11001 3405 11065
rect 3469 11001 3493 11065
rect 3557 11001 3581 11065
rect 3645 11001 3669 11065
rect 3733 11001 3757 11065
rect 3821 11001 3840 11065
rect 2944 10985 3840 11001
rect 2944 10921 2965 10985
rect 3029 10921 3053 10985
rect 3117 10921 3141 10985
rect 3205 10921 3229 10985
rect 3293 10921 3317 10985
rect 3381 10921 3405 10985
rect 3469 10921 3493 10985
rect 3557 10921 3581 10985
rect 3645 10921 3669 10985
rect 3733 10921 3757 10985
rect 3821 10921 3840 10985
rect 2944 10905 3840 10921
rect 2944 10841 2965 10905
rect 3029 10841 3053 10905
rect 3117 10841 3141 10905
rect 3205 10841 3229 10905
rect 3293 10841 3317 10905
rect 3381 10841 3405 10905
rect 3469 10841 3493 10905
rect 3557 10841 3581 10905
rect 3645 10841 3669 10905
rect 3733 10841 3757 10905
rect 3821 10841 3840 10905
rect 2944 10825 3840 10841
rect 2944 10761 2965 10825
rect 3029 10761 3053 10825
rect 3117 10761 3141 10825
rect 3205 10761 3229 10825
rect 3293 10761 3317 10825
rect 3381 10761 3405 10825
rect 3469 10761 3493 10825
rect 3557 10761 3581 10825
rect 3645 10761 3669 10825
rect 3733 10761 3757 10825
rect 3821 10761 3840 10825
rect 2944 10745 3840 10761
rect 2944 10681 2965 10745
rect 3029 10681 3053 10745
rect 3117 10681 3141 10745
rect 3205 10681 3229 10745
rect 3293 10681 3317 10745
rect 3381 10681 3405 10745
rect 3469 10681 3493 10745
rect 3557 10681 3581 10745
rect 3645 10681 3669 10745
rect 3733 10681 3757 10745
rect 3821 10681 3840 10745
rect 2944 10665 3840 10681
rect 2944 10601 2965 10665
rect 3029 10601 3053 10665
rect 3117 10601 3141 10665
rect 3205 10601 3229 10665
rect 3293 10601 3317 10665
rect 3381 10601 3405 10665
rect 3469 10601 3493 10665
rect 3557 10601 3581 10665
rect 3645 10601 3669 10665
rect 3733 10601 3757 10665
rect 3821 10601 3840 10665
rect 2944 10585 3840 10601
rect 2944 10521 2965 10585
rect 3029 10521 3053 10585
rect 3117 10521 3141 10585
rect 3205 10521 3229 10585
rect 3293 10521 3317 10585
rect 3381 10521 3405 10585
rect 3469 10521 3493 10585
rect 3557 10521 3581 10585
rect 3645 10521 3669 10585
rect 3733 10521 3757 10585
rect 3821 10521 3840 10585
rect 2944 10505 3840 10521
rect 2944 10441 2965 10505
rect 3029 10441 3053 10505
rect 3117 10441 3141 10505
rect 3205 10441 3229 10505
rect 3293 10441 3317 10505
rect 3381 10441 3405 10505
rect 3469 10441 3493 10505
rect 3557 10441 3581 10505
rect 3645 10441 3669 10505
rect 3733 10441 3757 10505
rect 3821 10441 3840 10505
rect 2944 10425 3840 10441
rect 2944 10361 2965 10425
rect 3029 10361 3053 10425
rect 3117 10361 3141 10425
rect 3205 10361 3229 10425
rect 3293 10361 3317 10425
rect 3381 10361 3405 10425
rect 3469 10361 3493 10425
rect 3557 10361 3581 10425
rect 3645 10361 3669 10425
rect 3733 10361 3757 10425
rect 3821 10361 3840 10425
rect 2944 10345 3840 10361
rect 2944 10281 2965 10345
rect 3029 10281 3053 10345
rect 3117 10281 3141 10345
rect 3205 10281 3229 10345
rect 3293 10281 3317 10345
rect 3381 10281 3405 10345
rect 3469 10281 3493 10345
rect 3557 10281 3581 10345
rect 3645 10281 3669 10345
rect 3733 10281 3757 10345
rect 3821 10281 3840 10345
rect 2944 10265 3840 10281
rect 2944 10201 2965 10265
rect 3029 10201 3053 10265
rect 3117 10201 3141 10265
rect 3205 10201 3229 10265
rect 3293 10201 3317 10265
rect 3381 10201 3405 10265
rect 3469 10201 3493 10265
rect 3557 10201 3581 10265
rect 3645 10201 3669 10265
rect 3733 10201 3757 10265
rect 3821 10201 3840 10265
rect 2944 10185 3840 10201
rect 2944 10121 2965 10185
rect 3029 10121 3053 10185
rect 3117 10121 3141 10185
rect 3205 10121 3229 10185
rect 3293 10121 3317 10185
rect 3381 10121 3405 10185
rect 3469 10121 3493 10185
rect 3557 10121 3581 10185
rect 3645 10121 3669 10185
rect 3733 10121 3757 10185
rect 3821 10121 3840 10185
rect 2944 10105 3840 10121
rect 2944 10041 2965 10105
rect 3029 10041 3053 10105
rect 3117 10041 3141 10105
rect 3205 10041 3229 10105
rect 3293 10041 3317 10105
rect 3381 10041 3405 10105
rect 3469 10041 3493 10105
rect 3557 10041 3581 10105
rect 3645 10041 3669 10105
rect 3733 10041 3757 10105
rect 3821 10041 3840 10105
rect 2944 10025 3840 10041
rect 2944 9961 2965 10025
rect 3029 9961 3053 10025
rect 3117 9961 3141 10025
rect 3205 9961 3229 10025
rect 3293 9961 3317 10025
rect 3381 9961 3405 10025
rect 3469 9961 3493 10025
rect 3557 9961 3581 10025
rect 3645 9961 3669 10025
rect 3733 9961 3757 10025
rect 3821 9961 3840 10025
rect 2944 9945 3840 9961
rect 2944 9881 2965 9945
rect 3029 9881 3053 9945
rect 3117 9881 3141 9945
rect 3205 9881 3229 9945
rect 3293 9881 3317 9945
rect 3381 9881 3405 9945
rect 3469 9881 3493 9945
rect 3557 9881 3581 9945
rect 3645 9881 3669 9945
rect 3733 9881 3757 9945
rect 3821 9881 3840 9945
rect 2944 9865 3840 9881
rect 2944 9801 2965 9865
rect 3029 9801 3053 9865
rect 3117 9801 3141 9865
rect 3205 9801 3229 9865
rect 3293 9801 3317 9865
rect 3381 9801 3405 9865
rect 3469 9801 3493 9865
rect 3557 9801 3581 9865
rect 3645 9801 3669 9865
rect 3733 9801 3757 9865
rect 3821 9801 3840 9865
rect 2944 9785 3840 9801
rect 2944 9721 2965 9785
rect 3029 9721 3053 9785
rect 3117 9721 3141 9785
rect 3205 9721 3229 9785
rect 3293 9721 3317 9785
rect 3381 9721 3405 9785
rect 3469 9721 3493 9785
rect 3557 9721 3581 9785
rect 3645 9721 3669 9785
rect 3733 9721 3757 9785
rect 3821 9721 3840 9785
rect 2944 9705 3840 9721
rect 2944 9641 2965 9705
rect 3029 9641 3053 9705
rect 3117 9641 3141 9705
rect 3205 9641 3229 9705
rect 3293 9641 3317 9705
rect 3381 9641 3405 9705
rect 3469 9641 3493 9705
rect 3557 9641 3581 9705
rect 3645 9641 3669 9705
rect 3733 9641 3757 9705
rect 3821 9641 3840 9705
rect 2944 9625 3840 9641
rect 2944 9561 2965 9625
rect 3029 9561 3053 9625
rect 3117 9561 3141 9625
rect 3205 9561 3229 9625
rect 3293 9561 3317 9625
rect 3381 9561 3405 9625
rect 3469 9561 3493 9625
rect 3557 9561 3581 9625
rect 3645 9561 3669 9625
rect 3733 9561 3757 9625
rect 3821 9561 3840 9625
rect 2944 9545 3840 9561
rect 2944 9481 2965 9545
rect 3029 9481 3053 9545
rect 3117 9481 3141 9545
rect 3205 9481 3229 9545
rect 3293 9481 3317 9545
rect 3381 9481 3405 9545
rect 3469 9481 3493 9545
rect 3557 9481 3581 9545
rect 3645 9481 3669 9545
rect 3733 9481 3757 9545
rect 3821 9481 3840 9545
rect 2944 9465 3840 9481
rect 2944 9401 2965 9465
rect 3029 9401 3053 9465
rect 3117 9401 3141 9465
rect 3205 9401 3229 9465
rect 3293 9401 3317 9465
rect 3381 9401 3405 9465
rect 3469 9401 3493 9465
rect 3557 9401 3581 9465
rect 3645 9401 3669 9465
rect 3733 9401 3757 9465
rect 3821 9401 3840 9465
rect 2944 9385 3840 9401
rect 2944 9321 2965 9385
rect 3029 9321 3053 9385
rect 3117 9321 3141 9385
rect 3205 9321 3229 9385
rect 3293 9321 3317 9385
rect 3381 9321 3405 9385
rect 3469 9321 3493 9385
rect 3557 9321 3581 9385
rect 3645 9321 3669 9385
rect 3733 9321 3757 9385
rect 3821 9321 3840 9385
rect 2944 9305 3840 9321
rect 2944 9241 2965 9305
rect 3029 9241 3053 9305
rect 3117 9241 3141 9305
rect 3205 9241 3229 9305
rect 3293 9241 3317 9305
rect 3381 9241 3405 9305
rect 3469 9241 3493 9305
rect 3557 9241 3581 9305
rect 3645 9241 3669 9305
rect 3733 9241 3757 9305
rect 3821 9241 3840 9305
rect 2944 9225 3840 9241
rect 2944 9161 2965 9225
rect 3029 9161 3053 9225
rect 3117 9161 3141 9225
rect 3205 9161 3229 9225
rect 3293 9161 3317 9225
rect 3381 9161 3405 9225
rect 3469 9161 3493 9225
rect 3557 9161 3581 9225
rect 3645 9161 3669 9225
rect 3733 9161 3757 9225
rect 3821 9161 3840 9225
rect 2944 9145 3840 9161
rect 2944 9081 2965 9145
rect 3029 9081 3053 9145
rect 3117 9081 3141 9145
rect 3205 9081 3229 9145
rect 3293 9081 3317 9145
rect 3381 9081 3405 9145
rect 3469 9081 3493 9145
rect 3557 9081 3581 9145
rect 3645 9081 3669 9145
rect 3733 9081 3757 9145
rect 3821 9081 3840 9145
rect 2944 9065 3840 9081
rect 2944 9001 2965 9065
rect 3029 9001 3053 9065
rect 3117 9001 3141 9065
rect 3205 9001 3229 9065
rect 3293 9001 3317 9065
rect 3381 9001 3405 9065
rect 3469 9001 3493 9065
rect 3557 9001 3581 9065
rect 3645 9001 3669 9065
rect 3733 9001 3757 9065
rect 3821 9001 3840 9065
rect 2944 8985 3840 9001
rect 2944 8921 2965 8985
rect 3029 8921 3053 8985
rect 3117 8921 3141 8985
rect 3205 8921 3229 8985
rect 3293 8921 3317 8985
rect 3381 8921 3405 8985
rect 3469 8921 3493 8985
rect 3557 8921 3581 8985
rect 3645 8921 3669 8985
rect 3733 8921 3757 8985
rect 3821 8921 3840 8985
rect 2944 8904 3840 8921
rect 2944 8840 2965 8904
rect 3029 8840 3053 8904
rect 3117 8840 3141 8904
rect 3205 8840 3229 8904
rect 3293 8840 3317 8904
rect 3381 8840 3405 8904
rect 3469 8840 3493 8904
rect 3557 8840 3581 8904
rect 3645 8840 3669 8904
rect 3733 8840 3757 8904
rect 3821 8840 3840 8904
rect 2944 8823 3840 8840
rect 2944 8759 2965 8823
rect 3029 8759 3053 8823
rect 3117 8759 3141 8823
rect 3205 8759 3229 8823
rect 3293 8759 3317 8823
rect 3381 8759 3405 8823
rect 3469 8759 3493 8823
rect 3557 8759 3581 8823
rect 3645 8759 3669 8823
rect 3733 8759 3757 8823
rect 3821 8759 3840 8823
rect 2944 8742 3840 8759
rect 2944 8678 2965 8742
rect 3029 8678 3053 8742
rect 3117 8678 3141 8742
rect 3205 8678 3229 8742
rect 3293 8678 3317 8742
rect 3381 8678 3405 8742
rect 3469 8678 3493 8742
rect 3557 8678 3581 8742
rect 3645 8678 3669 8742
rect 3733 8678 3757 8742
rect 3821 8678 3840 8742
rect 2944 8661 3840 8678
rect 2944 8597 2965 8661
rect 3029 8597 3053 8661
rect 3117 8597 3141 8661
rect 3205 8597 3229 8661
rect 3293 8597 3317 8661
rect 3381 8597 3405 8661
rect 3469 8597 3493 8661
rect 3557 8597 3581 8661
rect 3645 8597 3669 8661
rect 3733 8597 3757 8661
rect 3821 8597 3840 8661
rect 2944 8580 3840 8597
rect 2944 8516 2965 8580
rect 3029 8516 3053 8580
rect 3117 8516 3141 8580
rect 3205 8516 3229 8580
rect 3293 8516 3317 8580
rect 3381 8516 3405 8580
rect 3469 8516 3493 8580
rect 3557 8516 3581 8580
rect 3645 8516 3669 8580
rect 3733 8516 3757 8580
rect 3821 8516 3840 8580
rect 2944 8499 3840 8516
rect 2944 8435 2965 8499
rect 3029 8435 3053 8499
rect 3117 8435 3141 8499
rect 3205 8435 3229 8499
rect 3293 8435 3317 8499
rect 3381 8435 3405 8499
rect 3469 8435 3493 8499
rect 3557 8435 3581 8499
rect 3645 8435 3669 8499
rect 3733 8435 3757 8499
rect 3821 8435 3840 8499
rect 2944 8418 3840 8435
rect 2944 8354 2965 8418
rect 3029 8354 3053 8418
rect 3117 8354 3141 8418
rect 3205 8354 3229 8418
rect 3293 8354 3317 8418
rect 3381 8354 3405 8418
rect 3469 8354 3493 8418
rect 3557 8354 3581 8418
rect 3645 8354 3669 8418
rect 3733 8354 3757 8418
rect 3821 8354 3840 8418
rect 2944 8337 3840 8354
rect 2944 8273 2965 8337
rect 3029 8273 3053 8337
rect 3117 8273 3141 8337
rect 3205 8273 3229 8337
rect 3293 8273 3317 8337
rect 3381 8273 3405 8337
rect 3469 8273 3493 8337
rect 3557 8273 3581 8337
rect 3645 8273 3669 8337
rect 3733 8273 3757 8337
rect 3821 8273 3840 8337
rect 2944 8256 3840 8273
rect 2944 8192 2965 8256
rect 3029 8192 3053 8256
rect 3117 8192 3141 8256
rect 3205 8192 3229 8256
rect 3293 8192 3317 8256
rect 3381 8192 3405 8256
rect 3469 8192 3493 8256
rect 3557 8192 3581 8256
rect 3645 8192 3669 8256
rect 3733 8192 3757 8256
rect 3821 8192 3840 8256
rect 2944 8175 3840 8192
rect 2944 8111 2965 8175
rect 3029 8111 3053 8175
rect 3117 8111 3141 8175
rect 3205 8111 3229 8175
rect 3293 8111 3317 8175
rect 3381 8111 3405 8175
rect 3469 8111 3493 8175
rect 3557 8111 3581 8175
rect 3645 8111 3669 8175
rect 3733 8111 3757 8175
rect 3821 8111 3840 8175
rect 2944 8094 3840 8111
rect 2944 8030 2965 8094
rect 3029 8030 3053 8094
rect 3117 8030 3141 8094
rect 3205 8030 3229 8094
rect 3293 8030 3317 8094
rect 3381 8030 3405 8094
rect 3469 8030 3493 8094
rect 3557 8030 3581 8094
rect 3645 8030 3669 8094
rect 3733 8030 3757 8094
rect 3821 8030 3840 8094
rect 2944 8013 3840 8030
rect 2944 7949 2965 8013
rect 3029 7949 3053 8013
rect 3117 7949 3141 8013
rect 3205 7949 3229 8013
rect 3293 7949 3317 8013
rect 3381 7949 3405 8013
rect 3469 7949 3493 8013
rect 3557 7949 3581 8013
rect 3645 7949 3669 8013
rect 3733 7949 3757 8013
rect 3821 7949 3840 8013
rect 2944 7932 3840 7949
rect 2944 7868 2965 7932
rect 3029 7868 3053 7932
rect 3117 7868 3141 7932
rect 3205 7868 3229 7932
rect 3293 7868 3317 7932
rect 3381 7868 3405 7932
rect 3469 7868 3493 7932
rect 3557 7868 3581 7932
rect 3645 7868 3669 7932
rect 3733 7868 3757 7932
rect 3821 7868 3840 7932
rect 2944 7851 3840 7868
rect 2944 7787 2965 7851
rect 3029 7787 3053 7851
rect 3117 7787 3141 7851
rect 3205 7787 3229 7851
rect 3293 7787 3317 7851
rect 3381 7787 3405 7851
rect 3469 7787 3493 7851
rect 3557 7787 3581 7851
rect 3645 7787 3669 7851
rect 3733 7787 3757 7851
rect 3821 7787 3840 7851
rect 2944 7773 3840 7787
rect 2919 7119 3248 7124
rect 2919 7063 2924 7119
rect 2980 7063 3012 7119
rect 3068 7063 3100 7119
rect 3156 7063 3187 7119
rect 3243 7063 3248 7119
rect 2919 7058 3248 7063
rect 21051 4437 21940 7202
rect 20892 2090 20958 2095
rect 20892 2034 20897 2090
rect 20953 2034 20958 2090
rect 20892 2010 20958 2034
rect 20892 1954 20897 2010
rect 20953 1954 20958 2010
rect 20892 952 20958 1954
rect 20892 896 20897 952
rect 20953 896 20958 952
rect 20892 872 20958 896
rect 20892 816 20897 872
rect 20953 816 20958 872
rect 20892 811 20958 816
rect 21051 265 21779 4437
tri 21779 4276 21940 4437 nw
rect 23057 1708 23177 15878
rect 23619 5601 23685 15967
rect 23619 5545 23624 5601
rect 23680 5545 23685 5601
rect 23619 5521 23685 5545
rect 23619 5465 23624 5521
rect 23680 5465 23685 5521
rect 23619 5460 23685 5465
rect 27059 2990 27535 2996
rect 27059 2926 27060 2990
rect 27124 2926 27142 2990
rect 27206 2926 27224 2990
rect 27288 2926 27306 2990
rect 27370 2926 27388 2990
rect 27452 2926 27470 2990
rect 27534 2926 27535 2990
rect 27059 2908 27535 2926
rect 27059 2844 27060 2908
rect 27124 2844 27142 2908
rect 27206 2844 27224 2908
rect 27288 2844 27306 2908
rect 27370 2844 27388 2908
rect 27452 2844 27470 2908
rect 27534 2844 27535 2908
rect 27059 2826 27535 2844
rect 25153 2793 25219 2798
rect 25153 2737 25158 2793
rect 25214 2737 25219 2793
rect 25153 2713 25219 2737
rect 25153 2657 25158 2713
rect 25214 2657 25219 2713
rect 25153 2652 25219 2657
rect 27059 2762 27060 2826
rect 27124 2762 27142 2826
rect 27206 2762 27224 2826
rect 27288 2762 27306 2826
rect 27370 2762 27388 2826
rect 27452 2762 27470 2826
rect 27534 2762 27535 2826
rect 27059 2743 27535 2762
rect 27059 2679 27060 2743
rect 27124 2679 27142 2743
rect 27206 2679 27224 2743
rect 27288 2679 27306 2743
rect 27370 2679 27388 2743
rect 27452 2679 27470 2743
rect 27534 2679 27535 2743
rect 27059 2660 27535 2679
rect 27059 2596 27060 2660
rect 27124 2596 27142 2660
rect 27206 2596 27224 2660
rect 27288 2596 27306 2660
rect 27370 2596 27388 2660
rect 27452 2596 27470 2660
rect 27534 2596 27535 2660
rect 27059 2577 27535 2596
rect 27059 2513 27060 2577
rect 27124 2513 27142 2577
rect 27206 2513 27224 2577
rect 27288 2513 27306 2577
rect 27370 2513 27388 2577
rect 27452 2513 27470 2577
rect 27534 2513 27535 2577
rect 27059 2494 27535 2513
rect 27059 2430 27060 2494
rect 27124 2430 27142 2494
rect 27206 2430 27224 2494
rect 27288 2430 27306 2494
rect 27370 2430 27388 2494
rect 27452 2430 27470 2494
rect 27534 2430 27535 2494
rect 27059 2411 27535 2430
rect 27059 2347 27060 2411
rect 27124 2347 27142 2411
rect 27206 2347 27224 2411
rect 27288 2347 27306 2411
rect 27370 2347 27388 2411
rect 27452 2347 27470 2411
rect 27534 2347 27535 2411
rect 27059 2328 27535 2347
rect 27059 2264 27060 2328
rect 27124 2264 27142 2328
rect 27206 2264 27224 2328
rect 27288 2264 27306 2328
rect 27370 2264 27388 2328
rect 27452 2264 27470 2328
rect 27534 2264 27535 2328
rect 27059 2245 27535 2264
rect 27059 2181 27060 2245
rect 27124 2181 27142 2245
rect 27206 2181 27224 2245
rect 27288 2181 27306 2245
rect 27370 2181 27388 2245
rect 27452 2181 27470 2245
rect 27534 2181 27535 2245
rect 27059 2162 27535 2181
rect 27059 2098 27060 2162
rect 27124 2098 27142 2162
rect 27206 2098 27224 2162
rect 27288 2098 27306 2162
rect 27370 2098 27388 2162
rect 27452 2098 27470 2162
rect 27534 2098 27535 2162
rect 27059 2092 27535 2098
rect 23057 1652 23062 1708
rect 23118 1652 23177 1708
rect 23057 1628 23177 1652
rect 23057 1572 23062 1628
rect 23118 1572 23177 1628
rect 23057 1561 23177 1572
rect 21051 209 21070 265
rect 21126 209 21151 265
rect 21207 209 21231 265
rect 21287 209 21311 265
rect 21367 209 21391 265
rect 21447 209 21471 265
rect 21527 209 21551 265
rect 21607 209 21631 265
rect 21687 209 21711 265
rect 21767 209 21779 265
rect 21051 133 21779 209
rect 21051 77 21070 133
rect 21126 77 21151 133
rect 21207 77 21231 133
rect 21287 77 21311 133
rect 21367 77 21391 133
rect 21447 77 21471 133
rect 21527 77 21551 133
rect 21607 77 21631 133
rect 21687 77 21711 133
rect 21767 77 21779 133
rect 21051 70 21779 77
rect 24775 49 24841 118
rect 24901 49 24967 115
rect 25027 43 25093 109
rect 25279 52 25345 127
rect 25153 -269 25219 26
rect 26287 -17 26353 49
rect 26413 -17 26479 49
rect 26539 -17 26605 49
rect 26665 -17 26731 49
rect 26791 -17 26857 49
rect 26917 -17 26983 77
<< via3 >>
rect 23395 29948 23459 30012
rect 23513 29948 23577 30012
rect 23631 29948 23695 30012
rect 23395 29865 23459 29929
rect 23513 29865 23577 29929
rect 23631 29865 23695 29929
rect 23395 29782 23459 29846
rect 23513 29782 23577 29846
rect 23631 29782 23695 29846
rect 23395 29699 23459 29763
rect 23513 29699 23577 29763
rect 23631 29699 23695 29763
rect 23395 29616 23459 29680
rect 23513 29616 23577 29680
rect 23631 29616 23695 29680
rect 23395 29533 23459 29597
rect 23513 29533 23577 29597
rect 23631 29533 23695 29597
rect 23395 29450 23459 29514
rect 23513 29450 23577 29514
rect 23631 29450 23695 29514
rect 23395 29367 23459 29431
rect 23513 29367 23577 29431
rect 23631 29367 23695 29431
rect 23395 29284 23459 29348
rect 23513 29284 23577 29348
rect 23631 29284 23695 29348
rect 23395 29201 23459 29265
rect 23513 29201 23577 29265
rect 23631 29201 23695 29265
rect 23395 29118 23459 29182
rect 23513 29118 23577 29182
rect 23631 29118 23695 29182
rect 23395 29034 23459 29098
rect 23513 29034 23577 29098
rect 23631 29034 23695 29098
rect 23395 28950 23459 29014
rect 23513 28950 23577 29014
rect 23631 28950 23695 29014
rect 2965 12681 3029 12745
rect 3053 12681 3117 12745
rect 3141 12681 3205 12745
rect 3229 12681 3293 12745
rect 3317 12681 3381 12745
rect 3405 12681 3469 12745
rect 3493 12681 3557 12745
rect 3581 12681 3645 12745
rect 3669 12681 3733 12745
rect 3757 12681 3821 12745
rect 2965 12601 3029 12665
rect 3053 12601 3117 12665
rect 3141 12601 3205 12665
rect 3229 12601 3293 12665
rect 3317 12601 3381 12665
rect 3405 12601 3469 12665
rect 3493 12601 3557 12665
rect 3581 12601 3645 12665
rect 3669 12601 3733 12665
rect 3757 12601 3821 12665
rect 2965 12521 3029 12585
rect 3053 12521 3117 12585
rect 3141 12521 3205 12585
rect 3229 12521 3293 12585
rect 3317 12521 3381 12585
rect 3405 12521 3469 12585
rect 3493 12521 3557 12585
rect 3581 12521 3645 12585
rect 3669 12521 3733 12585
rect 3757 12521 3821 12585
rect 2965 12441 3029 12505
rect 3053 12441 3117 12505
rect 3141 12441 3205 12505
rect 3229 12441 3293 12505
rect 3317 12441 3381 12505
rect 3405 12441 3469 12505
rect 3493 12441 3557 12505
rect 3581 12441 3645 12505
rect 3669 12441 3733 12505
rect 3757 12441 3821 12505
rect 2965 12361 3029 12425
rect 3053 12361 3117 12425
rect 3141 12361 3205 12425
rect 3229 12361 3293 12425
rect 3317 12361 3381 12425
rect 3405 12361 3469 12425
rect 3493 12361 3557 12425
rect 3581 12361 3645 12425
rect 3669 12361 3733 12425
rect 3757 12361 3821 12425
rect 2965 12281 3029 12345
rect 3053 12281 3117 12345
rect 3141 12281 3205 12345
rect 3229 12281 3293 12345
rect 3317 12281 3381 12345
rect 3405 12281 3469 12345
rect 3493 12281 3557 12345
rect 3581 12281 3645 12345
rect 3669 12281 3733 12345
rect 3757 12281 3821 12345
rect 2965 12201 3029 12265
rect 3053 12201 3117 12265
rect 3141 12201 3205 12265
rect 3229 12201 3293 12265
rect 3317 12201 3381 12265
rect 3405 12201 3469 12265
rect 3493 12201 3557 12265
rect 3581 12201 3645 12265
rect 3669 12201 3733 12265
rect 3757 12201 3821 12265
rect 2965 12121 3029 12185
rect 3053 12121 3117 12185
rect 3141 12121 3205 12185
rect 3229 12121 3293 12185
rect 3317 12121 3381 12185
rect 3405 12121 3469 12185
rect 3493 12121 3557 12185
rect 3581 12121 3645 12185
rect 3669 12121 3733 12185
rect 3757 12121 3821 12185
rect 2965 12041 3029 12105
rect 3053 12041 3117 12105
rect 3141 12041 3205 12105
rect 3229 12041 3293 12105
rect 3317 12041 3381 12105
rect 3405 12041 3469 12105
rect 3493 12041 3557 12105
rect 3581 12041 3645 12105
rect 3669 12041 3733 12105
rect 3757 12041 3821 12105
rect 2965 11961 3029 12025
rect 3053 11961 3117 12025
rect 3141 11961 3205 12025
rect 3229 11961 3293 12025
rect 3317 11961 3381 12025
rect 3405 11961 3469 12025
rect 3493 11961 3557 12025
rect 3581 11961 3645 12025
rect 3669 11961 3733 12025
rect 3757 11961 3821 12025
rect 2965 11881 3029 11945
rect 3053 11881 3117 11945
rect 3141 11881 3205 11945
rect 3229 11881 3293 11945
rect 3317 11881 3381 11945
rect 3405 11881 3469 11945
rect 3493 11881 3557 11945
rect 3581 11881 3645 11945
rect 3669 11881 3733 11945
rect 3757 11881 3821 11945
rect 2965 11801 3029 11865
rect 3053 11801 3117 11865
rect 3141 11801 3205 11865
rect 3229 11801 3293 11865
rect 3317 11801 3381 11865
rect 3405 11801 3469 11865
rect 3493 11801 3557 11865
rect 3581 11801 3645 11865
rect 3669 11801 3733 11865
rect 3757 11801 3821 11865
rect 2965 11721 3029 11785
rect 3053 11721 3117 11785
rect 3141 11721 3205 11785
rect 3229 11721 3293 11785
rect 3317 11721 3381 11785
rect 3405 11721 3469 11785
rect 3493 11721 3557 11785
rect 3581 11721 3645 11785
rect 3669 11721 3733 11785
rect 3757 11721 3821 11785
rect 2965 11641 3029 11705
rect 3053 11641 3117 11705
rect 3141 11641 3205 11705
rect 3229 11641 3293 11705
rect 3317 11641 3381 11705
rect 3405 11641 3469 11705
rect 3493 11641 3557 11705
rect 3581 11641 3645 11705
rect 3669 11641 3733 11705
rect 3757 11641 3821 11705
rect 2965 11561 3029 11625
rect 3053 11561 3117 11625
rect 3141 11561 3205 11625
rect 3229 11561 3293 11625
rect 3317 11561 3381 11625
rect 3405 11561 3469 11625
rect 3493 11561 3557 11625
rect 3581 11561 3645 11625
rect 3669 11561 3733 11625
rect 3757 11561 3821 11625
rect 2965 11481 3029 11545
rect 3053 11481 3117 11545
rect 3141 11481 3205 11545
rect 3229 11481 3293 11545
rect 3317 11481 3381 11545
rect 3405 11481 3469 11545
rect 3493 11481 3557 11545
rect 3581 11481 3645 11545
rect 3669 11481 3733 11545
rect 3757 11481 3821 11545
rect 2965 11401 3029 11465
rect 3053 11401 3117 11465
rect 3141 11401 3205 11465
rect 3229 11401 3293 11465
rect 3317 11401 3381 11465
rect 3405 11401 3469 11465
rect 3493 11401 3557 11465
rect 3581 11401 3645 11465
rect 3669 11401 3733 11465
rect 3757 11401 3821 11465
rect 2965 11321 3029 11385
rect 3053 11321 3117 11385
rect 3141 11321 3205 11385
rect 3229 11321 3293 11385
rect 3317 11321 3381 11385
rect 3405 11321 3469 11385
rect 3493 11321 3557 11385
rect 3581 11321 3645 11385
rect 3669 11321 3733 11385
rect 3757 11321 3821 11385
rect 2965 11241 3029 11305
rect 3053 11241 3117 11305
rect 3141 11241 3205 11305
rect 3229 11241 3293 11305
rect 3317 11241 3381 11305
rect 3405 11241 3469 11305
rect 3493 11241 3557 11305
rect 3581 11241 3645 11305
rect 3669 11241 3733 11305
rect 3757 11241 3821 11305
rect 2965 11161 3029 11225
rect 3053 11161 3117 11225
rect 3141 11161 3205 11225
rect 3229 11161 3293 11225
rect 3317 11161 3381 11225
rect 3405 11161 3469 11225
rect 3493 11161 3557 11225
rect 3581 11161 3645 11225
rect 3669 11161 3733 11225
rect 3757 11161 3821 11225
rect 2965 11081 3029 11145
rect 3053 11081 3117 11145
rect 3141 11081 3205 11145
rect 3229 11081 3293 11145
rect 3317 11081 3381 11145
rect 3405 11081 3469 11145
rect 3493 11081 3557 11145
rect 3581 11081 3645 11145
rect 3669 11081 3733 11145
rect 3757 11081 3821 11145
rect 2965 11001 3029 11065
rect 3053 11001 3117 11065
rect 3141 11001 3205 11065
rect 3229 11001 3293 11065
rect 3317 11001 3381 11065
rect 3405 11001 3469 11065
rect 3493 11001 3557 11065
rect 3581 11001 3645 11065
rect 3669 11001 3733 11065
rect 3757 11001 3821 11065
rect 2965 10921 3029 10985
rect 3053 10921 3117 10985
rect 3141 10921 3205 10985
rect 3229 10921 3293 10985
rect 3317 10921 3381 10985
rect 3405 10921 3469 10985
rect 3493 10921 3557 10985
rect 3581 10921 3645 10985
rect 3669 10921 3733 10985
rect 3757 10921 3821 10985
rect 2965 10841 3029 10905
rect 3053 10841 3117 10905
rect 3141 10841 3205 10905
rect 3229 10841 3293 10905
rect 3317 10841 3381 10905
rect 3405 10841 3469 10905
rect 3493 10841 3557 10905
rect 3581 10841 3645 10905
rect 3669 10841 3733 10905
rect 3757 10841 3821 10905
rect 2965 10761 3029 10825
rect 3053 10761 3117 10825
rect 3141 10761 3205 10825
rect 3229 10761 3293 10825
rect 3317 10761 3381 10825
rect 3405 10761 3469 10825
rect 3493 10761 3557 10825
rect 3581 10761 3645 10825
rect 3669 10761 3733 10825
rect 3757 10761 3821 10825
rect 2965 10681 3029 10745
rect 3053 10681 3117 10745
rect 3141 10681 3205 10745
rect 3229 10681 3293 10745
rect 3317 10681 3381 10745
rect 3405 10681 3469 10745
rect 3493 10681 3557 10745
rect 3581 10681 3645 10745
rect 3669 10681 3733 10745
rect 3757 10681 3821 10745
rect 2965 10601 3029 10665
rect 3053 10601 3117 10665
rect 3141 10601 3205 10665
rect 3229 10601 3293 10665
rect 3317 10601 3381 10665
rect 3405 10601 3469 10665
rect 3493 10601 3557 10665
rect 3581 10601 3645 10665
rect 3669 10601 3733 10665
rect 3757 10601 3821 10665
rect 2965 10521 3029 10585
rect 3053 10521 3117 10585
rect 3141 10521 3205 10585
rect 3229 10521 3293 10585
rect 3317 10521 3381 10585
rect 3405 10521 3469 10585
rect 3493 10521 3557 10585
rect 3581 10521 3645 10585
rect 3669 10521 3733 10585
rect 3757 10521 3821 10585
rect 2965 10441 3029 10505
rect 3053 10441 3117 10505
rect 3141 10441 3205 10505
rect 3229 10441 3293 10505
rect 3317 10441 3381 10505
rect 3405 10441 3469 10505
rect 3493 10441 3557 10505
rect 3581 10441 3645 10505
rect 3669 10441 3733 10505
rect 3757 10441 3821 10505
rect 2965 10361 3029 10425
rect 3053 10361 3117 10425
rect 3141 10361 3205 10425
rect 3229 10361 3293 10425
rect 3317 10361 3381 10425
rect 3405 10361 3469 10425
rect 3493 10361 3557 10425
rect 3581 10361 3645 10425
rect 3669 10361 3733 10425
rect 3757 10361 3821 10425
rect 2965 10281 3029 10345
rect 3053 10281 3117 10345
rect 3141 10281 3205 10345
rect 3229 10281 3293 10345
rect 3317 10281 3381 10345
rect 3405 10281 3469 10345
rect 3493 10281 3557 10345
rect 3581 10281 3645 10345
rect 3669 10281 3733 10345
rect 3757 10281 3821 10345
rect 2965 10201 3029 10265
rect 3053 10201 3117 10265
rect 3141 10201 3205 10265
rect 3229 10201 3293 10265
rect 3317 10201 3381 10265
rect 3405 10201 3469 10265
rect 3493 10201 3557 10265
rect 3581 10201 3645 10265
rect 3669 10201 3733 10265
rect 3757 10201 3821 10265
rect 2965 10121 3029 10185
rect 3053 10121 3117 10185
rect 3141 10121 3205 10185
rect 3229 10121 3293 10185
rect 3317 10121 3381 10185
rect 3405 10121 3469 10185
rect 3493 10121 3557 10185
rect 3581 10121 3645 10185
rect 3669 10121 3733 10185
rect 3757 10121 3821 10185
rect 2965 10041 3029 10105
rect 3053 10041 3117 10105
rect 3141 10041 3205 10105
rect 3229 10041 3293 10105
rect 3317 10041 3381 10105
rect 3405 10041 3469 10105
rect 3493 10041 3557 10105
rect 3581 10041 3645 10105
rect 3669 10041 3733 10105
rect 3757 10041 3821 10105
rect 2965 9961 3029 10025
rect 3053 9961 3117 10025
rect 3141 9961 3205 10025
rect 3229 9961 3293 10025
rect 3317 9961 3381 10025
rect 3405 9961 3469 10025
rect 3493 9961 3557 10025
rect 3581 9961 3645 10025
rect 3669 9961 3733 10025
rect 3757 9961 3821 10025
rect 2965 9881 3029 9945
rect 3053 9881 3117 9945
rect 3141 9881 3205 9945
rect 3229 9881 3293 9945
rect 3317 9881 3381 9945
rect 3405 9881 3469 9945
rect 3493 9881 3557 9945
rect 3581 9881 3645 9945
rect 3669 9881 3733 9945
rect 3757 9881 3821 9945
rect 2965 9801 3029 9865
rect 3053 9801 3117 9865
rect 3141 9801 3205 9865
rect 3229 9801 3293 9865
rect 3317 9801 3381 9865
rect 3405 9801 3469 9865
rect 3493 9801 3557 9865
rect 3581 9801 3645 9865
rect 3669 9801 3733 9865
rect 3757 9801 3821 9865
rect 2965 9721 3029 9785
rect 3053 9721 3117 9785
rect 3141 9721 3205 9785
rect 3229 9721 3293 9785
rect 3317 9721 3381 9785
rect 3405 9721 3469 9785
rect 3493 9721 3557 9785
rect 3581 9721 3645 9785
rect 3669 9721 3733 9785
rect 3757 9721 3821 9785
rect 2965 9641 3029 9705
rect 3053 9641 3117 9705
rect 3141 9641 3205 9705
rect 3229 9641 3293 9705
rect 3317 9641 3381 9705
rect 3405 9641 3469 9705
rect 3493 9641 3557 9705
rect 3581 9641 3645 9705
rect 3669 9641 3733 9705
rect 3757 9641 3821 9705
rect 2965 9561 3029 9625
rect 3053 9561 3117 9625
rect 3141 9561 3205 9625
rect 3229 9561 3293 9625
rect 3317 9561 3381 9625
rect 3405 9561 3469 9625
rect 3493 9561 3557 9625
rect 3581 9561 3645 9625
rect 3669 9561 3733 9625
rect 3757 9561 3821 9625
rect 2965 9481 3029 9545
rect 3053 9481 3117 9545
rect 3141 9481 3205 9545
rect 3229 9481 3293 9545
rect 3317 9481 3381 9545
rect 3405 9481 3469 9545
rect 3493 9481 3557 9545
rect 3581 9481 3645 9545
rect 3669 9481 3733 9545
rect 3757 9481 3821 9545
rect 2965 9401 3029 9465
rect 3053 9401 3117 9465
rect 3141 9401 3205 9465
rect 3229 9401 3293 9465
rect 3317 9401 3381 9465
rect 3405 9401 3469 9465
rect 3493 9401 3557 9465
rect 3581 9401 3645 9465
rect 3669 9401 3733 9465
rect 3757 9401 3821 9465
rect 2965 9321 3029 9385
rect 3053 9321 3117 9385
rect 3141 9321 3205 9385
rect 3229 9321 3293 9385
rect 3317 9321 3381 9385
rect 3405 9321 3469 9385
rect 3493 9321 3557 9385
rect 3581 9321 3645 9385
rect 3669 9321 3733 9385
rect 3757 9321 3821 9385
rect 2965 9241 3029 9305
rect 3053 9241 3117 9305
rect 3141 9241 3205 9305
rect 3229 9241 3293 9305
rect 3317 9241 3381 9305
rect 3405 9241 3469 9305
rect 3493 9241 3557 9305
rect 3581 9241 3645 9305
rect 3669 9241 3733 9305
rect 3757 9241 3821 9305
rect 2965 9161 3029 9225
rect 3053 9161 3117 9225
rect 3141 9161 3205 9225
rect 3229 9161 3293 9225
rect 3317 9161 3381 9225
rect 3405 9161 3469 9225
rect 3493 9161 3557 9225
rect 3581 9161 3645 9225
rect 3669 9161 3733 9225
rect 3757 9161 3821 9225
rect 2965 9081 3029 9145
rect 3053 9081 3117 9145
rect 3141 9081 3205 9145
rect 3229 9081 3293 9145
rect 3317 9081 3381 9145
rect 3405 9081 3469 9145
rect 3493 9081 3557 9145
rect 3581 9081 3645 9145
rect 3669 9081 3733 9145
rect 3757 9081 3821 9145
rect 2965 9001 3029 9065
rect 3053 9001 3117 9065
rect 3141 9001 3205 9065
rect 3229 9001 3293 9065
rect 3317 9001 3381 9065
rect 3405 9001 3469 9065
rect 3493 9001 3557 9065
rect 3581 9001 3645 9065
rect 3669 9001 3733 9065
rect 3757 9001 3821 9065
rect 2965 8921 3029 8985
rect 3053 8921 3117 8985
rect 3141 8921 3205 8985
rect 3229 8921 3293 8985
rect 3317 8921 3381 8985
rect 3405 8921 3469 8985
rect 3493 8921 3557 8985
rect 3581 8921 3645 8985
rect 3669 8921 3733 8985
rect 3757 8921 3821 8985
rect 2965 8840 3029 8904
rect 3053 8840 3117 8904
rect 3141 8840 3205 8904
rect 3229 8840 3293 8904
rect 3317 8840 3381 8904
rect 3405 8840 3469 8904
rect 3493 8840 3557 8904
rect 3581 8840 3645 8904
rect 3669 8840 3733 8904
rect 3757 8840 3821 8904
rect 2965 8759 3029 8823
rect 3053 8759 3117 8823
rect 3141 8759 3205 8823
rect 3229 8759 3293 8823
rect 3317 8759 3381 8823
rect 3405 8759 3469 8823
rect 3493 8759 3557 8823
rect 3581 8759 3645 8823
rect 3669 8759 3733 8823
rect 3757 8759 3821 8823
rect 2965 8678 3029 8742
rect 3053 8678 3117 8742
rect 3141 8678 3205 8742
rect 3229 8678 3293 8742
rect 3317 8678 3381 8742
rect 3405 8678 3469 8742
rect 3493 8678 3557 8742
rect 3581 8678 3645 8742
rect 3669 8678 3733 8742
rect 3757 8678 3821 8742
rect 2965 8597 3029 8661
rect 3053 8597 3117 8661
rect 3141 8597 3205 8661
rect 3229 8597 3293 8661
rect 3317 8597 3381 8661
rect 3405 8597 3469 8661
rect 3493 8597 3557 8661
rect 3581 8597 3645 8661
rect 3669 8597 3733 8661
rect 3757 8597 3821 8661
rect 2965 8516 3029 8580
rect 3053 8516 3117 8580
rect 3141 8516 3205 8580
rect 3229 8516 3293 8580
rect 3317 8516 3381 8580
rect 3405 8516 3469 8580
rect 3493 8516 3557 8580
rect 3581 8516 3645 8580
rect 3669 8516 3733 8580
rect 3757 8516 3821 8580
rect 2965 8435 3029 8499
rect 3053 8435 3117 8499
rect 3141 8435 3205 8499
rect 3229 8435 3293 8499
rect 3317 8435 3381 8499
rect 3405 8435 3469 8499
rect 3493 8435 3557 8499
rect 3581 8435 3645 8499
rect 3669 8435 3733 8499
rect 3757 8435 3821 8499
rect 2965 8354 3029 8418
rect 3053 8354 3117 8418
rect 3141 8354 3205 8418
rect 3229 8354 3293 8418
rect 3317 8354 3381 8418
rect 3405 8354 3469 8418
rect 3493 8354 3557 8418
rect 3581 8354 3645 8418
rect 3669 8354 3733 8418
rect 3757 8354 3821 8418
rect 2965 8273 3029 8337
rect 3053 8273 3117 8337
rect 3141 8273 3205 8337
rect 3229 8273 3293 8337
rect 3317 8273 3381 8337
rect 3405 8273 3469 8337
rect 3493 8273 3557 8337
rect 3581 8273 3645 8337
rect 3669 8273 3733 8337
rect 3757 8273 3821 8337
rect 2965 8192 3029 8256
rect 3053 8192 3117 8256
rect 3141 8192 3205 8256
rect 3229 8192 3293 8256
rect 3317 8192 3381 8256
rect 3405 8192 3469 8256
rect 3493 8192 3557 8256
rect 3581 8192 3645 8256
rect 3669 8192 3733 8256
rect 3757 8192 3821 8256
rect 2965 8111 3029 8175
rect 3053 8111 3117 8175
rect 3141 8111 3205 8175
rect 3229 8111 3293 8175
rect 3317 8111 3381 8175
rect 3405 8111 3469 8175
rect 3493 8111 3557 8175
rect 3581 8111 3645 8175
rect 3669 8111 3733 8175
rect 3757 8111 3821 8175
rect 2965 8030 3029 8094
rect 3053 8030 3117 8094
rect 3141 8030 3205 8094
rect 3229 8030 3293 8094
rect 3317 8030 3381 8094
rect 3405 8030 3469 8094
rect 3493 8030 3557 8094
rect 3581 8030 3645 8094
rect 3669 8030 3733 8094
rect 3757 8030 3821 8094
rect 2965 7949 3029 8013
rect 3053 7949 3117 8013
rect 3141 7949 3205 8013
rect 3229 7949 3293 8013
rect 3317 7949 3381 8013
rect 3405 7949 3469 8013
rect 3493 7949 3557 8013
rect 3581 7949 3645 8013
rect 3669 7949 3733 8013
rect 3757 7949 3821 8013
rect 2965 7868 3029 7932
rect 3053 7868 3117 7932
rect 3141 7868 3205 7932
rect 3229 7868 3293 7932
rect 3317 7868 3381 7932
rect 3405 7868 3469 7932
rect 3493 7868 3557 7932
rect 3581 7868 3645 7932
rect 3669 7868 3733 7932
rect 3757 7868 3821 7932
rect 2965 7787 3029 7851
rect 3053 7787 3117 7851
rect 3141 7787 3205 7851
rect 3229 7787 3293 7851
rect 3317 7787 3381 7851
rect 3405 7787 3469 7851
rect 3493 7787 3557 7851
rect 3581 7787 3645 7851
rect 3669 7787 3733 7851
rect 3757 7787 3821 7851
rect 27060 2926 27124 2990
rect 27142 2926 27206 2990
rect 27224 2926 27288 2990
rect 27306 2926 27370 2990
rect 27388 2926 27452 2990
rect 27470 2926 27534 2990
rect 27060 2844 27124 2908
rect 27142 2844 27206 2908
rect 27224 2844 27288 2908
rect 27306 2844 27370 2908
rect 27388 2844 27452 2908
rect 27470 2844 27534 2908
rect 27060 2762 27124 2826
rect 27142 2762 27206 2826
rect 27224 2762 27288 2826
rect 27306 2762 27370 2826
rect 27388 2762 27452 2826
rect 27470 2762 27534 2826
rect 27060 2679 27124 2743
rect 27142 2679 27206 2743
rect 27224 2679 27288 2743
rect 27306 2679 27370 2743
rect 27388 2679 27452 2743
rect 27470 2679 27534 2743
rect 27060 2596 27124 2660
rect 27142 2596 27206 2660
rect 27224 2596 27288 2660
rect 27306 2596 27370 2660
rect 27388 2596 27452 2660
rect 27470 2596 27534 2660
rect 27060 2513 27124 2577
rect 27142 2513 27206 2577
rect 27224 2513 27288 2577
rect 27306 2513 27370 2577
rect 27388 2513 27452 2577
rect 27470 2513 27534 2577
rect 27060 2430 27124 2494
rect 27142 2430 27206 2494
rect 27224 2430 27288 2494
rect 27306 2430 27370 2494
rect 27388 2430 27452 2494
rect 27470 2430 27534 2494
rect 27060 2347 27124 2411
rect 27142 2347 27206 2411
rect 27224 2347 27288 2411
rect 27306 2347 27370 2411
rect 27388 2347 27452 2411
rect 27470 2347 27534 2411
rect 27060 2264 27124 2328
rect 27142 2264 27206 2328
rect 27224 2264 27288 2328
rect 27306 2264 27370 2328
rect 27388 2264 27452 2328
rect 27470 2264 27534 2328
rect 27060 2181 27124 2245
rect 27142 2181 27206 2245
rect 27224 2181 27288 2245
rect 27306 2181 27370 2245
rect 27388 2181 27452 2245
rect 27470 2181 27534 2245
rect 27060 2098 27124 2162
rect 27142 2098 27206 2162
rect 27224 2098 27288 2162
rect 27306 2098 27370 2162
rect 27388 2098 27452 2162
rect 27470 2098 27534 2162
<< metal4 >>
rect 6845 30419 7737 31355
rect 23394 30012 23696 30013
rect 23394 29948 23395 30012
rect 23459 29948 23513 30012
rect 23577 29948 23631 30012
rect 23695 29948 23696 30012
rect 23394 29929 23696 29948
rect 23394 29865 23395 29929
rect 23459 29865 23513 29929
rect 23577 29865 23631 29929
rect 23695 29865 23696 29929
rect 23394 29846 23696 29865
rect 23394 29782 23395 29846
rect 23459 29782 23513 29846
rect 23577 29782 23631 29846
rect 23695 29782 23696 29846
rect 23394 29763 23696 29782
rect 23394 29699 23395 29763
rect 23459 29699 23513 29763
rect 23577 29699 23631 29763
rect 23695 29699 23696 29763
rect 23394 29680 23696 29699
rect 23394 29616 23395 29680
rect 23459 29616 23513 29680
rect 23577 29616 23631 29680
rect 23695 29616 23696 29680
rect 23394 29597 23696 29616
rect 23394 29533 23395 29597
rect 23459 29533 23513 29597
rect 23577 29533 23631 29597
rect 23695 29533 23696 29597
rect 23394 29514 23696 29533
rect 23394 29450 23395 29514
rect 23459 29450 23513 29514
rect 23577 29450 23631 29514
rect 23695 29450 23696 29514
rect 23394 29431 23696 29450
rect 23394 29367 23395 29431
rect 23459 29367 23513 29431
rect 23577 29367 23631 29431
rect 23695 29367 23696 29431
rect 23394 29348 23696 29367
rect 23394 29284 23395 29348
rect 23459 29284 23513 29348
rect 23577 29284 23631 29348
rect 23695 29284 23696 29348
rect 23394 29265 23696 29284
rect 23394 29201 23395 29265
rect 23459 29201 23513 29265
rect 23577 29201 23631 29265
rect 23695 29201 23696 29265
rect 23394 29182 23696 29201
rect 23394 29118 23395 29182
rect 23459 29118 23513 29182
rect 23577 29118 23631 29182
rect 23695 29118 23696 29182
rect 23394 29098 23696 29118
rect 23394 29034 23395 29098
rect 23459 29034 23513 29098
rect 23577 29034 23631 29098
rect 23695 29034 23696 29098
rect 23394 29014 23696 29034
rect 23394 28950 23395 29014
rect 23459 28950 23513 29014
rect 23577 28950 23631 29014
rect 23695 28950 23696 29014
rect 23394 28949 23696 28950
rect 12354 14735 12837 15238
rect 2961 12745 3825 12746
rect 2961 12681 2965 12745
rect 3029 12681 3053 12745
rect 3117 12681 3141 12745
rect 3205 12681 3229 12745
rect 3293 12681 3317 12745
rect 3381 12681 3405 12745
rect 3469 12681 3493 12745
rect 3557 12681 3581 12745
rect 3645 12681 3669 12745
rect 3733 12681 3757 12745
rect 3821 12681 3825 12745
rect 2961 12665 3825 12681
rect 2961 12601 2965 12665
rect 3029 12601 3053 12665
rect 3117 12601 3141 12665
rect 3205 12601 3229 12665
rect 3293 12601 3317 12665
rect 3381 12601 3405 12665
rect 3469 12601 3493 12665
rect 3557 12601 3581 12665
rect 3645 12601 3669 12665
rect 3733 12601 3757 12665
rect 3821 12601 3825 12665
rect 2961 12585 3825 12601
rect 2961 12521 2965 12585
rect 3029 12521 3053 12585
rect 3117 12521 3141 12585
rect 3205 12521 3229 12585
rect 3293 12521 3317 12585
rect 3381 12521 3405 12585
rect 3469 12521 3493 12585
rect 3557 12521 3581 12585
rect 3645 12521 3669 12585
rect 3733 12521 3757 12585
rect 3821 12521 3825 12585
rect 2961 12505 3825 12521
rect 2961 12441 2965 12505
rect 3029 12441 3053 12505
rect 3117 12441 3141 12505
rect 3205 12441 3229 12505
rect 3293 12441 3317 12505
rect 3381 12441 3405 12505
rect 3469 12441 3493 12505
rect 3557 12441 3581 12505
rect 3645 12441 3669 12505
rect 3733 12441 3757 12505
rect 3821 12441 3825 12505
rect 2961 12425 3825 12441
rect 2961 12361 2965 12425
rect 3029 12361 3053 12425
rect 3117 12361 3141 12425
rect 3205 12361 3229 12425
rect 3293 12361 3317 12425
rect 3381 12361 3405 12425
rect 3469 12361 3493 12425
rect 3557 12361 3581 12425
rect 3645 12361 3669 12425
rect 3733 12361 3757 12425
rect 3821 12361 3825 12425
rect 2961 12345 3825 12361
rect 2961 12281 2965 12345
rect 3029 12281 3053 12345
rect 3117 12281 3141 12345
rect 3205 12281 3229 12345
rect 3293 12281 3317 12345
rect 3381 12281 3405 12345
rect 3469 12281 3493 12345
rect 3557 12281 3581 12345
rect 3645 12281 3669 12345
rect 3733 12281 3757 12345
rect 3821 12281 3825 12345
rect 2961 12265 3825 12281
rect 2961 12201 2965 12265
rect 3029 12201 3053 12265
rect 3117 12201 3141 12265
rect 3205 12201 3229 12265
rect 3293 12201 3317 12265
rect 3381 12201 3405 12265
rect 3469 12201 3493 12265
rect 3557 12201 3581 12265
rect 3645 12201 3669 12265
rect 3733 12201 3757 12265
rect 3821 12201 3825 12265
rect 2961 12185 3825 12201
rect 2961 12121 2965 12185
rect 3029 12121 3053 12185
rect 3117 12121 3141 12185
rect 3205 12121 3229 12185
rect 3293 12121 3317 12185
rect 3381 12121 3405 12185
rect 3469 12121 3493 12185
rect 3557 12121 3581 12185
rect 3645 12121 3669 12185
rect 3733 12121 3757 12185
rect 3821 12121 3825 12185
rect 2961 12105 3825 12121
rect 2961 12041 2965 12105
rect 3029 12041 3053 12105
rect 3117 12041 3141 12105
rect 3205 12041 3229 12105
rect 3293 12041 3317 12105
rect 3381 12041 3405 12105
rect 3469 12041 3493 12105
rect 3557 12041 3581 12105
rect 3645 12041 3669 12105
rect 3733 12041 3757 12105
rect 3821 12041 3825 12105
rect 2961 12025 3825 12041
rect 2961 11961 2965 12025
rect 3029 11961 3053 12025
rect 3117 11961 3141 12025
rect 3205 11961 3229 12025
rect 3293 11961 3317 12025
rect 3381 11961 3405 12025
rect 3469 11961 3493 12025
rect 3557 11961 3581 12025
rect 3645 11961 3669 12025
rect 3733 11961 3757 12025
rect 3821 11961 3825 12025
rect 2961 11945 3825 11961
rect 2961 11881 2965 11945
rect 3029 11881 3053 11945
rect 3117 11881 3141 11945
rect 3205 11881 3229 11945
rect 3293 11881 3317 11945
rect 3381 11881 3405 11945
rect 3469 11881 3493 11945
rect 3557 11881 3581 11945
rect 3645 11881 3669 11945
rect 3733 11881 3757 11945
rect 3821 11881 3825 11945
rect 2961 11865 3825 11881
rect 2961 11801 2965 11865
rect 3029 11801 3053 11865
rect 3117 11801 3141 11865
rect 3205 11801 3229 11865
rect 3293 11801 3317 11865
rect 3381 11801 3405 11865
rect 3469 11801 3493 11865
rect 3557 11801 3581 11865
rect 3645 11801 3669 11865
rect 3733 11801 3757 11865
rect 3821 11801 3825 11865
rect 2961 11785 3825 11801
rect 2961 11721 2965 11785
rect 3029 11721 3053 11785
rect 3117 11721 3141 11785
rect 3205 11721 3229 11785
rect 3293 11721 3317 11785
rect 3381 11721 3405 11785
rect 3469 11721 3493 11785
rect 3557 11721 3581 11785
rect 3645 11721 3669 11785
rect 3733 11721 3757 11785
rect 3821 11721 3825 11785
rect 2961 11705 3825 11721
rect 2961 11641 2965 11705
rect 3029 11641 3053 11705
rect 3117 11641 3141 11705
rect 3205 11641 3229 11705
rect 3293 11641 3317 11705
rect 3381 11641 3405 11705
rect 3469 11641 3493 11705
rect 3557 11641 3581 11705
rect 3645 11641 3669 11705
rect 3733 11641 3757 11705
rect 3821 11641 3825 11705
rect 2961 11625 3825 11641
rect 2961 11561 2965 11625
rect 3029 11561 3053 11625
rect 3117 11561 3141 11625
rect 3205 11561 3229 11625
rect 3293 11561 3317 11625
rect 3381 11561 3405 11625
rect 3469 11561 3493 11625
rect 3557 11561 3581 11625
rect 3645 11561 3669 11625
rect 3733 11561 3757 11625
rect 3821 11561 3825 11625
rect 2961 11545 3825 11561
rect 2961 11481 2965 11545
rect 3029 11481 3053 11545
rect 3117 11481 3141 11545
rect 3205 11481 3229 11545
rect 3293 11481 3317 11545
rect 3381 11481 3405 11545
rect 3469 11481 3493 11545
rect 3557 11481 3581 11545
rect 3645 11481 3669 11545
rect 3733 11481 3757 11545
rect 3821 11481 3825 11545
rect 2961 11465 3825 11481
rect 2961 11401 2965 11465
rect 3029 11401 3053 11465
rect 3117 11401 3141 11465
rect 3205 11401 3229 11465
rect 3293 11401 3317 11465
rect 3381 11401 3405 11465
rect 3469 11401 3493 11465
rect 3557 11401 3581 11465
rect 3645 11401 3669 11465
rect 3733 11401 3757 11465
rect 3821 11401 3825 11465
rect 2961 11385 3825 11401
rect 2961 11321 2965 11385
rect 3029 11321 3053 11385
rect 3117 11321 3141 11385
rect 3205 11321 3229 11385
rect 3293 11321 3317 11385
rect 3381 11321 3405 11385
rect 3469 11321 3493 11385
rect 3557 11321 3581 11385
rect 3645 11321 3669 11385
rect 3733 11321 3757 11385
rect 3821 11321 3825 11385
rect 2961 11305 3825 11321
rect 2961 11241 2965 11305
rect 3029 11241 3053 11305
rect 3117 11241 3141 11305
rect 3205 11241 3229 11305
rect 3293 11241 3317 11305
rect 3381 11241 3405 11305
rect 3469 11241 3493 11305
rect 3557 11241 3581 11305
rect 3645 11241 3669 11305
rect 3733 11241 3757 11305
rect 3821 11241 3825 11305
rect 2961 11225 3825 11241
rect 2961 11161 2965 11225
rect 3029 11161 3053 11225
rect 3117 11161 3141 11225
rect 3205 11161 3229 11225
rect 3293 11161 3317 11225
rect 3381 11161 3405 11225
rect 3469 11161 3493 11225
rect 3557 11161 3581 11225
rect 3645 11161 3669 11225
rect 3733 11161 3757 11225
rect 3821 11161 3825 11225
rect 2961 11145 3825 11161
rect 2961 11081 2965 11145
rect 3029 11081 3053 11145
rect 3117 11081 3141 11145
rect 3205 11081 3229 11145
rect 3293 11081 3317 11145
rect 3381 11081 3405 11145
rect 3469 11081 3493 11145
rect 3557 11081 3581 11145
rect 3645 11081 3669 11145
rect 3733 11081 3757 11145
rect 3821 11081 3825 11145
rect 2961 11065 3825 11081
rect 2961 11001 2965 11065
rect 3029 11001 3053 11065
rect 3117 11001 3141 11065
rect 3205 11001 3229 11065
rect 3293 11001 3317 11065
rect 3381 11001 3405 11065
rect 3469 11001 3493 11065
rect 3557 11001 3581 11065
rect 3645 11001 3669 11065
rect 3733 11001 3757 11065
rect 3821 11001 3825 11065
rect 2961 10985 3825 11001
rect 2961 10921 2965 10985
rect 3029 10921 3053 10985
rect 3117 10921 3141 10985
rect 3205 10921 3229 10985
rect 3293 10921 3317 10985
rect 3381 10921 3405 10985
rect 3469 10921 3493 10985
rect 3557 10921 3581 10985
rect 3645 10921 3669 10985
rect 3733 10921 3757 10985
rect 3821 10921 3825 10985
rect 2961 10905 3825 10921
rect 2961 10841 2965 10905
rect 3029 10841 3053 10905
rect 3117 10841 3141 10905
rect 3205 10841 3229 10905
rect 3293 10841 3317 10905
rect 3381 10841 3405 10905
rect 3469 10841 3493 10905
rect 3557 10841 3581 10905
rect 3645 10841 3669 10905
rect 3733 10841 3757 10905
rect 3821 10841 3825 10905
rect 2961 10825 3825 10841
rect 2961 10761 2965 10825
rect 3029 10761 3053 10825
rect 3117 10761 3141 10825
rect 3205 10761 3229 10825
rect 3293 10761 3317 10825
rect 3381 10761 3405 10825
rect 3469 10761 3493 10825
rect 3557 10761 3581 10825
rect 3645 10761 3669 10825
rect 3733 10761 3757 10825
rect 3821 10761 3825 10825
rect 2961 10745 3825 10761
rect 2961 10681 2965 10745
rect 3029 10681 3053 10745
rect 3117 10681 3141 10745
rect 3205 10681 3229 10745
rect 3293 10681 3317 10745
rect 3381 10681 3405 10745
rect 3469 10681 3493 10745
rect 3557 10681 3581 10745
rect 3645 10681 3669 10745
rect 3733 10681 3757 10745
rect 3821 10681 3825 10745
rect 2961 10665 3825 10681
rect 2961 10601 2965 10665
rect 3029 10601 3053 10665
rect 3117 10601 3141 10665
rect 3205 10601 3229 10665
rect 3293 10601 3317 10665
rect 3381 10601 3405 10665
rect 3469 10601 3493 10665
rect 3557 10601 3581 10665
rect 3645 10601 3669 10665
rect 3733 10601 3757 10665
rect 3821 10601 3825 10665
rect 2961 10585 3825 10601
rect 2961 10521 2965 10585
rect 3029 10521 3053 10585
rect 3117 10521 3141 10585
rect 3205 10521 3229 10585
rect 3293 10521 3317 10585
rect 3381 10521 3405 10585
rect 3469 10521 3493 10585
rect 3557 10521 3581 10585
rect 3645 10521 3669 10585
rect 3733 10521 3757 10585
rect 3821 10521 3825 10585
rect 2961 10505 3825 10521
rect 2961 10441 2965 10505
rect 3029 10441 3053 10505
rect 3117 10441 3141 10505
rect 3205 10441 3229 10505
rect 3293 10441 3317 10505
rect 3381 10441 3405 10505
rect 3469 10441 3493 10505
rect 3557 10441 3581 10505
rect 3645 10441 3669 10505
rect 3733 10441 3757 10505
rect 3821 10441 3825 10505
rect 2961 10425 3825 10441
rect 2961 10361 2965 10425
rect 3029 10361 3053 10425
rect 3117 10361 3141 10425
rect 3205 10361 3229 10425
rect 3293 10361 3317 10425
rect 3381 10361 3405 10425
rect 3469 10361 3493 10425
rect 3557 10361 3581 10425
rect 3645 10361 3669 10425
rect 3733 10361 3757 10425
rect 3821 10361 3825 10425
rect 2961 10345 3825 10361
rect 2961 10281 2965 10345
rect 3029 10281 3053 10345
rect 3117 10281 3141 10345
rect 3205 10281 3229 10345
rect 3293 10281 3317 10345
rect 3381 10281 3405 10345
rect 3469 10281 3493 10345
rect 3557 10281 3581 10345
rect 3645 10281 3669 10345
rect 3733 10281 3757 10345
rect 3821 10281 3825 10345
rect 2961 10265 3825 10281
rect 2961 10201 2965 10265
rect 3029 10201 3053 10265
rect 3117 10201 3141 10265
rect 3205 10201 3229 10265
rect 3293 10201 3317 10265
rect 3381 10201 3405 10265
rect 3469 10201 3493 10265
rect 3557 10201 3581 10265
rect 3645 10201 3669 10265
rect 3733 10201 3757 10265
rect 3821 10201 3825 10265
rect 2961 10185 3825 10201
rect 2961 10121 2965 10185
rect 3029 10121 3053 10185
rect 3117 10121 3141 10185
rect 3205 10121 3229 10185
rect 3293 10121 3317 10185
rect 3381 10121 3405 10185
rect 3469 10121 3493 10185
rect 3557 10121 3581 10185
rect 3645 10121 3669 10185
rect 3733 10121 3757 10185
rect 3821 10121 3825 10185
rect 2961 10105 3825 10121
rect 2961 10041 2965 10105
rect 3029 10041 3053 10105
rect 3117 10041 3141 10105
rect 3205 10041 3229 10105
rect 3293 10041 3317 10105
rect 3381 10041 3405 10105
rect 3469 10041 3493 10105
rect 3557 10041 3581 10105
rect 3645 10041 3669 10105
rect 3733 10041 3757 10105
rect 3821 10041 3825 10105
rect 2961 10025 3825 10041
rect 2961 9961 2965 10025
rect 3029 9961 3053 10025
rect 3117 9961 3141 10025
rect 3205 9961 3229 10025
rect 3293 9961 3317 10025
rect 3381 9961 3405 10025
rect 3469 9961 3493 10025
rect 3557 9961 3581 10025
rect 3645 9961 3669 10025
rect 3733 9961 3757 10025
rect 3821 9961 3825 10025
rect 2961 9945 3825 9961
rect 2961 9881 2965 9945
rect 3029 9881 3053 9945
rect 3117 9881 3141 9945
rect 3205 9881 3229 9945
rect 3293 9881 3317 9945
rect 3381 9881 3405 9945
rect 3469 9881 3493 9945
rect 3557 9881 3581 9945
rect 3645 9881 3669 9945
rect 3733 9881 3757 9945
rect 3821 9881 3825 9945
rect 2961 9865 3825 9881
rect 2961 9801 2965 9865
rect 3029 9801 3053 9865
rect 3117 9801 3141 9865
rect 3205 9801 3229 9865
rect 3293 9801 3317 9865
rect 3381 9801 3405 9865
rect 3469 9801 3493 9865
rect 3557 9801 3581 9865
rect 3645 9801 3669 9865
rect 3733 9801 3757 9865
rect 3821 9801 3825 9865
rect 2961 9785 3825 9801
rect 2961 9721 2965 9785
rect 3029 9721 3053 9785
rect 3117 9721 3141 9785
rect 3205 9721 3229 9785
rect 3293 9721 3317 9785
rect 3381 9721 3405 9785
rect 3469 9721 3493 9785
rect 3557 9721 3581 9785
rect 3645 9721 3669 9785
rect 3733 9721 3757 9785
rect 3821 9721 3825 9785
rect 2961 9705 3825 9721
rect 2961 9641 2965 9705
rect 3029 9641 3053 9705
rect 3117 9641 3141 9705
rect 3205 9641 3229 9705
rect 3293 9641 3317 9705
rect 3381 9641 3405 9705
rect 3469 9641 3493 9705
rect 3557 9641 3581 9705
rect 3645 9641 3669 9705
rect 3733 9641 3757 9705
rect 3821 9641 3825 9705
rect 2961 9625 3825 9641
rect 16141 9637 17244 10662
rect 2961 9561 2965 9625
rect 3029 9561 3053 9625
rect 3117 9561 3141 9625
rect 3205 9561 3229 9625
rect 3293 9561 3317 9625
rect 3381 9561 3405 9625
rect 3469 9561 3493 9625
rect 3557 9561 3581 9625
rect 3645 9561 3669 9625
rect 3733 9561 3757 9625
rect 3821 9561 3825 9625
rect 2961 9545 3825 9561
rect 2961 9481 2965 9545
rect 3029 9481 3053 9545
rect 3117 9481 3141 9545
rect 3205 9481 3229 9545
rect 3293 9481 3317 9545
rect 3381 9481 3405 9545
rect 3469 9481 3493 9545
rect 3557 9481 3581 9545
rect 3645 9481 3669 9545
rect 3733 9481 3757 9545
rect 3821 9481 3825 9545
rect 2961 9465 3825 9481
rect 2961 9401 2965 9465
rect 3029 9401 3053 9465
rect 3117 9401 3141 9465
rect 3205 9401 3229 9465
rect 3293 9401 3317 9465
rect 3381 9401 3405 9465
rect 3469 9401 3493 9465
rect 3557 9401 3581 9465
rect 3645 9401 3669 9465
rect 3733 9401 3757 9465
rect 3821 9401 3825 9465
rect 2961 9385 3825 9401
rect 2961 9321 2965 9385
rect 3029 9321 3053 9385
rect 3117 9321 3141 9385
rect 3205 9321 3229 9385
rect 3293 9321 3317 9385
rect 3381 9321 3405 9385
rect 3469 9321 3493 9385
rect 3557 9321 3581 9385
rect 3645 9321 3669 9385
rect 3733 9321 3757 9385
rect 3821 9321 3825 9385
rect 2961 9305 3825 9321
rect 2961 9241 2965 9305
rect 3029 9241 3053 9305
rect 3117 9241 3141 9305
rect 3205 9241 3229 9305
rect 3293 9241 3317 9305
rect 3381 9241 3405 9305
rect 3469 9241 3493 9305
rect 3557 9241 3581 9305
rect 3645 9241 3669 9305
rect 3733 9241 3757 9305
rect 3821 9241 3825 9305
rect 2961 9225 3825 9241
rect 2961 9161 2965 9225
rect 3029 9161 3053 9225
rect 3117 9161 3141 9225
rect 3205 9161 3229 9225
rect 3293 9161 3317 9225
rect 3381 9161 3405 9225
rect 3469 9161 3493 9225
rect 3557 9161 3581 9225
rect 3645 9161 3669 9225
rect 3733 9161 3757 9225
rect 3821 9161 3825 9225
rect 2961 9145 3825 9161
rect 2961 9081 2965 9145
rect 3029 9081 3053 9145
rect 3117 9081 3141 9145
rect 3205 9081 3229 9145
rect 3293 9081 3317 9145
rect 3381 9081 3405 9145
rect 3469 9081 3493 9145
rect 3557 9081 3581 9145
rect 3645 9081 3669 9145
rect 3733 9081 3757 9145
rect 3821 9081 3825 9145
rect 2961 9065 3825 9081
rect 2961 9001 2965 9065
rect 3029 9001 3053 9065
rect 3117 9001 3141 9065
rect 3205 9001 3229 9065
rect 3293 9001 3317 9065
rect 3381 9001 3405 9065
rect 3469 9001 3493 9065
rect 3557 9001 3581 9065
rect 3645 9001 3669 9065
rect 3733 9001 3757 9065
rect 3821 9001 3825 9065
rect 2961 8985 3825 9001
rect 2961 8921 2965 8985
rect 3029 8921 3053 8985
rect 3117 8921 3141 8985
rect 3205 8921 3229 8985
rect 3293 8921 3317 8985
rect 3381 8921 3405 8985
rect 3469 8921 3493 8985
rect 3557 8921 3581 8985
rect 3645 8921 3669 8985
rect 3733 8921 3757 8985
rect 3821 8921 3825 8985
rect 2961 8904 3825 8921
rect 2961 8840 2965 8904
rect 3029 8840 3053 8904
rect 3117 8840 3141 8904
rect 3205 8840 3229 8904
rect 3293 8840 3317 8904
rect 3381 8840 3405 8904
rect 3469 8840 3493 8904
rect 3557 8840 3581 8904
rect 3645 8840 3669 8904
rect 3733 8840 3757 8904
rect 3821 8840 3825 8904
rect 2961 8823 3825 8840
rect 2961 8759 2965 8823
rect 3029 8759 3053 8823
rect 3117 8759 3141 8823
rect 3205 8759 3229 8823
rect 3293 8759 3317 8823
rect 3381 8759 3405 8823
rect 3469 8759 3493 8823
rect 3557 8759 3581 8823
rect 3645 8759 3669 8823
rect 3733 8759 3757 8823
rect 3821 8759 3825 8823
rect 2961 8742 3825 8759
rect 2961 8678 2965 8742
rect 3029 8678 3053 8742
rect 3117 8678 3141 8742
rect 3205 8678 3229 8742
rect 3293 8678 3317 8742
rect 3381 8678 3405 8742
rect 3469 8678 3493 8742
rect 3557 8678 3581 8742
rect 3645 8678 3669 8742
rect 3733 8678 3757 8742
rect 3821 8678 3825 8742
rect 2961 8661 3825 8678
rect 2961 8597 2965 8661
rect 3029 8597 3053 8661
rect 3117 8597 3141 8661
rect 3205 8597 3229 8661
rect 3293 8597 3317 8661
rect 3381 8597 3405 8661
rect 3469 8597 3493 8661
rect 3557 8597 3581 8661
rect 3645 8597 3669 8661
rect 3733 8597 3757 8661
rect 3821 8597 3825 8661
rect 2961 8580 3825 8597
rect 2961 8516 2965 8580
rect 3029 8516 3053 8580
rect 3117 8516 3141 8580
rect 3205 8516 3229 8580
rect 3293 8516 3317 8580
rect 3381 8516 3405 8580
rect 3469 8516 3493 8580
rect 3557 8516 3581 8580
rect 3645 8516 3669 8580
rect 3733 8516 3757 8580
rect 3821 8516 3825 8580
rect 2961 8499 3825 8516
rect 2961 8435 2965 8499
rect 3029 8435 3053 8499
rect 3117 8435 3141 8499
rect 3205 8435 3229 8499
rect 3293 8435 3317 8499
rect 3381 8435 3405 8499
rect 3469 8435 3493 8499
rect 3557 8435 3581 8499
rect 3645 8435 3669 8499
rect 3733 8435 3757 8499
rect 3821 8435 3825 8499
rect 2961 8418 3825 8435
rect 2961 8354 2965 8418
rect 3029 8354 3053 8418
rect 3117 8354 3141 8418
rect 3205 8354 3229 8418
rect 3293 8354 3317 8418
rect 3381 8354 3405 8418
rect 3469 8354 3493 8418
rect 3557 8354 3581 8418
rect 3645 8354 3669 8418
rect 3733 8354 3757 8418
rect 3821 8354 3825 8418
rect 2961 8337 3825 8354
rect 2961 8273 2965 8337
rect 3029 8273 3053 8337
rect 3117 8273 3141 8337
rect 3205 8273 3229 8337
rect 3293 8273 3317 8337
rect 3381 8273 3405 8337
rect 3469 8273 3493 8337
rect 3557 8273 3581 8337
rect 3645 8273 3669 8337
rect 3733 8273 3757 8337
rect 3821 8273 3825 8337
rect 2961 8256 3825 8273
rect 2961 8192 2965 8256
rect 3029 8192 3053 8256
rect 3117 8192 3141 8256
rect 3205 8192 3229 8256
rect 3293 8192 3317 8256
rect 3381 8192 3405 8256
rect 3469 8192 3493 8256
rect 3557 8192 3581 8256
rect 3645 8192 3669 8256
rect 3733 8192 3757 8256
rect 3821 8192 3825 8256
rect 2961 8175 3825 8192
rect 2961 8111 2965 8175
rect 3029 8111 3053 8175
rect 3117 8111 3141 8175
rect 3205 8111 3229 8175
rect 3293 8111 3317 8175
rect 3381 8111 3405 8175
rect 3469 8111 3493 8175
rect 3557 8111 3581 8175
rect 3645 8111 3669 8175
rect 3733 8111 3757 8175
rect 3821 8111 3825 8175
rect 2961 8094 3825 8111
rect 2961 8030 2965 8094
rect 3029 8030 3053 8094
rect 3117 8030 3141 8094
rect 3205 8030 3229 8094
rect 3293 8030 3317 8094
rect 3381 8030 3405 8094
rect 3469 8030 3493 8094
rect 3557 8030 3581 8094
rect 3645 8030 3669 8094
rect 3733 8030 3757 8094
rect 3821 8030 3825 8094
rect 2961 8013 3825 8030
rect 2961 7949 2965 8013
rect 3029 7949 3053 8013
rect 3117 7949 3141 8013
rect 3205 7949 3229 8013
rect 3293 7949 3317 8013
rect 3381 7949 3405 8013
rect 3469 7949 3493 8013
rect 3557 7949 3581 8013
rect 3645 7949 3669 8013
rect 3733 7949 3757 8013
rect 3821 7949 3825 8013
rect 2961 7932 3825 7949
rect 2961 7868 2965 7932
rect 3029 7868 3053 7932
rect 3117 7868 3141 7932
rect 3205 7868 3229 7932
rect 3293 7868 3317 7932
rect 3381 7868 3405 7932
rect 3469 7868 3493 7932
rect 3557 7868 3581 7932
rect 3645 7868 3669 7932
rect 3733 7868 3757 7932
rect 3821 7868 3825 7932
rect 2961 7851 3825 7868
rect 2961 7787 2965 7851
rect 3029 7787 3053 7851
rect 3117 7787 3141 7851
rect 3205 7787 3229 7851
rect 3293 7787 3317 7851
rect 3381 7787 3405 7851
rect 3469 7787 3493 7851
rect 3557 7787 3581 7851
rect 3645 7787 3669 7851
rect 3733 7787 3757 7851
rect 3821 7787 3825 7851
rect 2961 7786 3825 7787
rect 27058 2990 27536 2991
rect 27058 2926 27060 2990
rect 27124 2926 27142 2990
rect 27206 2926 27224 2990
rect 27288 2926 27306 2990
rect 27370 2926 27388 2990
rect 27452 2926 27470 2990
rect 27534 2926 27536 2990
rect 27058 2908 27536 2926
rect 27058 2844 27060 2908
rect 27124 2844 27142 2908
rect 27206 2844 27224 2908
rect 27288 2844 27306 2908
rect 27370 2844 27388 2908
rect 27452 2844 27470 2908
rect 27534 2844 27536 2908
rect 27058 2826 27536 2844
rect 27058 2762 27060 2826
rect 27124 2762 27142 2826
rect 27206 2762 27224 2826
rect 27288 2762 27306 2826
rect 27370 2762 27388 2826
rect 27452 2762 27470 2826
rect 27534 2762 27536 2826
rect 27058 2743 27536 2762
rect 27058 2679 27060 2743
rect 27124 2679 27142 2743
rect 27206 2679 27224 2743
rect 27288 2679 27306 2743
rect 27370 2679 27388 2743
rect 27452 2679 27470 2743
rect 27534 2679 27536 2743
rect 27058 2660 27536 2679
rect 27058 2596 27060 2660
rect 27124 2596 27142 2660
rect 27206 2596 27224 2660
rect 27288 2596 27306 2660
rect 27370 2596 27388 2660
rect 27452 2596 27470 2660
rect 27534 2596 27536 2660
rect 27058 2577 27536 2596
rect 27058 2513 27060 2577
rect 27124 2513 27142 2577
rect 27206 2513 27224 2577
rect 27288 2513 27306 2577
rect 27370 2513 27388 2577
rect 27452 2513 27470 2577
rect 27534 2513 27536 2577
rect 27058 2494 27536 2513
rect 27058 2430 27060 2494
rect 27124 2430 27142 2494
rect 27206 2430 27224 2494
rect 27288 2430 27306 2494
rect 27370 2430 27388 2494
rect 27452 2430 27470 2494
rect 27534 2430 27536 2494
rect 27058 2411 27536 2430
rect 27058 2347 27060 2411
rect 27124 2347 27142 2411
rect 27206 2347 27224 2411
rect 27288 2347 27306 2411
rect 27370 2347 27388 2411
rect 27452 2347 27470 2411
rect 27534 2347 27536 2411
rect 27058 2328 27536 2347
rect 27058 2264 27060 2328
rect 27124 2264 27142 2328
rect 27206 2264 27224 2328
rect 27288 2264 27306 2328
rect 27370 2264 27388 2328
rect 27452 2264 27470 2328
rect 27534 2264 27536 2328
rect 27058 2245 27536 2264
rect 27058 2181 27060 2245
rect 27124 2181 27142 2245
rect 27206 2181 27224 2245
rect 27288 2181 27306 2245
rect 27370 2181 27388 2245
rect 27452 2181 27470 2245
rect 27534 2181 27536 2245
rect 27058 2162 27536 2181
rect 27058 2098 27060 2162
rect 27124 2098 27142 2162
rect 27206 2098 27224 2162
rect 27288 2098 27306 2162
rect 27370 2098 27388 2162
rect 27452 2098 27470 2162
rect 27534 2098 27536 2162
rect 27058 2097 27536 2098
use sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix_0
timestamp 1648127584
transform 1 0 0 0 1 0
box 206 -5849 28170 33916
use sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix_0
timestamp 1648127584
transform 1 0 1013 0 1 6483
box -877 -6624 27197 26120
<< labels >>
flabel metal4 s 16141 9637 17244 10662 3 FreeSans 200 0 0 0 VDDIO
port 1 nsew
flabel metal4 s 6845 30419 7737 31355 3 FreeSans 200 0 0 0 VSSIO
port 2 nsew
flabel metal4 s 12354 14735 12837 15238 3 FreeSans 200 0 0 0 PAD
port 3 nsew
flabel metal3 s 26917 -17 26983 77 3 FreeSans 200 90 0 0 DM_H[0]
port 4 nsew
flabel metal3 s 26791 -17 26857 49 3 FreeSans 200 90 0 0 DM_H[1]
port 5 nsew
flabel metal3 s 26665 -17 26731 49 3 FreeSans 200 90 0 0 DM_H[2]
port 6 nsew
flabel metal3 s 26539 -17 26605 49 3 FreeSans 200 90 0 0 DM_H_N[0]
port 7 nsew
flabel metal3 s 26413 -17 26479 49 3 FreeSans 200 90 0 0 DM_H_N[1]
port 8 nsew
flabel metal3 s 26287 -17 26353 49 3 FreeSans 200 90 0 0 DM_H_N[2]
port 9 nsew
flabel metal3 s 25279 52 25345 127 3 FreeSans 200 0 0 0 HLD_I_H_N
port 10 nsew
flabel metal3 s 24901 49 24967 115 3 FreeSans 200 90 0 0 OE_N
port 11 nsew
flabel metal3 s 24775 49 24841 118 3 FreeSans 200 90 0 0 OUT
port 12 nsew
flabel metal3 s 2174 27784 2228 27844 3 FreeSans 200 90 0 0 SLEW_CTL_H[0]
port 13 nsew
flabel metal3 s 1429 27806 1489 27866 3 FreeSans 200 90 0 0 SLEW_CTL_H[1]
port 14 nsew
flabel metal3 s 1309 27806 1369 27866 3 FreeSans 200 90 0 0 SLEW_CTL_H_N[0]
port 15 nsew
flabel metal3 s 1189 27807 1249 27867 3 FreeSans 200 90 0 0 SLEW_CTL_H_N[1]
port 16 nsew
flabel metal3 s 25027 43 25093 109 3 FreeSans 200 90 0 0 SLOW
port 17 nsew
flabel metal3 s 27651 32483 27999 32585 3 FreeSans 200 0 0 0 VCCD
port 18 nsew
flabel metal3 s 17953 28367 18013 28427 3 FreeSans 520 90 0 0 NGA_PAD_VPMP_H
port 19 nsew
flabel metal3 s 18098 28362 18158 28422 3 FreeSans 520 90 0 0 NGB_PAD_VPMP_H
port 20 nsew
flabel metal2 s 2536 12352 2588 12430 3 FreeSans 200 0 0 0 PU_CSD_H
port 21 nsew
flabel metal2 s 3533 14228 3585 14268 3 FreeSans 200 0 0 0 PGHS_H
port 22 nsew
flabel metal1 s 23083 1691 23154 1780 3 FreeSans 200 0 0 0 HLD_I_OVR_H
port 23 nsew
flabel metal1 s 12691 771 12752 803 3 FreeSans 200 0 0 0 OD_I_H_N
port 24 nsew
flabel metal1 s 4286 26662 4411 26737 3 FreeSans 200 0 0 0 PD_CSD_H
port 25 nsew
flabel metal1 s 22371 1902 22619 2181 3 FreeSans 200 0 0 0 VPWR_KA
port 26 nsew
flabel metal1 s 1982 7609 2123 7747 3 FreeSans 200 0 0 0 VSSD
port 27 nsew
flabel metal1 s 6437 17954 6539 18043 3 FreeSans 200 0 0 0 VSSIO_AMX
port 28 nsew
flabel metal1 s 25592 15812 25711 15930 3 FreeSans 200 0 0 0 TIE_HI_ESD
port 29 nsew
flabel metal1 s 18580 27001 18626 27046 3 FreeSans 200 90 0 0 TIE_LO_ESD
port 30 nsew
flabel metal1 s 10043 14120 10107 14152 3 FreeSans 200 0 0 0 PUG_H[5]
port 31 nsew
flabel metal1 s 8397 13471 8437 13503 3 FreeSans 200 0 0 0 PUG_H[6]
port 32 nsew
flabel metal1 s 10741 11936 10936 12030 3 FreeSans 200 0 0 0 VDDIO_AMX
port 33 nsew
flabel metal1 s 2382 8577 2692 8746 3 FreeSans 200 0 0 0 VPB_DRVR
port 34 nsew
flabel comment s 2955 32848 2955 32848 0 FreeSans 800 0 0 0 VDDIO
<< properties >>
string GDS_END 46640978
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 46558308
<< end >>
