magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< metal3 >>
rect 11966 18573 14932 18592
rect 11966 18347 12211 18573
rect 12243 18539 12283 18573
rect 12324 18539 12364 18573
rect 12405 18539 12445 18573
rect 12486 18539 12526 18573
rect 12568 18539 12608 18573
rect 12650 18539 12690 18573
rect 12732 18539 12772 18573
rect 12814 18539 12854 18573
rect 12896 18539 12936 18573
rect 12978 18539 13018 18573
rect 13060 18539 13100 18573
rect 13142 18539 13182 18573
rect 13224 18539 13264 18573
rect 13306 18539 13346 18573
rect 13388 18539 13428 18573
rect 13470 18539 13510 18573
rect 13552 18539 13592 18573
rect 13634 18539 13674 18573
rect 13716 18539 13756 18573
rect 13798 18539 13838 18573
rect 13880 18539 13920 18573
rect 13962 18539 14002 18573
rect 14044 18539 14084 18573
rect 14126 18539 14166 18573
rect 14208 18539 14248 18573
rect 14290 18539 14330 18573
rect 14372 18539 14412 18573
rect 14454 18539 14494 18573
rect 14536 18539 14576 18573
rect 14618 18539 14658 18573
rect 14700 18539 14740 18573
rect 14782 18539 14822 18573
rect 14864 18539 14904 18573
rect 12231 18493 12295 18509
rect 12312 18493 12376 18509
rect 12393 18493 12457 18509
rect 12474 18493 12538 18509
rect 12556 18493 12620 18509
rect 12638 18493 12702 18509
rect 12720 18493 12784 18509
rect 12802 18493 12866 18509
rect 12884 18493 12948 18509
rect 12966 18493 13030 18509
rect 13048 18493 13112 18509
rect 13130 18493 13194 18509
rect 13212 18493 13276 18509
rect 13294 18493 13358 18509
rect 13376 18493 13440 18509
rect 13458 18493 13522 18509
rect 13540 18493 13604 18509
rect 13622 18493 13686 18509
rect 13704 18493 13768 18509
rect 13786 18493 13850 18509
rect 13868 18493 13932 18509
rect 13950 18493 14014 18509
rect 14032 18493 14096 18509
rect 14114 18493 14178 18509
rect 14196 18493 14260 18509
rect 14278 18493 14342 18509
rect 14360 18493 14424 18509
rect 14442 18493 14506 18509
rect 14524 18493 14588 18509
rect 14606 18493 14670 18509
rect 14688 18493 14752 18509
rect 14770 18493 14834 18509
rect 14852 18493 14916 18509
rect 12231 18445 12291 18493
rect 12231 18363 12291 18427
rect 11788 18169 11966 18347
rect 11979 18277 12043 18341
rect 12135 18277 12199 18341
rect 12231 18281 12291 18345
rect 11979 18191 12043 18255
rect 11530 17911 11788 18169
rect 11803 18099 11867 18163
rect 11885 18099 11949 18163
rect 11967 18099 12031 18163
rect 11803 18013 11867 18077
rect 11803 17927 11867 17991
rect 11283 17664 11530 17911
rect 11547 17841 11611 17905
rect 11703 17841 11767 17905
rect 11803 17841 11867 17905
rect 11547 17757 11610 17821
rect 11547 17674 11610 17738
rect 11027 17408 11283 17664
rect 11286 17563 11350 17627
rect 11368 17584 11432 17627
rect 11450 17584 11514 17627
rect 11532 17584 11596 17627
rect 11286 17482 11350 17546
rect 10742 17123 11027 17408
rect 11039 17338 11103 17402
rect 11187 17338 11251 17402
rect 11286 17401 11350 17465
rect 11286 17328 11350 17384
rect 11039 17250 11103 17314
rect 11039 17163 11103 17227
rect 10481 16862 10742 17123
rect 10765 17053 10829 17117
rect 10861 17053 10925 17117
rect 10957 17053 11021 17117
rect 11053 17053 11107 17117
rect 10765 16960 10822 17024
rect 10765 16867 10822 16931
rect 10152 16533 10481 16862
rect 10498 16792 10562 16856
rect 10656 16792 10720 16856
rect 10765 16782 10822 16838
rect 10498 16682 10561 16746
rect 10498 16613 10561 16636
rect 10498 16572 10562 16613
rect 10656 16572 10720 16613
rect 10765 16590 10829 16613
rect 10861 16590 10925 16613
rect 10957 16590 11021 16613
rect 11053 16590 11117 16613
rect 11149 16590 11213 16613
rect 11286 16599 11350 16613
rect 11368 16599 11432 16613
rect 11450 16599 11514 16613
rect 11532 16599 11596 16613
rect 11614 16599 11678 16613
rect 11696 16599 11760 16613
rect 11778 16599 11842 16613
rect 11860 16599 11924 16613
rect 11942 16599 12006 16613
rect 12024 16599 12088 16613
rect 12106 16599 12170 16613
rect 12231 16559 12295 16613
rect 12312 16559 12376 16613
rect 12393 16559 12457 16613
rect 12474 16559 12538 16613
rect 12556 16559 12620 16613
rect 12638 16559 12702 16613
rect 12720 16559 12784 16613
rect 12802 16559 12866 16613
rect 12884 16559 12948 16613
rect 12966 16559 13030 16613
rect 13048 16559 13112 16613
rect 13130 16559 13194 16613
rect 13212 16559 13276 16613
rect 13294 16559 13358 16613
rect 13376 16559 13440 16613
rect 13458 16559 13522 16613
rect 13540 16559 13604 16613
rect 13622 16559 13686 16613
rect 13704 16559 13768 16613
rect 13786 16559 13850 16613
rect 13868 16559 13932 16613
rect 13950 16559 14014 16613
rect 14032 16559 14096 16613
rect 14114 16559 14178 16613
rect 14196 16559 14260 16613
rect 14278 16559 14342 16613
rect 14360 16559 14424 16613
rect 14442 16559 14506 16613
rect 14524 16559 14588 16613
rect 14606 16559 14670 16613
rect 14688 16559 14752 16613
rect 14770 16559 14834 16613
rect 14852 16559 14916 16613
rect 10152 13607 14932 16533
rect 10151 12418 14931 13306
rect 120 3558 4900 4486
rect 10151 3558 14931 4486
<< obsm3 >>
rect 119 18427 11886 18591
rect 119 18249 11708 18427
rect 119 17991 11450 18249
rect 12291 18267 14932 18493
rect 119 17744 11203 17991
rect 12046 18089 14932 18267
rect 119 17488 10947 17744
rect 11868 17831 14932 18089
rect 119 17203 10662 17488
rect 11610 17584 14932 17831
rect 119 16942 10401 17203
rect 11363 17328 14932 17584
rect 119 13527 10072 16942
rect 11107 17043 14932 17328
rect 10822 16782 14932 17043
rect 10561 16613 14932 16782
rect 119 13386 14932 13527
rect 119 12418 10071 13386
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 18591 254 18600
rect 0 18527 281 18591
rect 299 18527 363 18591
rect 381 18527 445 18591
rect 463 18527 527 18591
rect 545 18527 609 18591
rect 627 18527 691 18591
rect 709 18527 773 18591
rect 791 18527 855 18591
rect 873 18527 937 18591
rect 955 18527 1019 18591
rect 1037 18527 1101 18591
rect 1119 18527 1183 18591
rect 1201 18527 1265 18591
rect 1283 18527 1347 18591
rect 1365 18527 1429 18591
rect 1447 18527 1511 18591
rect 1529 18527 1593 18591
rect 1611 18527 1675 18591
rect 1693 18527 1757 18591
rect 1775 18527 1839 18591
rect 1857 18527 1921 18591
rect 1939 18527 2003 18591
rect 2021 18527 2085 18591
rect 2103 18527 2167 18591
rect 2185 18527 2249 18591
rect 2267 18527 2331 18591
rect 2349 18527 2413 18591
rect 2431 18527 2495 18591
rect 2513 18527 2577 18591
rect 2594 18527 2658 18591
rect 2675 18527 2739 18591
rect 2756 18527 2820 18591
rect 0 18509 254 18527
rect 14746 18509 15000 18600
rect 0 18445 281 18509
rect 299 18445 363 18509
rect 381 18445 445 18509
rect 463 18445 527 18509
rect 545 18445 609 18509
rect 627 18445 691 18509
rect 709 18445 773 18509
rect 791 18445 855 18509
rect 873 18445 937 18509
rect 955 18445 1019 18509
rect 1037 18445 1101 18509
rect 1119 18445 1183 18509
rect 1201 18445 1265 18509
rect 1283 18445 1347 18509
rect 1365 18445 1429 18509
rect 1447 18445 1511 18509
rect 1529 18445 1593 18509
rect 1611 18445 1675 18509
rect 1693 18445 1757 18509
rect 1775 18445 1839 18509
rect 1857 18445 1921 18509
rect 1939 18445 2003 18509
rect 2021 18445 2085 18509
rect 2103 18445 2167 18509
rect 2185 18445 2249 18509
rect 2267 18445 2331 18509
rect 2349 18445 2413 18509
rect 2431 18445 2495 18509
rect 2513 18445 2577 18509
rect 2594 18445 2658 18509
rect 2675 18445 2739 18509
rect 2756 18445 2820 18509
rect 12231 18445 12295 18509
rect 12312 18445 12376 18509
rect 12393 18445 12457 18509
rect 12474 18445 12538 18509
rect 12556 18445 12620 18509
rect 12638 18445 12702 18509
rect 12720 18445 12784 18509
rect 12802 18445 12866 18509
rect 12884 18445 12948 18509
rect 12966 18445 13030 18509
rect 13048 18445 13112 18509
rect 13130 18445 13194 18509
rect 13212 18445 13276 18509
rect 13294 18445 13358 18509
rect 13376 18445 13440 18509
rect 13458 18445 13522 18509
rect 13540 18445 13604 18509
rect 13622 18445 13686 18509
rect 13704 18445 13768 18509
rect 13786 18445 13850 18509
rect 13868 18445 13932 18509
rect 13950 18445 14014 18509
rect 14032 18445 14096 18509
rect 14114 18445 14178 18509
rect 14196 18445 14260 18509
rect 14278 18445 14342 18509
rect 14360 18445 14424 18509
rect 14442 18445 14506 18509
rect 14524 18445 14588 18509
rect 14606 18445 14670 18509
rect 14688 18445 15000 18509
rect 0 18427 254 18445
rect 14746 18427 15000 18445
rect 0 18363 281 18427
rect 299 18363 363 18427
rect 381 18363 445 18427
rect 463 18363 527 18427
rect 545 18363 609 18427
rect 627 18363 691 18427
rect 709 18363 773 18427
rect 791 18363 855 18427
rect 873 18363 937 18427
rect 955 18363 1019 18427
rect 1037 18363 1101 18427
rect 1119 18363 1183 18427
rect 1201 18363 1265 18427
rect 1283 18363 1347 18427
rect 1365 18363 1429 18427
rect 1447 18363 1511 18427
rect 1529 18363 1593 18427
rect 1611 18363 1675 18427
rect 1693 18363 1757 18427
rect 1775 18363 1839 18427
rect 1857 18363 1921 18427
rect 1939 18363 2003 18427
rect 2021 18363 2085 18427
rect 2103 18363 2167 18427
rect 2185 18363 2249 18427
rect 2267 18363 2331 18427
rect 2349 18363 2413 18427
rect 2431 18363 2495 18427
rect 2513 18363 2577 18427
rect 2594 18363 2658 18427
rect 2675 18363 2739 18427
rect 2756 18363 2820 18427
rect 0 18345 254 18363
rect 0 18281 281 18345
rect 299 18281 363 18345
rect 381 18281 445 18345
rect 463 18281 527 18345
rect 545 18281 609 18345
rect 627 18281 691 18345
rect 709 18281 773 18345
rect 791 18281 855 18345
rect 873 18281 937 18345
rect 955 18281 1019 18345
rect 1037 18281 1101 18345
rect 1119 18281 1183 18345
rect 1201 18281 1265 18345
rect 1283 18281 1347 18345
rect 1365 18281 1429 18345
rect 1447 18281 1511 18345
rect 1529 18281 1593 18345
rect 1611 18281 1675 18345
rect 1693 18281 1757 18345
rect 1775 18281 1839 18345
rect 1857 18281 1921 18345
rect 1939 18281 2003 18345
rect 2021 18281 2085 18345
rect 2103 18281 2167 18345
rect 2185 18281 2249 18345
rect 2267 18281 2331 18345
rect 2349 18281 2413 18345
rect 2431 18281 2495 18345
rect 2513 18281 2577 18345
rect 2594 18281 2658 18345
rect 2675 18281 2739 18345
rect 2756 18281 2820 18345
rect 0 18263 254 18281
rect 0 18199 281 18263
rect 299 18199 363 18263
rect 381 18199 445 18263
rect 463 18199 527 18263
rect 545 18199 609 18263
rect 627 18199 691 18263
rect 709 18199 773 18263
rect 791 18199 855 18263
rect 873 18199 937 18263
rect 955 18199 1019 18263
rect 1037 18199 1101 18263
rect 1119 18199 1183 18263
rect 1201 18199 1265 18263
rect 1283 18199 1347 18263
rect 1365 18199 1429 18263
rect 1447 18199 1511 18263
rect 1529 18199 1593 18263
rect 1611 18199 1675 18263
rect 1693 18199 1757 18263
rect 1775 18199 1839 18263
rect 1857 18199 1921 18263
rect 1939 18199 2003 18263
rect 2021 18199 2085 18263
rect 2103 18199 2167 18263
rect 2185 18199 2249 18263
rect 2267 18199 2331 18263
rect 2349 18199 2413 18263
rect 2431 18199 2495 18263
rect 2513 18199 2577 18263
rect 2594 18199 2658 18263
rect 2675 18199 2739 18263
rect 2756 18199 2820 18263
rect 0 18181 254 18199
rect 2851 18190 3073 18342
rect 12231 18363 12295 18427
rect 12312 18363 12376 18427
rect 12393 18363 12457 18427
rect 12474 18363 12538 18427
rect 12556 18363 12620 18427
rect 12638 18363 12702 18427
rect 12720 18363 12784 18427
rect 12802 18363 12866 18427
rect 12884 18363 12948 18427
rect 12966 18363 13030 18427
rect 13048 18363 13112 18427
rect 13130 18363 13194 18427
rect 13212 18363 13276 18427
rect 13294 18363 13358 18427
rect 13376 18363 13440 18427
rect 13458 18363 13522 18427
rect 13540 18363 13604 18427
rect 13622 18363 13686 18427
rect 13704 18363 13768 18427
rect 13786 18363 13850 18427
rect 13868 18363 13932 18427
rect 13950 18363 14014 18427
rect 14032 18363 14096 18427
rect 14114 18363 14178 18427
rect 14196 18363 14260 18427
rect 14278 18363 14342 18427
rect 14360 18363 14424 18427
rect 14442 18363 14506 18427
rect 14524 18363 14588 18427
rect 14606 18363 14670 18427
rect 14688 18363 15000 18427
rect 14746 18345 15000 18363
rect 0 18117 281 18181
rect 299 18117 363 18181
rect 381 18117 445 18181
rect 463 18117 527 18181
rect 545 18117 609 18181
rect 627 18117 691 18181
rect 709 18117 773 18181
rect 791 18117 855 18181
rect 873 18117 937 18181
rect 955 18117 1019 18181
rect 1037 18117 1101 18181
rect 1119 18117 1183 18181
rect 1201 18117 1265 18181
rect 1283 18117 1347 18181
rect 1365 18117 1429 18181
rect 1447 18117 1511 18181
rect 1529 18117 1593 18181
rect 1611 18117 1675 18181
rect 1693 18117 1757 18181
rect 1775 18117 1839 18181
rect 1857 18117 1921 18181
rect 1939 18117 2003 18181
rect 2021 18117 2085 18181
rect 2103 18117 2167 18181
rect 2185 18117 2249 18181
rect 2267 18117 2331 18181
rect 2349 18117 2413 18181
rect 2431 18117 2495 18181
rect 2513 18117 2577 18181
rect 2594 18117 2658 18181
rect 2675 18117 2739 18181
rect 2756 18117 2820 18181
rect 0 18099 254 18117
rect 0 18035 281 18099
rect 299 18035 363 18099
rect 381 18035 445 18099
rect 463 18035 527 18099
rect 545 18035 609 18099
rect 627 18035 691 18099
rect 709 18035 773 18099
rect 791 18035 855 18099
rect 873 18035 937 18099
rect 955 18035 1019 18099
rect 1037 18035 1101 18099
rect 1119 18035 1183 18099
rect 1201 18035 1265 18099
rect 1283 18035 1347 18099
rect 1365 18035 1429 18099
rect 1447 18035 1511 18099
rect 1529 18035 1593 18099
rect 1611 18035 1675 18099
rect 1693 18035 1757 18099
rect 1775 18035 1839 18099
rect 1857 18035 1921 18099
rect 1939 18035 2003 18099
rect 2021 18035 2085 18099
rect 2103 18035 2167 18099
rect 2185 18035 2249 18099
rect 2267 18035 2331 18099
rect 2349 18035 2413 18099
rect 2431 18035 2495 18099
rect 2513 18035 2577 18099
rect 2594 18035 2658 18099
rect 2675 18035 2739 18099
rect 2756 18035 2820 18099
rect 0 18017 254 18035
rect 0 17953 281 18017
rect 299 17953 363 18017
rect 381 17953 445 18017
rect 463 17953 527 18017
rect 545 17953 609 18017
rect 627 17953 691 18017
rect 709 17953 773 18017
rect 791 17953 855 18017
rect 873 17953 937 18017
rect 955 17953 1019 18017
rect 1037 17953 1101 18017
rect 1119 17953 1183 18017
rect 1201 17953 1265 18017
rect 1283 17953 1347 18017
rect 1365 17953 1429 18017
rect 1447 17953 1511 18017
rect 1529 17953 1593 18017
rect 1611 17953 1675 18017
rect 1693 17953 1757 18017
rect 1775 17953 1839 18017
rect 1857 17953 1921 18017
rect 1939 17953 2003 18017
rect 2021 17953 2085 18017
rect 2103 17953 2167 18017
rect 2185 17953 2249 18017
rect 2267 17953 2331 18017
rect 2349 17953 2413 18017
rect 2431 17953 2495 18017
rect 2513 17953 2577 18017
rect 2594 17953 2658 18017
rect 2675 17953 2739 18017
rect 2756 17953 2820 18017
rect 0 17935 254 17953
rect 0 17871 281 17935
rect 299 17871 363 17935
rect 381 17871 445 17935
rect 463 17871 527 17935
rect 545 17871 609 17935
rect 627 17871 691 17935
rect 709 17871 773 17935
rect 791 17871 855 17935
rect 873 17871 937 17935
rect 955 17871 1019 17935
rect 1037 17871 1101 17935
rect 1119 17871 1183 17935
rect 1201 17871 1265 17935
rect 1283 17871 1347 17935
rect 1365 17871 1429 17935
rect 1447 17871 1511 17935
rect 1529 17871 1593 17935
rect 1611 17871 1675 17935
rect 1693 17871 1757 17935
rect 1775 17871 1839 17935
rect 1857 17871 1921 17935
rect 1939 17871 2003 17935
rect 2021 17871 2085 17935
rect 2103 17871 2167 17935
rect 2185 17871 2249 17935
rect 2267 17871 2331 17935
rect 2349 17871 2413 17935
rect 2431 17871 2495 17935
rect 2513 17871 2577 17935
rect 2594 17871 2658 17935
rect 2675 17871 2739 17935
rect 2756 17871 2820 17935
rect 0 17853 254 17871
rect 0 17789 281 17853
rect 299 17789 363 17853
rect 381 17789 445 17853
rect 463 17789 527 17853
rect 545 17789 609 17853
rect 627 17789 691 17853
rect 709 17789 773 17853
rect 791 17789 855 17853
rect 873 17789 937 17853
rect 955 17789 1019 17853
rect 1037 17789 1101 17853
rect 1119 17789 1183 17853
rect 1201 17789 1265 17853
rect 1283 17789 1347 17853
rect 1365 17789 1429 17853
rect 1447 17789 1511 17853
rect 1529 17789 1593 17853
rect 1611 17789 1675 17853
rect 1693 17789 1757 17853
rect 1775 17789 1839 17853
rect 1857 17789 1921 17853
rect 1939 17789 2003 17853
rect 2021 17789 2085 17853
rect 2103 17789 2167 17853
rect 2185 17789 2249 17853
rect 2267 17789 2331 17853
rect 2349 17789 2413 17853
rect 2431 17789 2495 17853
rect 2513 17789 2577 17853
rect 2594 17789 2658 17853
rect 2675 17789 2739 17853
rect 2756 17789 2820 17853
rect 0 17771 254 17789
rect 0 17707 281 17771
rect 299 17707 363 17771
rect 381 17707 445 17771
rect 463 17707 527 17771
rect 545 17707 609 17771
rect 627 17707 691 17771
rect 709 17707 773 17771
rect 791 17707 855 17771
rect 873 17707 937 17771
rect 955 17707 1019 17771
rect 1037 17707 1101 17771
rect 1119 17707 1183 17771
rect 1201 17707 1265 17771
rect 1283 17707 1347 17771
rect 1365 17707 1429 17771
rect 1447 17707 1511 17771
rect 1529 17707 1593 17771
rect 1611 17707 1675 17771
rect 1693 17707 1757 17771
rect 1775 17707 1839 17771
rect 1857 17707 1921 17771
rect 1939 17707 2003 17771
rect 2021 17707 2085 17771
rect 2103 17707 2167 17771
rect 2185 17707 2249 17771
rect 2267 17707 2331 17771
rect 2349 17707 2413 17771
rect 2431 17707 2495 17771
rect 2513 17707 2577 17771
rect 2594 17707 2658 17771
rect 2675 17707 2739 17771
rect 2756 17707 2820 17771
rect 0 17689 254 17707
rect 0 17625 281 17689
rect 299 17625 363 17689
rect 381 17625 445 17689
rect 463 17625 527 17689
rect 545 17625 609 17689
rect 627 17625 691 17689
rect 709 17625 773 17689
rect 791 17625 855 17689
rect 873 17625 937 17689
rect 955 17625 1019 17689
rect 1037 17625 1101 17689
rect 1119 17625 1183 17689
rect 1201 17625 1265 17689
rect 1283 17625 1347 17689
rect 1365 17625 1429 17689
rect 1447 17625 1511 17689
rect 1529 17625 1593 17689
rect 1611 17625 1675 17689
rect 1693 17625 1757 17689
rect 1775 17625 1839 17689
rect 1857 17625 1921 17689
rect 1939 17625 2003 17689
rect 2021 17625 2085 17689
rect 2103 17625 2167 17689
rect 2185 17625 2249 17689
rect 2267 17625 2331 17689
rect 2349 17625 2413 17689
rect 2431 17625 2495 17689
rect 2513 17625 2577 17689
rect 2594 17625 2658 17689
rect 2675 17625 2739 17689
rect 2756 17625 2820 17689
rect 2854 17669 3250 18164
rect 11978 18190 12200 18342
rect 12231 18281 12295 18345
rect 12312 18281 12376 18345
rect 12393 18281 12457 18345
rect 12474 18281 12538 18345
rect 12556 18281 12620 18345
rect 12638 18281 12702 18345
rect 12720 18281 12784 18345
rect 12802 18281 12866 18345
rect 12884 18281 12948 18345
rect 12966 18281 13030 18345
rect 13048 18281 13112 18345
rect 13130 18281 13194 18345
rect 13212 18281 13276 18345
rect 13294 18281 13358 18345
rect 13376 18281 13440 18345
rect 13458 18281 13522 18345
rect 13540 18281 13604 18345
rect 13622 18281 13686 18345
rect 13704 18281 13768 18345
rect 13786 18281 13850 18345
rect 13868 18281 13932 18345
rect 13950 18281 14014 18345
rect 14032 18281 14096 18345
rect 14114 18281 14178 18345
rect 14196 18281 14260 18345
rect 14278 18281 14342 18345
rect 14360 18281 14424 18345
rect 14442 18281 14506 18345
rect 14524 18281 14588 18345
rect 14606 18281 14670 18345
rect 14688 18281 15000 18345
rect 14746 18263 15000 18281
rect 12231 18199 12295 18263
rect 12312 18199 12376 18263
rect 12393 18199 12457 18263
rect 12474 18199 12538 18263
rect 12556 18199 12620 18263
rect 12638 18199 12702 18263
rect 12720 18199 12784 18263
rect 12802 18199 12866 18263
rect 12884 18199 12948 18263
rect 12966 18199 13030 18263
rect 13048 18199 13112 18263
rect 13130 18199 13194 18263
rect 13212 18199 13276 18263
rect 13294 18199 13358 18263
rect 13376 18199 13440 18263
rect 13458 18199 13522 18263
rect 13540 18199 13604 18263
rect 13622 18199 13686 18263
rect 13704 18199 13768 18263
rect 13786 18199 13850 18263
rect 13868 18199 13932 18263
rect 13950 18199 14014 18263
rect 14032 18199 14096 18263
rect 14114 18199 14178 18263
rect 14196 18199 14260 18263
rect 14278 18199 14342 18263
rect 14360 18199 14424 18263
rect 14442 18199 14506 18263
rect 14524 18199 14588 18263
rect 14606 18199 14670 18263
rect 14688 18199 15000 18263
rect 14746 18181 15000 18199
rect 3283 17673 3505 17906
rect 0 17607 254 17625
rect 0 17543 281 17607
rect 299 17543 363 17607
rect 381 17543 445 17607
rect 463 17543 527 17607
rect 545 17543 609 17607
rect 627 17543 691 17607
rect 709 17543 773 17607
rect 791 17543 855 17607
rect 873 17543 937 17607
rect 955 17543 1019 17607
rect 1037 17543 1101 17607
rect 1119 17543 1183 17607
rect 1201 17543 1265 17607
rect 1283 17543 1347 17607
rect 1365 17543 1429 17607
rect 1447 17543 1511 17607
rect 1529 17543 1593 17607
rect 1611 17543 1675 17607
rect 1693 17543 1757 17607
rect 1775 17543 1839 17607
rect 1857 17543 1921 17607
rect 1939 17543 2003 17607
rect 2021 17543 2085 17607
rect 2103 17543 2167 17607
rect 2185 17543 2249 17607
rect 2267 17543 2331 17607
rect 2349 17543 2413 17607
rect 2431 17543 2495 17607
rect 2513 17543 2577 17607
rect 2594 17543 2658 17607
rect 2675 17543 2739 17607
rect 2756 17543 2820 17607
rect 0 17525 254 17543
rect 0 17461 281 17525
rect 299 17461 363 17525
rect 381 17461 445 17525
rect 463 17461 527 17525
rect 545 17461 609 17525
rect 627 17461 691 17525
rect 709 17461 773 17525
rect 791 17461 855 17525
rect 873 17461 937 17525
rect 955 17461 1019 17525
rect 1037 17461 1101 17525
rect 1119 17461 1183 17525
rect 1201 17461 1265 17525
rect 1283 17461 1347 17525
rect 1365 17461 1429 17525
rect 1447 17461 1511 17525
rect 1529 17461 1593 17525
rect 1611 17461 1675 17525
rect 1693 17461 1757 17525
rect 1775 17461 1839 17525
rect 1857 17461 1921 17525
rect 1939 17461 2003 17525
rect 2021 17461 2085 17525
rect 2103 17461 2167 17525
rect 2185 17461 2249 17525
rect 2267 17461 2331 17525
rect 2349 17461 2413 17525
rect 2431 17461 2495 17525
rect 2513 17461 2577 17525
rect 2594 17461 2658 17525
rect 2675 17461 2739 17525
rect 2756 17461 2820 17525
rect 0 17443 254 17461
rect 0 17379 281 17443
rect 299 17379 363 17443
rect 381 17379 445 17443
rect 463 17379 527 17443
rect 545 17379 609 17443
rect 627 17379 691 17443
rect 709 17379 773 17443
rect 791 17379 855 17443
rect 873 17379 937 17443
rect 955 17379 1019 17443
rect 1037 17379 1101 17443
rect 1119 17379 1183 17443
rect 1201 17379 1265 17443
rect 1283 17379 1347 17443
rect 1365 17379 1429 17443
rect 1447 17379 1511 17443
rect 1529 17379 1593 17443
rect 1611 17379 1675 17443
rect 1693 17379 1757 17443
rect 1775 17379 1839 17443
rect 1857 17379 1921 17443
rect 1939 17379 2003 17443
rect 2021 17379 2085 17443
rect 2103 17379 2167 17443
rect 2185 17379 2249 17443
rect 2267 17379 2331 17443
rect 2349 17379 2413 17443
rect 2431 17379 2495 17443
rect 2513 17379 2577 17443
rect 2594 17379 2658 17443
rect 2675 17379 2739 17443
rect 2756 17379 2820 17443
rect 0 17361 254 17379
rect 0 17297 281 17361
rect 299 17297 363 17361
rect 381 17297 445 17361
rect 463 17297 527 17361
rect 545 17297 609 17361
rect 627 17297 691 17361
rect 709 17297 773 17361
rect 791 17297 855 17361
rect 873 17297 937 17361
rect 955 17297 1019 17361
rect 1037 17297 1101 17361
rect 1119 17297 1183 17361
rect 1201 17297 1265 17361
rect 1283 17297 1347 17361
rect 1365 17297 1429 17361
rect 1447 17297 1511 17361
rect 1529 17297 1593 17361
rect 1611 17297 1675 17361
rect 1693 17297 1757 17361
rect 1775 17297 1839 17361
rect 1857 17297 1921 17361
rect 1939 17297 2003 17361
rect 2021 17297 2085 17361
rect 2103 17297 2167 17361
rect 2185 17297 2249 17361
rect 2267 17297 2331 17361
rect 2349 17297 2413 17361
rect 2431 17297 2495 17361
rect 2513 17297 2577 17361
rect 2594 17297 2658 17361
rect 2675 17297 2739 17361
rect 2756 17297 2820 17361
rect 0 17279 254 17297
rect 0 17215 281 17279
rect 299 17215 363 17279
rect 381 17215 445 17279
rect 463 17215 527 17279
rect 545 17215 609 17279
rect 627 17215 691 17279
rect 709 17215 773 17279
rect 791 17215 855 17279
rect 873 17215 937 17279
rect 955 17215 1019 17279
rect 1037 17215 1101 17279
rect 1119 17215 1183 17279
rect 1201 17215 1265 17279
rect 1283 17215 1347 17279
rect 1365 17215 1429 17279
rect 1447 17215 1511 17279
rect 1529 17215 1593 17279
rect 1611 17215 1675 17279
rect 1693 17215 1757 17279
rect 1775 17215 1839 17279
rect 1857 17215 1921 17279
rect 1939 17215 2003 17279
rect 2021 17215 2085 17279
rect 2103 17215 2167 17279
rect 2185 17215 2249 17279
rect 2267 17215 2331 17279
rect 2349 17215 2413 17279
rect 2431 17215 2495 17279
rect 2513 17215 2577 17279
rect 2594 17215 2658 17279
rect 2675 17215 2739 17279
rect 2756 17215 2820 17279
rect 0 17197 254 17215
rect 0 17133 281 17197
rect 299 17133 363 17197
rect 381 17133 445 17197
rect 463 17133 527 17197
rect 545 17133 609 17197
rect 627 17133 691 17197
rect 709 17133 773 17197
rect 791 17133 855 17197
rect 873 17133 937 17197
rect 955 17133 1019 17197
rect 1037 17133 1101 17197
rect 1119 17133 1183 17197
rect 1201 17133 1265 17197
rect 1283 17133 1347 17197
rect 1365 17133 1429 17197
rect 1447 17133 1511 17197
rect 1529 17133 1593 17197
rect 1611 17133 1675 17197
rect 1693 17133 1757 17197
rect 1775 17133 1839 17197
rect 1857 17133 1921 17197
rect 1939 17133 2003 17197
rect 2021 17133 2085 17197
rect 2103 17133 2167 17197
rect 2185 17133 2249 17197
rect 2267 17133 2331 17197
rect 2349 17133 2413 17197
rect 2431 17133 2495 17197
rect 2513 17133 2577 17197
rect 2594 17133 2658 17197
rect 2675 17133 2739 17197
rect 2756 17133 2820 17197
rect 0 17115 254 17133
rect 0 17051 281 17115
rect 299 17051 363 17115
rect 381 17051 445 17115
rect 463 17051 527 17115
rect 545 17051 609 17115
rect 627 17051 691 17115
rect 709 17051 773 17115
rect 791 17051 855 17115
rect 873 17051 937 17115
rect 955 17051 1019 17115
rect 1037 17051 1101 17115
rect 1119 17051 1183 17115
rect 1201 17051 1265 17115
rect 1283 17051 1347 17115
rect 1365 17051 1429 17115
rect 1447 17051 1511 17115
rect 1529 17051 1593 17115
rect 1611 17051 1675 17115
rect 1693 17051 1757 17115
rect 1775 17051 1839 17115
rect 1857 17051 1921 17115
rect 1939 17051 2003 17115
rect 2021 17051 2085 17115
rect 2103 17051 2167 17115
rect 2185 17051 2249 17115
rect 2267 17051 2331 17115
rect 2349 17051 2413 17115
rect 2431 17051 2495 17115
rect 2513 17051 2577 17115
rect 2594 17051 2658 17115
rect 2675 17051 2739 17115
rect 2756 17051 2820 17115
rect 0 17033 254 17051
rect 0 16969 281 17033
rect 299 16969 363 17033
rect 381 16969 445 17033
rect 463 16969 527 17033
rect 545 16969 609 17033
rect 627 16969 691 17033
rect 709 16969 773 17033
rect 791 16969 855 17033
rect 873 16969 937 17033
rect 955 16969 1019 17033
rect 1037 16969 1101 17033
rect 1119 16969 1183 17033
rect 1201 16969 1265 17033
rect 1283 16969 1347 17033
rect 1365 16969 1429 17033
rect 1447 16969 1511 17033
rect 1529 16969 1593 17033
rect 1611 16969 1675 17033
rect 1693 16969 1757 17033
rect 1775 16969 1839 17033
rect 1857 16969 1921 17033
rect 1939 16969 2003 17033
rect 2021 16969 2085 17033
rect 2103 16969 2167 17033
rect 2185 16969 2249 17033
rect 2267 16969 2331 17033
rect 2349 16969 2413 17033
rect 2431 16969 2495 17033
rect 2513 16969 2577 17033
rect 2594 16969 2658 17033
rect 2675 16969 2739 17033
rect 2756 16969 2820 17033
rect 0 16951 254 16969
rect 0 16887 281 16951
rect 299 16887 363 16951
rect 381 16887 445 16951
rect 463 16887 527 16951
rect 545 16887 609 16951
rect 627 16887 691 16951
rect 709 16887 773 16951
rect 791 16887 855 16951
rect 873 16887 937 16951
rect 955 16887 1019 16951
rect 1037 16887 1101 16951
rect 1119 16887 1183 16951
rect 1201 16887 1265 16951
rect 1283 16887 1347 16951
rect 1365 16887 1429 16951
rect 1447 16887 1511 16951
rect 1529 16887 1593 16951
rect 1611 16887 1675 16951
rect 1693 16887 1757 16951
rect 1775 16887 1839 16951
rect 1857 16887 1921 16951
rect 1939 16887 2003 16951
rect 2021 16887 2085 16951
rect 2103 16887 2167 16951
rect 2185 16887 2249 16951
rect 2267 16887 2331 16951
rect 2349 16887 2413 16951
rect 2431 16887 2495 16951
rect 2513 16887 2577 16951
rect 2594 16887 2658 16951
rect 2675 16887 2739 16951
rect 2756 16887 2820 16951
rect 0 16869 254 16887
rect 0 16805 281 16869
rect 299 16805 363 16869
rect 381 16805 445 16869
rect 463 16805 527 16869
rect 545 16805 609 16869
rect 627 16805 691 16869
rect 709 16805 773 16869
rect 791 16805 855 16869
rect 873 16805 937 16869
rect 955 16805 1019 16869
rect 1037 16805 1101 16869
rect 1119 16805 1183 16869
rect 1201 16805 1265 16869
rect 1283 16805 1347 16869
rect 1365 16805 1429 16869
rect 1447 16805 1511 16869
rect 1529 16805 1593 16869
rect 1611 16805 1675 16869
rect 1693 16805 1757 16869
rect 1775 16805 1839 16869
rect 1857 16805 1921 16869
rect 1939 16805 2003 16869
rect 2021 16805 2085 16869
rect 2103 16805 2167 16869
rect 2185 16805 2249 16869
rect 2267 16805 2331 16869
rect 2349 16805 2413 16869
rect 2431 16805 2495 16869
rect 2513 16805 2577 16869
rect 2594 16805 2658 16869
rect 2675 16805 2739 16869
rect 2756 16805 2820 16869
rect 0 16787 254 16805
rect 0 16723 281 16787
rect 299 16723 363 16787
rect 381 16723 445 16787
rect 463 16723 527 16787
rect 545 16723 609 16787
rect 627 16723 691 16787
rect 709 16723 773 16787
rect 791 16723 855 16787
rect 873 16723 937 16787
rect 955 16723 1019 16787
rect 1037 16723 1101 16787
rect 1119 16723 1183 16787
rect 1201 16723 1265 16787
rect 1283 16723 1347 16787
rect 1365 16723 1429 16787
rect 1447 16723 1511 16787
rect 1529 16723 1593 16787
rect 1611 16723 1675 16787
rect 1693 16723 1757 16787
rect 1775 16723 1839 16787
rect 1857 16723 1921 16787
rect 1939 16723 2003 16787
rect 2021 16723 2085 16787
rect 2103 16723 2167 16787
rect 2185 16723 2249 16787
rect 2267 16723 2331 16787
rect 2349 16723 2413 16787
rect 2431 16723 2495 16787
rect 2513 16723 2577 16787
rect 2594 16723 2658 16787
rect 2675 16723 2739 16787
rect 2756 16723 2820 16787
rect 0 16705 254 16723
rect 0 16641 281 16705
rect 299 16641 363 16705
rect 381 16641 445 16705
rect 463 16641 527 16705
rect 545 16641 609 16705
rect 627 16641 691 16705
rect 709 16641 773 16705
rect 791 16641 855 16705
rect 873 16641 937 16705
rect 955 16641 1019 16705
rect 1037 16641 1101 16705
rect 1119 16641 1183 16705
rect 1201 16641 1265 16705
rect 1283 16641 1347 16705
rect 1365 16641 1429 16705
rect 1447 16641 1511 16705
rect 1529 16641 1593 16705
rect 1611 16641 1675 16705
rect 1693 16641 1757 16705
rect 1775 16641 1839 16705
rect 1857 16641 1921 16705
rect 1939 16641 2003 16705
rect 2021 16641 2085 16705
rect 2103 16641 2167 16705
rect 2185 16641 2249 16705
rect 2267 16641 2331 16705
rect 2349 16641 2413 16705
rect 2431 16641 2495 16705
rect 2513 16641 2577 16705
rect 2594 16641 2658 16705
rect 2675 16641 2739 16705
rect 2756 16641 2820 16705
rect 0 16623 254 16641
rect 0 16559 281 16623
rect 299 16559 363 16623
rect 381 16559 445 16623
rect 463 16559 527 16623
rect 545 16559 609 16623
rect 627 16559 691 16623
rect 709 16559 773 16623
rect 791 16559 855 16623
rect 873 16559 937 16623
rect 955 16559 1019 16623
rect 1037 16559 1101 16623
rect 1119 16559 1183 16623
rect 1201 16559 1265 16623
rect 1283 16559 1347 16623
rect 1365 16559 1429 16623
rect 1447 16559 1511 16623
rect 1529 16559 1593 16623
rect 1611 16559 1675 16623
rect 1693 16559 1757 16623
rect 1775 16559 1839 16623
rect 1857 16559 1921 16623
rect 1939 16559 2003 16623
rect 2021 16559 2085 16623
rect 2103 16559 2167 16623
rect 2185 16559 2249 16623
rect 2267 16559 2331 16623
rect 2349 16559 2413 16623
rect 2431 16559 2495 16623
rect 2513 16559 2577 16623
rect 2594 16559 2658 16623
rect 2675 16559 2739 16623
rect 2756 16559 2820 16623
rect 2875 16598 3771 17628
rect 11546 17673 11768 17906
rect 11801 17669 12197 18164
rect 12231 18117 12295 18181
rect 12312 18117 12376 18181
rect 12393 18117 12457 18181
rect 12474 18117 12538 18181
rect 12556 18117 12620 18181
rect 12638 18117 12702 18181
rect 12720 18117 12784 18181
rect 12802 18117 12866 18181
rect 12884 18117 12948 18181
rect 12966 18117 13030 18181
rect 13048 18117 13112 18181
rect 13130 18117 13194 18181
rect 13212 18117 13276 18181
rect 13294 18117 13358 18181
rect 13376 18117 13440 18181
rect 13458 18117 13522 18181
rect 13540 18117 13604 18181
rect 13622 18117 13686 18181
rect 13704 18117 13768 18181
rect 13786 18117 13850 18181
rect 13868 18117 13932 18181
rect 13950 18117 14014 18181
rect 14032 18117 14096 18181
rect 14114 18117 14178 18181
rect 14196 18117 14260 18181
rect 14278 18117 14342 18181
rect 14360 18117 14424 18181
rect 14442 18117 14506 18181
rect 14524 18117 14588 18181
rect 14606 18117 14670 18181
rect 14688 18117 15000 18181
rect 14746 18099 15000 18117
rect 12231 18035 12295 18099
rect 12312 18035 12376 18099
rect 12393 18035 12457 18099
rect 12474 18035 12538 18099
rect 12556 18035 12620 18099
rect 12638 18035 12702 18099
rect 12720 18035 12784 18099
rect 12802 18035 12866 18099
rect 12884 18035 12948 18099
rect 12966 18035 13030 18099
rect 13048 18035 13112 18099
rect 13130 18035 13194 18099
rect 13212 18035 13276 18099
rect 13294 18035 13358 18099
rect 13376 18035 13440 18099
rect 13458 18035 13522 18099
rect 13540 18035 13604 18099
rect 13622 18035 13686 18099
rect 13704 18035 13768 18099
rect 13786 18035 13850 18099
rect 13868 18035 13932 18099
rect 13950 18035 14014 18099
rect 14032 18035 14096 18099
rect 14114 18035 14178 18099
rect 14196 18035 14260 18099
rect 14278 18035 14342 18099
rect 14360 18035 14424 18099
rect 14442 18035 14506 18099
rect 14524 18035 14588 18099
rect 14606 18035 14670 18099
rect 14688 18035 15000 18099
rect 14746 18017 15000 18035
rect 12231 17953 12295 18017
rect 12312 17953 12376 18017
rect 12393 17953 12457 18017
rect 12474 17953 12538 18017
rect 12556 17953 12620 18017
rect 12638 17953 12702 18017
rect 12720 17953 12784 18017
rect 12802 17953 12866 18017
rect 12884 17953 12948 18017
rect 12966 17953 13030 18017
rect 13048 17953 13112 18017
rect 13130 17953 13194 18017
rect 13212 17953 13276 18017
rect 13294 17953 13358 18017
rect 13376 17953 13440 18017
rect 13458 17953 13522 18017
rect 13540 17953 13604 18017
rect 13622 17953 13686 18017
rect 13704 17953 13768 18017
rect 13786 17953 13850 18017
rect 13868 17953 13932 18017
rect 13950 17953 14014 18017
rect 14032 17953 14096 18017
rect 14114 17953 14178 18017
rect 14196 17953 14260 18017
rect 14278 17953 14342 18017
rect 14360 17953 14424 18017
rect 14442 17953 14506 18017
rect 14524 17953 14588 18017
rect 14606 17953 14670 18017
rect 14688 17953 15000 18017
rect 14746 17935 15000 17953
rect 12231 17871 12295 17935
rect 12312 17871 12376 17935
rect 12393 17871 12457 17935
rect 12474 17871 12538 17935
rect 12556 17871 12620 17935
rect 12638 17871 12702 17935
rect 12720 17871 12784 17935
rect 12802 17871 12866 17935
rect 12884 17871 12948 17935
rect 12966 17871 13030 17935
rect 13048 17871 13112 17935
rect 13130 17871 13194 17935
rect 13212 17871 13276 17935
rect 13294 17871 13358 17935
rect 13376 17871 13440 17935
rect 13458 17871 13522 17935
rect 13540 17871 13604 17935
rect 13622 17871 13686 17935
rect 13704 17871 13768 17935
rect 13786 17871 13850 17935
rect 13868 17871 13932 17935
rect 13950 17871 14014 17935
rect 14032 17871 14096 17935
rect 14114 17871 14178 17935
rect 14196 17871 14260 17935
rect 14278 17871 14342 17935
rect 14360 17871 14424 17935
rect 14442 17871 14506 17935
rect 14524 17871 14588 17935
rect 14606 17871 14670 17935
rect 14688 17871 15000 17935
rect 14746 17853 15000 17871
rect 12231 17789 12295 17853
rect 12312 17789 12376 17853
rect 12393 17789 12457 17853
rect 12474 17789 12538 17853
rect 12556 17789 12620 17853
rect 12638 17789 12702 17853
rect 12720 17789 12784 17853
rect 12802 17789 12866 17853
rect 12884 17789 12948 17853
rect 12966 17789 13030 17853
rect 13048 17789 13112 17853
rect 13130 17789 13194 17853
rect 13212 17789 13276 17853
rect 13294 17789 13358 17853
rect 13376 17789 13440 17853
rect 13458 17789 13522 17853
rect 13540 17789 13604 17853
rect 13622 17789 13686 17853
rect 13704 17789 13768 17853
rect 13786 17789 13850 17853
rect 13868 17789 13932 17853
rect 13950 17789 14014 17853
rect 14032 17789 14096 17853
rect 14114 17789 14178 17853
rect 14196 17789 14260 17853
rect 14278 17789 14342 17853
rect 14360 17789 14424 17853
rect 14442 17789 14506 17853
rect 14524 17789 14588 17853
rect 14606 17789 14670 17853
rect 14688 17789 15000 17853
rect 14746 17771 15000 17789
rect 12231 17707 12295 17771
rect 12312 17707 12376 17771
rect 12393 17707 12457 17771
rect 12474 17707 12538 17771
rect 12556 17707 12620 17771
rect 12638 17707 12702 17771
rect 12720 17707 12784 17771
rect 12802 17707 12866 17771
rect 12884 17707 12948 17771
rect 12966 17707 13030 17771
rect 13048 17707 13112 17771
rect 13130 17707 13194 17771
rect 13212 17707 13276 17771
rect 13294 17707 13358 17771
rect 13376 17707 13440 17771
rect 13458 17707 13522 17771
rect 13540 17707 13604 17771
rect 13622 17707 13686 17771
rect 13704 17707 13768 17771
rect 13786 17707 13850 17771
rect 13868 17707 13932 17771
rect 13950 17707 14014 17771
rect 14032 17707 14096 17771
rect 14114 17707 14178 17771
rect 14196 17707 14260 17771
rect 14278 17707 14342 17771
rect 14360 17707 14424 17771
rect 14442 17707 14506 17771
rect 14524 17707 14588 17771
rect 14606 17707 14670 17771
rect 14688 17707 15000 17771
rect 14746 17689 15000 17707
rect 3799 17162 4013 17403
rect 3834 16589 4290 17118
rect 11038 17162 11252 17403
rect 4330 16571 4554 16857
rect 0 16524 254 16559
rect 10497 16571 10721 16857
rect 10761 16589 11217 17118
rect 11280 16598 12176 17628
rect 12231 17625 12295 17689
rect 12312 17625 12376 17689
rect 12393 17625 12457 17689
rect 12474 17625 12538 17689
rect 12556 17625 12620 17689
rect 12638 17625 12702 17689
rect 12720 17625 12784 17689
rect 12802 17625 12866 17689
rect 12884 17625 12948 17689
rect 12966 17625 13030 17689
rect 13048 17625 13112 17689
rect 13130 17625 13194 17689
rect 13212 17625 13276 17689
rect 13294 17625 13358 17689
rect 13376 17625 13440 17689
rect 13458 17625 13522 17689
rect 13540 17625 13604 17689
rect 13622 17625 13686 17689
rect 13704 17625 13768 17689
rect 13786 17625 13850 17689
rect 13868 17625 13932 17689
rect 13950 17625 14014 17689
rect 14032 17625 14096 17689
rect 14114 17625 14178 17689
rect 14196 17625 14260 17689
rect 14278 17625 14342 17689
rect 14360 17625 14424 17689
rect 14442 17625 14506 17689
rect 14524 17625 14588 17689
rect 14606 17625 14670 17689
rect 14688 17625 15000 17689
rect 14746 17607 15000 17625
rect 12231 17543 12295 17607
rect 12312 17543 12376 17607
rect 12393 17543 12457 17607
rect 12474 17543 12538 17607
rect 12556 17543 12620 17607
rect 12638 17543 12702 17607
rect 12720 17543 12784 17607
rect 12802 17543 12866 17607
rect 12884 17543 12948 17607
rect 12966 17543 13030 17607
rect 13048 17543 13112 17607
rect 13130 17543 13194 17607
rect 13212 17543 13276 17607
rect 13294 17543 13358 17607
rect 13376 17543 13440 17607
rect 13458 17543 13522 17607
rect 13540 17543 13604 17607
rect 13622 17543 13686 17607
rect 13704 17543 13768 17607
rect 13786 17543 13850 17607
rect 13868 17543 13932 17607
rect 13950 17543 14014 17607
rect 14032 17543 14096 17607
rect 14114 17543 14178 17607
rect 14196 17543 14260 17607
rect 14278 17543 14342 17607
rect 14360 17543 14424 17607
rect 14442 17543 14506 17607
rect 14524 17543 14588 17607
rect 14606 17543 14670 17607
rect 14688 17543 15000 17607
rect 14746 17525 15000 17543
rect 12231 17461 12295 17525
rect 12312 17461 12376 17525
rect 12393 17461 12457 17525
rect 12474 17461 12538 17525
rect 12556 17461 12620 17525
rect 12638 17461 12702 17525
rect 12720 17461 12784 17525
rect 12802 17461 12866 17525
rect 12884 17461 12948 17525
rect 12966 17461 13030 17525
rect 13048 17461 13112 17525
rect 13130 17461 13194 17525
rect 13212 17461 13276 17525
rect 13294 17461 13358 17525
rect 13376 17461 13440 17525
rect 13458 17461 13522 17525
rect 13540 17461 13604 17525
rect 13622 17461 13686 17525
rect 13704 17461 13768 17525
rect 13786 17461 13850 17525
rect 13868 17461 13932 17525
rect 13950 17461 14014 17525
rect 14032 17461 14096 17525
rect 14114 17461 14178 17525
rect 14196 17461 14260 17525
rect 14278 17461 14342 17525
rect 14360 17461 14424 17525
rect 14442 17461 14506 17525
rect 14524 17461 14588 17525
rect 14606 17461 14670 17525
rect 14688 17461 15000 17525
rect 14746 17443 15000 17461
rect 12231 17379 12295 17443
rect 12312 17379 12376 17443
rect 12393 17379 12457 17443
rect 12474 17379 12538 17443
rect 12556 17379 12620 17443
rect 12638 17379 12702 17443
rect 12720 17379 12784 17443
rect 12802 17379 12866 17443
rect 12884 17379 12948 17443
rect 12966 17379 13030 17443
rect 13048 17379 13112 17443
rect 13130 17379 13194 17443
rect 13212 17379 13276 17443
rect 13294 17379 13358 17443
rect 13376 17379 13440 17443
rect 13458 17379 13522 17443
rect 13540 17379 13604 17443
rect 13622 17379 13686 17443
rect 13704 17379 13768 17443
rect 13786 17379 13850 17443
rect 13868 17379 13932 17443
rect 13950 17379 14014 17443
rect 14032 17379 14096 17443
rect 14114 17379 14178 17443
rect 14196 17379 14260 17443
rect 14278 17379 14342 17443
rect 14360 17379 14424 17443
rect 14442 17379 14506 17443
rect 14524 17379 14588 17443
rect 14606 17379 14670 17443
rect 14688 17379 15000 17443
rect 14746 17361 15000 17379
rect 12231 17297 12295 17361
rect 12312 17297 12376 17361
rect 12393 17297 12457 17361
rect 12474 17297 12538 17361
rect 12556 17297 12620 17361
rect 12638 17297 12702 17361
rect 12720 17297 12784 17361
rect 12802 17297 12866 17361
rect 12884 17297 12948 17361
rect 12966 17297 13030 17361
rect 13048 17297 13112 17361
rect 13130 17297 13194 17361
rect 13212 17297 13276 17361
rect 13294 17297 13358 17361
rect 13376 17297 13440 17361
rect 13458 17297 13522 17361
rect 13540 17297 13604 17361
rect 13622 17297 13686 17361
rect 13704 17297 13768 17361
rect 13786 17297 13850 17361
rect 13868 17297 13932 17361
rect 13950 17297 14014 17361
rect 14032 17297 14096 17361
rect 14114 17297 14178 17361
rect 14196 17297 14260 17361
rect 14278 17297 14342 17361
rect 14360 17297 14424 17361
rect 14442 17297 14506 17361
rect 14524 17297 14588 17361
rect 14606 17297 14670 17361
rect 14688 17297 15000 17361
rect 14746 17279 15000 17297
rect 12231 17215 12295 17279
rect 12312 17215 12376 17279
rect 12393 17215 12457 17279
rect 12474 17215 12538 17279
rect 12556 17215 12620 17279
rect 12638 17215 12702 17279
rect 12720 17215 12784 17279
rect 12802 17215 12866 17279
rect 12884 17215 12948 17279
rect 12966 17215 13030 17279
rect 13048 17215 13112 17279
rect 13130 17215 13194 17279
rect 13212 17215 13276 17279
rect 13294 17215 13358 17279
rect 13376 17215 13440 17279
rect 13458 17215 13522 17279
rect 13540 17215 13604 17279
rect 13622 17215 13686 17279
rect 13704 17215 13768 17279
rect 13786 17215 13850 17279
rect 13868 17215 13932 17279
rect 13950 17215 14014 17279
rect 14032 17215 14096 17279
rect 14114 17215 14178 17279
rect 14196 17215 14260 17279
rect 14278 17215 14342 17279
rect 14360 17215 14424 17279
rect 14442 17215 14506 17279
rect 14524 17215 14588 17279
rect 14606 17215 14670 17279
rect 14688 17215 15000 17279
rect 14746 17197 15000 17215
rect 12231 17133 12295 17197
rect 12312 17133 12376 17197
rect 12393 17133 12457 17197
rect 12474 17133 12538 17197
rect 12556 17133 12620 17197
rect 12638 17133 12702 17197
rect 12720 17133 12784 17197
rect 12802 17133 12866 17197
rect 12884 17133 12948 17197
rect 12966 17133 13030 17197
rect 13048 17133 13112 17197
rect 13130 17133 13194 17197
rect 13212 17133 13276 17197
rect 13294 17133 13358 17197
rect 13376 17133 13440 17197
rect 13458 17133 13522 17197
rect 13540 17133 13604 17197
rect 13622 17133 13686 17197
rect 13704 17133 13768 17197
rect 13786 17133 13850 17197
rect 13868 17133 13932 17197
rect 13950 17133 14014 17197
rect 14032 17133 14096 17197
rect 14114 17133 14178 17197
rect 14196 17133 14260 17197
rect 14278 17133 14342 17197
rect 14360 17133 14424 17197
rect 14442 17133 14506 17197
rect 14524 17133 14588 17197
rect 14606 17133 14670 17197
rect 14688 17133 15000 17197
rect 14746 17115 15000 17133
rect 12231 17051 12295 17115
rect 12312 17051 12376 17115
rect 12393 17051 12457 17115
rect 12474 17051 12538 17115
rect 12556 17051 12620 17115
rect 12638 17051 12702 17115
rect 12720 17051 12784 17115
rect 12802 17051 12866 17115
rect 12884 17051 12948 17115
rect 12966 17051 13030 17115
rect 13048 17051 13112 17115
rect 13130 17051 13194 17115
rect 13212 17051 13276 17115
rect 13294 17051 13358 17115
rect 13376 17051 13440 17115
rect 13458 17051 13522 17115
rect 13540 17051 13604 17115
rect 13622 17051 13686 17115
rect 13704 17051 13768 17115
rect 13786 17051 13850 17115
rect 13868 17051 13932 17115
rect 13950 17051 14014 17115
rect 14032 17051 14096 17115
rect 14114 17051 14178 17115
rect 14196 17051 14260 17115
rect 14278 17051 14342 17115
rect 14360 17051 14424 17115
rect 14442 17051 14506 17115
rect 14524 17051 14588 17115
rect 14606 17051 14670 17115
rect 14688 17051 15000 17115
rect 14746 17033 15000 17051
rect 12231 16969 12295 17033
rect 12312 16969 12376 17033
rect 12393 16969 12457 17033
rect 12474 16969 12538 17033
rect 12556 16969 12620 17033
rect 12638 16969 12702 17033
rect 12720 16969 12784 17033
rect 12802 16969 12866 17033
rect 12884 16969 12948 17033
rect 12966 16969 13030 17033
rect 13048 16969 13112 17033
rect 13130 16969 13194 17033
rect 13212 16969 13276 17033
rect 13294 16969 13358 17033
rect 13376 16969 13440 17033
rect 13458 16969 13522 17033
rect 13540 16969 13604 17033
rect 13622 16969 13686 17033
rect 13704 16969 13768 17033
rect 13786 16969 13850 17033
rect 13868 16969 13932 17033
rect 13950 16969 14014 17033
rect 14032 16969 14096 17033
rect 14114 16969 14178 17033
rect 14196 16969 14260 17033
rect 14278 16969 14342 17033
rect 14360 16969 14424 17033
rect 14442 16969 14506 17033
rect 14524 16969 14588 17033
rect 14606 16969 14670 17033
rect 14688 16969 15000 17033
rect 14746 16951 15000 16969
rect 12231 16887 12295 16951
rect 12312 16887 12376 16951
rect 12393 16887 12457 16951
rect 12474 16887 12538 16951
rect 12556 16887 12620 16951
rect 12638 16887 12702 16951
rect 12720 16887 12784 16951
rect 12802 16887 12866 16951
rect 12884 16887 12948 16951
rect 12966 16887 13030 16951
rect 13048 16887 13112 16951
rect 13130 16887 13194 16951
rect 13212 16887 13276 16951
rect 13294 16887 13358 16951
rect 13376 16887 13440 16951
rect 13458 16887 13522 16951
rect 13540 16887 13604 16951
rect 13622 16887 13686 16951
rect 13704 16887 13768 16951
rect 13786 16887 13850 16951
rect 13868 16887 13932 16951
rect 13950 16887 14014 16951
rect 14032 16887 14096 16951
rect 14114 16887 14178 16951
rect 14196 16887 14260 16951
rect 14278 16887 14342 16951
rect 14360 16887 14424 16951
rect 14442 16887 14506 16951
rect 14524 16887 14588 16951
rect 14606 16887 14670 16951
rect 14688 16887 15000 16951
rect 14746 16869 15000 16887
rect 12231 16805 12295 16869
rect 12312 16805 12376 16869
rect 12393 16805 12457 16869
rect 12474 16805 12538 16869
rect 12556 16805 12620 16869
rect 12638 16805 12702 16869
rect 12720 16805 12784 16869
rect 12802 16805 12866 16869
rect 12884 16805 12948 16869
rect 12966 16805 13030 16869
rect 13048 16805 13112 16869
rect 13130 16805 13194 16869
rect 13212 16805 13276 16869
rect 13294 16805 13358 16869
rect 13376 16805 13440 16869
rect 13458 16805 13522 16869
rect 13540 16805 13604 16869
rect 13622 16805 13686 16869
rect 13704 16805 13768 16869
rect 13786 16805 13850 16869
rect 13868 16805 13932 16869
rect 13950 16805 14014 16869
rect 14032 16805 14096 16869
rect 14114 16805 14178 16869
rect 14196 16805 14260 16869
rect 14278 16805 14342 16869
rect 14360 16805 14424 16869
rect 14442 16805 14506 16869
rect 14524 16805 14588 16869
rect 14606 16805 14670 16869
rect 14688 16805 15000 16869
rect 14746 16787 15000 16805
rect 12231 16723 12295 16787
rect 12312 16723 12376 16787
rect 12393 16723 12457 16787
rect 12474 16723 12538 16787
rect 12556 16723 12620 16787
rect 12638 16723 12702 16787
rect 12720 16723 12784 16787
rect 12802 16723 12866 16787
rect 12884 16723 12948 16787
rect 12966 16723 13030 16787
rect 13048 16723 13112 16787
rect 13130 16723 13194 16787
rect 13212 16723 13276 16787
rect 13294 16723 13358 16787
rect 13376 16723 13440 16787
rect 13458 16723 13522 16787
rect 13540 16723 13604 16787
rect 13622 16723 13686 16787
rect 13704 16723 13768 16787
rect 13786 16723 13850 16787
rect 13868 16723 13932 16787
rect 13950 16723 14014 16787
rect 14032 16723 14096 16787
rect 14114 16723 14178 16787
rect 14196 16723 14260 16787
rect 14278 16723 14342 16787
rect 14360 16723 14424 16787
rect 14442 16723 14506 16787
rect 14524 16723 14588 16787
rect 14606 16723 14670 16787
rect 14688 16723 15000 16787
rect 14746 16705 15000 16723
rect 12231 16641 12295 16705
rect 12312 16641 12376 16705
rect 12393 16641 12457 16705
rect 12474 16641 12538 16705
rect 12556 16641 12620 16705
rect 12638 16641 12702 16705
rect 12720 16641 12784 16705
rect 12802 16641 12866 16705
rect 12884 16641 12948 16705
rect 12966 16641 13030 16705
rect 13048 16641 13112 16705
rect 13130 16641 13194 16705
rect 13212 16641 13276 16705
rect 13294 16641 13358 16705
rect 13376 16641 13440 16705
rect 13458 16641 13522 16705
rect 13540 16641 13604 16705
rect 13622 16641 13686 16705
rect 13704 16641 13768 16705
rect 13786 16641 13850 16705
rect 13868 16641 13932 16705
rect 13950 16641 14014 16705
rect 14032 16641 14096 16705
rect 14114 16641 14178 16705
rect 14196 16641 14260 16705
rect 14278 16641 14342 16705
rect 14360 16641 14424 16705
rect 14442 16641 14506 16705
rect 14524 16641 14588 16705
rect 14606 16641 14670 16705
rect 14688 16641 15000 16705
rect 14746 16623 15000 16641
rect 12231 16559 12295 16623
rect 12312 16559 12376 16623
rect 12393 16559 12457 16623
rect 12474 16559 12538 16623
rect 12556 16559 12620 16623
rect 12638 16559 12702 16623
rect 12720 16559 12784 16623
rect 12802 16559 12866 16623
rect 12884 16559 12948 16623
rect 12966 16559 13030 16623
rect 13048 16559 13112 16623
rect 13130 16559 13194 16623
rect 13212 16559 13276 16623
rect 13294 16559 13358 16623
rect 13376 16559 13440 16623
rect 13458 16559 13522 16623
rect 13540 16559 13604 16623
rect 13622 16559 13686 16623
rect 13704 16559 13768 16623
rect 13786 16559 13850 16623
rect 13868 16559 13932 16623
rect 13950 16559 14014 16623
rect 14032 16559 14096 16623
rect 14114 16559 14178 16623
rect 14196 16559 14260 16623
rect 14278 16559 14342 16623
rect 14360 16559 14424 16623
rect 14442 16559 14506 16623
rect 14524 16559 14588 16623
rect 14606 16559 14670 16623
rect 14688 16559 15000 16623
rect 0 16460 301 16524
rect 317 16460 381 16524
rect 397 16460 461 16524
rect 477 16460 541 16524
rect 557 16460 621 16524
rect 637 16460 701 16524
rect 717 16460 781 16524
rect 797 16460 861 16524
rect 877 16460 941 16524
rect 957 16460 1021 16524
rect 1037 16460 1101 16524
rect 1117 16460 1181 16524
rect 1197 16460 1261 16524
rect 1277 16460 1341 16524
rect 1357 16460 1421 16524
rect 1437 16460 1501 16524
rect 1517 16460 1581 16524
rect 1597 16460 1661 16524
rect 1677 16460 1741 16524
rect 1757 16460 1821 16524
rect 1837 16460 1901 16524
rect 1917 16460 1981 16524
rect 1997 16460 2061 16524
rect 2077 16460 2141 16524
rect 2157 16460 2221 16524
rect 2237 16460 2301 16524
rect 2317 16460 2381 16524
rect 2397 16460 2461 16524
rect 2477 16460 2541 16524
rect 2557 16460 2621 16524
rect 2637 16460 2701 16524
rect 2717 16460 2781 16524
rect 2797 16460 2861 16524
rect 2877 16460 2941 16524
rect 2957 16460 3021 16524
rect 3037 16460 3101 16524
rect 3117 16460 3181 16524
rect 3197 16460 3261 16524
rect 3277 16460 3341 16524
rect 3357 16460 3421 16524
rect 3437 16460 3501 16524
rect 3517 16460 3581 16524
rect 3597 16460 3661 16524
rect 3677 16460 3741 16524
rect 3757 16460 3821 16524
rect 3837 16460 3901 16524
rect 3917 16460 3981 16524
rect 3997 16460 4061 16524
rect 4077 16460 4141 16524
rect 4157 16460 4221 16524
rect 4237 16460 4301 16524
rect 4317 16460 4381 16524
rect 4397 16460 4461 16524
rect 4477 16460 4541 16524
rect 4557 16460 4621 16524
rect 4637 16460 4701 16524
rect 4717 16460 4781 16524
rect 4797 16460 4861 16524
rect 0 16443 254 16460
rect 0 16379 301 16443
rect 317 16379 381 16443
rect 397 16379 461 16443
rect 477 16379 541 16443
rect 557 16379 621 16443
rect 637 16379 701 16443
rect 717 16379 781 16443
rect 797 16379 861 16443
rect 877 16379 941 16443
rect 957 16379 1021 16443
rect 1037 16379 1101 16443
rect 1117 16379 1181 16443
rect 1197 16379 1261 16443
rect 1277 16379 1341 16443
rect 1357 16379 1421 16443
rect 1437 16379 1501 16443
rect 1517 16379 1581 16443
rect 1597 16379 1661 16443
rect 1677 16379 1741 16443
rect 1757 16379 1821 16443
rect 1837 16379 1901 16443
rect 1917 16379 1981 16443
rect 1997 16379 2061 16443
rect 2077 16379 2141 16443
rect 2157 16379 2221 16443
rect 2237 16379 2301 16443
rect 2317 16379 2381 16443
rect 2397 16379 2461 16443
rect 2477 16379 2541 16443
rect 2557 16379 2621 16443
rect 2637 16379 2701 16443
rect 2717 16379 2781 16443
rect 2797 16379 2861 16443
rect 2877 16379 2941 16443
rect 2957 16379 3021 16443
rect 3037 16379 3101 16443
rect 3117 16379 3181 16443
rect 3197 16379 3261 16443
rect 3277 16379 3341 16443
rect 3357 16379 3421 16443
rect 3437 16379 3501 16443
rect 3517 16379 3581 16443
rect 3597 16379 3661 16443
rect 3677 16379 3741 16443
rect 3757 16379 3821 16443
rect 3837 16379 3901 16443
rect 3917 16379 3981 16443
rect 3997 16379 4061 16443
rect 4077 16379 4141 16443
rect 4157 16379 4221 16443
rect 4237 16379 4301 16443
rect 4317 16379 4381 16443
rect 4397 16379 4461 16443
rect 4477 16379 4541 16443
rect 4557 16379 4621 16443
rect 4637 16379 4701 16443
rect 4717 16379 4781 16443
rect 4797 16379 4861 16443
rect 0 16362 254 16379
rect 0 16298 301 16362
rect 317 16298 381 16362
rect 397 16298 461 16362
rect 477 16298 541 16362
rect 557 16298 621 16362
rect 637 16298 701 16362
rect 717 16298 781 16362
rect 797 16298 861 16362
rect 877 16298 941 16362
rect 957 16298 1021 16362
rect 1037 16298 1101 16362
rect 1117 16298 1181 16362
rect 1197 16298 1261 16362
rect 1277 16298 1341 16362
rect 1357 16298 1421 16362
rect 1437 16298 1501 16362
rect 1517 16298 1581 16362
rect 1597 16298 1661 16362
rect 1677 16298 1741 16362
rect 1757 16298 1821 16362
rect 1837 16298 1901 16362
rect 1917 16298 1981 16362
rect 1997 16298 2061 16362
rect 2077 16298 2141 16362
rect 2157 16298 2221 16362
rect 2237 16298 2301 16362
rect 2317 16298 2381 16362
rect 2397 16298 2461 16362
rect 2477 16298 2541 16362
rect 2557 16298 2621 16362
rect 2637 16298 2701 16362
rect 2717 16298 2781 16362
rect 2797 16298 2861 16362
rect 2877 16298 2941 16362
rect 2957 16298 3021 16362
rect 3037 16298 3101 16362
rect 3117 16298 3181 16362
rect 3197 16298 3261 16362
rect 3277 16298 3341 16362
rect 3357 16298 3421 16362
rect 3437 16298 3501 16362
rect 3517 16298 3581 16362
rect 3597 16298 3661 16362
rect 3677 16298 3741 16362
rect 3757 16298 3821 16362
rect 3837 16298 3901 16362
rect 3917 16298 3981 16362
rect 3997 16298 4061 16362
rect 4077 16298 4141 16362
rect 4157 16298 4221 16362
rect 4237 16298 4301 16362
rect 4317 16298 4381 16362
rect 4397 16298 4461 16362
rect 4477 16298 4541 16362
rect 4557 16298 4621 16362
rect 4637 16298 4701 16362
rect 4717 16298 4781 16362
rect 4797 16298 4861 16362
rect 0 16281 254 16298
rect 0 16217 301 16281
rect 317 16217 381 16281
rect 397 16217 461 16281
rect 477 16217 541 16281
rect 557 16217 621 16281
rect 637 16217 701 16281
rect 717 16217 781 16281
rect 797 16217 861 16281
rect 877 16217 941 16281
rect 957 16217 1021 16281
rect 1037 16217 1101 16281
rect 1117 16217 1181 16281
rect 1197 16217 1261 16281
rect 1277 16217 1341 16281
rect 1357 16217 1421 16281
rect 1437 16217 1501 16281
rect 1517 16217 1581 16281
rect 1597 16217 1661 16281
rect 1677 16217 1741 16281
rect 1757 16217 1821 16281
rect 1837 16217 1901 16281
rect 1917 16217 1981 16281
rect 1997 16217 2061 16281
rect 2077 16217 2141 16281
rect 2157 16217 2221 16281
rect 2237 16217 2301 16281
rect 2317 16217 2381 16281
rect 2397 16217 2461 16281
rect 2477 16217 2541 16281
rect 2557 16217 2621 16281
rect 2637 16217 2701 16281
rect 2717 16217 2781 16281
rect 2797 16217 2861 16281
rect 2877 16217 2941 16281
rect 2957 16217 3021 16281
rect 3037 16217 3101 16281
rect 3117 16217 3181 16281
rect 3197 16217 3261 16281
rect 3277 16217 3341 16281
rect 3357 16217 3421 16281
rect 3437 16217 3501 16281
rect 3517 16217 3581 16281
rect 3597 16217 3661 16281
rect 3677 16217 3741 16281
rect 3757 16217 3821 16281
rect 3837 16217 3901 16281
rect 3917 16217 3981 16281
rect 3997 16217 4061 16281
rect 4077 16217 4141 16281
rect 4157 16217 4221 16281
rect 4237 16217 4301 16281
rect 4317 16217 4381 16281
rect 4397 16217 4461 16281
rect 4477 16217 4541 16281
rect 4557 16217 4621 16281
rect 4637 16217 4701 16281
rect 4717 16217 4781 16281
rect 4797 16217 4861 16281
rect 0 16200 254 16217
rect 0 16136 301 16200
rect 317 16136 381 16200
rect 397 16136 461 16200
rect 477 16136 541 16200
rect 557 16136 621 16200
rect 637 16136 701 16200
rect 717 16136 781 16200
rect 797 16136 861 16200
rect 877 16136 941 16200
rect 957 16136 1021 16200
rect 1037 16136 1101 16200
rect 1117 16136 1181 16200
rect 1197 16136 1261 16200
rect 1277 16136 1341 16200
rect 1357 16136 1421 16200
rect 1437 16136 1501 16200
rect 1517 16136 1581 16200
rect 1597 16136 1661 16200
rect 1677 16136 1741 16200
rect 1757 16136 1821 16200
rect 1837 16136 1901 16200
rect 1917 16136 1981 16200
rect 1997 16136 2061 16200
rect 2077 16136 2141 16200
rect 2157 16136 2221 16200
rect 2237 16136 2301 16200
rect 2317 16136 2381 16200
rect 2397 16136 2461 16200
rect 2477 16136 2541 16200
rect 2557 16136 2621 16200
rect 2637 16136 2701 16200
rect 2717 16136 2781 16200
rect 2797 16136 2861 16200
rect 2877 16136 2941 16200
rect 2957 16136 3021 16200
rect 3037 16136 3101 16200
rect 3117 16136 3181 16200
rect 3197 16136 3261 16200
rect 3277 16136 3341 16200
rect 3357 16136 3421 16200
rect 3437 16136 3501 16200
rect 3517 16136 3581 16200
rect 3597 16136 3661 16200
rect 3677 16136 3741 16200
rect 3757 16136 3821 16200
rect 3837 16136 3901 16200
rect 3917 16136 3981 16200
rect 3997 16136 4061 16200
rect 4077 16136 4141 16200
rect 4157 16136 4221 16200
rect 4237 16136 4301 16200
rect 4317 16136 4381 16200
rect 4397 16136 4461 16200
rect 4477 16136 4541 16200
rect 4557 16136 4621 16200
rect 4637 16136 4701 16200
rect 4717 16136 4781 16200
rect 4797 16136 4861 16200
rect 0 16119 254 16136
rect 0 16055 301 16119
rect 317 16055 381 16119
rect 397 16055 461 16119
rect 477 16055 541 16119
rect 557 16055 621 16119
rect 637 16055 701 16119
rect 717 16055 781 16119
rect 797 16055 861 16119
rect 877 16055 941 16119
rect 957 16055 1021 16119
rect 1037 16055 1101 16119
rect 1117 16055 1181 16119
rect 1197 16055 1261 16119
rect 1277 16055 1341 16119
rect 1357 16055 1421 16119
rect 1437 16055 1501 16119
rect 1517 16055 1581 16119
rect 1597 16055 1661 16119
rect 1677 16055 1741 16119
rect 1757 16055 1821 16119
rect 1837 16055 1901 16119
rect 1917 16055 1981 16119
rect 1997 16055 2061 16119
rect 2077 16055 2141 16119
rect 2157 16055 2221 16119
rect 2237 16055 2301 16119
rect 2317 16055 2381 16119
rect 2397 16055 2461 16119
rect 2477 16055 2541 16119
rect 2557 16055 2621 16119
rect 2637 16055 2701 16119
rect 2717 16055 2781 16119
rect 2797 16055 2861 16119
rect 2877 16055 2941 16119
rect 2957 16055 3021 16119
rect 3037 16055 3101 16119
rect 3117 16055 3181 16119
rect 3197 16055 3261 16119
rect 3277 16055 3341 16119
rect 3357 16055 3421 16119
rect 3437 16055 3501 16119
rect 3517 16055 3581 16119
rect 3597 16055 3661 16119
rect 3677 16055 3741 16119
rect 3757 16055 3821 16119
rect 3837 16055 3901 16119
rect 3917 16055 3981 16119
rect 3997 16055 4061 16119
rect 4077 16055 4141 16119
rect 4157 16055 4221 16119
rect 4237 16055 4301 16119
rect 4317 16055 4381 16119
rect 4397 16055 4461 16119
rect 4477 16055 4541 16119
rect 4557 16055 4621 16119
rect 4637 16055 4701 16119
rect 4717 16055 4781 16119
rect 4797 16055 4861 16119
rect 0 16038 254 16055
rect 0 15974 301 16038
rect 317 15974 381 16038
rect 397 15974 461 16038
rect 477 15974 541 16038
rect 557 15974 621 16038
rect 637 15974 701 16038
rect 717 15974 781 16038
rect 797 15974 861 16038
rect 877 15974 941 16038
rect 957 15974 1021 16038
rect 1037 15974 1101 16038
rect 1117 15974 1181 16038
rect 1197 15974 1261 16038
rect 1277 15974 1341 16038
rect 1357 15974 1421 16038
rect 1437 15974 1501 16038
rect 1517 15974 1581 16038
rect 1597 15974 1661 16038
rect 1677 15974 1741 16038
rect 1757 15974 1821 16038
rect 1837 15974 1901 16038
rect 1917 15974 1981 16038
rect 1997 15974 2061 16038
rect 2077 15974 2141 16038
rect 2157 15974 2221 16038
rect 2237 15974 2301 16038
rect 2317 15974 2381 16038
rect 2397 15974 2461 16038
rect 2477 15974 2541 16038
rect 2557 15974 2621 16038
rect 2637 15974 2701 16038
rect 2717 15974 2781 16038
rect 2797 15974 2861 16038
rect 2877 15974 2941 16038
rect 2957 15974 3021 16038
rect 3037 15974 3101 16038
rect 3117 15974 3181 16038
rect 3197 15974 3261 16038
rect 3277 15974 3341 16038
rect 3357 15974 3421 16038
rect 3437 15974 3501 16038
rect 3517 15974 3581 16038
rect 3597 15974 3661 16038
rect 3677 15974 3741 16038
rect 3757 15974 3821 16038
rect 3837 15974 3901 16038
rect 3917 15974 3981 16038
rect 3997 15974 4061 16038
rect 4077 15974 4141 16038
rect 4157 15974 4221 16038
rect 4237 15974 4301 16038
rect 4317 15974 4381 16038
rect 4397 15974 4461 16038
rect 4477 15974 4541 16038
rect 4557 15974 4621 16038
rect 4637 15974 4701 16038
rect 4717 15974 4781 16038
rect 4797 15974 4861 16038
rect 0 15957 254 15974
rect 0 15893 301 15957
rect 317 15893 381 15957
rect 397 15893 461 15957
rect 477 15893 541 15957
rect 557 15893 621 15957
rect 637 15893 701 15957
rect 717 15893 781 15957
rect 797 15893 861 15957
rect 877 15893 941 15957
rect 957 15893 1021 15957
rect 1037 15893 1101 15957
rect 1117 15893 1181 15957
rect 1197 15893 1261 15957
rect 1277 15893 1341 15957
rect 1357 15893 1421 15957
rect 1437 15893 1501 15957
rect 1517 15893 1581 15957
rect 1597 15893 1661 15957
rect 1677 15893 1741 15957
rect 1757 15893 1821 15957
rect 1837 15893 1901 15957
rect 1917 15893 1981 15957
rect 1997 15893 2061 15957
rect 2077 15893 2141 15957
rect 2157 15893 2221 15957
rect 2237 15893 2301 15957
rect 2317 15893 2381 15957
rect 2397 15893 2461 15957
rect 2477 15893 2541 15957
rect 2557 15893 2621 15957
rect 2637 15893 2701 15957
rect 2717 15893 2781 15957
rect 2797 15893 2861 15957
rect 2877 15893 2941 15957
rect 2957 15893 3021 15957
rect 3037 15893 3101 15957
rect 3117 15893 3181 15957
rect 3197 15893 3261 15957
rect 3277 15893 3341 15957
rect 3357 15893 3421 15957
rect 3437 15893 3501 15957
rect 3517 15893 3581 15957
rect 3597 15893 3661 15957
rect 3677 15893 3741 15957
rect 3757 15893 3821 15957
rect 3837 15893 3901 15957
rect 3917 15893 3981 15957
rect 3997 15893 4061 15957
rect 4077 15893 4141 15957
rect 4157 15893 4221 15957
rect 4237 15893 4301 15957
rect 4317 15893 4381 15957
rect 4397 15893 4461 15957
rect 4477 15893 4541 15957
rect 4557 15893 4621 15957
rect 4637 15893 4701 15957
rect 4717 15893 4781 15957
rect 4797 15893 4861 15957
rect 0 15876 254 15893
rect 0 15812 301 15876
rect 317 15812 381 15876
rect 397 15812 461 15876
rect 477 15812 541 15876
rect 557 15812 621 15876
rect 637 15812 701 15876
rect 717 15812 781 15876
rect 797 15812 861 15876
rect 877 15812 941 15876
rect 957 15812 1021 15876
rect 1037 15812 1101 15876
rect 1117 15812 1181 15876
rect 1197 15812 1261 15876
rect 1277 15812 1341 15876
rect 1357 15812 1421 15876
rect 1437 15812 1501 15876
rect 1517 15812 1581 15876
rect 1597 15812 1661 15876
rect 1677 15812 1741 15876
rect 1757 15812 1821 15876
rect 1837 15812 1901 15876
rect 1917 15812 1981 15876
rect 1997 15812 2061 15876
rect 2077 15812 2141 15876
rect 2157 15812 2221 15876
rect 2237 15812 2301 15876
rect 2317 15812 2381 15876
rect 2397 15812 2461 15876
rect 2477 15812 2541 15876
rect 2557 15812 2621 15876
rect 2637 15812 2701 15876
rect 2717 15812 2781 15876
rect 2797 15812 2861 15876
rect 2877 15812 2941 15876
rect 2957 15812 3021 15876
rect 3037 15812 3101 15876
rect 3117 15812 3181 15876
rect 3197 15812 3261 15876
rect 3277 15812 3341 15876
rect 3357 15812 3421 15876
rect 3437 15812 3501 15876
rect 3517 15812 3581 15876
rect 3597 15812 3661 15876
rect 3677 15812 3741 15876
rect 3757 15812 3821 15876
rect 3837 15812 3901 15876
rect 3917 15812 3981 15876
rect 3997 15812 4061 15876
rect 4077 15812 4141 15876
rect 4157 15812 4221 15876
rect 4237 15812 4301 15876
rect 4317 15812 4381 15876
rect 4397 15812 4461 15876
rect 4477 15812 4541 15876
rect 4557 15812 4621 15876
rect 4637 15812 4701 15876
rect 4717 15812 4781 15876
rect 4797 15812 4861 15876
rect 0 15795 254 15812
rect 0 15731 301 15795
rect 317 15731 381 15795
rect 397 15731 461 15795
rect 477 15731 541 15795
rect 557 15731 621 15795
rect 637 15731 701 15795
rect 717 15731 781 15795
rect 797 15731 861 15795
rect 877 15731 941 15795
rect 957 15731 1021 15795
rect 1037 15731 1101 15795
rect 1117 15731 1181 15795
rect 1197 15731 1261 15795
rect 1277 15731 1341 15795
rect 1357 15731 1421 15795
rect 1437 15731 1501 15795
rect 1517 15731 1581 15795
rect 1597 15731 1661 15795
rect 1677 15731 1741 15795
rect 1757 15731 1821 15795
rect 1837 15731 1901 15795
rect 1917 15731 1981 15795
rect 1997 15731 2061 15795
rect 2077 15731 2141 15795
rect 2157 15731 2221 15795
rect 2237 15731 2301 15795
rect 2317 15731 2381 15795
rect 2397 15731 2461 15795
rect 2477 15731 2541 15795
rect 2557 15731 2621 15795
rect 2637 15731 2701 15795
rect 2717 15731 2781 15795
rect 2797 15731 2861 15795
rect 2877 15731 2941 15795
rect 2957 15731 3021 15795
rect 3037 15731 3101 15795
rect 3117 15731 3181 15795
rect 3197 15731 3261 15795
rect 3277 15731 3341 15795
rect 3357 15731 3421 15795
rect 3437 15731 3501 15795
rect 3517 15731 3581 15795
rect 3597 15731 3661 15795
rect 3677 15731 3741 15795
rect 3757 15731 3821 15795
rect 3837 15731 3901 15795
rect 3917 15731 3981 15795
rect 3997 15731 4061 15795
rect 4077 15731 4141 15795
rect 4157 15731 4221 15795
rect 4237 15731 4301 15795
rect 4317 15731 4381 15795
rect 4397 15731 4461 15795
rect 4477 15731 4541 15795
rect 4557 15731 4621 15795
rect 4637 15731 4701 15795
rect 4717 15731 4781 15795
rect 4797 15731 4861 15795
rect 0 15714 254 15731
rect 0 15650 301 15714
rect 317 15650 381 15714
rect 397 15650 461 15714
rect 477 15650 541 15714
rect 557 15650 621 15714
rect 637 15650 701 15714
rect 717 15650 781 15714
rect 797 15650 861 15714
rect 877 15650 941 15714
rect 957 15650 1021 15714
rect 1037 15650 1101 15714
rect 1117 15650 1181 15714
rect 1197 15650 1261 15714
rect 1277 15650 1341 15714
rect 1357 15650 1421 15714
rect 1437 15650 1501 15714
rect 1517 15650 1581 15714
rect 1597 15650 1661 15714
rect 1677 15650 1741 15714
rect 1757 15650 1821 15714
rect 1837 15650 1901 15714
rect 1917 15650 1981 15714
rect 1997 15650 2061 15714
rect 2077 15650 2141 15714
rect 2157 15650 2221 15714
rect 2237 15650 2301 15714
rect 2317 15650 2381 15714
rect 2397 15650 2461 15714
rect 2477 15650 2541 15714
rect 2557 15650 2621 15714
rect 2637 15650 2701 15714
rect 2717 15650 2781 15714
rect 2797 15650 2861 15714
rect 2877 15650 2941 15714
rect 2957 15650 3021 15714
rect 3037 15650 3101 15714
rect 3117 15650 3181 15714
rect 3197 15650 3261 15714
rect 3277 15650 3341 15714
rect 3357 15650 3421 15714
rect 3437 15650 3501 15714
rect 3517 15650 3581 15714
rect 3597 15650 3661 15714
rect 3677 15650 3741 15714
rect 3757 15650 3821 15714
rect 3837 15650 3901 15714
rect 3917 15650 3981 15714
rect 3997 15650 4061 15714
rect 4077 15650 4141 15714
rect 4157 15650 4221 15714
rect 4237 15650 4301 15714
rect 4317 15650 4381 15714
rect 4397 15650 4461 15714
rect 4477 15650 4541 15714
rect 4557 15650 4621 15714
rect 4637 15650 4701 15714
rect 4717 15650 4781 15714
rect 4797 15650 4861 15714
rect 0 15633 254 15650
rect 0 15569 301 15633
rect 317 15569 381 15633
rect 397 15569 461 15633
rect 477 15569 541 15633
rect 557 15569 621 15633
rect 637 15569 701 15633
rect 717 15569 781 15633
rect 797 15569 861 15633
rect 877 15569 941 15633
rect 957 15569 1021 15633
rect 1037 15569 1101 15633
rect 1117 15569 1181 15633
rect 1197 15569 1261 15633
rect 1277 15569 1341 15633
rect 1357 15569 1421 15633
rect 1437 15569 1501 15633
rect 1517 15569 1581 15633
rect 1597 15569 1661 15633
rect 1677 15569 1741 15633
rect 1757 15569 1821 15633
rect 1837 15569 1901 15633
rect 1917 15569 1981 15633
rect 1997 15569 2061 15633
rect 2077 15569 2141 15633
rect 2157 15569 2221 15633
rect 2237 15569 2301 15633
rect 2317 15569 2381 15633
rect 2397 15569 2461 15633
rect 2477 15569 2541 15633
rect 2557 15569 2621 15633
rect 2637 15569 2701 15633
rect 2717 15569 2781 15633
rect 2797 15569 2861 15633
rect 2877 15569 2941 15633
rect 2957 15569 3021 15633
rect 3037 15569 3101 15633
rect 3117 15569 3181 15633
rect 3197 15569 3261 15633
rect 3277 15569 3341 15633
rect 3357 15569 3421 15633
rect 3437 15569 3501 15633
rect 3517 15569 3581 15633
rect 3597 15569 3661 15633
rect 3677 15569 3741 15633
rect 3757 15569 3821 15633
rect 3837 15569 3901 15633
rect 3917 15569 3981 15633
rect 3997 15569 4061 15633
rect 4077 15569 4141 15633
rect 4157 15569 4221 15633
rect 4237 15569 4301 15633
rect 4317 15569 4381 15633
rect 4397 15569 4461 15633
rect 4477 15569 4541 15633
rect 4557 15569 4621 15633
rect 4637 15569 4701 15633
rect 4717 15569 4781 15633
rect 4797 15569 4861 15633
rect 0 15552 254 15569
rect 0 15488 301 15552
rect 317 15488 381 15552
rect 397 15488 461 15552
rect 477 15488 541 15552
rect 557 15488 621 15552
rect 637 15488 701 15552
rect 717 15488 781 15552
rect 797 15488 861 15552
rect 877 15488 941 15552
rect 957 15488 1021 15552
rect 1037 15488 1101 15552
rect 1117 15488 1181 15552
rect 1197 15488 1261 15552
rect 1277 15488 1341 15552
rect 1357 15488 1421 15552
rect 1437 15488 1501 15552
rect 1517 15488 1581 15552
rect 1597 15488 1661 15552
rect 1677 15488 1741 15552
rect 1757 15488 1821 15552
rect 1837 15488 1901 15552
rect 1917 15488 1981 15552
rect 1997 15488 2061 15552
rect 2077 15488 2141 15552
rect 2157 15488 2221 15552
rect 2237 15488 2301 15552
rect 2317 15488 2381 15552
rect 2397 15488 2461 15552
rect 2477 15488 2541 15552
rect 2557 15488 2621 15552
rect 2637 15488 2701 15552
rect 2717 15488 2781 15552
rect 2797 15488 2861 15552
rect 2877 15488 2941 15552
rect 2957 15488 3021 15552
rect 3037 15488 3101 15552
rect 3117 15488 3181 15552
rect 3197 15488 3261 15552
rect 3277 15488 3341 15552
rect 3357 15488 3421 15552
rect 3437 15488 3501 15552
rect 3517 15488 3581 15552
rect 3597 15488 3661 15552
rect 3677 15488 3741 15552
rect 3757 15488 3821 15552
rect 3837 15488 3901 15552
rect 3917 15488 3981 15552
rect 3997 15488 4061 15552
rect 4077 15488 4141 15552
rect 4157 15488 4221 15552
rect 4237 15488 4301 15552
rect 4317 15488 4381 15552
rect 4397 15488 4461 15552
rect 4477 15488 4541 15552
rect 4557 15488 4621 15552
rect 4637 15488 4701 15552
rect 4717 15488 4781 15552
rect 4797 15488 4861 15552
rect 0 15471 254 15488
rect 0 15407 301 15471
rect 317 15407 381 15471
rect 397 15407 461 15471
rect 477 15407 541 15471
rect 557 15407 621 15471
rect 637 15407 701 15471
rect 717 15407 781 15471
rect 797 15407 861 15471
rect 877 15407 941 15471
rect 957 15407 1021 15471
rect 1037 15407 1101 15471
rect 1117 15407 1181 15471
rect 1197 15407 1261 15471
rect 1277 15407 1341 15471
rect 1357 15407 1421 15471
rect 1437 15407 1501 15471
rect 1517 15407 1581 15471
rect 1597 15407 1661 15471
rect 1677 15407 1741 15471
rect 1757 15407 1821 15471
rect 1837 15407 1901 15471
rect 1917 15407 1981 15471
rect 1997 15407 2061 15471
rect 2077 15407 2141 15471
rect 2157 15407 2221 15471
rect 2237 15407 2301 15471
rect 2317 15407 2381 15471
rect 2397 15407 2461 15471
rect 2477 15407 2541 15471
rect 2557 15407 2621 15471
rect 2637 15407 2701 15471
rect 2717 15407 2781 15471
rect 2797 15407 2861 15471
rect 2877 15407 2941 15471
rect 2957 15407 3021 15471
rect 3037 15407 3101 15471
rect 3117 15407 3181 15471
rect 3197 15407 3261 15471
rect 3277 15407 3341 15471
rect 3357 15407 3421 15471
rect 3437 15407 3501 15471
rect 3517 15407 3581 15471
rect 3597 15407 3661 15471
rect 3677 15407 3741 15471
rect 3757 15407 3821 15471
rect 3837 15407 3901 15471
rect 3917 15407 3981 15471
rect 3997 15407 4061 15471
rect 4077 15407 4141 15471
rect 4157 15407 4221 15471
rect 4237 15407 4301 15471
rect 4317 15407 4381 15471
rect 4397 15407 4461 15471
rect 4477 15407 4541 15471
rect 4557 15407 4621 15471
rect 4637 15407 4701 15471
rect 4717 15407 4781 15471
rect 4797 15407 4861 15471
rect 0 15390 254 15407
rect 0 15326 301 15390
rect 317 15326 381 15390
rect 397 15326 461 15390
rect 477 15326 541 15390
rect 557 15326 621 15390
rect 637 15326 701 15390
rect 717 15326 781 15390
rect 797 15326 861 15390
rect 877 15326 941 15390
rect 957 15326 1021 15390
rect 1037 15326 1101 15390
rect 1117 15326 1181 15390
rect 1197 15326 1261 15390
rect 1277 15326 1341 15390
rect 1357 15326 1421 15390
rect 1437 15326 1501 15390
rect 1517 15326 1581 15390
rect 1597 15326 1661 15390
rect 1677 15326 1741 15390
rect 1757 15326 1821 15390
rect 1837 15326 1901 15390
rect 1917 15326 1981 15390
rect 1997 15326 2061 15390
rect 2077 15326 2141 15390
rect 2157 15326 2221 15390
rect 2237 15326 2301 15390
rect 2317 15326 2381 15390
rect 2397 15326 2461 15390
rect 2477 15326 2541 15390
rect 2557 15326 2621 15390
rect 2637 15326 2701 15390
rect 2717 15326 2781 15390
rect 2797 15326 2861 15390
rect 2877 15326 2941 15390
rect 2957 15326 3021 15390
rect 3037 15326 3101 15390
rect 3117 15326 3181 15390
rect 3197 15326 3261 15390
rect 3277 15326 3341 15390
rect 3357 15326 3421 15390
rect 3437 15326 3501 15390
rect 3517 15326 3581 15390
rect 3597 15326 3661 15390
rect 3677 15326 3741 15390
rect 3757 15326 3821 15390
rect 3837 15326 3901 15390
rect 3917 15326 3981 15390
rect 3997 15326 4061 15390
rect 4077 15326 4141 15390
rect 4157 15326 4221 15390
rect 4237 15326 4301 15390
rect 4317 15326 4381 15390
rect 4397 15326 4461 15390
rect 4477 15326 4541 15390
rect 4557 15326 4621 15390
rect 4637 15326 4701 15390
rect 4717 15326 4781 15390
rect 4797 15326 4861 15390
rect 0 15309 254 15326
rect 0 15245 301 15309
rect 317 15245 381 15309
rect 397 15245 461 15309
rect 477 15245 541 15309
rect 557 15245 621 15309
rect 637 15245 701 15309
rect 717 15245 781 15309
rect 797 15245 861 15309
rect 877 15245 941 15309
rect 957 15245 1021 15309
rect 1037 15245 1101 15309
rect 1117 15245 1181 15309
rect 1197 15245 1261 15309
rect 1277 15245 1341 15309
rect 1357 15245 1421 15309
rect 1437 15245 1501 15309
rect 1517 15245 1581 15309
rect 1597 15245 1661 15309
rect 1677 15245 1741 15309
rect 1757 15245 1821 15309
rect 1837 15245 1901 15309
rect 1917 15245 1981 15309
rect 1997 15245 2061 15309
rect 2077 15245 2141 15309
rect 2157 15245 2221 15309
rect 2237 15245 2301 15309
rect 2317 15245 2381 15309
rect 2397 15245 2461 15309
rect 2477 15245 2541 15309
rect 2557 15245 2621 15309
rect 2637 15245 2701 15309
rect 2717 15245 2781 15309
rect 2797 15245 2861 15309
rect 2877 15245 2941 15309
rect 2957 15245 3021 15309
rect 3037 15245 3101 15309
rect 3117 15245 3181 15309
rect 3197 15245 3261 15309
rect 3277 15245 3341 15309
rect 3357 15245 3421 15309
rect 3437 15245 3501 15309
rect 3517 15245 3581 15309
rect 3597 15245 3661 15309
rect 3677 15245 3741 15309
rect 3757 15245 3821 15309
rect 3837 15245 3901 15309
rect 3917 15245 3981 15309
rect 3997 15245 4061 15309
rect 4077 15245 4141 15309
rect 4157 15245 4221 15309
rect 4237 15245 4301 15309
rect 4317 15245 4381 15309
rect 4397 15245 4461 15309
rect 4477 15245 4541 15309
rect 4557 15245 4621 15309
rect 4637 15245 4701 15309
rect 4717 15245 4781 15309
rect 4797 15245 4861 15309
rect 0 15228 254 15245
rect 0 15164 301 15228
rect 317 15164 381 15228
rect 397 15164 461 15228
rect 477 15164 541 15228
rect 557 15164 621 15228
rect 637 15164 701 15228
rect 717 15164 781 15228
rect 797 15164 861 15228
rect 877 15164 941 15228
rect 957 15164 1021 15228
rect 1037 15164 1101 15228
rect 1117 15164 1181 15228
rect 1197 15164 1261 15228
rect 1277 15164 1341 15228
rect 1357 15164 1421 15228
rect 1437 15164 1501 15228
rect 1517 15164 1581 15228
rect 1597 15164 1661 15228
rect 1677 15164 1741 15228
rect 1757 15164 1821 15228
rect 1837 15164 1901 15228
rect 1917 15164 1981 15228
rect 1997 15164 2061 15228
rect 2077 15164 2141 15228
rect 2157 15164 2221 15228
rect 2237 15164 2301 15228
rect 2317 15164 2381 15228
rect 2397 15164 2461 15228
rect 2477 15164 2541 15228
rect 2557 15164 2621 15228
rect 2637 15164 2701 15228
rect 2717 15164 2781 15228
rect 2797 15164 2861 15228
rect 2877 15164 2941 15228
rect 2957 15164 3021 15228
rect 3037 15164 3101 15228
rect 3117 15164 3181 15228
rect 3197 15164 3261 15228
rect 3277 15164 3341 15228
rect 3357 15164 3421 15228
rect 3437 15164 3501 15228
rect 3517 15164 3581 15228
rect 3597 15164 3661 15228
rect 3677 15164 3741 15228
rect 3757 15164 3821 15228
rect 3837 15164 3901 15228
rect 3917 15164 3981 15228
rect 3997 15164 4061 15228
rect 4077 15164 4141 15228
rect 4157 15164 4221 15228
rect 4237 15164 4301 15228
rect 4317 15164 4381 15228
rect 4397 15164 4461 15228
rect 4477 15164 4541 15228
rect 4557 15164 4621 15228
rect 4637 15164 4701 15228
rect 4717 15164 4781 15228
rect 4797 15164 4861 15228
rect 0 15147 254 15164
rect 0 15083 301 15147
rect 317 15083 381 15147
rect 397 15083 461 15147
rect 477 15083 541 15147
rect 557 15083 621 15147
rect 637 15083 701 15147
rect 717 15083 781 15147
rect 797 15083 861 15147
rect 877 15083 941 15147
rect 957 15083 1021 15147
rect 1037 15083 1101 15147
rect 1117 15083 1181 15147
rect 1197 15083 1261 15147
rect 1277 15083 1341 15147
rect 1357 15083 1421 15147
rect 1437 15083 1501 15147
rect 1517 15083 1581 15147
rect 1597 15083 1661 15147
rect 1677 15083 1741 15147
rect 1757 15083 1821 15147
rect 1837 15083 1901 15147
rect 1917 15083 1981 15147
rect 1997 15083 2061 15147
rect 2077 15083 2141 15147
rect 2157 15083 2221 15147
rect 2237 15083 2301 15147
rect 2317 15083 2381 15147
rect 2397 15083 2461 15147
rect 2477 15083 2541 15147
rect 2557 15083 2621 15147
rect 2637 15083 2701 15147
rect 2717 15083 2781 15147
rect 2797 15083 2861 15147
rect 2877 15083 2941 15147
rect 2957 15083 3021 15147
rect 3037 15083 3101 15147
rect 3117 15083 3181 15147
rect 3197 15083 3261 15147
rect 3277 15083 3341 15147
rect 3357 15083 3421 15147
rect 3437 15083 3501 15147
rect 3517 15083 3581 15147
rect 3597 15083 3661 15147
rect 3677 15083 3741 15147
rect 3757 15083 3821 15147
rect 3837 15083 3901 15147
rect 3917 15083 3981 15147
rect 3997 15083 4061 15147
rect 4077 15083 4141 15147
rect 4157 15083 4221 15147
rect 4237 15083 4301 15147
rect 4317 15083 4381 15147
rect 4397 15083 4461 15147
rect 4477 15083 4541 15147
rect 4557 15083 4621 15147
rect 4637 15083 4701 15147
rect 4717 15083 4781 15147
rect 4797 15083 4861 15147
rect 0 15066 254 15083
rect 0 15002 301 15066
rect 317 15002 381 15066
rect 397 15002 461 15066
rect 477 15002 541 15066
rect 557 15002 621 15066
rect 637 15002 701 15066
rect 717 15002 781 15066
rect 797 15002 861 15066
rect 877 15002 941 15066
rect 957 15002 1021 15066
rect 1037 15002 1101 15066
rect 1117 15002 1181 15066
rect 1197 15002 1261 15066
rect 1277 15002 1341 15066
rect 1357 15002 1421 15066
rect 1437 15002 1501 15066
rect 1517 15002 1581 15066
rect 1597 15002 1661 15066
rect 1677 15002 1741 15066
rect 1757 15002 1821 15066
rect 1837 15002 1901 15066
rect 1917 15002 1981 15066
rect 1997 15002 2061 15066
rect 2077 15002 2141 15066
rect 2157 15002 2221 15066
rect 2237 15002 2301 15066
rect 2317 15002 2381 15066
rect 2397 15002 2461 15066
rect 2477 15002 2541 15066
rect 2557 15002 2621 15066
rect 2637 15002 2701 15066
rect 2717 15002 2781 15066
rect 2797 15002 2861 15066
rect 2877 15002 2941 15066
rect 2957 15002 3021 15066
rect 3037 15002 3101 15066
rect 3117 15002 3181 15066
rect 3197 15002 3261 15066
rect 3277 15002 3341 15066
rect 3357 15002 3421 15066
rect 3437 15002 3501 15066
rect 3517 15002 3581 15066
rect 3597 15002 3661 15066
rect 3677 15002 3741 15066
rect 3757 15002 3821 15066
rect 3837 15002 3901 15066
rect 3917 15002 3981 15066
rect 3997 15002 4061 15066
rect 4077 15002 4141 15066
rect 4157 15002 4221 15066
rect 4237 15002 4301 15066
rect 4317 15002 4381 15066
rect 4397 15002 4461 15066
rect 4477 15002 4541 15066
rect 4557 15002 4621 15066
rect 4637 15002 4701 15066
rect 4717 15002 4781 15066
rect 4797 15002 4861 15066
rect 0 14985 254 15002
rect 0 14921 301 14985
rect 317 14921 381 14985
rect 397 14921 461 14985
rect 477 14921 541 14985
rect 557 14921 621 14985
rect 637 14921 701 14985
rect 717 14921 781 14985
rect 797 14921 861 14985
rect 877 14921 941 14985
rect 957 14921 1021 14985
rect 1037 14921 1101 14985
rect 1117 14921 1181 14985
rect 1197 14921 1261 14985
rect 1277 14921 1341 14985
rect 1357 14921 1421 14985
rect 1437 14921 1501 14985
rect 1517 14921 1581 14985
rect 1597 14921 1661 14985
rect 1677 14921 1741 14985
rect 1757 14921 1821 14985
rect 1837 14921 1901 14985
rect 1917 14921 1981 14985
rect 1997 14921 2061 14985
rect 2077 14921 2141 14985
rect 2157 14921 2221 14985
rect 2237 14921 2301 14985
rect 2317 14921 2381 14985
rect 2397 14921 2461 14985
rect 2477 14921 2541 14985
rect 2557 14921 2621 14985
rect 2637 14921 2701 14985
rect 2717 14921 2781 14985
rect 2797 14921 2861 14985
rect 2877 14921 2941 14985
rect 2957 14921 3021 14985
rect 3037 14921 3101 14985
rect 3117 14921 3181 14985
rect 3197 14921 3261 14985
rect 3277 14921 3341 14985
rect 3357 14921 3421 14985
rect 3437 14921 3501 14985
rect 3517 14921 3581 14985
rect 3597 14921 3661 14985
rect 3677 14921 3741 14985
rect 3757 14921 3821 14985
rect 3837 14921 3901 14985
rect 3917 14921 3981 14985
rect 3997 14921 4061 14985
rect 4077 14921 4141 14985
rect 4157 14921 4221 14985
rect 4237 14921 4301 14985
rect 4317 14921 4381 14985
rect 4397 14921 4461 14985
rect 4477 14921 4541 14985
rect 4557 14921 4621 14985
rect 4637 14921 4701 14985
rect 4717 14921 4781 14985
rect 4797 14921 4861 14985
rect 0 14904 254 14921
rect 0 14840 301 14904
rect 317 14840 381 14904
rect 397 14840 461 14904
rect 477 14840 541 14904
rect 557 14840 621 14904
rect 637 14840 701 14904
rect 717 14840 781 14904
rect 797 14840 861 14904
rect 877 14840 941 14904
rect 957 14840 1021 14904
rect 1037 14840 1101 14904
rect 1117 14840 1181 14904
rect 1197 14840 1261 14904
rect 1277 14840 1341 14904
rect 1357 14840 1421 14904
rect 1437 14840 1501 14904
rect 1517 14840 1581 14904
rect 1597 14840 1661 14904
rect 1677 14840 1741 14904
rect 1757 14840 1821 14904
rect 1837 14840 1901 14904
rect 1917 14840 1981 14904
rect 1997 14840 2061 14904
rect 2077 14840 2141 14904
rect 2157 14840 2221 14904
rect 2237 14840 2301 14904
rect 2317 14840 2381 14904
rect 2397 14840 2461 14904
rect 2477 14840 2541 14904
rect 2557 14840 2621 14904
rect 2637 14840 2701 14904
rect 2717 14840 2781 14904
rect 2797 14840 2861 14904
rect 2877 14840 2941 14904
rect 2957 14840 3021 14904
rect 3037 14840 3101 14904
rect 3117 14840 3181 14904
rect 3197 14840 3261 14904
rect 3277 14840 3341 14904
rect 3357 14840 3421 14904
rect 3437 14840 3501 14904
rect 3517 14840 3581 14904
rect 3597 14840 3661 14904
rect 3677 14840 3741 14904
rect 3757 14840 3821 14904
rect 3837 14840 3901 14904
rect 3917 14840 3981 14904
rect 3997 14840 4061 14904
rect 4077 14840 4141 14904
rect 4157 14840 4221 14904
rect 4237 14840 4301 14904
rect 4317 14840 4381 14904
rect 4397 14840 4461 14904
rect 4477 14840 4541 14904
rect 4557 14840 4621 14904
rect 4637 14840 4701 14904
rect 4717 14840 4781 14904
rect 4797 14840 4861 14904
rect 0 14823 254 14840
rect 0 14759 301 14823
rect 317 14759 381 14823
rect 397 14759 461 14823
rect 477 14759 541 14823
rect 557 14759 621 14823
rect 637 14759 701 14823
rect 717 14759 781 14823
rect 797 14759 861 14823
rect 877 14759 941 14823
rect 957 14759 1021 14823
rect 1037 14759 1101 14823
rect 1117 14759 1181 14823
rect 1197 14759 1261 14823
rect 1277 14759 1341 14823
rect 1357 14759 1421 14823
rect 1437 14759 1501 14823
rect 1517 14759 1581 14823
rect 1597 14759 1661 14823
rect 1677 14759 1741 14823
rect 1757 14759 1821 14823
rect 1837 14759 1901 14823
rect 1917 14759 1981 14823
rect 1997 14759 2061 14823
rect 2077 14759 2141 14823
rect 2157 14759 2221 14823
rect 2237 14759 2301 14823
rect 2317 14759 2381 14823
rect 2397 14759 2461 14823
rect 2477 14759 2541 14823
rect 2557 14759 2621 14823
rect 2637 14759 2701 14823
rect 2717 14759 2781 14823
rect 2797 14759 2861 14823
rect 2877 14759 2941 14823
rect 2957 14759 3021 14823
rect 3037 14759 3101 14823
rect 3117 14759 3181 14823
rect 3197 14759 3261 14823
rect 3277 14759 3341 14823
rect 3357 14759 3421 14823
rect 3437 14759 3501 14823
rect 3517 14759 3581 14823
rect 3597 14759 3661 14823
rect 3677 14759 3741 14823
rect 3757 14759 3821 14823
rect 3837 14759 3901 14823
rect 3917 14759 3981 14823
rect 3997 14759 4061 14823
rect 4077 14759 4141 14823
rect 4157 14759 4221 14823
rect 4237 14759 4301 14823
rect 4317 14759 4381 14823
rect 4397 14759 4461 14823
rect 4477 14759 4541 14823
rect 4557 14759 4621 14823
rect 4637 14759 4701 14823
rect 4717 14759 4781 14823
rect 4797 14759 4861 14823
rect 0 14742 254 14759
rect 0 14678 301 14742
rect 317 14678 381 14742
rect 397 14678 461 14742
rect 477 14678 541 14742
rect 557 14678 621 14742
rect 637 14678 701 14742
rect 717 14678 781 14742
rect 797 14678 861 14742
rect 877 14678 941 14742
rect 957 14678 1021 14742
rect 1037 14678 1101 14742
rect 1117 14678 1181 14742
rect 1197 14678 1261 14742
rect 1277 14678 1341 14742
rect 1357 14678 1421 14742
rect 1437 14678 1501 14742
rect 1517 14678 1581 14742
rect 1597 14678 1661 14742
rect 1677 14678 1741 14742
rect 1757 14678 1821 14742
rect 1837 14678 1901 14742
rect 1917 14678 1981 14742
rect 1997 14678 2061 14742
rect 2077 14678 2141 14742
rect 2157 14678 2221 14742
rect 2237 14678 2301 14742
rect 2317 14678 2381 14742
rect 2397 14678 2461 14742
rect 2477 14678 2541 14742
rect 2557 14678 2621 14742
rect 2637 14678 2701 14742
rect 2717 14678 2781 14742
rect 2797 14678 2861 14742
rect 2877 14678 2941 14742
rect 2957 14678 3021 14742
rect 3037 14678 3101 14742
rect 3117 14678 3181 14742
rect 3197 14678 3261 14742
rect 3277 14678 3341 14742
rect 3357 14678 3421 14742
rect 3437 14678 3501 14742
rect 3517 14678 3581 14742
rect 3597 14678 3661 14742
rect 3677 14678 3741 14742
rect 3757 14678 3821 14742
rect 3837 14678 3901 14742
rect 3917 14678 3981 14742
rect 3997 14678 4061 14742
rect 4077 14678 4141 14742
rect 4157 14678 4221 14742
rect 4237 14678 4301 14742
rect 4317 14678 4381 14742
rect 4397 14678 4461 14742
rect 4477 14678 4541 14742
rect 4557 14678 4621 14742
rect 4637 14678 4701 14742
rect 4717 14678 4781 14742
rect 4797 14678 4861 14742
rect 0 14661 254 14678
rect 0 14597 301 14661
rect 317 14597 381 14661
rect 397 14597 461 14661
rect 477 14597 541 14661
rect 557 14597 621 14661
rect 637 14597 701 14661
rect 717 14597 781 14661
rect 797 14597 861 14661
rect 877 14597 941 14661
rect 957 14597 1021 14661
rect 1037 14597 1101 14661
rect 1117 14597 1181 14661
rect 1197 14597 1261 14661
rect 1277 14597 1341 14661
rect 1357 14597 1421 14661
rect 1437 14597 1501 14661
rect 1517 14597 1581 14661
rect 1597 14597 1661 14661
rect 1677 14597 1741 14661
rect 1757 14597 1821 14661
rect 1837 14597 1901 14661
rect 1917 14597 1981 14661
rect 1997 14597 2061 14661
rect 2077 14597 2141 14661
rect 2157 14597 2221 14661
rect 2237 14597 2301 14661
rect 2317 14597 2381 14661
rect 2397 14597 2461 14661
rect 2477 14597 2541 14661
rect 2557 14597 2621 14661
rect 2637 14597 2701 14661
rect 2717 14597 2781 14661
rect 2797 14597 2861 14661
rect 2877 14597 2941 14661
rect 2957 14597 3021 14661
rect 3037 14597 3101 14661
rect 3117 14597 3181 14661
rect 3197 14597 3261 14661
rect 3277 14597 3341 14661
rect 3357 14597 3421 14661
rect 3437 14597 3501 14661
rect 3517 14597 3581 14661
rect 3597 14597 3661 14661
rect 3677 14597 3741 14661
rect 3757 14597 3821 14661
rect 3837 14597 3901 14661
rect 3917 14597 3981 14661
rect 3997 14597 4061 14661
rect 4077 14597 4141 14661
rect 4157 14597 4221 14661
rect 4237 14597 4301 14661
rect 4317 14597 4381 14661
rect 4397 14597 4461 14661
rect 4477 14597 4541 14661
rect 4557 14597 4621 14661
rect 4637 14597 4701 14661
rect 4717 14597 4781 14661
rect 4797 14597 4861 14661
rect 0 14579 254 14597
rect 0 14515 301 14579
rect 317 14515 381 14579
rect 397 14515 461 14579
rect 477 14515 541 14579
rect 557 14515 621 14579
rect 637 14515 701 14579
rect 717 14515 781 14579
rect 797 14515 861 14579
rect 877 14515 941 14579
rect 957 14515 1021 14579
rect 1037 14515 1101 14579
rect 1117 14515 1181 14579
rect 1197 14515 1261 14579
rect 1277 14515 1341 14579
rect 1357 14515 1421 14579
rect 1437 14515 1501 14579
rect 1517 14515 1581 14579
rect 1597 14515 1661 14579
rect 1677 14515 1741 14579
rect 1757 14515 1821 14579
rect 1837 14515 1901 14579
rect 1917 14515 1981 14579
rect 1997 14515 2061 14579
rect 2077 14515 2141 14579
rect 2157 14515 2221 14579
rect 2237 14515 2301 14579
rect 2317 14515 2381 14579
rect 2397 14515 2461 14579
rect 2477 14515 2541 14579
rect 2557 14515 2621 14579
rect 2637 14515 2701 14579
rect 2717 14515 2781 14579
rect 2797 14515 2861 14579
rect 2877 14515 2941 14579
rect 2957 14515 3021 14579
rect 3037 14515 3101 14579
rect 3117 14515 3181 14579
rect 3197 14515 3261 14579
rect 3277 14515 3341 14579
rect 3357 14515 3421 14579
rect 3437 14515 3501 14579
rect 3517 14515 3581 14579
rect 3597 14515 3661 14579
rect 3677 14515 3741 14579
rect 3757 14515 3821 14579
rect 3837 14515 3901 14579
rect 3917 14515 3981 14579
rect 3997 14515 4061 14579
rect 4077 14515 4141 14579
rect 4157 14515 4221 14579
rect 4237 14515 4301 14579
rect 4317 14515 4381 14579
rect 4397 14515 4461 14579
rect 4477 14515 4541 14579
rect 4557 14515 4621 14579
rect 4637 14515 4701 14579
rect 4717 14515 4781 14579
rect 4797 14515 4861 14579
rect 0 14497 254 14515
rect 0 14433 301 14497
rect 317 14433 381 14497
rect 397 14433 461 14497
rect 477 14433 541 14497
rect 557 14433 621 14497
rect 637 14433 701 14497
rect 717 14433 781 14497
rect 797 14433 861 14497
rect 877 14433 941 14497
rect 957 14433 1021 14497
rect 1037 14433 1101 14497
rect 1117 14433 1181 14497
rect 1197 14433 1261 14497
rect 1277 14433 1341 14497
rect 1357 14433 1421 14497
rect 1437 14433 1501 14497
rect 1517 14433 1581 14497
rect 1597 14433 1661 14497
rect 1677 14433 1741 14497
rect 1757 14433 1821 14497
rect 1837 14433 1901 14497
rect 1917 14433 1981 14497
rect 1997 14433 2061 14497
rect 2077 14433 2141 14497
rect 2157 14433 2221 14497
rect 2237 14433 2301 14497
rect 2317 14433 2381 14497
rect 2397 14433 2461 14497
rect 2477 14433 2541 14497
rect 2557 14433 2621 14497
rect 2637 14433 2701 14497
rect 2717 14433 2781 14497
rect 2797 14433 2861 14497
rect 2877 14433 2941 14497
rect 2957 14433 3021 14497
rect 3037 14433 3101 14497
rect 3117 14433 3181 14497
rect 3197 14433 3261 14497
rect 3277 14433 3341 14497
rect 3357 14433 3421 14497
rect 3437 14433 3501 14497
rect 3517 14433 3581 14497
rect 3597 14433 3661 14497
rect 3677 14433 3741 14497
rect 3757 14433 3821 14497
rect 3837 14433 3901 14497
rect 3917 14433 3981 14497
rect 3997 14433 4061 14497
rect 4077 14433 4141 14497
rect 4157 14433 4221 14497
rect 4237 14433 4301 14497
rect 4317 14433 4381 14497
rect 4397 14433 4461 14497
rect 4477 14433 4541 14497
rect 4557 14433 4621 14497
rect 4637 14433 4701 14497
rect 4717 14433 4781 14497
rect 4797 14433 4861 14497
rect 0 14415 254 14433
rect 0 14351 301 14415
rect 317 14351 381 14415
rect 397 14351 461 14415
rect 477 14351 541 14415
rect 557 14351 621 14415
rect 637 14351 701 14415
rect 717 14351 781 14415
rect 797 14351 861 14415
rect 877 14351 941 14415
rect 957 14351 1021 14415
rect 1037 14351 1101 14415
rect 1117 14351 1181 14415
rect 1197 14351 1261 14415
rect 1277 14351 1341 14415
rect 1357 14351 1421 14415
rect 1437 14351 1501 14415
rect 1517 14351 1581 14415
rect 1597 14351 1661 14415
rect 1677 14351 1741 14415
rect 1757 14351 1821 14415
rect 1837 14351 1901 14415
rect 1917 14351 1981 14415
rect 1997 14351 2061 14415
rect 2077 14351 2141 14415
rect 2157 14351 2221 14415
rect 2237 14351 2301 14415
rect 2317 14351 2381 14415
rect 2397 14351 2461 14415
rect 2477 14351 2541 14415
rect 2557 14351 2621 14415
rect 2637 14351 2701 14415
rect 2717 14351 2781 14415
rect 2797 14351 2861 14415
rect 2877 14351 2941 14415
rect 2957 14351 3021 14415
rect 3037 14351 3101 14415
rect 3117 14351 3181 14415
rect 3197 14351 3261 14415
rect 3277 14351 3341 14415
rect 3357 14351 3421 14415
rect 3437 14351 3501 14415
rect 3517 14351 3581 14415
rect 3597 14351 3661 14415
rect 3677 14351 3741 14415
rect 3757 14351 3821 14415
rect 3837 14351 3901 14415
rect 3917 14351 3981 14415
rect 3997 14351 4061 14415
rect 4077 14351 4141 14415
rect 4157 14351 4221 14415
rect 4237 14351 4301 14415
rect 4317 14351 4381 14415
rect 4397 14351 4461 14415
rect 4477 14351 4541 14415
rect 4557 14351 4621 14415
rect 4637 14351 4701 14415
rect 4717 14351 4781 14415
rect 4797 14351 4861 14415
rect 0 14333 254 14351
rect 0 14269 301 14333
rect 317 14269 381 14333
rect 397 14269 461 14333
rect 477 14269 541 14333
rect 557 14269 621 14333
rect 637 14269 701 14333
rect 717 14269 781 14333
rect 797 14269 861 14333
rect 877 14269 941 14333
rect 957 14269 1021 14333
rect 1037 14269 1101 14333
rect 1117 14269 1181 14333
rect 1197 14269 1261 14333
rect 1277 14269 1341 14333
rect 1357 14269 1421 14333
rect 1437 14269 1501 14333
rect 1517 14269 1581 14333
rect 1597 14269 1661 14333
rect 1677 14269 1741 14333
rect 1757 14269 1821 14333
rect 1837 14269 1901 14333
rect 1917 14269 1981 14333
rect 1997 14269 2061 14333
rect 2077 14269 2141 14333
rect 2157 14269 2221 14333
rect 2237 14269 2301 14333
rect 2317 14269 2381 14333
rect 2397 14269 2461 14333
rect 2477 14269 2541 14333
rect 2557 14269 2621 14333
rect 2637 14269 2701 14333
rect 2717 14269 2781 14333
rect 2797 14269 2861 14333
rect 2877 14269 2941 14333
rect 2957 14269 3021 14333
rect 3037 14269 3101 14333
rect 3117 14269 3181 14333
rect 3197 14269 3261 14333
rect 3277 14269 3341 14333
rect 3357 14269 3421 14333
rect 3437 14269 3501 14333
rect 3517 14269 3581 14333
rect 3597 14269 3661 14333
rect 3677 14269 3741 14333
rect 3757 14269 3821 14333
rect 3837 14269 3901 14333
rect 3917 14269 3981 14333
rect 3997 14269 4061 14333
rect 4077 14269 4141 14333
rect 4157 14269 4221 14333
rect 4237 14269 4301 14333
rect 4317 14269 4381 14333
rect 4397 14269 4461 14333
rect 4477 14269 4541 14333
rect 4557 14269 4621 14333
rect 4637 14269 4701 14333
rect 4717 14269 4781 14333
rect 4797 14269 4861 14333
rect 0 14251 254 14269
rect 0 14187 301 14251
rect 317 14187 381 14251
rect 397 14187 461 14251
rect 477 14187 541 14251
rect 557 14187 621 14251
rect 637 14187 701 14251
rect 717 14187 781 14251
rect 797 14187 861 14251
rect 877 14187 941 14251
rect 957 14187 1021 14251
rect 1037 14187 1101 14251
rect 1117 14187 1181 14251
rect 1197 14187 1261 14251
rect 1277 14187 1341 14251
rect 1357 14187 1421 14251
rect 1437 14187 1501 14251
rect 1517 14187 1581 14251
rect 1597 14187 1661 14251
rect 1677 14187 1741 14251
rect 1757 14187 1821 14251
rect 1837 14187 1901 14251
rect 1917 14187 1981 14251
rect 1997 14187 2061 14251
rect 2077 14187 2141 14251
rect 2157 14187 2221 14251
rect 2237 14187 2301 14251
rect 2317 14187 2381 14251
rect 2397 14187 2461 14251
rect 2477 14187 2541 14251
rect 2557 14187 2621 14251
rect 2637 14187 2701 14251
rect 2717 14187 2781 14251
rect 2797 14187 2861 14251
rect 2877 14187 2941 14251
rect 2957 14187 3021 14251
rect 3037 14187 3101 14251
rect 3117 14187 3181 14251
rect 3197 14187 3261 14251
rect 3277 14187 3341 14251
rect 3357 14187 3421 14251
rect 3437 14187 3501 14251
rect 3517 14187 3581 14251
rect 3597 14187 3661 14251
rect 3677 14187 3741 14251
rect 3757 14187 3821 14251
rect 3837 14187 3901 14251
rect 3917 14187 3981 14251
rect 3997 14187 4061 14251
rect 4077 14187 4141 14251
rect 4157 14187 4221 14251
rect 4237 14187 4301 14251
rect 4317 14187 4381 14251
rect 4397 14187 4461 14251
rect 4477 14187 4541 14251
rect 4557 14187 4621 14251
rect 4637 14187 4701 14251
rect 4717 14187 4781 14251
rect 4797 14187 4861 14251
rect 0 14169 254 14187
rect 0 14105 301 14169
rect 317 14105 381 14169
rect 397 14105 461 14169
rect 477 14105 541 14169
rect 557 14105 621 14169
rect 637 14105 701 14169
rect 717 14105 781 14169
rect 797 14105 861 14169
rect 877 14105 941 14169
rect 957 14105 1021 14169
rect 1037 14105 1101 14169
rect 1117 14105 1181 14169
rect 1197 14105 1261 14169
rect 1277 14105 1341 14169
rect 1357 14105 1421 14169
rect 1437 14105 1501 14169
rect 1517 14105 1581 14169
rect 1597 14105 1661 14169
rect 1677 14105 1741 14169
rect 1757 14105 1821 14169
rect 1837 14105 1901 14169
rect 1917 14105 1981 14169
rect 1997 14105 2061 14169
rect 2077 14105 2141 14169
rect 2157 14105 2221 14169
rect 2237 14105 2301 14169
rect 2317 14105 2381 14169
rect 2397 14105 2461 14169
rect 2477 14105 2541 14169
rect 2557 14105 2621 14169
rect 2637 14105 2701 14169
rect 2717 14105 2781 14169
rect 2797 14105 2861 14169
rect 2877 14105 2941 14169
rect 2957 14105 3021 14169
rect 3037 14105 3101 14169
rect 3117 14105 3181 14169
rect 3197 14105 3261 14169
rect 3277 14105 3341 14169
rect 3357 14105 3421 14169
rect 3437 14105 3501 14169
rect 3517 14105 3581 14169
rect 3597 14105 3661 14169
rect 3677 14105 3741 14169
rect 3757 14105 3821 14169
rect 3837 14105 3901 14169
rect 3917 14105 3981 14169
rect 3997 14105 4061 14169
rect 4077 14105 4141 14169
rect 4157 14105 4221 14169
rect 4237 14105 4301 14169
rect 4317 14105 4381 14169
rect 4397 14105 4461 14169
rect 4477 14105 4541 14169
rect 4557 14105 4621 14169
rect 4637 14105 4701 14169
rect 4717 14105 4781 14169
rect 4797 14105 4861 14169
rect 0 14087 254 14105
rect 0 14023 301 14087
rect 317 14023 381 14087
rect 397 14023 461 14087
rect 477 14023 541 14087
rect 557 14023 621 14087
rect 637 14023 701 14087
rect 717 14023 781 14087
rect 797 14023 861 14087
rect 877 14023 941 14087
rect 957 14023 1021 14087
rect 1037 14023 1101 14087
rect 1117 14023 1181 14087
rect 1197 14023 1261 14087
rect 1277 14023 1341 14087
rect 1357 14023 1421 14087
rect 1437 14023 1501 14087
rect 1517 14023 1581 14087
rect 1597 14023 1661 14087
rect 1677 14023 1741 14087
rect 1757 14023 1821 14087
rect 1837 14023 1901 14087
rect 1917 14023 1981 14087
rect 1997 14023 2061 14087
rect 2077 14023 2141 14087
rect 2157 14023 2221 14087
rect 2237 14023 2301 14087
rect 2317 14023 2381 14087
rect 2397 14023 2461 14087
rect 2477 14023 2541 14087
rect 2557 14023 2621 14087
rect 2637 14023 2701 14087
rect 2717 14023 2781 14087
rect 2797 14023 2861 14087
rect 2877 14023 2941 14087
rect 2957 14023 3021 14087
rect 3037 14023 3101 14087
rect 3117 14023 3181 14087
rect 3197 14023 3261 14087
rect 3277 14023 3341 14087
rect 3357 14023 3421 14087
rect 3437 14023 3501 14087
rect 3517 14023 3581 14087
rect 3597 14023 3661 14087
rect 3677 14023 3741 14087
rect 3757 14023 3821 14087
rect 3837 14023 3901 14087
rect 3917 14023 3981 14087
rect 3997 14023 4061 14087
rect 4077 14023 4141 14087
rect 4157 14023 4221 14087
rect 4237 14023 4301 14087
rect 4317 14023 4381 14087
rect 4397 14023 4461 14087
rect 4477 14023 4541 14087
rect 4557 14023 4621 14087
rect 4637 14023 4701 14087
rect 4717 14023 4781 14087
rect 4797 14023 4861 14087
rect 0 14005 254 14023
rect 0 13941 301 14005
rect 317 13941 381 14005
rect 397 13941 461 14005
rect 477 13941 541 14005
rect 557 13941 621 14005
rect 637 13941 701 14005
rect 717 13941 781 14005
rect 797 13941 861 14005
rect 877 13941 941 14005
rect 957 13941 1021 14005
rect 1037 13941 1101 14005
rect 1117 13941 1181 14005
rect 1197 13941 1261 14005
rect 1277 13941 1341 14005
rect 1357 13941 1421 14005
rect 1437 13941 1501 14005
rect 1517 13941 1581 14005
rect 1597 13941 1661 14005
rect 1677 13941 1741 14005
rect 1757 13941 1821 14005
rect 1837 13941 1901 14005
rect 1917 13941 1981 14005
rect 1997 13941 2061 14005
rect 2077 13941 2141 14005
rect 2157 13941 2221 14005
rect 2237 13941 2301 14005
rect 2317 13941 2381 14005
rect 2397 13941 2461 14005
rect 2477 13941 2541 14005
rect 2557 13941 2621 14005
rect 2637 13941 2701 14005
rect 2717 13941 2781 14005
rect 2797 13941 2861 14005
rect 2877 13941 2941 14005
rect 2957 13941 3021 14005
rect 3037 13941 3101 14005
rect 3117 13941 3181 14005
rect 3197 13941 3261 14005
rect 3277 13941 3341 14005
rect 3357 13941 3421 14005
rect 3437 13941 3501 14005
rect 3517 13941 3581 14005
rect 3597 13941 3661 14005
rect 3677 13941 3741 14005
rect 3757 13941 3821 14005
rect 3837 13941 3901 14005
rect 3917 13941 3981 14005
rect 3997 13941 4061 14005
rect 4077 13941 4141 14005
rect 4157 13941 4221 14005
rect 4237 13941 4301 14005
rect 4317 13941 4381 14005
rect 4397 13941 4461 14005
rect 4477 13941 4541 14005
rect 4557 13941 4621 14005
rect 4637 13941 4701 14005
rect 4717 13941 4781 14005
rect 4797 13941 4861 14005
rect 0 13923 254 13941
rect 0 13859 301 13923
rect 317 13859 381 13923
rect 397 13859 461 13923
rect 477 13859 541 13923
rect 557 13859 621 13923
rect 637 13859 701 13923
rect 717 13859 781 13923
rect 797 13859 861 13923
rect 877 13859 941 13923
rect 957 13859 1021 13923
rect 1037 13859 1101 13923
rect 1117 13859 1181 13923
rect 1197 13859 1261 13923
rect 1277 13859 1341 13923
rect 1357 13859 1421 13923
rect 1437 13859 1501 13923
rect 1517 13859 1581 13923
rect 1597 13859 1661 13923
rect 1677 13859 1741 13923
rect 1757 13859 1821 13923
rect 1837 13859 1901 13923
rect 1917 13859 1981 13923
rect 1997 13859 2061 13923
rect 2077 13859 2141 13923
rect 2157 13859 2221 13923
rect 2237 13859 2301 13923
rect 2317 13859 2381 13923
rect 2397 13859 2461 13923
rect 2477 13859 2541 13923
rect 2557 13859 2621 13923
rect 2637 13859 2701 13923
rect 2717 13859 2781 13923
rect 2797 13859 2861 13923
rect 2877 13859 2941 13923
rect 2957 13859 3021 13923
rect 3037 13859 3101 13923
rect 3117 13859 3181 13923
rect 3197 13859 3261 13923
rect 3277 13859 3341 13923
rect 3357 13859 3421 13923
rect 3437 13859 3501 13923
rect 3517 13859 3581 13923
rect 3597 13859 3661 13923
rect 3677 13859 3741 13923
rect 3757 13859 3821 13923
rect 3837 13859 3901 13923
rect 3917 13859 3981 13923
rect 3997 13859 4061 13923
rect 4077 13859 4141 13923
rect 4157 13859 4221 13923
rect 4237 13859 4301 13923
rect 4317 13859 4381 13923
rect 4397 13859 4461 13923
rect 4477 13859 4541 13923
rect 4557 13859 4621 13923
rect 4637 13859 4701 13923
rect 4717 13859 4781 13923
rect 4797 13859 4861 13923
rect 0 13841 254 13859
rect 0 13777 301 13841
rect 317 13777 381 13841
rect 397 13777 461 13841
rect 477 13777 541 13841
rect 557 13777 621 13841
rect 637 13777 701 13841
rect 717 13777 781 13841
rect 797 13777 861 13841
rect 877 13777 941 13841
rect 957 13777 1021 13841
rect 1037 13777 1101 13841
rect 1117 13777 1181 13841
rect 1197 13777 1261 13841
rect 1277 13777 1341 13841
rect 1357 13777 1421 13841
rect 1437 13777 1501 13841
rect 1517 13777 1581 13841
rect 1597 13777 1661 13841
rect 1677 13777 1741 13841
rect 1757 13777 1821 13841
rect 1837 13777 1901 13841
rect 1917 13777 1981 13841
rect 1997 13777 2061 13841
rect 2077 13777 2141 13841
rect 2157 13777 2221 13841
rect 2237 13777 2301 13841
rect 2317 13777 2381 13841
rect 2397 13777 2461 13841
rect 2477 13777 2541 13841
rect 2557 13777 2621 13841
rect 2637 13777 2701 13841
rect 2717 13777 2781 13841
rect 2797 13777 2861 13841
rect 2877 13777 2941 13841
rect 2957 13777 3021 13841
rect 3037 13777 3101 13841
rect 3117 13777 3181 13841
rect 3197 13777 3261 13841
rect 3277 13777 3341 13841
rect 3357 13777 3421 13841
rect 3437 13777 3501 13841
rect 3517 13777 3581 13841
rect 3597 13777 3661 13841
rect 3677 13777 3741 13841
rect 3757 13777 3821 13841
rect 3837 13777 3901 13841
rect 3917 13777 3981 13841
rect 3997 13777 4061 13841
rect 4077 13777 4141 13841
rect 4157 13777 4221 13841
rect 4237 13777 4301 13841
rect 4317 13777 4381 13841
rect 4397 13777 4461 13841
rect 4477 13777 4541 13841
rect 4557 13777 4621 13841
rect 4637 13777 4701 13841
rect 4717 13777 4781 13841
rect 4797 13777 4861 13841
rect 0 13759 254 13777
rect 0 13695 301 13759
rect 317 13695 381 13759
rect 397 13695 461 13759
rect 477 13695 541 13759
rect 557 13695 621 13759
rect 637 13695 701 13759
rect 717 13695 781 13759
rect 797 13695 861 13759
rect 877 13695 941 13759
rect 957 13695 1021 13759
rect 1037 13695 1101 13759
rect 1117 13695 1181 13759
rect 1197 13695 1261 13759
rect 1277 13695 1341 13759
rect 1357 13695 1421 13759
rect 1437 13695 1501 13759
rect 1517 13695 1581 13759
rect 1597 13695 1661 13759
rect 1677 13695 1741 13759
rect 1757 13695 1821 13759
rect 1837 13695 1901 13759
rect 1917 13695 1981 13759
rect 1997 13695 2061 13759
rect 2077 13695 2141 13759
rect 2157 13695 2221 13759
rect 2237 13695 2301 13759
rect 2317 13695 2381 13759
rect 2397 13695 2461 13759
rect 2477 13695 2541 13759
rect 2557 13695 2621 13759
rect 2637 13695 2701 13759
rect 2717 13695 2781 13759
rect 2797 13695 2861 13759
rect 2877 13695 2941 13759
rect 2957 13695 3021 13759
rect 3037 13695 3101 13759
rect 3117 13695 3181 13759
rect 3197 13695 3261 13759
rect 3277 13695 3341 13759
rect 3357 13695 3421 13759
rect 3437 13695 3501 13759
rect 3517 13695 3581 13759
rect 3597 13695 3661 13759
rect 3677 13695 3741 13759
rect 3757 13695 3821 13759
rect 3837 13695 3901 13759
rect 3917 13695 3981 13759
rect 3997 13695 4061 13759
rect 4077 13695 4141 13759
rect 4157 13695 4221 13759
rect 4237 13695 4301 13759
rect 4317 13695 4381 13759
rect 4397 13695 4461 13759
rect 4477 13695 4541 13759
rect 4557 13695 4621 13759
rect 4637 13695 4701 13759
rect 4717 13695 4781 13759
rect 4797 13695 4861 13759
rect 0 13677 254 13695
rect 0 13613 301 13677
rect 317 13613 381 13677
rect 397 13613 461 13677
rect 477 13613 541 13677
rect 557 13613 621 13677
rect 637 13613 701 13677
rect 717 13613 781 13677
rect 797 13613 861 13677
rect 877 13613 941 13677
rect 957 13613 1021 13677
rect 1037 13613 1101 13677
rect 1117 13613 1181 13677
rect 1197 13613 1261 13677
rect 1277 13613 1341 13677
rect 1357 13613 1421 13677
rect 1437 13613 1501 13677
rect 1517 13613 1581 13677
rect 1597 13613 1661 13677
rect 1677 13613 1741 13677
rect 1757 13613 1821 13677
rect 1837 13613 1901 13677
rect 1917 13613 1981 13677
rect 1997 13613 2061 13677
rect 2077 13613 2141 13677
rect 2157 13613 2221 13677
rect 2237 13613 2301 13677
rect 2317 13613 2381 13677
rect 2397 13613 2461 13677
rect 2477 13613 2541 13677
rect 2557 13613 2621 13677
rect 2637 13613 2701 13677
rect 2717 13613 2781 13677
rect 2797 13613 2861 13677
rect 2877 13613 2941 13677
rect 2957 13613 3021 13677
rect 3037 13613 3101 13677
rect 3117 13613 3181 13677
rect 3197 13613 3261 13677
rect 3277 13613 3341 13677
rect 3357 13613 3421 13677
rect 3437 13613 3501 13677
rect 3517 13613 3581 13677
rect 3597 13613 3661 13677
rect 3677 13613 3741 13677
rect 3757 13613 3821 13677
rect 3837 13613 3901 13677
rect 3917 13613 3981 13677
rect 3997 13613 4061 13677
rect 4077 13613 4141 13677
rect 4157 13613 4221 13677
rect 4237 13613 4301 13677
rect 4317 13613 4381 13677
rect 4397 13613 4461 13677
rect 4477 13613 4541 13677
rect 4557 13613 4621 13677
rect 4637 13613 4701 13677
rect 4717 13613 4781 13677
rect 4797 13613 4861 13677
rect 0 13607 254 13613
rect 14746 13607 15000 16559
rect 0 13304 254 13307
rect 0 13240 271 13304
rect 288 13240 352 13304
rect 369 13240 433 13304
rect 450 13240 514 13304
rect 531 13240 595 13304
rect 612 13240 676 13304
rect 693 13240 757 13304
rect 774 13240 838 13304
rect 855 13240 919 13304
rect 936 13240 1000 13304
rect 1017 13240 1081 13304
rect 1098 13240 1162 13304
rect 1179 13240 1243 13304
rect 1260 13240 1324 13304
rect 1341 13240 1405 13304
rect 1422 13240 1486 13304
rect 1503 13240 1567 13304
rect 1584 13240 1648 13304
rect 1665 13240 1729 13304
rect 1746 13240 1810 13304
rect 1827 13240 1891 13304
rect 1908 13240 1972 13304
rect 1989 13240 2053 13304
rect 2070 13240 2134 13304
rect 2151 13240 2215 13304
rect 2232 13240 2296 13304
rect 2313 13240 2377 13304
rect 2394 13240 2458 13304
rect 2475 13240 2539 13304
rect 2556 13240 2620 13304
rect 2637 13240 2701 13304
rect 2718 13240 2782 13304
rect 2799 13240 2863 13304
rect 2880 13240 2944 13304
rect 2961 13240 3025 13304
rect 3042 13240 3106 13304
rect 3123 13240 3187 13304
rect 3204 13240 3268 13304
rect 3285 13240 3349 13304
rect 3366 13240 3430 13304
rect 3447 13240 3511 13304
rect 3528 13240 3592 13304
rect 3609 13240 3673 13304
rect 3690 13240 3754 13304
rect 3771 13240 3835 13304
rect 3852 13240 3916 13304
rect 3933 13240 3997 13304
rect 4014 13240 4078 13304
rect 4095 13240 4159 13304
rect 4176 13240 4240 13304
rect 4257 13240 4321 13304
rect 4338 13240 4402 13304
rect 4420 13240 4484 13304
rect 4502 13240 4566 13304
rect 4584 13240 4648 13304
rect 4666 13240 4730 13304
rect 4748 13240 4812 13304
rect 4830 13240 4894 13304
rect 0 13222 254 13240
rect 0 13158 271 13222
rect 288 13158 352 13222
rect 369 13158 433 13222
rect 450 13158 514 13222
rect 531 13158 595 13222
rect 612 13158 676 13222
rect 693 13158 757 13222
rect 774 13158 838 13222
rect 855 13158 919 13222
rect 936 13158 1000 13222
rect 1017 13158 1081 13222
rect 1098 13158 1162 13222
rect 1179 13158 1243 13222
rect 1260 13158 1324 13222
rect 1341 13158 1405 13222
rect 1422 13158 1486 13222
rect 1503 13158 1567 13222
rect 1584 13158 1648 13222
rect 1665 13158 1729 13222
rect 1746 13158 1810 13222
rect 1827 13158 1891 13222
rect 1908 13158 1972 13222
rect 1989 13158 2053 13222
rect 2070 13158 2134 13222
rect 2151 13158 2215 13222
rect 2232 13158 2296 13222
rect 2313 13158 2377 13222
rect 2394 13158 2458 13222
rect 2475 13158 2539 13222
rect 2556 13158 2620 13222
rect 2637 13158 2701 13222
rect 2718 13158 2782 13222
rect 2799 13158 2863 13222
rect 2880 13158 2944 13222
rect 2961 13158 3025 13222
rect 3042 13158 3106 13222
rect 3123 13158 3187 13222
rect 3204 13158 3268 13222
rect 3285 13158 3349 13222
rect 3366 13158 3430 13222
rect 3447 13158 3511 13222
rect 3528 13158 3592 13222
rect 3609 13158 3673 13222
rect 3690 13158 3754 13222
rect 3771 13158 3835 13222
rect 3852 13158 3916 13222
rect 3933 13158 3997 13222
rect 4014 13158 4078 13222
rect 4095 13158 4159 13222
rect 4176 13158 4240 13222
rect 4257 13158 4321 13222
rect 4338 13158 4402 13222
rect 4420 13158 4484 13222
rect 4502 13158 4566 13222
rect 4584 13158 4648 13222
rect 4666 13158 4730 13222
rect 4748 13158 4812 13222
rect 4830 13158 4894 13222
rect 0 13140 254 13158
rect 0 13076 271 13140
rect 288 13076 352 13140
rect 369 13076 433 13140
rect 450 13076 514 13140
rect 531 13076 595 13140
rect 612 13076 676 13140
rect 693 13076 757 13140
rect 774 13076 838 13140
rect 855 13076 919 13140
rect 936 13076 1000 13140
rect 1017 13076 1081 13140
rect 1098 13076 1162 13140
rect 1179 13076 1243 13140
rect 1260 13076 1324 13140
rect 1341 13076 1405 13140
rect 1422 13076 1486 13140
rect 1503 13076 1567 13140
rect 1584 13076 1648 13140
rect 1665 13076 1729 13140
rect 1746 13076 1810 13140
rect 1827 13076 1891 13140
rect 1908 13076 1972 13140
rect 1989 13076 2053 13140
rect 2070 13076 2134 13140
rect 2151 13076 2215 13140
rect 2232 13076 2296 13140
rect 2313 13076 2377 13140
rect 2394 13076 2458 13140
rect 2475 13076 2539 13140
rect 2556 13076 2620 13140
rect 2637 13076 2701 13140
rect 2718 13076 2782 13140
rect 2799 13076 2863 13140
rect 2880 13076 2944 13140
rect 2961 13076 3025 13140
rect 3042 13076 3106 13140
rect 3123 13076 3187 13140
rect 3204 13076 3268 13140
rect 3285 13076 3349 13140
rect 3366 13076 3430 13140
rect 3447 13076 3511 13140
rect 3528 13076 3592 13140
rect 3609 13076 3673 13140
rect 3690 13076 3754 13140
rect 3771 13076 3835 13140
rect 3852 13076 3916 13140
rect 3933 13076 3997 13140
rect 4014 13076 4078 13140
rect 4095 13076 4159 13140
rect 4176 13076 4240 13140
rect 4257 13076 4321 13140
rect 4338 13076 4402 13140
rect 4420 13076 4484 13140
rect 4502 13076 4566 13140
rect 4584 13076 4648 13140
rect 4666 13076 4730 13140
rect 4748 13076 4812 13140
rect 4830 13076 4894 13140
rect 0 13058 254 13076
rect 0 12994 271 13058
rect 288 12994 352 13058
rect 369 12994 433 13058
rect 450 12994 514 13058
rect 531 12994 595 13058
rect 612 12994 676 13058
rect 693 12994 757 13058
rect 774 12994 838 13058
rect 855 12994 919 13058
rect 936 12994 1000 13058
rect 1017 12994 1081 13058
rect 1098 12994 1162 13058
rect 1179 12994 1243 13058
rect 1260 12994 1324 13058
rect 1341 12994 1405 13058
rect 1422 12994 1486 13058
rect 1503 12994 1567 13058
rect 1584 12994 1648 13058
rect 1665 12994 1729 13058
rect 1746 12994 1810 13058
rect 1827 12994 1891 13058
rect 1908 12994 1972 13058
rect 1989 12994 2053 13058
rect 2070 12994 2134 13058
rect 2151 12994 2215 13058
rect 2232 12994 2296 13058
rect 2313 12994 2377 13058
rect 2394 12994 2458 13058
rect 2475 12994 2539 13058
rect 2556 12994 2620 13058
rect 2637 12994 2701 13058
rect 2718 12994 2782 13058
rect 2799 12994 2863 13058
rect 2880 12994 2944 13058
rect 2961 12994 3025 13058
rect 3042 12994 3106 13058
rect 3123 12994 3187 13058
rect 3204 12994 3268 13058
rect 3285 12994 3349 13058
rect 3366 12994 3430 13058
rect 3447 12994 3511 13058
rect 3528 12994 3592 13058
rect 3609 12994 3673 13058
rect 3690 12994 3754 13058
rect 3771 12994 3835 13058
rect 3852 12994 3916 13058
rect 3933 12994 3997 13058
rect 4014 12994 4078 13058
rect 4095 12994 4159 13058
rect 4176 12994 4240 13058
rect 4257 12994 4321 13058
rect 4338 12994 4402 13058
rect 4420 12994 4484 13058
rect 4502 12994 4566 13058
rect 4584 12994 4648 13058
rect 4666 12994 4730 13058
rect 4748 12994 4812 13058
rect 4830 12994 4894 13058
rect 0 12976 254 12994
rect 0 12912 271 12976
rect 288 12912 352 12976
rect 369 12912 433 12976
rect 450 12912 514 12976
rect 531 12912 595 12976
rect 612 12912 676 12976
rect 693 12912 757 12976
rect 774 12912 838 12976
rect 855 12912 919 12976
rect 936 12912 1000 12976
rect 1017 12912 1081 12976
rect 1098 12912 1162 12976
rect 1179 12912 1243 12976
rect 1260 12912 1324 12976
rect 1341 12912 1405 12976
rect 1422 12912 1486 12976
rect 1503 12912 1567 12976
rect 1584 12912 1648 12976
rect 1665 12912 1729 12976
rect 1746 12912 1810 12976
rect 1827 12912 1891 12976
rect 1908 12912 1972 12976
rect 1989 12912 2053 12976
rect 2070 12912 2134 12976
rect 2151 12912 2215 12976
rect 2232 12912 2296 12976
rect 2313 12912 2377 12976
rect 2394 12912 2458 12976
rect 2475 12912 2539 12976
rect 2556 12912 2620 12976
rect 2637 12912 2701 12976
rect 2718 12912 2782 12976
rect 2799 12912 2863 12976
rect 2880 12912 2944 12976
rect 2961 12912 3025 12976
rect 3042 12912 3106 12976
rect 3123 12912 3187 12976
rect 3204 12912 3268 12976
rect 3285 12912 3349 12976
rect 3366 12912 3430 12976
rect 3447 12912 3511 12976
rect 3528 12912 3592 12976
rect 3609 12912 3673 12976
rect 3690 12912 3754 12976
rect 3771 12912 3835 12976
rect 3852 12912 3916 12976
rect 3933 12912 3997 12976
rect 4014 12912 4078 12976
rect 4095 12912 4159 12976
rect 4176 12912 4240 12976
rect 4257 12912 4321 12976
rect 4338 12912 4402 12976
rect 4420 12912 4484 12976
rect 4502 12912 4566 12976
rect 4584 12912 4648 12976
rect 4666 12912 4730 12976
rect 4748 12912 4812 12976
rect 4830 12912 4894 12976
rect 0 12894 254 12912
rect 0 12830 271 12894
rect 288 12830 352 12894
rect 369 12830 433 12894
rect 450 12830 514 12894
rect 531 12830 595 12894
rect 612 12830 676 12894
rect 693 12830 757 12894
rect 774 12830 838 12894
rect 855 12830 919 12894
rect 936 12830 1000 12894
rect 1017 12830 1081 12894
rect 1098 12830 1162 12894
rect 1179 12830 1243 12894
rect 1260 12830 1324 12894
rect 1341 12830 1405 12894
rect 1422 12830 1486 12894
rect 1503 12830 1567 12894
rect 1584 12830 1648 12894
rect 1665 12830 1729 12894
rect 1746 12830 1810 12894
rect 1827 12830 1891 12894
rect 1908 12830 1972 12894
rect 1989 12830 2053 12894
rect 2070 12830 2134 12894
rect 2151 12830 2215 12894
rect 2232 12830 2296 12894
rect 2313 12830 2377 12894
rect 2394 12830 2458 12894
rect 2475 12830 2539 12894
rect 2556 12830 2620 12894
rect 2637 12830 2701 12894
rect 2718 12830 2782 12894
rect 2799 12830 2863 12894
rect 2880 12830 2944 12894
rect 2961 12830 3025 12894
rect 3042 12830 3106 12894
rect 3123 12830 3187 12894
rect 3204 12830 3268 12894
rect 3285 12830 3349 12894
rect 3366 12830 3430 12894
rect 3447 12830 3511 12894
rect 3528 12830 3592 12894
rect 3609 12830 3673 12894
rect 3690 12830 3754 12894
rect 3771 12830 3835 12894
rect 3852 12830 3916 12894
rect 3933 12830 3997 12894
rect 4014 12830 4078 12894
rect 4095 12830 4159 12894
rect 4176 12830 4240 12894
rect 4257 12830 4321 12894
rect 4338 12830 4402 12894
rect 4420 12830 4484 12894
rect 4502 12830 4566 12894
rect 4584 12830 4648 12894
rect 4666 12830 4730 12894
rect 4748 12830 4812 12894
rect 4830 12830 4894 12894
rect 0 12812 254 12830
rect 0 12748 271 12812
rect 288 12748 352 12812
rect 369 12748 433 12812
rect 450 12748 514 12812
rect 531 12748 595 12812
rect 612 12748 676 12812
rect 693 12748 757 12812
rect 774 12748 838 12812
rect 855 12748 919 12812
rect 936 12748 1000 12812
rect 1017 12748 1081 12812
rect 1098 12748 1162 12812
rect 1179 12748 1243 12812
rect 1260 12748 1324 12812
rect 1341 12748 1405 12812
rect 1422 12748 1486 12812
rect 1503 12748 1567 12812
rect 1584 12748 1648 12812
rect 1665 12748 1729 12812
rect 1746 12748 1810 12812
rect 1827 12748 1891 12812
rect 1908 12748 1972 12812
rect 1989 12748 2053 12812
rect 2070 12748 2134 12812
rect 2151 12748 2215 12812
rect 2232 12748 2296 12812
rect 2313 12748 2377 12812
rect 2394 12748 2458 12812
rect 2475 12748 2539 12812
rect 2556 12748 2620 12812
rect 2637 12748 2701 12812
rect 2718 12748 2782 12812
rect 2799 12748 2863 12812
rect 2880 12748 2944 12812
rect 2961 12748 3025 12812
rect 3042 12748 3106 12812
rect 3123 12748 3187 12812
rect 3204 12748 3268 12812
rect 3285 12748 3349 12812
rect 3366 12748 3430 12812
rect 3447 12748 3511 12812
rect 3528 12748 3592 12812
rect 3609 12748 3673 12812
rect 3690 12748 3754 12812
rect 3771 12748 3835 12812
rect 3852 12748 3916 12812
rect 3933 12748 3997 12812
rect 4014 12748 4078 12812
rect 4095 12748 4159 12812
rect 4176 12748 4240 12812
rect 4257 12748 4321 12812
rect 4338 12748 4402 12812
rect 4420 12748 4484 12812
rect 4502 12748 4566 12812
rect 4584 12748 4648 12812
rect 4666 12748 4730 12812
rect 4748 12748 4812 12812
rect 4830 12748 4894 12812
rect 0 12730 254 12748
rect 0 12666 271 12730
rect 288 12666 352 12730
rect 369 12666 433 12730
rect 450 12666 514 12730
rect 531 12666 595 12730
rect 612 12666 676 12730
rect 693 12666 757 12730
rect 774 12666 838 12730
rect 855 12666 919 12730
rect 936 12666 1000 12730
rect 1017 12666 1081 12730
rect 1098 12666 1162 12730
rect 1179 12666 1243 12730
rect 1260 12666 1324 12730
rect 1341 12666 1405 12730
rect 1422 12666 1486 12730
rect 1503 12666 1567 12730
rect 1584 12666 1648 12730
rect 1665 12666 1729 12730
rect 1746 12666 1810 12730
rect 1827 12666 1891 12730
rect 1908 12666 1972 12730
rect 1989 12666 2053 12730
rect 2070 12666 2134 12730
rect 2151 12666 2215 12730
rect 2232 12666 2296 12730
rect 2313 12666 2377 12730
rect 2394 12666 2458 12730
rect 2475 12666 2539 12730
rect 2556 12666 2620 12730
rect 2637 12666 2701 12730
rect 2718 12666 2782 12730
rect 2799 12666 2863 12730
rect 2880 12666 2944 12730
rect 2961 12666 3025 12730
rect 3042 12666 3106 12730
rect 3123 12666 3187 12730
rect 3204 12666 3268 12730
rect 3285 12666 3349 12730
rect 3366 12666 3430 12730
rect 3447 12666 3511 12730
rect 3528 12666 3592 12730
rect 3609 12666 3673 12730
rect 3690 12666 3754 12730
rect 3771 12666 3835 12730
rect 3852 12666 3916 12730
rect 3933 12666 3997 12730
rect 4014 12666 4078 12730
rect 4095 12666 4159 12730
rect 4176 12666 4240 12730
rect 4257 12666 4321 12730
rect 4338 12666 4402 12730
rect 4420 12666 4484 12730
rect 4502 12666 4566 12730
rect 4584 12666 4648 12730
rect 4666 12666 4730 12730
rect 4748 12666 4812 12730
rect 4830 12666 4894 12730
rect 0 12648 254 12666
rect 0 12584 271 12648
rect 288 12584 352 12648
rect 369 12584 433 12648
rect 450 12584 514 12648
rect 531 12584 595 12648
rect 612 12584 676 12648
rect 693 12584 757 12648
rect 774 12584 838 12648
rect 855 12584 919 12648
rect 936 12584 1000 12648
rect 1017 12584 1081 12648
rect 1098 12584 1162 12648
rect 1179 12584 1243 12648
rect 1260 12584 1324 12648
rect 1341 12584 1405 12648
rect 1422 12584 1486 12648
rect 1503 12584 1567 12648
rect 1584 12584 1648 12648
rect 1665 12584 1729 12648
rect 1746 12584 1810 12648
rect 1827 12584 1891 12648
rect 1908 12584 1972 12648
rect 1989 12584 2053 12648
rect 2070 12584 2134 12648
rect 2151 12584 2215 12648
rect 2232 12584 2296 12648
rect 2313 12584 2377 12648
rect 2394 12584 2458 12648
rect 2475 12584 2539 12648
rect 2556 12584 2620 12648
rect 2637 12584 2701 12648
rect 2718 12584 2782 12648
rect 2799 12584 2863 12648
rect 2880 12584 2944 12648
rect 2961 12584 3025 12648
rect 3042 12584 3106 12648
rect 3123 12584 3187 12648
rect 3204 12584 3268 12648
rect 3285 12584 3349 12648
rect 3366 12584 3430 12648
rect 3447 12584 3511 12648
rect 3528 12584 3592 12648
rect 3609 12584 3673 12648
rect 3690 12584 3754 12648
rect 3771 12584 3835 12648
rect 3852 12584 3916 12648
rect 3933 12584 3997 12648
rect 4014 12584 4078 12648
rect 4095 12584 4159 12648
rect 4176 12584 4240 12648
rect 4257 12584 4321 12648
rect 4338 12584 4402 12648
rect 4420 12584 4484 12648
rect 4502 12584 4566 12648
rect 4584 12584 4648 12648
rect 4666 12584 4730 12648
rect 4748 12584 4812 12648
rect 4830 12584 4894 12648
rect 0 12566 254 12584
rect 0 12502 271 12566
rect 288 12502 352 12566
rect 369 12502 433 12566
rect 450 12502 514 12566
rect 531 12502 595 12566
rect 612 12502 676 12566
rect 693 12502 757 12566
rect 774 12502 838 12566
rect 855 12502 919 12566
rect 936 12502 1000 12566
rect 1017 12502 1081 12566
rect 1098 12502 1162 12566
rect 1179 12502 1243 12566
rect 1260 12502 1324 12566
rect 1341 12502 1405 12566
rect 1422 12502 1486 12566
rect 1503 12502 1567 12566
rect 1584 12502 1648 12566
rect 1665 12502 1729 12566
rect 1746 12502 1810 12566
rect 1827 12502 1891 12566
rect 1908 12502 1972 12566
rect 1989 12502 2053 12566
rect 2070 12502 2134 12566
rect 2151 12502 2215 12566
rect 2232 12502 2296 12566
rect 2313 12502 2377 12566
rect 2394 12502 2458 12566
rect 2475 12502 2539 12566
rect 2556 12502 2620 12566
rect 2637 12502 2701 12566
rect 2718 12502 2782 12566
rect 2799 12502 2863 12566
rect 2880 12502 2944 12566
rect 2961 12502 3025 12566
rect 3042 12502 3106 12566
rect 3123 12502 3187 12566
rect 3204 12502 3268 12566
rect 3285 12502 3349 12566
rect 3366 12502 3430 12566
rect 3447 12502 3511 12566
rect 3528 12502 3592 12566
rect 3609 12502 3673 12566
rect 3690 12502 3754 12566
rect 3771 12502 3835 12566
rect 3852 12502 3916 12566
rect 3933 12502 3997 12566
rect 4014 12502 4078 12566
rect 4095 12502 4159 12566
rect 4176 12502 4240 12566
rect 4257 12502 4321 12566
rect 4338 12502 4402 12566
rect 4420 12502 4484 12566
rect 4502 12502 4566 12566
rect 4584 12502 4648 12566
rect 4666 12502 4730 12566
rect 4748 12502 4812 12566
rect 4830 12502 4894 12566
rect 0 12484 254 12502
rect 0 12420 271 12484
rect 288 12420 352 12484
rect 369 12420 433 12484
rect 450 12420 514 12484
rect 531 12420 595 12484
rect 612 12420 676 12484
rect 693 12420 757 12484
rect 774 12420 838 12484
rect 855 12420 919 12484
rect 936 12420 1000 12484
rect 1017 12420 1081 12484
rect 1098 12420 1162 12484
rect 1179 12420 1243 12484
rect 1260 12420 1324 12484
rect 1341 12420 1405 12484
rect 1422 12420 1486 12484
rect 1503 12420 1567 12484
rect 1584 12420 1648 12484
rect 1665 12420 1729 12484
rect 1746 12420 1810 12484
rect 1827 12420 1891 12484
rect 1908 12420 1972 12484
rect 1989 12420 2053 12484
rect 2070 12420 2134 12484
rect 2151 12420 2215 12484
rect 2232 12420 2296 12484
rect 2313 12420 2377 12484
rect 2394 12420 2458 12484
rect 2475 12420 2539 12484
rect 2556 12420 2620 12484
rect 2637 12420 2701 12484
rect 2718 12420 2782 12484
rect 2799 12420 2863 12484
rect 2880 12420 2944 12484
rect 2961 12420 3025 12484
rect 3042 12420 3106 12484
rect 3123 12420 3187 12484
rect 3204 12420 3268 12484
rect 3285 12420 3349 12484
rect 3366 12420 3430 12484
rect 3447 12420 3511 12484
rect 3528 12420 3592 12484
rect 3609 12420 3673 12484
rect 3690 12420 3754 12484
rect 3771 12420 3835 12484
rect 3852 12420 3916 12484
rect 3933 12420 3997 12484
rect 4014 12420 4078 12484
rect 4095 12420 4159 12484
rect 4176 12420 4240 12484
rect 4257 12420 4321 12484
rect 4338 12420 4402 12484
rect 4420 12420 4484 12484
rect 4502 12420 4566 12484
rect 4584 12420 4648 12484
rect 4666 12420 4730 12484
rect 4748 12420 4812 12484
rect 4830 12420 4894 12484
rect 0 12417 254 12420
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 18591 14666 18680
rect 363 18527 381 18591
rect 445 18527 463 18591
rect 527 18527 545 18591
rect 609 18527 627 18591
rect 691 18527 709 18591
rect 773 18527 791 18591
rect 855 18527 873 18591
rect 937 18527 955 18591
rect 1019 18527 1037 18591
rect 1101 18527 1119 18591
rect 1183 18527 1201 18591
rect 1265 18527 1283 18591
rect 1347 18527 1365 18591
rect 1429 18527 1447 18591
rect 1511 18527 1529 18591
rect 1593 18527 1611 18591
rect 1675 18527 1693 18591
rect 1757 18527 1775 18591
rect 1839 18527 1857 18591
rect 1921 18527 1939 18591
rect 2003 18527 2021 18591
rect 2085 18527 2103 18591
rect 2167 18527 2185 18591
rect 2249 18527 2267 18591
rect 2331 18527 2349 18591
rect 2413 18527 2431 18591
rect 2495 18527 2513 18591
rect 2577 18527 2594 18591
rect 2658 18527 2675 18591
rect 2739 18527 2756 18591
rect 2820 18527 14666 18591
rect 334 18509 14666 18527
rect 363 18445 381 18509
rect 445 18445 463 18509
rect 527 18445 545 18509
rect 609 18445 627 18509
rect 691 18445 709 18509
rect 773 18445 791 18509
rect 855 18445 873 18509
rect 937 18445 955 18509
rect 1019 18445 1037 18509
rect 1101 18445 1119 18509
rect 1183 18445 1201 18509
rect 1265 18445 1283 18509
rect 1347 18445 1365 18509
rect 1429 18445 1447 18509
rect 1511 18445 1529 18509
rect 1593 18445 1611 18509
rect 1675 18445 1693 18509
rect 1757 18445 1775 18509
rect 1839 18445 1857 18509
rect 1921 18445 1939 18509
rect 2003 18445 2021 18509
rect 2085 18445 2103 18509
rect 2167 18445 2185 18509
rect 2249 18445 2267 18509
rect 2331 18445 2349 18509
rect 2413 18445 2431 18509
rect 2495 18445 2513 18509
rect 2577 18445 2594 18509
rect 2658 18445 2675 18509
rect 2739 18445 2756 18509
rect 2820 18445 12231 18509
rect 12295 18445 12312 18509
rect 12376 18445 12393 18509
rect 12457 18445 12474 18509
rect 12538 18445 12556 18509
rect 12620 18445 12638 18509
rect 12702 18445 12720 18509
rect 12784 18445 12802 18509
rect 12866 18445 12884 18509
rect 12948 18445 12966 18509
rect 13030 18445 13048 18509
rect 13112 18445 13130 18509
rect 13194 18445 13212 18509
rect 13276 18445 13294 18509
rect 13358 18445 13376 18509
rect 13440 18445 13458 18509
rect 13522 18445 13540 18509
rect 13604 18445 13622 18509
rect 13686 18445 13704 18509
rect 13768 18445 13786 18509
rect 13850 18445 13868 18509
rect 13932 18445 13950 18509
rect 14014 18445 14032 18509
rect 14096 18445 14114 18509
rect 14178 18445 14196 18509
rect 14260 18445 14278 18509
rect 14342 18445 14360 18509
rect 14424 18445 14442 18509
rect 14506 18445 14524 18509
rect 14588 18445 14606 18509
rect 334 18427 14666 18445
rect 363 18363 381 18427
rect 445 18363 463 18427
rect 527 18363 545 18427
rect 609 18363 627 18427
rect 691 18363 709 18427
rect 773 18363 791 18427
rect 855 18363 873 18427
rect 937 18363 955 18427
rect 1019 18363 1037 18427
rect 1101 18363 1119 18427
rect 1183 18363 1201 18427
rect 1265 18363 1283 18427
rect 1347 18363 1365 18427
rect 1429 18363 1447 18427
rect 1511 18363 1529 18427
rect 1593 18363 1611 18427
rect 1675 18363 1693 18427
rect 1757 18363 1775 18427
rect 1839 18363 1857 18427
rect 1921 18363 1939 18427
rect 2003 18363 2021 18427
rect 2085 18363 2103 18427
rect 2167 18363 2185 18427
rect 2249 18363 2267 18427
rect 2331 18363 2349 18427
rect 2413 18363 2431 18427
rect 2495 18363 2513 18427
rect 2577 18363 2594 18427
rect 2658 18363 2675 18427
rect 2739 18363 2756 18427
rect 2820 18422 12231 18427
rect 334 18345 2771 18363
rect 363 18281 381 18345
rect 445 18281 463 18345
rect 527 18281 545 18345
rect 609 18281 627 18345
rect 691 18281 709 18345
rect 773 18281 791 18345
rect 855 18281 873 18345
rect 937 18281 955 18345
rect 1019 18281 1037 18345
rect 1101 18281 1119 18345
rect 1183 18281 1201 18345
rect 1265 18281 1283 18345
rect 1347 18281 1365 18345
rect 1429 18281 1447 18345
rect 1511 18281 1529 18345
rect 1593 18281 1611 18345
rect 1675 18281 1693 18345
rect 1757 18281 1775 18345
rect 1839 18281 1857 18345
rect 1921 18281 1939 18345
rect 2003 18281 2021 18345
rect 2085 18281 2103 18345
rect 2167 18281 2185 18345
rect 2249 18281 2267 18345
rect 2331 18281 2349 18345
rect 2413 18281 2431 18345
rect 2495 18281 2513 18345
rect 2577 18281 2594 18345
rect 2658 18281 2675 18345
rect 2739 18281 2756 18345
rect 334 18263 2771 18281
rect 363 18199 381 18263
rect 445 18199 463 18263
rect 527 18199 545 18263
rect 609 18199 627 18263
rect 691 18199 709 18263
rect 773 18199 791 18263
rect 855 18199 873 18263
rect 937 18199 955 18263
rect 1019 18199 1037 18263
rect 1101 18199 1119 18263
rect 1183 18199 1201 18263
rect 1265 18199 1283 18263
rect 1347 18199 1365 18263
rect 1429 18199 1447 18263
rect 1511 18199 1529 18263
rect 1593 18199 1611 18263
rect 1675 18199 1693 18263
rect 1757 18199 1775 18263
rect 1839 18199 1857 18263
rect 1921 18199 1939 18263
rect 2003 18199 2021 18263
rect 2085 18199 2103 18263
rect 2167 18199 2185 18263
rect 2249 18199 2267 18263
rect 2331 18199 2349 18263
rect 2413 18199 2431 18263
rect 2495 18199 2513 18263
rect 2577 18199 2594 18263
rect 2658 18199 2675 18263
rect 2739 18199 2756 18263
rect 334 18181 2771 18199
rect 3153 18244 11898 18422
rect 12295 18363 12312 18427
rect 12376 18363 12393 18427
rect 12457 18363 12474 18427
rect 12538 18363 12556 18427
rect 12620 18363 12638 18427
rect 12702 18363 12720 18427
rect 12784 18363 12802 18427
rect 12866 18363 12884 18427
rect 12948 18363 12966 18427
rect 13030 18363 13048 18427
rect 13112 18363 13130 18427
rect 13194 18363 13212 18427
rect 13276 18363 13294 18427
rect 13358 18363 13376 18427
rect 13440 18363 13458 18427
rect 13522 18363 13540 18427
rect 13604 18363 13622 18427
rect 13686 18363 13704 18427
rect 13768 18363 13786 18427
rect 13850 18363 13868 18427
rect 13932 18363 13950 18427
rect 14014 18363 14032 18427
rect 14096 18363 14114 18427
rect 14178 18363 14196 18427
rect 14260 18363 14278 18427
rect 14342 18363 14360 18427
rect 14424 18363 14442 18427
rect 14506 18363 14524 18427
rect 14588 18363 14606 18427
rect 12280 18345 14666 18363
rect 363 18117 381 18181
rect 445 18117 463 18181
rect 527 18117 545 18181
rect 609 18117 627 18181
rect 691 18117 709 18181
rect 773 18117 791 18181
rect 855 18117 873 18181
rect 937 18117 955 18181
rect 1019 18117 1037 18181
rect 1101 18117 1119 18181
rect 1183 18117 1201 18181
rect 1265 18117 1283 18181
rect 1347 18117 1365 18181
rect 1429 18117 1447 18181
rect 1511 18117 1529 18181
rect 1593 18117 1611 18181
rect 1675 18117 1693 18181
rect 1757 18117 1775 18181
rect 1839 18117 1857 18181
rect 1921 18117 1939 18181
rect 2003 18117 2021 18181
rect 2085 18117 2103 18181
rect 2167 18117 2185 18181
rect 2249 18117 2267 18181
rect 2331 18117 2349 18181
rect 2413 18117 2431 18181
rect 2495 18117 2513 18181
rect 2577 18117 2594 18181
rect 2658 18117 2675 18181
rect 2739 18117 2756 18181
rect 334 18110 2771 18117
rect 334 18099 2774 18110
rect 363 18035 381 18099
rect 445 18035 463 18099
rect 527 18035 545 18099
rect 609 18035 627 18099
rect 691 18035 709 18099
rect 773 18035 791 18099
rect 855 18035 873 18099
rect 937 18035 955 18099
rect 1019 18035 1037 18099
rect 1101 18035 1119 18099
rect 1183 18035 1201 18099
rect 1265 18035 1283 18099
rect 1347 18035 1365 18099
rect 1429 18035 1447 18099
rect 1511 18035 1529 18099
rect 1593 18035 1611 18099
rect 1675 18035 1693 18099
rect 1757 18035 1775 18099
rect 1839 18035 1857 18099
rect 1921 18035 1939 18099
rect 2003 18035 2021 18099
rect 2085 18035 2103 18099
rect 2167 18035 2185 18099
rect 2249 18035 2267 18099
rect 2331 18035 2349 18099
rect 2413 18035 2431 18099
rect 2495 18035 2513 18099
rect 2577 18035 2594 18099
rect 2658 18035 2675 18099
rect 2739 18035 2756 18099
rect 334 18017 2774 18035
rect 363 17953 381 18017
rect 445 17953 463 18017
rect 527 17953 545 18017
rect 609 17953 627 18017
rect 691 17953 709 18017
rect 773 17953 791 18017
rect 855 17953 873 18017
rect 937 17953 955 18017
rect 1019 17953 1037 18017
rect 1101 17953 1119 18017
rect 1183 17953 1201 18017
rect 1265 17953 1283 18017
rect 1347 17953 1365 18017
rect 1429 17953 1447 18017
rect 1511 17953 1529 18017
rect 1593 17953 1611 18017
rect 1675 17953 1693 18017
rect 1757 17953 1775 18017
rect 1839 17953 1857 18017
rect 1921 17953 1939 18017
rect 2003 17953 2021 18017
rect 2085 17953 2103 18017
rect 2167 17953 2185 18017
rect 2249 17953 2267 18017
rect 2331 17953 2349 18017
rect 2413 17953 2431 18017
rect 2495 17953 2513 18017
rect 2577 17953 2594 18017
rect 2658 17953 2675 18017
rect 2739 17953 2756 18017
rect 334 17935 2774 17953
rect 363 17871 381 17935
rect 445 17871 463 17935
rect 527 17871 545 17935
rect 609 17871 627 17935
rect 691 17871 709 17935
rect 773 17871 791 17935
rect 855 17871 873 17935
rect 937 17871 955 17935
rect 1019 17871 1037 17935
rect 1101 17871 1119 17935
rect 1183 17871 1201 17935
rect 1265 17871 1283 17935
rect 1347 17871 1365 17935
rect 1429 17871 1447 17935
rect 1511 17871 1529 17935
rect 1593 17871 1611 17935
rect 1675 17871 1693 17935
rect 1757 17871 1775 17935
rect 1839 17871 1857 17935
rect 1921 17871 1939 17935
rect 2003 17871 2021 17935
rect 2085 17871 2103 17935
rect 2167 17871 2185 17935
rect 2249 17871 2267 17935
rect 2331 17871 2349 17935
rect 2413 17871 2431 17935
rect 2495 17871 2513 17935
rect 2577 17871 2594 17935
rect 2658 17871 2675 17935
rect 2739 17871 2756 17935
rect 334 17853 2774 17871
rect 363 17789 381 17853
rect 445 17789 463 17853
rect 527 17789 545 17853
rect 609 17789 627 17853
rect 691 17789 709 17853
rect 773 17789 791 17853
rect 855 17789 873 17853
rect 937 17789 955 17853
rect 1019 17789 1037 17853
rect 1101 17789 1119 17853
rect 1183 17789 1201 17853
rect 1265 17789 1283 17853
rect 1347 17789 1365 17853
rect 1429 17789 1447 17853
rect 1511 17789 1529 17853
rect 1593 17789 1611 17853
rect 1675 17789 1693 17853
rect 1757 17789 1775 17853
rect 1839 17789 1857 17853
rect 1921 17789 1939 17853
rect 2003 17789 2021 17853
rect 2085 17789 2103 17853
rect 2167 17789 2185 17853
rect 2249 17789 2267 17853
rect 2331 17789 2349 17853
rect 2413 17789 2431 17853
rect 2495 17789 2513 17853
rect 2577 17789 2594 17853
rect 2658 17789 2675 17853
rect 2739 17789 2756 17853
rect 334 17771 2774 17789
rect 363 17707 381 17771
rect 445 17707 463 17771
rect 527 17707 545 17771
rect 609 17707 627 17771
rect 691 17707 709 17771
rect 773 17707 791 17771
rect 855 17707 873 17771
rect 937 17707 955 17771
rect 1019 17707 1037 17771
rect 1101 17707 1119 17771
rect 1183 17707 1201 17771
rect 1265 17707 1283 17771
rect 1347 17707 1365 17771
rect 1429 17707 1447 17771
rect 1511 17707 1529 17771
rect 1593 17707 1611 17771
rect 1675 17707 1693 17771
rect 1757 17707 1775 17771
rect 1839 17707 1857 17771
rect 1921 17707 1939 17771
rect 2003 17707 2021 17771
rect 2085 17707 2103 17771
rect 2167 17707 2185 17771
rect 2249 17707 2267 17771
rect 2331 17707 2349 17771
rect 2413 17707 2431 17771
rect 2495 17707 2513 17771
rect 2577 17707 2594 17771
rect 2658 17707 2675 17771
rect 2739 17707 2756 17771
rect 334 17689 2774 17707
rect 363 17625 381 17689
rect 445 17625 463 17689
rect 527 17625 545 17689
rect 609 17625 627 17689
rect 691 17625 709 17689
rect 773 17625 791 17689
rect 855 17625 873 17689
rect 937 17625 955 17689
rect 1019 17625 1037 17689
rect 1101 17625 1119 17689
rect 1183 17625 1201 17689
rect 1265 17625 1283 17689
rect 1347 17625 1365 17689
rect 1429 17625 1447 17689
rect 1511 17625 1529 17689
rect 1593 17625 1611 17689
rect 1675 17625 1693 17689
rect 1757 17625 1775 17689
rect 1839 17625 1857 17689
rect 1921 17625 1939 17689
rect 2003 17625 2021 17689
rect 2085 17625 2103 17689
rect 2167 17625 2185 17689
rect 2249 17625 2267 17689
rect 2331 17625 2349 17689
rect 2413 17625 2431 17689
rect 2495 17625 2513 17689
rect 2577 17625 2594 17689
rect 2658 17625 2675 17689
rect 2739 17625 2756 17689
rect 3330 17986 11721 18244
rect 12295 18281 12312 18345
rect 12376 18281 12393 18345
rect 12457 18281 12474 18345
rect 12538 18281 12556 18345
rect 12620 18281 12638 18345
rect 12702 18281 12720 18345
rect 12784 18281 12802 18345
rect 12866 18281 12884 18345
rect 12948 18281 12966 18345
rect 13030 18281 13048 18345
rect 13112 18281 13130 18345
rect 13194 18281 13212 18345
rect 13276 18281 13294 18345
rect 13358 18281 13376 18345
rect 13440 18281 13458 18345
rect 13522 18281 13540 18345
rect 13604 18281 13622 18345
rect 13686 18281 13704 18345
rect 13768 18281 13786 18345
rect 13850 18281 13868 18345
rect 13932 18281 13950 18345
rect 14014 18281 14032 18345
rect 14096 18281 14114 18345
rect 14178 18281 14196 18345
rect 14260 18281 14278 18345
rect 14342 18281 14360 18345
rect 14424 18281 14442 18345
rect 14506 18281 14524 18345
rect 14588 18281 14606 18345
rect 12280 18263 14666 18281
rect 12295 18199 12312 18263
rect 12376 18199 12393 18263
rect 12457 18199 12474 18263
rect 12538 18199 12556 18263
rect 12620 18199 12638 18263
rect 12702 18199 12720 18263
rect 12784 18199 12802 18263
rect 12866 18199 12884 18263
rect 12948 18199 12966 18263
rect 13030 18199 13048 18263
rect 13112 18199 13130 18263
rect 13194 18199 13212 18263
rect 13276 18199 13294 18263
rect 13358 18199 13376 18263
rect 13440 18199 13458 18263
rect 13522 18199 13540 18263
rect 13604 18199 13622 18263
rect 13686 18199 13704 18263
rect 13768 18199 13786 18263
rect 13850 18199 13868 18263
rect 13932 18199 13950 18263
rect 14014 18199 14032 18263
rect 14096 18199 14114 18263
rect 14178 18199 14196 18263
rect 14260 18199 14278 18263
rect 14342 18199 14360 18263
rect 14424 18199 14442 18263
rect 14506 18199 14524 18263
rect 14588 18199 14606 18263
rect 12280 18181 14666 18199
rect 3585 17708 11466 17986
rect 334 17607 2774 17625
rect 363 17543 381 17607
rect 445 17543 463 17607
rect 527 17543 545 17607
rect 609 17543 627 17607
rect 691 17543 709 17607
rect 773 17543 791 17607
rect 855 17543 873 17607
rect 937 17543 955 17607
rect 1019 17543 1037 17607
rect 1101 17543 1119 17607
rect 1183 17543 1201 17607
rect 1265 17543 1283 17607
rect 1347 17543 1365 17607
rect 1429 17543 1447 17607
rect 1511 17543 1529 17607
rect 1593 17543 1611 17607
rect 1675 17543 1693 17607
rect 1757 17543 1775 17607
rect 1839 17543 1857 17607
rect 1921 17543 1939 17607
rect 2003 17543 2021 17607
rect 2085 17543 2103 17607
rect 2167 17543 2185 17607
rect 2249 17543 2267 17607
rect 2331 17543 2349 17607
rect 2413 17543 2431 17607
rect 2495 17543 2513 17607
rect 2577 17543 2594 17607
rect 2658 17543 2675 17607
rect 2739 17543 2756 17607
rect 334 17525 2795 17543
rect 363 17461 381 17525
rect 445 17461 463 17525
rect 527 17461 545 17525
rect 609 17461 627 17525
rect 691 17461 709 17525
rect 773 17461 791 17525
rect 855 17461 873 17525
rect 937 17461 955 17525
rect 1019 17461 1037 17525
rect 1101 17461 1119 17525
rect 1183 17461 1201 17525
rect 1265 17461 1283 17525
rect 1347 17461 1365 17525
rect 1429 17461 1447 17525
rect 1511 17461 1529 17525
rect 1593 17461 1611 17525
rect 1675 17461 1693 17525
rect 1757 17461 1775 17525
rect 1839 17461 1857 17525
rect 1921 17461 1939 17525
rect 2003 17461 2021 17525
rect 2085 17461 2103 17525
rect 2167 17461 2185 17525
rect 2249 17461 2267 17525
rect 2331 17461 2349 17525
rect 2413 17461 2431 17525
rect 2495 17461 2513 17525
rect 2577 17461 2594 17525
rect 2658 17461 2675 17525
rect 2739 17461 2756 17525
rect 334 17443 2795 17461
rect 363 17379 381 17443
rect 445 17379 463 17443
rect 527 17379 545 17443
rect 609 17379 627 17443
rect 691 17379 709 17443
rect 773 17379 791 17443
rect 855 17379 873 17443
rect 937 17379 955 17443
rect 1019 17379 1037 17443
rect 1101 17379 1119 17443
rect 1183 17379 1201 17443
rect 1265 17379 1283 17443
rect 1347 17379 1365 17443
rect 1429 17379 1447 17443
rect 1511 17379 1529 17443
rect 1593 17379 1611 17443
rect 1675 17379 1693 17443
rect 1757 17379 1775 17443
rect 1839 17379 1857 17443
rect 1921 17379 1939 17443
rect 2003 17379 2021 17443
rect 2085 17379 2103 17443
rect 2167 17379 2185 17443
rect 2249 17379 2267 17443
rect 2331 17379 2349 17443
rect 2413 17379 2431 17443
rect 2495 17379 2513 17443
rect 2577 17379 2594 17443
rect 2658 17379 2675 17443
rect 2739 17379 2756 17443
rect 334 17361 2795 17379
rect 363 17297 381 17361
rect 445 17297 463 17361
rect 527 17297 545 17361
rect 609 17297 627 17361
rect 691 17297 709 17361
rect 773 17297 791 17361
rect 855 17297 873 17361
rect 937 17297 955 17361
rect 1019 17297 1037 17361
rect 1101 17297 1119 17361
rect 1183 17297 1201 17361
rect 1265 17297 1283 17361
rect 1347 17297 1365 17361
rect 1429 17297 1447 17361
rect 1511 17297 1529 17361
rect 1593 17297 1611 17361
rect 1675 17297 1693 17361
rect 1757 17297 1775 17361
rect 1839 17297 1857 17361
rect 1921 17297 1939 17361
rect 2003 17297 2021 17361
rect 2085 17297 2103 17361
rect 2167 17297 2185 17361
rect 2249 17297 2267 17361
rect 2331 17297 2349 17361
rect 2413 17297 2431 17361
rect 2495 17297 2513 17361
rect 2577 17297 2594 17361
rect 2658 17297 2675 17361
rect 2739 17297 2756 17361
rect 334 17279 2795 17297
rect 363 17215 381 17279
rect 445 17215 463 17279
rect 527 17215 545 17279
rect 609 17215 627 17279
rect 691 17215 709 17279
rect 773 17215 791 17279
rect 855 17215 873 17279
rect 937 17215 955 17279
rect 1019 17215 1037 17279
rect 1101 17215 1119 17279
rect 1183 17215 1201 17279
rect 1265 17215 1283 17279
rect 1347 17215 1365 17279
rect 1429 17215 1447 17279
rect 1511 17215 1529 17279
rect 1593 17215 1611 17279
rect 1675 17215 1693 17279
rect 1757 17215 1775 17279
rect 1839 17215 1857 17279
rect 1921 17215 1939 17279
rect 2003 17215 2021 17279
rect 2085 17215 2103 17279
rect 2167 17215 2185 17279
rect 2249 17215 2267 17279
rect 2331 17215 2349 17279
rect 2413 17215 2431 17279
rect 2495 17215 2513 17279
rect 2577 17215 2594 17279
rect 2658 17215 2675 17279
rect 2739 17215 2756 17279
rect 334 17197 2795 17215
rect 363 17133 381 17197
rect 445 17133 463 17197
rect 527 17133 545 17197
rect 609 17133 627 17197
rect 691 17133 709 17197
rect 773 17133 791 17197
rect 855 17133 873 17197
rect 937 17133 955 17197
rect 1019 17133 1037 17197
rect 1101 17133 1119 17197
rect 1183 17133 1201 17197
rect 1265 17133 1283 17197
rect 1347 17133 1365 17197
rect 1429 17133 1447 17197
rect 1511 17133 1529 17197
rect 1593 17133 1611 17197
rect 1675 17133 1693 17197
rect 1757 17133 1775 17197
rect 1839 17133 1857 17197
rect 1921 17133 1939 17197
rect 2003 17133 2021 17197
rect 2085 17133 2103 17197
rect 2167 17133 2185 17197
rect 2249 17133 2267 17197
rect 2331 17133 2349 17197
rect 2413 17133 2431 17197
rect 2495 17133 2513 17197
rect 2577 17133 2594 17197
rect 2658 17133 2675 17197
rect 2739 17133 2756 17197
rect 334 17115 2795 17133
rect 363 17051 381 17115
rect 445 17051 463 17115
rect 527 17051 545 17115
rect 609 17051 627 17115
rect 691 17051 709 17115
rect 773 17051 791 17115
rect 855 17051 873 17115
rect 937 17051 955 17115
rect 1019 17051 1037 17115
rect 1101 17051 1119 17115
rect 1183 17051 1201 17115
rect 1265 17051 1283 17115
rect 1347 17051 1365 17115
rect 1429 17051 1447 17115
rect 1511 17051 1529 17115
rect 1593 17051 1611 17115
rect 1675 17051 1693 17115
rect 1757 17051 1775 17115
rect 1839 17051 1857 17115
rect 1921 17051 1939 17115
rect 2003 17051 2021 17115
rect 2085 17051 2103 17115
rect 2167 17051 2185 17115
rect 2249 17051 2267 17115
rect 2331 17051 2349 17115
rect 2413 17051 2431 17115
rect 2495 17051 2513 17115
rect 2577 17051 2594 17115
rect 2658 17051 2675 17115
rect 2739 17051 2756 17115
rect 334 17033 2795 17051
rect 363 16969 381 17033
rect 445 16969 463 17033
rect 527 16969 545 17033
rect 609 16969 627 17033
rect 691 16969 709 17033
rect 773 16969 791 17033
rect 855 16969 873 17033
rect 937 16969 955 17033
rect 1019 16969 1037 17033
rect 1101 16969 1119 17033
rect 1183 16969 1201 17033
rect 1265 16969 1283 17033
rect 1347 16969 1365 17033
rect 1429 16969 1447 17033
rect 1511 16969 1529 17033
rect 1593 16969 1611 17033
rect 1675 16969 1693 17033
rect 1757 16969 1775 17033
rect 1839 16969 1857 17033
rect 1921 16969 1939 17033
rect 2003 16969 2021 17033
rect 2085 16969 2103 17033
rect 2167 16969 2185 17033
rect 2249 16969 2267 17033
rect 2331 16969 2349 17033
rect 2413 16969 2431 17033
rect 2495 16969 2513 17033
rect 2577 16969 2594 17033
rect 2658 16969 2675 17033
rect 2739 16969 2756 17033
rect 334 16951 2795 16969
rect 363 16887 381 16951
rect 445 16887 463 16951
rect 527 16887 545 16951
rect 609 16887 627 16951
rect 691 16887 709 16951
rect 773 16887 791 16951
rect 855 16887 873 16951
rect 937 16887 955 16951
rect 1019 16887 1037 16951
rect 1101 16887 1119 16951
rect 1183 16887 1201 16951
rect 1265 16887 1283 16951
rect 1347 16887 1365 16951
rect 1429 16887 1447 16951
rect 1511 16887 1529 16951
rect 1593 16887 1611 16951
rect 1675 16887 1693 16951
rect 1757 16887 1775 16951
rect 1839 16887 1857 16951
rect 1921 16887 1939 16951
rect 2003 16887 2021 16951
rect 2085 16887 2103 16951
rect 2167 16887 2185 16951
rect 2249 16887 2267 16951
rect 2331 16887 2349 16951
rect 2413 16887 2431 16951
rect 2495 16887 2513 16951
rect 2577 16887 2594 16951
rect 2658 16887 2675 16951
rect 2739 16887 2756 16951
rect 334 16869 2795 16887
rect 363 16805 381 16869
rect 445 16805 463 16869
rect 527 16805 545 16869
rect 609 16805 627 16869
rect 691 16805 709 16869
rect 773 16805 791 16869
rect 855 16805 873 16869
rect 937 16805 955 16869
rect 1019 16805 1037 16869
rect 1101 16805 1119 16869
rect 1183 16805 1201 16869
rect 1265 16805 1283 16869
rect 1347 16805 1365 16869
rect 1429 16805 1447 16869
rect 1511 16805 1529 16869
rect 1593 16805 1611 16869
rect 1675 16805 1693 16869
rect 1757 16805 1775 16869
rect 1839 16805 1857 16869
rect 1921 16805 1939 16869
rect 2003 16805 2021 16869
rect 2085 16805 2103 16869
rect 2167 16805 2185 16869
rect 2249 16805 2267 16869
rect 2331 16805 2349 16869
rect 2413 16805 2431 16869
rect 2495 16805 2513 16869
rect 2577 16805 2594 16869
rect 2658 16805 2675 16869
rect 2739 16805 2756 16869
rect 334 16787 2795 16805
rect 363 16723 381 16787
rect 445 16723 463 16787
rect 527 16723 545 16787
rect 609 16723 627 16787
rect 691 16723 709 16787
rect 773 16723 791 16787
rect 855 16723 873 16787
rect 937 16723 955 16787
rect 1019 16723 1037 16787
rect 1101 16723 1119 16787
rect 1183 16723 1201 16787
rect 1265 16723 1283 16787
rect 1347 16723 1365 16787
rect 1429 16723 1447 16787
rect 1511 16723 1529 16787
rect 1593 16723 1611 16787
rect 1675 16723 1693 16787
rect 1757 16723 1775 16787
rect 1839 16723 1857 16787
rect 1921 16723 1939 16787
rect 2003 16723 2021 16787
rect 2085 16723 2103 16787
rect 2167 16723 2185 16787
rect 2249 16723 2267 16787
rect 2331 16723 2349 16787
rect 2413 16723 2431 16787
rect 2495 16723 2513 16787
rect 2577 16723 2594 16787
rect 2658 16723 2675 16787
rect 2739 16723 2756 16787
rect 334 16705 2795 16723
rect 363 16641 381 16705
rect 445 16641 463 16705
rect 527 16641 545 16705
rect 609 16641 627 16705
rect 691 16641 709 16705
rect 773 16641 791 16705
rect 855 16641 873 16705
rect 937 16641 955 16705
rect 1019 16641 1037 16705
rect 1101 16641 1119 16705
rect 1183 16641 1201 16705
rect 1265 16641 1283 16705
rect 1347 16641 1365 16705
rect 1429 16641 1447 16705
rect 1511 16641 1529 16705
rect 1593 16641 1611 16705
rect 1675 16641 1693 16705
rect 1757 16641 1775 16705
rect 1839 16641 1857 16705
rect 1921 16641 1939 16705
rect 2003 16641 2021 16705
rect 2085 16641 2103 16705
rect 2167 16641 2185 16705
rect 2249 16641 2267 16705
rect 2331 16641 2349 16705
rect 2413 16641 2431 16705
rect 2495 16641 2513 16705
rect 2577 16641 2594 16705
rect 2658 16641 2675 16705
rect 2739 16641 2756 16705
rect 334 16623 2795 16641
rect 363 16559 381 16623
rect 445 16559 463 16623
rect 527 16559 545 16623
rect 609 16559 627 16623
rect 691 16559 709 16623
rect 773 16559 791 16623
rect 855 16559 873 16623
rect 937 16559 955 16623
rect 1019 16559 1037 16623
rect 1101 16559 1119 16623
rect 1183 16559 1201 16623
rect 1265 16559 1283 16623
rect 1347 16559 1365 16623
rect 1429 16559 1447 16623
rect 1511 16559 1529 16623
rect 1593 16559 1611 16623
rect 1675 16559 1693 16623
rect 1757 16559 1775 16623
rect 1839 16559 1857 16623
rect 1921 16559 1939 16623
rect 2003 16559 2021 16623
rect 2085 16559 2103 16623
rect 2167 16559 2185 16623
rect 2249 16559 2267 16623
rect 2331 16559 2349 16623
rect 2413 16559 2431 16623
rect 2495 16559 2513 16623
rect 2577 16559 2594 16623
rect 2658 16559 2675 16623
rect 2739 16559 2756 16623
rect 3851 17483 11200 17708
rect 12295 18117 12312 18181
rect 12376 18117 12393 18181
rect 12457 18117 12474 18181
rect 12538 18117 12556 18181
rect 12620 18117 12638 18181
rect 12702 18117 12720 18181
rect 12784 18117 12802 18181
rect 12866 18117 12884 18181
rect 12948 18117 12966 18181
rect 13030 18117 13048 18181
rect 13112 18117 13130 18181
rect 13194 18117 13212 18181
rect 13276 18117 13294 18181
rect 13358 18117 13376 18181
rect 13440 18117 13458 18181
rect 13522 18117 13540 18181
rect 13604 18117 13622 18181
rect 13686 18117 13704 18181
rect 13768 18117 13786 18181
rect 13850 18117 13868 18181
rect 13932 18117 13950 18181
rect 14014 18117 14032 18181
rect 14096 18117 14114 18181
rect 14178 18117 14196 18181
rect 14260 18117 14278 18181
rect 14342 18117 14360 18181
rect 14424 18117 14442 18181
rect 14506 18117 14524 18181
rect 14588 18117 14606 18181
rect 12280 18110 14666 18117
rect 12277 18099 14666 18110
rect 12295 18035 12312 18099
rect 12376 18035 12393 18099
rect 12457 18035 12474 18099
rect 12538 18035 12556 18099
rect 12620 18035 12638 18099
rect 12702 18035 12720 18099
rect 12784 18035 12802 18099
rect 12866 18035 12884 18099
rect 12948 18035 12966 18099
rect 13030 18035 13048 18099
rect 13112 18035 13130 18099
rect 13194 18035 13212 18099
rect 13276 18035 13294 18099
rect 13358 18035 13376 18099
rect 13440 18035 13458 18099
rect 13522 18035 13540 18099
rect 13604 18035 13622 18099
rect 13686 18035 13704 18099
rect 13768 18035 13786 18099
rect 13850 18035 13868 18099
rect 13932 18035 13950 18099
rect 14014 18035 14032 18099
rect 14096 18035 14114 18099
rect 14178 18035 14196 18099
rect 14260 18035 14278 18099
rect 14342 18035 14360 18099
rect 14424 18035 14442 18099
rect 14506 18035 14524 18099
rect 14588 18035 14606 18099
rect 12277 18017 14666 18035
rect 12295 17953 12312 18017
rect 12376 17953 12393 18017
rect 12457 17953 12474 18017
rect 12538 17953 12556 18017
rect 12620 17953 12638 18017
rect 12702 17953 12720 18017
rect 12784 17953 12802 18017
rect 12866 17953 12884 18017
rect 12948 17953 12966 18017
rect 13030 17953 13048 18017
rect 13112 17953 13130 18017
rect 13194 17953 13212 18017
rect 13276 17953 13294 18017
rect 13358 17953 13376 18017
rect 13440 17953 13458 18017
rect 13522 17953 13540 18017
rect 13604 17953 13622 18017
rect 13686 17953 13704 18017
rect 13768 17953 13786 18017
rect 13850 17953 13868 18017
rect 13932 17953 13950 18017
rect 14014 17953 14032 18017
rect 14096 17953 14114 18017
rect 14178 17953 14196 18017
rect 14260 17953 14278 18017
rect 14342 17953 14360 18017
rect 14424 17953 14442 18017
rect 14506 17953 14524 18017
rect 14588 17953 14606 18017
rect 12277 17935 14666 17953
rect 12295 17871 12312 17935
rect 12376 17871 12393 17935
rect 12457 17871 12474 17935
rect 12538 17871 12556 17935
rect 12620 17871 12638 17935
rect 12702 17871 12720 17935
rect 12784 17871 12802 17935
rect 12866 17871 12884 17935
rect 12948 17871 12966 17935
rect 13030 17871 13048 17935
rect 13112 17871 13130 17935
rect 13194 17871 13212 17935
rect 13276 17871 13294 17935
rect 13358 17871 13376 17935
rect 13440 17871 13458 17935
rect 13522 17871 13540 17935
rect 13604 17871 13622 17935
rect 13686 17871 13704 17935
rect 13768 17871 13786 17935
rect 13850 17871 13868 17935
rect 13932 17871 13950 17935
rect 14014 17871 14032 17935
rect 14096 17871 14114 17935
rect 14178 17871 14196 17935
rect 14260 17871 14278 17935
rect 14342 17871 14360 17935
rect 14424 17871 14442 17935
rect 14506 17871 14524 17935
rect 14588 17871 14606 17935
rect 12277 17853 14666 17871
rect 12295 17789 12312 17853
rect 12376 17789 12393 17853
rect 12457 17789 12474 17853
rect 12538 17789 12556 17853
rect 12620 17789 12638 17853
rect 12702 17789 12720 17853
rect 12784 17789 12802 17853
rect 12866 17789 12884 17853
rect 12948 17789 12966 17853
rect 13030 17789 13048 17853
rect 13112 17789 13130 17853
rect 13194 17789 13212 17853
rect 13276 17789 13294 17853
rect 13358 17789 13376 17853
rect 13440 17789 13458 17853
rect 13522 17789 13540 17853
rect 13604 17789 13622 17853
rect 13686 17789 13704 17853
rect 13768 17789 13786 17853
rect 13850 17789 13868 17853
rect 13932 17789 13950 17853
rect 14014 17789 14032 17853
rect 14096 17789 14114 17853
rect 14178 17789 14196 17853
rect 14260 17789 14278 17853
rect 14342 17789 14360 17853
rect 14424 17789 14442 17853
rect 14506 17789 14524 17853
rect 14588 17789 14606 17853
rect 12277 17771 14666 17789
rect 12295 17707 12312 17771
rect 12376 17707 12393 17771
rect 12457 17707 12474 17771
rect 12538 17707 12556 17771
rect 12620 17707 12638 17771
rect 12702 17707 12720 17771
rect 12784 17707 12802 17771
rect 12866 17707 12884 17771
rect 12948 17707 12966 17771
rect 13030 17707 13048 17771
rect 13112 17707 13130 17771
rect 13194 17707 13212 17771
rect 13276 17707 13294 17771
rect 13358 17707 13376 17771
rect 13440 17707 13458 17771
rect 13522 17707 13540 17771
rect 13604 17707 13622 17771
rect 13686 17707 13704 17771
rect 13768 17707 13786 17771
rect 13850 17707 13868 17771
rect 13932 17707 13950 17771
rect 14014 17707 14032 17771
rect 14096 17707 14114 17771
rect 14178 17707 14196 17771
rect 14260 17707 14278 17771
rect 14342 17707 14360 17771
rect 14424 17707 14442 17771
rect 14506 17707 14524 17771
rect 14588 17707 14606 17771
rect 12277 17689 14666 17707
rect 4093 17198 10958 17483
rect 4370 16937 10681 17198
rect 334 16524 2795 16559
rect 4634 16524 10417 16937
rect 12295 17625 12312 17689
rect 12376 17625 12393 17689
rect 12457 17625 12474 17689
rect 12538 17625 12556 17689
rect 12620 17625 12638 17689
rect 12702 17625 12720 17689
rect 12784 17625 12802 17689
rect 12866 17625 12884 17689
rect 12948 17625 12966 17689
rect 13030 17625 13048 17689
rect 13112 17625 13130 17689
rect 13194 17625 13212 17689
rect 13276 17625 13294 17689
rect 13358 17625 13376 17689
rect 13440 17625 13458 17689
rect 13522 17625 13540 17689
rect 13604 17625 13622 17689
rect 13686 17625 13704 17689
rect 13768 17625 13786 17689
rect 13850 17625 13868 17689
rect 13932 17625 13950 17689
rect 14014 17625 14032 17689
rect 14096 17625 14114 17689
rect 14178 17625 14196 17689
rect 14260 17625 14278 17689
rect 14342 17625 14360 17689
rect 14424 17625 14442 17689
rect 14506 17625 14524 17689
rect 14588 17625 14606 17689
rect 12277 17607 14666 17625
rect 12295 17543 12312 17607
rect 12376 17543 12393 17607
rect 12457 17543 12474 17607
rect 12538 17543 12556 17607
rect 12620 17543 12638 17607
rect 12702 17543 12720 17607
rect 12784 17543 12802 17607
rect 12866 17543 12884 17607
rect 12948 17543 12966 17607
rect 13030 17543 13048 17607
rect 13112 17543 13130 17607
rect 13194 17543 13212 17607
rect 13276 17543 13294 17607
rect 13358 17543 13376 17607
rect 13440 17543 13458 17607
rect 13522 17543 13540 17607
rect 13604 17543 13622 17607
rect 13686 17543 13704 17607
rect 13768 17543 13786 17607
rect 13850 17543 13868 17607
rect 13932 17543 13950 17607
rect 14014 17543 14032 17607
rect 14096 17543 14114 17607
rect 14178 17543 14196 17607
rect 14260 17543 14278 17607
rect 14342 17543 14360 17607
rect 14424 17543 14442 17607
rect 14506 17543 14524 17607
rect 14588 17543 14606 17607
rect 12256 17525 14666 17543
rect 12295 17461 12312 17525
rect 12376 17461 12393 17525
rect 12457 17461 12474 17525
rect 12538 17461 12556 17525
rect 12620 17461 12638 17525
rect 12702 17461 12720 17525
rect 12784 17461 12802 17525
rect 12866 17461 12884 17525
rect 12948 17461 12966 17525
rect 13030 17461 13048 17525
rect 13112 17461 13130 17525
rect 13194 17461 13212 17525
rect 13276 17461 13294 17525
rect 13358 17461 13376 17525
rect 13440 17461 13458 17525
rect 13522 17461 13540 17525
rect 13604 17461 13622 17525
rect 13686 17461 13704 17525
rect 13768 17461 13786 17525
rect 13850 17461 13868 17525
rect 13932 17461 13950 17525
rect 14014 17461 14032 17525
rect 14096 17461 14114 17525
rect 14178 17461 14196 17525
rect 14260 17461 14278 17525
rect 14342 17461 14360 17525
rect 14424 17461 14442 17525
rect 14506 17461 14524 17525
rect 14588 17461 14606 17525
rect 12256 17443 14666 17461
rect 12295 17379 12312 17443
rect 12376 17379 12393 17443
rect 12457 17379 12474 17443
rect 12538 17379 12556 17443
rect 12620 17379 12638 17443
rect 12702 17379 12720 17443
rect 12784 17379 12802 17443
rect 12866 17379 12884 17443
rect 12948 17379 12966 17443
rect 13030 17379 13048 17443
rect 13112 17379 13130 17443
rect 13194 17379 13212 17443
rect 13276 17379 13294 17443
rect 13358 17379 13376 17443
rect 13440 17379 13458 17443
rect 13522 17379 13540 17443
rect 13604 17379 13622 17443
rect 13686 17379 13704 17443
rect 13768 17379 13786 17443
rect 13850 17379 13868 17443
rect 13932 17379 13950 17443
rect 14014 17379 14032 17443
rect 14096 17379 14114 17443
rect 14178 17379 14196 17443
rect 14260 17379 14278 17443
rect 14342 17379 14360 17443
rect 14424 17379 14442 17443
rect 14506 17379 14524 17443
rect 14588 17379 14606 17443
rect 12256 17361 14666 17379
rect 12295 17297 12312 17361
rect 12376 17297 12393 17361
rect 12457 17297 12474 17361
rect 12538 17297 12556 17361
rect 12620 17297 12638 17361
rect 12702 17297 12720 17361
rect 12784 17297 12802 17361
rect 12866 17297 12884 17361
rect 12948 17297 12966 17361
rect 13030 17297 13048 17361
rect 13112 17297 13130 17361
rect 13194 17297 13212 17361
rect 13276 17297 13294 17361
rect 13358 17297 13376 17361
rect 13440 17297 13458 17361
rect 13522 17297 13540 17361
rect 13604 17297 13622 17361
rect 13686 17297 13704 17361
rect 13768 17297 13786 17361
rect 13850 17297 13868 17361
rect 13932 17297 13950 17361
rect 14014 17297 14032 17361
rect 14096 17297 14114 17361
rect 14178 17297 14196 17361
rect 14260 17297 14278 17361
rect 14342 17297 14360 17361
rect 14424 17297 14442 17361
rect 14506 17297 14524 17361
rect 14588 17297 14606 17361
rect 12256 17279 14666 17297
rect 12295 17215 12312 17279
rect 12376 17215 12393 17279
rect 12457 17215 12474 17279
rect 12538 17215 12556 17279
rect 12620 17215 12638 17279
rect 12702 17215 12720 17279
rect 12784 17215 12802 17279
rect 12866 17215 12884 17279
rect 12948 17215 12966 17279
rect 13030 17215 13048 17279
rect 13112 17215 13130 17279
rect 13194 17215 13212 17279
rect 13276 17215 13294 17279
rect 13358 17215 13376 17279
rect 13440 17215 13458 17279
rect 13522 17215 13540 17279
rect 13604 17215 13622 17279
rect 13686 17215 13704 17279
rect 13768 17215 13786 17279
rect 13850 17215 13868 17279
rect 13932 17215 13950 17279
rect 14014 17215 14032 17279
rect 14096 17215 14114 17279
rect 14178 17215 14196 17279
rect 14260 17215 14278 17279
rect 14342 17215 14360 17279
rect 14424 17215 14442 17279
rect 14506 17215 14524 17279
rect 14588 17215 14606 17279
rect 12256 17197 14666 17215
rect 12295 17133 12312 17197
rect 12376 17133 12393 17197
rect 12457 17133 12474 17197
rect 12538 17133 12556 17197
rect 12620 17133 12638 17197
rect 12702 17133 12720 17197
rect 12784 17133 12802 17197
rect 12866 17133 12884 17197
rect 12948 17133 12966 17197
rect 13030 17133 13048 17197
rect 13112 17133 13130 17197
rect 13194 17133 13212 17197
rect 13276 17133 13294 17197
rect 13358 17133 13376 17197
rect 13440 17133 13458 17197
rect 13522 17133 13540 17197
rect 13604 17133 13622 17197
rect 13686 17133 13704 17197
rect 13768 17133 13786 17197
rect 13850 17133 13868 17197
rect 13932 17133 13950 17197
rect 14014 17133 14032 17197
rect 14096 17133 14114 17197
rect 14178 17133 14196 17197
rect 14260 17133 14278 17197
rect 14342 17133 14360 17197
rect 14424 17133 14442 17197
rect 14506 17133 14524 17197
rect 14588 17133 14606 17197
rect 12256 17115 14666 17133
rect 12295 17051 12312 17115
rect 12376 17051 12393 17115
rect 12457 17051 12474 17115
rect 12538 17051 12556 17115
rect 12620 17051 12638 17115
rect 12702 17051 12720 17115
rect 12784 17051 12802 17115
rect 12866 17051 12884 17115
rect 12948 17051 12966 17115
rect 13030 17051 13048 17115
rect 13112 17051 13130 17115
rect 13194 17051 13212 17115
rect 13276 17051 13294 17115
rect 13358 17051 13376 17115
rect 13440 17051 13458 17115
rect 13522 17051 13540 17115
rect 13604 17051 13622 17115
rect 13686 17051 13704 17115
rect 13768 17051 13786 17115
rect 13850 17051 13868 17115
rect 13932 17051 13950 17115
rect 14014 17051 14032 17115
rect 14096 17051 14114 17115
rect 14178 17051 14196 17115
rect 14260 17051 14278 17115
rect 14342 17051 14360 17115
rect 14424 17051 14442 17115
rect 14506 17051 14524 17115
rect 14588 17051 14606 17115
rect 12256 17033 14666 17051
rect 12295 16969 12312 17033
rect 12376 16969 12393 17033
rect 12457 16969 12474 17033
rect 12538 16969 12556 17033
rect 12620 16969 12638 17033
rect 12702 16969 12720 17033
rect 12784 16969 12802 17033
rect 12866 16969 12884 17033
rect 12948 16969 12966 17033
rect 13030 16969 13048 17033
rect 13112 16969 13130 17033
rect 13194 16969 13212 17033
rect 13276 16969 13294 17033
rect 13358 16969 13376 17033
rect 13440 16969 13458 17033
rect 13522 16969 13540 17033
rect 13604 16969 13622 17033
rect 13686 16969 13704 17033
rect 13768 16969 13786 17033
rect 13850 16969 13868 17033
rect 13932 16969 13950 17033
rect 14014 16969 14032 17033
rect 14096 16969 14114 17033
rect 14178 16969 14196 17033
rect 14260 16969 14278 17033
rect 14342 16969 14360 17033
rect 14424 16969 14442 17033
rect 14506 16969 14524 17033
rect 14588 16969 14606 17033
rect 12256 16951 14666 16969
rect 12295 16887 12312 16951
rect 12376 16887 12393 16951
rect 12457 16887 12474 16951
rect 12538 16887 12556 16951
rect 12620 16887 12638 16951
rect 12702 16887 12720 16951
rect 12784 16887 12802 16951
rect 12866 16887 12884 16951
rect 12948 16887 12966 16951
rect 13030 16887 13048 16951
rect 13112 16887 13130 16951
rect 13194 16887 13212 16951
rect 13276 16887 13294 16951
rect 13358 16887 13376 16951
rect 13440 16887 13458 16951
rect 13522 16887 13540 16951
rect 13604 16887 13622 16951
rect 13686 16887 13704 16951
rect 13768 16887 13786 16951
rect 13850 16887 13868 16951
rect 13932 16887 13950 16951
rect 14014 16887 14032 16951
rect 14096 16887 14114 16951
rect 14178 16887 14196 16951
rect 14260 16887 14278 16951
rect 14342 16887 14360 16951
rect 14424 16887 14442 16951
rect 14506 16887 14524 16951
rect 14588 16887 14606 16951
rect 12256 16869 14666 16887
rect 12295 16805 12312 16869
rect 12376 16805 12393 16869
rect 12457 16805 12474 16869
rect 12538 16805 12556 16869
rect 12620 16805 12638 16869
rect 12702 16805 12720 16869
rect 12784 16805 12802 16869
rect 12866 16805 12884 16869
rect 12948 16805 12966 16869
rect 13030 16805 13048 16869
rect 13112 16805 13130 16869
rect 13194 16805 13212 16869
rect 13276 16805 13294 16869
rect 13358 16805 13376 16869
rect 13440 16805 13458 16869
rect 13522 16805 13540 16869
rect 13604 16805 13622 16869
rect 13686 16805 13704 16869
rect 13768 16805 13786 16869
rect 13850 16805 13868 16869
rect 13932 16805 13950 16869
rect 14014 16805 14032 16869
rect 14096 16805 14114 16869
rect 14178 16805 14196 16869
rect 14260 16805 14278 16869
rect 14342 16805 14360 16869
rect 14424 16805 14442 16869
rect 14506 16805 14524 16869
rect 14588 16805 14606 16869
rect 12256 16787 14666 16805
rect 12295 16723 12312 16787
rect 12376 16723 12393 16787
rect 12457 16723 12474 16787
rect 12538 16723 12556 16787
rect 12620 16723 12638 16787
rect 12702 16723 12720 16787
rect 12784 16723 12802 16787
rect 12866 16723 12884 16787
rect 12948 16723 12966 16787
rect 13030 16723 13048 16787
rect 13112 16723 13130 16787
rect 13194 16723 13212 16787
rect 13276 16723 13294 16787
rect 13358 16723 13376 16787
rect 13440 16723 13458 16787
rect 13522 16723 13540 16787
rect 13604 16723 13622 16787
rect 13686 16723 13704 16787
rect 13768 16723 13786 16787
rect 13850 16723 13868 16787
rect 13932 16723 13950 16787
rect 14014 16723 14032 16787
rect 14096 16723 14114 16787
rect 14178 16723 14196 16787
rect 14260 16723 14278 16787
rect 14342 16723 14360 16787
rect 14424 16723 14442 16787
rect 14506 16723 14524 16787
rect 14588 16723 14606 16787
rect 12256 16705 14666 16723
rect 12295 16641 12312 16705
rect 12376 16641 12393 16705
rect 12457 16641 12474 16705
rect 12538 16641 12556 16705
rect 12620 16641 12638 16705
rect 12702 16641 12720 16705
rect 12784 16641 12802 16705
rect 12866 16641 12884 16705
rect 12948 16641 12966 16705
rect 13030 16641 13048 16705
rect 13112 16641 13130 16705
rect 13194 16641 13212 16705
rect 13276 16641 13294 16705
rect 13358 16641 13376 16705
rect 13440 16641 13458 16705
rect 13522 16641 13540 16705
rect 13604 16641 13622 16705
rect 13686 16641 13704 16705
rect 13768 16641 13786 16705
rect 13850 16641 13868 16705
rect 13932 16641 13950 16705
rect 14014 16641 14032 16705
rect 14096 16641 14114 16705
rect 14178 16641 14196 16705
rect 14260 16641 14278 16705
rect 14342 16641 14360 16705
rect 14424 16641 14442 16705
rect 14506 16641 14524 16705
rect 14588 16641 14606 16705
rect 12256 16623 14666 16641
rect 12295 16559 12312 16623
rect 12376 16559 12393 16623
rect 12457 16559 12474 16623
rect 12538 16559 12556 16623
rect 12620 16559 12638 16623
rect 12702 16559 12720 16623
rect 12784 16559 12802 16623
rect 12866 16559 12884 16623
rect 12948 16559 12966 16623
rect 13030 16559 13048 16623
rect 13112 16559 13130 16623
rect 13194 16559 13212 16623
rect 13276 16559 13294 16623
rect 13358 16559 13376 16623
rect 13440 16559 13458 16623
rect 13522 16559 13540 16623
rect 13604 16559 13622 16623
rect 13686 16559 13704 16623
rect 13768 16559 13786 16623
rect 13850 16559 13868 16623
rect 13932 16559 13950 16623
rect 14014 16559 14032 16623
rect 14096 16559 14114 16623
rect 14178 16559 14196 16623
rect 14260 16559 14278 16623
rect 14342 16559 14360 16623
rect 14424 16559 14442 16623
rect 14506 16559 14524 16623
rect 14588 16559 14606 16623
rect 381 16460 397 16524
rect 461 16460 477 16524
rect 541 16460 557 16524
rect 621 16460 637 16524
rect 701 16460 717 16524
rect 781 16460 797 16524
rect 861 16460 877 16524
rect 941 16460 957 16524
rect 1021 16460 1037 16524
rect 1101 16460 1117 16524
rect 1181 16460 1197 16524
rect 1261 16460 1277 16524
rect 1341 16460 1357 16524
rect 1421 16460 1437 16524
rect 1501 16460 1517 16524
rect 1581 16460 1597 16524
rect 1661 16460 1677 16524
rect 1741 16460 1757 16524
rect 1821 16460 1837 16524
rect 1901 16460 1917 16524
rect 1981 16460 1997 16524
rect 2061 16460 2077 16524
rect 2141 16460 2157 16524
rect 2221 16460 2237 16524
rect 2301 16460 2317 16524
rect 2381 16460 2397 16524
rect 2461 16460 2477 16524
rect 2541 16460 2557 16524
rect 2621 16460 2637 16524
rect 2701 16460 2717 16524
rect 2781 16518 2795 16524
rect 2781 16460 2797 16518
rect 2861 16460 2877 16518
rect 2941 16460 2957 16518
rect 3021 16460 3037 16518
rect 3101 16460 3117 16518
rect 3181 16460 3197 16518
rect 3261 16460 3277 16518
rect 3341 16460 3357 16518
rect 3421 16460 3437 16518
rect 3501 16460 3517 16518
rect 3581 16460 3597 16518
rect 3661 16460 3677 16518
rect 3741 16509 3754 16518
rect 3741 16460 3757 16509
rect 3821 16460 3837 16509
rect 3901 16460 3917 16509
rect 3981 16460 3997 16509
rect 4061 16460 4077 16509
rect 4141 16460 4157 16509
rect 4221 16460 4237 16509
rect 4301 16460 4317 16491
rect 4381 16460 4397 16491
rect 4461 16460 4477 16491
rect 4541 16460 4557 16491
rect 4634 16491 4637 16524
rect 4621 16460 4637 16491
rect 4701 16460 4717 16524
rect 4781 16460 4797 16524
rect 4861 16491 10417 16524
rect 12256 16518 14666 16559
rect 11297 16509 14666 16518
rect 10801 16491 14666 16509
rect 4861 16460 14666 16491
rect 334 16443 14666 16460
rect 381 16379 397 16443
rect 461 16379 477 16443
rect 541 16379 557 16443
rect 621 16379 637 16443
rect 701 16379 717 16443
rect 781 16379 797 16443
rect 861 16379 877 16443
rect 941 16379 957 16443
rect 1021 16379 1037 16443
rect 1101 16379 1117 16443
rect 1181 16379 1197 16443
rect 1261 16379 1277 16443
rect 1341 16379 1357 16443
rect 1421 16379 1437 16443
rect 1501 16379 1517 16443
rect 1581 16379 1597 16443
rect 1661 16379 1677 16443
rect 1741 16379 1757 16443
rect 1821 16379 1837 16443
rect 1901 16379 1917 16443
rect 1981 16379 1997 16443
rect 2061 16379 2077 16443
rect 2141 16379 2157 16443
rect 2221 16379 2237 16443
rect 2301 16379 2317 16443
rect 2381 16379 2397 16443
rect 2461 16379 2477 16443
rect 2541 16379 2557 16443
rect 2621 16379 2637 16443
rect 2701 16379 2717 16443
rect 2781 16379 2797 16443
rect 2861 16379 2877 16443
rect 2941 16379 2957 16443
rect 3021 16379 3037 16443
rect 3101 16379 3117 16443
rect 3181 16379 3197 16443
rect 3261 16379 3277 16443
rect 3341 16379 3357 16443
rect 3421 16379 3437 16443
rect 3501 16379 3517 16443
rect 3581 16379 3597 16443
rect 3661 16379 3677 16443
rect 3741 16379 3757 16443
rect 3821 16379 3837 16443
rect 3901 16379 3917 16443
rect 3981 16379 3997 16443
rect 4061 16379 4077 16443
rect 4141 16379 4157 16443
rect 4221 16379 4237 16443
rect 4301 16379 4317 16443
rect 4381 16379 4397 16443
rect 4461 16379 4477 16443
rect 4541 16379 4557 16443
rect 4621 16379 4637 16443
rect 4701 16379 4717 16443
rect 4781 16379 4797 16443
rect 4861 16379 14666 16443
rect 334 16362 14666 16379
rect 381 16298 397 16362
rect 461 16298 477 16362
rect 541 16298 557 16362
rect 621 16298 637 16362
rect 701 16298 717 16362
rect 781 16298 797 16362
rect 861 16298 877 16362
rect 941 16298 957 16362
rect 1021 16298 1037 16362
rect 1101 16298 1117 16362
rect 1181 16298 1197 16362
rect 1261 16298 1277 16362
rect 1341 16298 1357 16362
rect 1421 16298 1437 16362
rect 1501 16298 1517 16362
rect 1581 16298 1597 16362
rect 1661 16298 1677 16362
rect 1741 16298 1757 16362
rect 1821 16298 1837 16362
rect 1901 16298 1917 16362
rect 1981 16298 1997 16362
rect 2061 16298 2077 16362
rect 2141 16298 2157 16362
rect 2221 16298 2237 16362
rect 2301 16298 2317 16362
rect 2381 16298 2397 16362
rect 2461 16298 2477 16362
rect 2541 16298 2557 16362
rect 2621 16298 2637 16362
rect 2701 16298 2717 16362
rect 2781 16298 2797 16362
rect 2861 16298 2877 16362
rect 2941 16298 2957 16362
rect 3021 16298 3037 16362
rect 3101 16298 3117 16362
rect 3181 16298 3197 16362
rect 3261 16298 3277 16362
rect 3341 16298 3357 16362
rect 3421 16298 3437 16362
rect 3501 16298 3517 16362
rect 3581 16298 3597 16362
rect 3661 16298 3677 16362
rect 3741 16298 3757 16362
rect 3821 16298 3837 16362
rect 3901 16298 3917 16362
rect 3981 16298 3997 16362
rect 4061 16298 4077 16362
rect 4141 16298 4157 16362
rect 4221 16298 4237 16362
rect 4301 16298 4317 16362
rect 4381 16298 4397 16362
rect 4461 16298 4477 16362
rect 4541 16298 4557 16362
rect 4621 16298 4637 16362
rect 4701 16298 4717 16362
rect 4781 16298 4797 16362
rect 4861 16298 14666 16362
rect 334 16281 14666 16298
rect 381 16217 397 16281
rect 461 16217 477 16281
rect 541 16217 557 16281
rect 621 16217 637 16281
rect 701 16217 717 16281
rect 781 16217 797 16281
rect 861 16217 877 16281
rect 941 16217 957 16281
rect 1021 16217 1037 16281
rect 1101 16217 1117 16281
rect 1181 16217 1197 16281
rect 1261 16217 1277 16281
rect 1341 16217 1357 16281
rect 1421 16217 1437 16281
rect 1501 16217 1517 16281
rect 1581 16217 1597 16281
rect 1661 16217 1677 16281
rect 1741 16217 1757 16281
rect 1821 16217 1837 16281
rect 1901 16217 1917 16281
rect 1981 16217 1997 16281
rect 2061 16217 2077 16281
rect 2141 16217 2157 16281
rect 2221 16217 2237 16281
rect 2301 16217 2317 16281
rect 2381 16217 2397 16281
rect 2461 16217 2477 16281
rect 2541 16217 2557 16281
rect 2621 16217 2637 16281
rect 2701 16217 2717 16281
rect 2781 16217 2797 16281
rect 2861 16217 2877 16281
rect 2941 16217 2957 16281
rect 3021 16217 3037 16281
rect 3101 16217 3117 16281
rect 3181 16217 3197 16281
rect 3261 16217 3277 16281
rect 3341 16217 3357 16281
rect 3421 16217 3437 16281
rect 3501 16217 3517 16281
rect 3581 16217 3597 16281
rect 3661 16217 3677 16281
rect 3741 16217 3757 16281
rect 3821 16217 3837 16281
rect 3901 16217 3917 16281
rect 3981 16217 3997 16281
rect 4061 16217 4077 16281
rect 4141 16217 4157 16281
rect 4221 16217 4237 16281
rect 4301 16217 4317 16281
rect 4381 16217 4397 16281
rect 4461 16217 4477 16281
rect 4541 16217 4557 16281
rect 4621 16217 4637 16281
rect 4701 16217 4717 16281
rect 4781 16217 4797 16281
rect 4861 16217 14666 16281
rect 334 16200 14666 16217
rect 381 16136 397 16200
rect 461 16136 477 16200
rect 541 16136 557 16200
rect 621 16136 637 16200
rect 701 16136 717 16200
rect 781 16136 797 16200
rect 861 16136 877 16200
rect 941 16136 957 16200
rect 1021 16136 1037 16200
rect 1101 16136 1117 16200
rect 1181 16136 1197 16200
rect 1261 16136 1277 16200
rect 1341 16136 1357 16200
rect 1421 16136 1437 16200
rect 1501 16136 1517 16200
rect 1581 16136 1597 16200
rect 1661 16136 1677 16200
rect 1741 16136 1757 16200
rect 1821 16136 1837 16200
rect 1901 16136 1917 16200
rect 1981 16136 1997 16200
rect 2061 16136 2077 16200
rect 2141 16136 2157 16200
rect 2221 16136 2237 16200
rect 2301 16136 2317 16200
rect 2381 16136 2397 16200
rect 2461 16136 2477 16200
rect 2541 16136 2557 16200
rect 2621 16136 2637 16200
rect 2701 16136 2717 16200
rect 2781 16136 2797 16200
rect 2861 16136 2877 16200
rect 2941 16136 2957 16200
rect 3021 16136 3037 16200
rect 3101 16136 3117 16200
rect 3181 16136 3197 16200
rect 3261 16136 3277 16200
rect 3341 16136 3357 16200
rect 3421 16136 3437 16200
rect 3501 16136 3517 16200
rect 3581 16136 3597 16200
rect 3661 16136 3677 16200
rect 3741 16136 3757 16200
rect 3821 16136 3837 16200
rect 3901 16136 3917 16200
rect 3981 16136 3997 16200
rect 4061 16136 4077 16200
rect 4141 16136 4157 16200
rect 4221 16136 4237 16200
rect 4301 16136 4317 16200
rect 4381 16136 4397 16200
rect 4461 16136 4477 16200
rect 4541 16136 4557 16200
rect 4621 16136 4637 16200
rect 4701 16136 4717 16200
rect 4781 16136 4797 16200
rect 4861 16136 14666 16200
rect 334 16119 14666 16136
rect 381 16055 397 16119
rect 461 16055 477 16119
rect 541 16055 557 16119
rect 621 16055 637 16119
rect 701 16055 717 16119
rect 781 16055 797 16119
rect 861 16055 877 16119
rect 941 16055 957 16119
rect 1021 16055 1037 16119
rect 1101 16055 1117 16119
rect 1181 16055 1197 16119
rect 1261 16055 1277 16119
rect 1341 16055 1357 16119
rect 1421 16055 1437 16119
rect 1501 16055 1517 16119
rect 1581 16055 1597 16119
rect 1661 16055 1677 16119
rect 1741 16055 1757 16119
rect 1821 16055 1837 16119
rect 1901 16055 1917 16119
rect 1981 16055 1997 16119
rect 2061 16055 2077 16119
rect 2141 16055 2157 16119
rect 2221 16055 2237 16119
rect 2301 16055 2317 16119
rect 2381 16055 2397 16119
rect 2461 16055 2477 16119
rect 2541 16055 2557 16119
rect 2621 16055 2637 16119
rect 2701 16055 2717 16119
rect 2781 16055 2797 16119
rect 2861 16055 2877 16119
rect 2941 16055 2957 16119
rect 3021 16055 3037 16119
rect 3101 16055 3117 16119
rect 3181 16055 3197 16119
rect 3261 16055 3277 16119
rect 3341 16055 3357 16119
rect 3421 16055 3437 16119
rect 3501 16055 3517 16119
rect 3581 16055 3597 16119
rect 3661 16055 3677 16119
rect 3741 16055 3757 16119
rect 3821 16055 3837 16119
rect 3901 16055 3917 16119
rect 3981 16055 3997 16119
rect 4061 16055 4077 16119
rect 4141 16055 4157 16119
rect 4221 16055 4237 16119
rect 4301 16055 4317 16119
rect 4381 16055 4397 16119
rect 4461 16055 4477 16119
rect 4541 16055 4557 16119
rect 4621 16055 4637 16119
rect 4701 16055 4717 16119
rect 4781 16055 4797 16119
rect 4861 16055 14666 16119
rect 334 16038 14666 16055
rect 381 15974 397 16038
rect 461 15974 477 16038
rect 541 15974 557 16038
rect 621 15974 637 16038
rect 701 15974 717 16038
rect 781 15974 797 16038
rect 861 15974 877 16038
rect 941 15974 957 16038
rect 1021 15974 1037 16038
rect 1101 15974 1117 16038
rect 1181 15974 1197 16038
rect 1261 15974 1277 16038
rect 1341 15974 1357 16038
rect 1421 15974 1437 16038
rect 1501 15974 1517 16038
rect 1581 15974 1597 16038
rect 1661 15974 1677 16038
rect 1741 15974 1757 16038
rect 1821 15974 1837 16038
rect 1901 15974 1917 16038
rect 1981 15974 1997 16038
rect 2061 15974 2077 16038
rect 2141 15974 2157 16038
rect 2221 15974 2237 16038
rect 2301 15974 2317 16038
rect 2381 15974 2397 16038
rect 2461 15974 2477 16038
rect 2541 15974 2557 16038
rect 2621 15974 2637 16038
rect 2701 15974 2717 16038
rect 2781 15974 2797 16038
rect 2861 15974 2877 16038
rect 2941 15974 2957 16038
rect 3021 15974 3037 16038
rect 3101 15974 3117 16038
rect 3181 15974 3197 16038
rect 3261 15974 3277 16038
rect 3341 15974 3357 16038
rect 3421 15974 3437 16038
rect 3501 15974 3517 16038
rect 3581 15974 3597 16038
rect 3661 15974 3677 16038
rect 3741 15974 3757 16038
rect 3821 15974 3837 16038
rect 3901 15974 3917 16038
rect 3981 15974 3997 16038
rect 4061 15974 4077 16038
rect 4141 15974 4157 16038
rect 4221 15974 4237 16038
rect 4301 15974 4317 16038
rect 4381 15974 4397 16038
rect 4461 15974 4477 16038
rect 4541 15974 4557 16038
rect 4621 15974 4637 16038
rect 4701 15974 4717 16038
rect 4781 15974 4797 16038
rect 4861 15974 14666 16038
rect 334 15957 14666 15974
rect 381 15893 397 15957
rect 461 15893 477 15957
rect 541 15893 557 15957
rect 621 15893 637 15957
rect 701 15893 717 15957
rect 781 15893 797 15957
rect 861 15893 877 15957
rect 941 15893 957 15957
rect 1021 15893 1037 15957
rect 1101 15893 1117 15957
rect 1181 15893 1197 15957
rect 1261 15893 1277 15957
rect 1341 15893 1357 15957
rect 1421 15893 1437 15957
rect 1501 15893 1517 15957
rect 1581 15893 1597 15957
rect 1661 15893 1677 15957
rect 1741 15893 1757 15957
rect 1821 15893 1837 15957
rect 1901 15893 1917 15957
rect 1981 15893 1997 15957
rect 2061 15893 2077 15957
rect 2141 15893 2157 15957
rect 2221 15893 2237 15957
rect 2301 15893 2317 15957
rect 2381 15893 2397 15957
rect 2461 15893 2477 15957
rect 2541 15893 2557 15957
rect 2621 15893 2637 15957
rect 2701 15893 2717 15957
rect 2781 15893 2797 15957
rect 2861 15893 2877 15957
rect 2941 15893 2957 15957
rect 3021 15893 3037 15957
rect 3101 15893 3117 15957
rect 3181 15893 3197 15957
rect 3261 15893 3277 15957
rect 3341 15893 3357 15957
rect 3421 15893 3437 15957
rect 3501 15893 3517 15957
rect 3581 15893 3597 15957
rect 3661 15893 3677 15957
rect 3741 15893 3757 15957
rect 3821 15893 3837 15957
rect 3901 15893 3917 15957
rect 3981 15893 3997 15957
rect 4061 15893 4077 15957
rect 4141 15893 4157 15957
rect 4221 15893 4237 15957
rect 4301 15893 4317 15957
rect 4381 15893 4397 15957
rect 4461 15893 4477 15957
rect 4541 15893 4557 15957
rect 4621 15893 4637 15957
rect 4701 15893 4717 15957
rect 4781 15893 4797 15957
rect 4861 15893 14666 15957
rect 334 15876 14666 15893
rect 381 15812 397 15876
rect 461 15812 477 15876
rect 541 15812 557 15876
rect 621 15812 637 15876
rect 701 15812 717 15876
rect 781 15812 797 15876
rect 861 15812 877 15876
rect 941 15812 957 15876
rect 1021 15812 1037 15876
rect 1101 15812 1117 15876
rect 1181 15812 1197 15876
rect 1261 15812 1277 15876
rect 1341 15812 1357 15876
rect 1421 15812 1437 15876
rect 1501 15812 1517 15876
rect 1581 15812 1597 15876
rect 1661 15812 1677 15876
rect 1741 15812 1757 15876
rect 1821 15812 1837 15876
rect 1901 15812 1917 15876
rect 1981 15812 1997 15876
rect 2061 15812 2077 15876
rect 2141 15812 2157 15876
rect 2221 15812 2237 15876
rect 2301 15812 2317 15876
rect 2381 15812 2397 15876
rect 2461 15812 2477 15876
rect 2541 15812 2557 15876
rect 2621 15812 2637 15876
rect 2701 15812 2717 15876
rect 2781 15812 2797 15876
rect 2861 15812 2877 15876
rect 2941 15812 2957 15876
rect 3021 15812 3037 15876
rect 3101 15812 3117 15876
rect 3181 15812 3197 15876
rect 3261 15812 3277 15876
rect 3341 15812 3357 15876
rect 3421 15812 3437 15876
rect 3501 15812 3517 15876
rect 3581 15812 3597 15876
rect 3661 15812 3677 15876
rect 3741 15812 3757 15876
rect 3821 15812 3837 15876
rect 3901 15812 3917 15876
rect 3981 15812 3997 15876
rect 4061 15812 4077 15876
rect 4141 15812 4157 15876
rect 4221 15812 4237 15876
rect 4301 15812 4317 15876
rect 4381 15812 4397 15876
rect 4461 15812 4477 15876
rect 4541 15812 4557 15876
rect 4621 15812 4637 15876
rect 4701 15812 4717 15876
rect 4781 15812 4797 15876
rect 4861 15812 14666 15876
rect 334 15795 14666 15812
rect 381 15731 397 15795
rect 461 15731 477 15795
rect 541 15731 557 15795
rect 621 15731 637 15795
rect 701 15731 717 15795
rect 781 15731 797 15795
rect 861 15731 877 15795
rect 941 15731 957 15795
rect 1021 15731 1037 15795
rect 1101 15731 1117 15795
rect 1181 15731 1197 15795
rect 1261 15731 1277 15795
rect 1341 15731 1357 15795
rect 1421 15731 1437 15795
rect 1501 15731 1517 15795
rect 1581 15731 1597 15795
rect 1661 15731 1677 15795
rect 1741 15731 1757 15795
rect 1821 15731 1837 15795
rect 1901 15731 1917 15795
rect 1981 15731 1997 15795
rect 2061 15731 2077 15795
rect 2141 15731 2157 15795
rect 2221 15731 2237 15795
rect 2301 15731 2317 15795
rect 2381 15731 2397 15795
rect 2461 15731 2477 15795
rect 2541 15731 2557 15795
rect 2621 15731 2637 15795
rect 2701 15731 2717 15795
rect 2781 15731 2797 15795
rect 2861 15731 2877 15795
rect 2941 15731 2957 15795
rect 3021 15731 3037 15795
rect 3101 15731 3117 15795
rect 3181 15731 3197 15795
rect 3261 15731 3277 15795
rect 3341 15731 3357 15795
rect 3421 15731 3437 15795
rect 3501 15731 3517 15795
rect 3581 15731 3597 15795
rect 3661 15731 3677 15795
rect 3741 15731 3757 15795
rect 3821 15731 3837 15795
rect 3901 15731 3917 15795
rect 3981 15731 3997 15795
rect 4061 15731 4077 15795
rect 4141 15731 4157 15795
rect 4221 15731 4237 15795
rect 4301 15731 4317 15795
rect 4381 15731 4397 15795
rect 4461 15731 4477 15795
rect 4541 15731 4557 15795
rect 4621 15731 4637 15795
rect 4701 15731 4717 15795
rect 4781 15731 4797 15795
rect 4861 15731 14666 15795
rect 334 15714 14666 15731
rect 381 15650 397 15714
rect 461 15650 477 15714
rect 541 15650 557 15714
rect 621 15650 637 15714
rect 701 15650 717 15714
rect 781 15650 797 15714
rect 861 15650 877 15714
rect 941 15650 957 15714
rect 1021 15650 1037 15714
rect 1101 15650 1117 15714
rect 1181 15650 1197 15714
rect 1261 15650 1277 15714
rect 1341 15650 1357 15714
rect 1421 15650 1437 15714
rect 1501 15650 1517 15714
rect 1581 15650 1597 15714
rect 1661 15650 1677 15714
rect 1741 15650 1757 15714
rect 1821 15650 1837 15714
rect 1901 15650 1917 15714
rect 1981 15650 1997 15714
rect 2061 15650 2077 15714
rect 2141 15650 2157 15714
rect 2221 15650 2237 15714
rect 2301 15650 2317 15714
rect 2381 15650 2397 15714
rect 2461 15650 2477 15714
rect 2541 15650 2557 15714
rect 2621 15650 2637 15714
rect 2701 15650 2717 15714
rect 2781 15650 2797 15714
rect 2861 15650 2877 15714
rect 2941 15650 2957 15714
rect 3021 15650 3037 15714
rect 3101 15650 3117 15714
rect 3181 15650 3197 15714
rect 3261 15650 3277 15714
rect 3341 15650 3357 15714
rect 3421 15650 3437 15714
rect 3501 15650 3517 15714
rect 3581 15650 3597 15714
rect 3661 15650 3677 15714
rect 3741 15650 3757 15714
rect 3821 15650 3837 15714
rect 3901 15650 3917 15714
rect 3981 15650 3997 15714
rect 4061 15650 4077 15714
rect 4141 15650 4157 15714
rect 4221 15650 4237 15714
rect 4301 15650 4317 15714
rect 4381 15650 4397 15714
rect 4461 15650 4477 15714
rect 4541 15650 4557 15714
rect 4621 15650 4637 15714
rect 4701 15650 4717 15714
rect 4781 15650 4797 15714
rect 4861 15650 14666 15714
rect 334 15633 14666 15650
rect 381 15569 397 15633
rect 461 15569 477 15633
rect 541 15569 557 15633
rect 621 15569 637 15633
rect 701 15569 717 15633
rect 781 15569 797 15633
rect 861 15569 877 15633
rect 941 15569 957 15633
rect 1021 15569 1037 15633
rect 1101 15569 1117 15633
rect 1181 15569 1197 15633
rect 1261 15569 1277 15633
rect 1341 15569 1357 15633
rect 1421 15569 1437 15633
rect 1501 15569 1517 15633
rect 1581 15569 1597 15633
rect 1661 15569 1677 15633
rect 1741 15569 1757 15633
rect 1821 15569 1837 15633
rect 1901 15569 1917 15633
rect 1981 15569 1997 15633
rect 2061 15569 2077 15633
rect 2141 15569 2157 15633
rect 2221 15569 2237 15633
rect 2301 15569 2317 15633
rect 2381 15569 2397 15633
rect 2461 15569 2477 15633
rect 2541 15569 2557 15633
rect 2621 15569 2637 15633
rect 2701 15569 2717 15633
rect 2781 15569 2797 15633
rect 2861 15569 2877 15633
rect 2941 15569 2957 15633
rect 3021 15569 3037 15633
rect 3101 15569 3117 15633
rect 3181 15569 3197 15633
rect 3261 15569 3277 15633
rect 3341 15569 3357 15633
rect 3421 15569 3437 15633
rect 3501 15569 3517 15633
rect 3581 15569 3597 15633
rect 3661 15569 3677 15633
rect 3741 15569 3757 15633
rect 3821 15569 3837 15633
rect 3901 15569 3917 15633
rect 3981 15569 3997 15633
rect 4061 15569 4077 15633
rect 4141 15569 4157 15633
rect 4221 15569 4237 15633
rect 4301 15569 4317 15633
rect 4381 15569 4397 15633
rect 4461 15569 4477 15633
rect 4541 15569 4557 15633
rect 4621 15569 4637 15633
rect 4701 15569 4717 15633
rect 4781 15569 4797 15633
rect 4861 15569 14666 15633
rect 334 15552 14666 15569
rect 381 15488 397 15552
rect 461 15488 477 15552
rect 541 15488 557 15552
rect 621 15488 637 15552
rect 701 15488 717 15552
rect 781 15488 797 15552
rect 861 15488 877 15552
rect 941 15488 957 15552
rect 1021 15488 1037 15552
rect 1101 15488 1117 15552
rect 1181 15488 1197 15552
rect 1261 15488 1277 15552
rect 1341 15488 1357 15552
rect 1421 15488 1437 15552
rect 1501 15488 1517 15552
rect 1581 15488 1597 15552
rect 1661 15488 1677 15552
rect 1741 15488 1757 15552
rect 1821 15488 1837 15552
rect 1901 15488 1917 15552
rect 1981 15488 1997 15552
rect 2061 15488 2077 15552
rect 2141 15488 2157 15552
rect 2221 15488 2237 15552
rect 2301 15488 2317 15552
rect 2381 15488 2397 15552
rect 2461 15488 2477 15552
rect 2541 15488 2557 15552
rect 2621 15488 2637 15552
rect 2701 15488 2717 15552
rect 2781 15488 2797 15552
rect 2861 15488 2877 15552
rect 2941 15488 2957 15552
rect 3021 15488 3037 15552
rect 3101 15488 3117 15552
rect 3181 15488 3197 15552
rect 3261 15488 3277 15552
rect 3341 15488 3357 15552
rect 3421 15488 3437 15552
rect 3501 15488 3517 15552
rect 3581 15488 3597 15552
rect 3661 15488 3677 15552
rect 3741 15488 3757 15552
rect 3821 15488 3837 15552
rect 3901 15488 3917 15552
rect 3981 15488 3997 15552
rect 4061 15488 4077 15552
rect 4141 15488 4157 15552
rect 4221 15488 4237 15552
rect 4301 15488 4317 15552
rect 4381 15488 4397 15552
rect 4461 15488 4477 15552
rect 4541 15488 4557 15552
rect 4621 15488 4637 15552
rect 4701 15488 4717 15552
rect 4781 15488 4797 15552
rect 4861 15488 14666 15552
rect 334 15471 14666 15488
rect 381 15407 397 15471
rect 461 15407 477 15471
rect 541 15407 557 15471
rect 621 15407 637 15471
rect 701 15407 717 15471
rect 781 15407 797 15471
rect 861 15407 877 15471
rect 941 15407 957 15471
rect 1021 15407 1037 15471
rect 1101 15407 1117 15471
rect 1181 15407 1197 15471
rect 1261 15407 1277 15471
rect 1341 15407 1357 15471
rect 1421 15407 1437 15471
rect 1501 15407 1517 15471
rect 1581 15407 1597 15471
rect 1661 15407 1677 15471
rect 1741 15407 1757 15471
rect 1821 15407 1837 15471
rect 1901 15407 1917 15471
rect 1981 15407 1997 15471
rect 2061 15407 2077 15471
rect 2141 15407 2157 15471
rect 2221 15407 2237 15471
rect 2301 15407 2317 15471
rect 2381 15407 2397 15471
rect 2461 15407 2477 15471
rect 2541 15407 2557 15471
rect 2621 15407 2637 15471
rect 2701 15407 2717 15471
rect 2781 15407 2797 15471
rect 2861 15407 2877 15471
rect 2941 15407 2957 15471
rect 3021 15407 3037 15471
rect 3101 15407 3117 15471
rect 3181 15407 3197 15471
rect 3261 15407 3277 15471
rect 3341 15407 3357 15471
rect 3421 15407 3437 15471
rect 3501 15407 3517 15471
rect 3581 15407 3597 15471
rect 3661 15407 3677 15471
rect 3741 15407 3757 15471
rect 3821 15407 3837 15471
rect 3901 15407 3917 15471
rect 3981 15407 3997 15471
rect 4061 15407 4077 15471
rect 4141 15407 4157 15471
rect 4221 15407 4237 15471
rect 4301 15407 4317 15471
rect 4381 15407 4397 15471
rect 4461 15407 4477 15471
rect 4541 15407 4557 15471
rect 4621 15407 4637 15471
rect 4701 15407 4717 15471
rect 4781 15407 4797 15471
rect 4861 15407 14666 15471
rect 334 15390 14666 15407
rect 381 15326 397 15390
rect 461 15326 477 15390
rect 541 15326 557 15390
rect 621 15326 637 15390
rect 701 15326 717 15390
rect 781 15326 797 15390
rect 861 15326 877 15390
rect 941 15326 957 15390
rect 1021 15326 1037 15390
rect 1101 15326 1117 15390
rect 1181 15326 1197 15390
rect 1261 15326 1277 15390
rect 1341 15326 1357 15390
rect 1421 15326 1437 15390
rect 1501 15326 1517 15390
rect 1581 15326 1597 15390
rect 1661 15326 1677 15390
rect 1741 15326 1757 15390
rect 1821 15326 1837 15390
rect 1901 15326 1917 15390
rect 1981 15326 1997 15390
rect 2061 15326 2077 15390
rect 2141 15326 2157 15390
rect 2221 15326 2237 15390
rect 2301 15326 2317 15390
rect 2381 15326 2397 15390
rect 2461 15326 2477 15390
rect 2541 15326 2557 15390
rect 2621 15326 2637 15390
rect 2701 15326 2717 15390
rect 2781 15326 2797 15390
rect 2861 15326 2877 15390
rect 2941 15326 2957 15390
rect 3021 15326 3037 15390
rect 3101 15326 3117 15390
rect 3181 15326 3197 15390
rect 3261 15326 3277 15390
rect 3341 15326 3357 15390
rect 3421 15326 3437 15390
rect 3501 15326 3517 15390
rect 3581 15326 3597 15390
rect 3661 15326 3677 15390
rect 3741 15326 3757 15390
rect 3821 15326 3837 15390
rect 3901 15326 3917 15390
rect 3981 15326 3997 15390
rect 4061 15326 4077 15390
rect 4141 15326 4157 15390
rect 4221 15326 4237 15390
rect 4301 15326 4317 15390
rect 4381 15326 4397 15390
rect 4461 15326 4477 15390
rect 4541 15326 4557 15390
rect 4621 15326 4637 15390
rect 4701 15326 4717 15390
rect 4781 15326 4797 15390
rect 4861 15326 14666 15390
rect 334 15309 14666 15326
rect 381 15245 397 15309
rect 461 15245 477 15309
rect 541 15245 557 15309
rect 621 15245 637 15309
rect 701 15245 717 15309
rect 781 15245 797 15309
rect 861 15245 877 15309
rect 941 15245 957 15309
rect 1021 15245 1037 15309
rect 1101 15245 1117 15309
rect 1181 15245 1197 15309
rect 1261 15245 1277 15309
rect 1341 15245 1357 15309
rect 1421 15245 1437 15309
rect 1501 15245 1517 15309
rect 1581 15245 1597 15309
rect 1661 15245 1677 15309
rect 1741 15245 1757 15309
rect 1821 15245 1837 15309
rect 1901 15245 1917 15309
rect 1981 15245 1997 15309
rect 2061 15245 2077 15309
rect 2141 15245 2157 15309
rect 2221 15245 2237 15309
rect 2301 15245 2317 15309
rect 2381 15245 2397 15309
rect 2461 15245 2477 15309
rect 2541 15245 2557 15309
rect 2621 15245 2637 15309
rect 2701 15245 2717 15309
rect 2781 15245 2797 15309
rect 2861 15245 2877 15309
rect 2941 15245 2957 15309
rect 3021 15245 3037 15309
rect 3101 15245 3117 15309
rect 3181 15245 3197 15309
rect 3261 15245 3277 15309
rect 3341 15245 3357 15309
rect 3421 15245 3437 15309
rect 3501 15245 3517 15309
rect 3581 15245 3597 15309
rect 3661 15245 3677 15309
rect 3741 15245 3757 15309
rect 3821 15245 3837 15309
rect 3901 15245 3917 15309
rect 3981 15245 3997 15309
rect 4061 15245 4077 15309
rect 4141 15245 4157 15309
rect 4221 15245 4237 15309
rect 4301 15245 4317 15309
rect 4381 15245 4397 15309
rect 4461 15245 4477 15309
rect 4541 15245 4557 15309
rect 4621 15245 4637 15309
rect 4701 15245 4717 15309
rect 4781 15245 4797 15309
rect 4861 15245 14666 15309
rect 334 15228 14666 15245
rect 381 15164 397 15228
rect 461 15164 477 15228
rect 541 15164 557 15228
rect 621 15164 637 15228
rect 701 15164 717 15228
rect 781 15164 797 15228
rect 861 15164 877 15228
rect 941 15164 957 15228
rect 1021 15164 1037 15228
rect 1101 15164 1117 15228
rect 1181 15164 1197 15228
rect 1261 15164 1277 15228
rect 1341 15164 1357 15228
rect 1421 15164 1437 15228
rect 1501 15164 1517 15228
rect 1581 15164 1597 15228
rect 1661 15164 1677 15228
rect 1741 15164 1757 15228
rect 1821 15164 1837 15228
rect 1901 15164 1917 15228
rect 1981 15164 1997 15228
rect 2061 15164 2077 15228
rect 2141 15164 2157 15228
rect 2221 15164 2237 15228
rect 2301 15164 2317 15228
rect 2381 15164 2397 15228
rect 2461 15164 2477 15228
rect 2541 15164 2557 15228
rect 2621 15164 2637 15228
rect 2701 15164 2717 15228
rect 2781 15164 2797 15228
rect 2861 15164 2877 15228
rect 2941 15164 2957 15228
rect 3021 15164 3037 15228
rect 3101 15164 3117 15228
rect 3181 15164 3197 15228
rect 3261 15164 3277 15228
rect 3341 15164 3357 15228
rect 3421 15164 3437 15228
rect 3501 15164 3517 15228
rect 3581 15164 3597 15228
rect 3661 15164 3677 15228
rect 3741 15164 3757 15228
rect 3821 15164 3837 15228
rect 3901 15164 3917 15228
rect 3981 15164 3997 15228
rect 4061 15164 4077 15228
rect 4141 15164 4157 15228
rect 4221 15164 4237 15228
rect 4301 15164 4317 15228
rect 4381 15164 4397 15228
rect 4461 15164 4477 15228
rect 4541 15164 4557 15228
rect 4621 15164 4637 15228
rect 4701 15164 4717 15228
rect 4781 15164 4797 15228
rect 4861 15164 14666 15228
rect 334 15147 14666 15164
rect 381 15083 397 15147
rect 461 15083 477 15147
rect 541 15083 557 15147
rect 621 15083 637 15147
rect 701 15083 717 15147
rect 781 15083 797 15147
rect 861 15083 877 15147
rect 941 15083 957 15147
rect 1021 15083 1037 15147
rect 1101 15083 1117 15147
rect 1181 15083 1197 15147
rect 1261 15083 1277 15147
rect 1341 15083 1357 15147
rect 1421 15083 1437 15147
rect 1501 15083 1517 15147
rect 1581 15083 1597 15147
rect 1661 15083 1677 15147
rect 1741 15083 1757 15147
rect 1821 15083 1837 15147
rect 1901 15083 1917 15147
rect 1981 15083 1997 15147
rect 2061 15083 2077 15147
rect 2141 15083 2157 15147
rect 2221 15083 2237 15147
rect 2301 15083 2317 15147
rect 2381 15083 2397 15147
rect 2461 15083 2477 15147
rect 2541 15083 2557 15147
rect 2621 15083 2637 15147
rect 2701 15083 2717 15147
rect 2781 15083 2797 15147
rect 2861 15083 2877 15147
rect 2941 15083 2957 15147
rect 3021 15083 3037 15147
rect 3101 15083 3117 15147
rect 3181 15083 3197 15147
rect 3261 15083 3277 15147
rect 3341 15083 3357 15147
rect 3421 15083 3437 15147
rect 3501 15083 3517 15147
rect 3581 15083 3597 15147
rect 3661 15083 3677 15147
rect 3741 15083 3757 15147
rect 3821 15083 3837 15147
rect 3901 15083 3917 15147
rect 3981 15083 3997 15147
rect 4061 15083 4077 15147
rect 4141 15083 4157 15147
rect 4221 15083 4237 15147
rect 4301 15083 4317 15147
rect 4381 15083 4397 15147
rect 4461 15083 4477 15147
rect 4541 15083 4557 15147
rect 4621 15083 4637 15147
rect 4701 15083 4717 15147
rect 4781 15083 4797 15147
rect 4861 15083 14666 15147
rect 334 15066 14666 15083
rect 381 15002 397 15066
rect 461 15002 477 15066
rect 541 15002 557 15066
rect 621 15002 637 15066
rect 701 15002 717 15066
rect 781 15002 797 15066
rect 861 15002 877 15066
rect 941 15002 957 15066
rect 1021 15002 1037 15066
rect 1101 15002 1117 15066
rect 1181 15002 1197 15066
rect 1261 15002 1277 15066
rect 1341 15002 1357 15066
rect 1421 15002 1437 15066
rect 1501 15002 1517 15066
rect 1581 15002 1597 15066
rect 1661 15002 1677 15066
rect 1741 15002 1757 15066
rect 1821 15002 1837 15066
rect 1901 15002 1917 15066
rect 1981 15002 1997 15066
rect 2061 15002 2077 15066
rect 2141 15002 2157 15066
rect 2221 15002 2237 15066
rect 2301 15002 2317 15066
rect 2381 15002 2397 15066
rect 2461 15002 2477 15066
rect 2541 15002 2557 15066
rect 2621 15002 2637 15066
rect 2701 15002 2717 15066
rect 2781 15002 2797 15066
rect 2861 15002 2877 15066
rect 2941 15002 2957 15066
rect 3021 15002 3037 15066
rect 3101 15002 3117 15066
rect 3181 15002 3197 15066
rect 3261 15002 3277 15066
rect 3341 15002 3357 15066
rect 3421 15002 3437 15066
rect 3501 15002 3517 15066
rect 3581 15002 3597 15066
rect 3661 15002 3677 15066
rect 3741 15002 3757 15066
rect 3821 15002 3837 15066
rect 3901 15002 3917 15066
rect 3981 15002 3997 15066
rect 4061 15002 4077 15066
rect 4141 15002 4157 15066
rect 4221 15002 4237 15066
rect 4301 15002 4317 15066
rect 4381 15002 4397 15066
rect 4461 15002 4477 15066
rect 4541 15002 4557 15066
rect 4621 15002 4637 15066
rect 4701 15002 4717 15066
rect 4781 15002 4797 15066
rect 4861 15002 14666 15066
rect 334 14985 14666 15002
rect 381 14921 397 14985
rect 461 14921 477 14985
rect 541 14921 557 14985
rect 621 14921 637 14985
rect 701 14921 717 14985
rect 781 14921 797 14985
rect 861 14921 877 14985
rect 941 14921 957 14985
rect 1021 14921 1037 14985
rect 1101 14921 1117 14985
rect 1181 14921 1197 14985
rect 1261 14921 1277 14985
rect 1341 14921 1357 14985
rect 1421 14921 1437 14985
rect 1501 14921 1517 14985
rect 1581 14921 1597 14985
rect 1661 14921 1677 14985
rect 1741 14921 1757 14985
rect 1821 14921 1837 14985
rect 1901 14921 1917 14985
rect 1981 14921 1997 14985
rect 2061 14921 2077 14985
rect 2141 14921 2157 14985
rect 2221 14921 2237 14985
rect 2301 14921 2317 14985
rect 2381 14921 2397 14985
rect 2461 14921 2477 14985
rect 2541 14921 2557 14985
rect 2621 14921 2637 14985
rect 2701 14921 2717 14985
rect 2781 14921 2797 14985
rect 2861 14921 2877 14985
rect 2941 14921 2957 14985
rect 3021 14921 3037 14985
rect 3101 14921 3117 14985
rect 3181 14921 3197 14985
rect 3261 14921 3277 14985
rect 3341 14921 3357 14985
rect 3421 14921 3437 14985
rect 3501 14921 3517 14985
rect 3581 14921 3597 14985
rect 3661 14921 3677 14985
rect 3741 14921 3757 14985
rect 3821 14921 3837 14985
rect 3901 14921 3917 14985
rect 3981 14921 3997 14985
rect 4061 14921 4077 14985
rect 4141 14921 4157 14985
rect 4221 14921 4237 14985
rect 4301 14921 4317 14985
rect 4381 14921 4397 14985
rect 4461 14921 4477 14985
rect 4541 14921 4557 14985
rect 4621 14921 4637 14985
rect 4701 14921 4717 14985
rect 4781 14921 4797 14985
rect 4861 14921 14666 14985
rect 334 14904 14666 14921
rect 381 14840 397 14904
rect 461 14840 477 14904
rect 541 14840 557 14904
rect 621 14840 637 14904
rect 701 14840 717 14904
rect 781 14840 797 14904
rect 861 14840 877 14904
rect 941 14840 957 14904
rect 1021 14840 1037 14904
rect 1101 14840 1117 14904
rect 1181 14840 1197 14904
rect 1261 14840 1277 14904
rect 1341 14840 1357 14904
rect 1421 14840 1437 14904
rect 1501 14840 1517 14904
rect 1581 14840 1597 14904
rect 1661 14840 1677 14904
rect 1741 14840 1757 14904
rect 1821 14840 1837 14904
rect 1901 14840 1917 14904
rect 1981 14840 1997 14904
rect 2061 14840 2077 14904
rect 2141 14840 2157 14904
rect 2221 14840 2237 14904
rect 2301 14840 2317 14904
rect 2381 14840 2397 14904
rect 2461 14840 2477 14904
rect 2541 14840 2557 14904
rect 2621 14840 2637 14904
rect 2701 14840 2717 14904
rect 2781 14840 2797 14904
rect 2861 14840 2877 14904
rect 2941 14840 2957 14904
rect 3021 14840 3037 14904
rect 3101 14840 3117 14904
rect 3181 14840 3197 14904
rect 3261 14840 3277 14904
rect 3341 14840 3357 14904
rect 3421 14840 3437 14904
rect 3501 14840 3517 14904
rect 3581 14840 3597 14904
rect 3661 14840 3677 14904
rect 3741 14840 3757 14904
rect 3821 14840 3837 14904
rect 3901 14840 3917 14904
rect 3981 14840 3997 14904
rect 4061 14840 4077 14904
rect 4141 14840 4157 14904
rect 4221 14840 4237 14904
rect 4301 14840 4317 14904
rect 4381 14840 4397 14904
rect 4461 14840 4477 14904
rect 4541 14840 4557 14904
rect 4621 14840 4637 14904
rect 4701 14840 4717 14904
rect 4781 14840 4797 14904
rect 4861 14840 14666 14904
rect 334 14823 14666 14840
rect 381 14759 397 14823
rect 461 14759 477 14823
rect 541 14759 557 14823
rect 621 14759 637 14823
rect 701 14759 717 14823
rect 781 14759 797 14823
rect 861 14759 877 14823
rect 941 14759 957 14823
rect 1021 14759 1037 14823
rect 1101 14759 1117 14823
rect 1181 14759 1197 14823
rect 1261 14759 1277 14823
rect 1341 14759 1357 14823
rect 1421 14759 1437 14823
rect 1501 14759 1517 14823
rect 1581 14759 1597 14823
rect 1661 14759 1677 14823
rect 1741 14759 1757 14823
rect 1821 14759 1837 14823
rect 1901 14759 1917 14823
rect 1981 14759 1997 14823
rect 2061 14759 2077 14823
rect 2141 14759 2157 14823
rect 2221 14759 2237 14823
rect 2301 14759 2317 14823
rect 2381 14759 2397 14823
rect 2461 14759 2477 14823
rect 2541 14759 2557 14823
rect 2621 14759 2637 14823
rect 2701 14759 2717 14823
rect 2781 14759 2797 14823
rect 2861 14759 2877 14823
rect 2941 14759 2957 14823
rect 3021 14759 3037 14823
rect 3101 14759 3117 14823
rect 3181 14759 3197 14823
rect 3261 14759 3277 14823
rect 3341 14759 3357 14823
rect 3421 14759 3437 14823
rect 3501 14759 3517 14823
rect 3581 14759 3597 14823
rect 3661 14759 3677 14823
rect 3741 14759 3757 14823
rect 3821 14759 3837 14823
rect 3901 14759 3917 14823
rect 3981 14759 3997 14823
rect 4061 14759 4077 14823
rect 4141 14759 4157 14823
rect 4221 14759 4237 14823
rect 4301 14759 4317 14823
rect 4381 14759 4397 14823
rect 4461 14759 4477 14823
rect 4541 14759 4557 14823
rect 4621 14759 4637 14823
rect 4701 14759 4717 14823
rect 4781 14759 4797 14823
rect 4861 14759 14666 14823
rect 334 14742 14666 14759
rect 381 14678 397 14742
rect 461 14678 477 14742
rect 541 14678 557 14742
rect 621 14678 637 14742
rect 701 14678 717 14742
rect 781 14678 797 14742
rect 861 14678 877 14742
rect 941 14678 957 14742
rect 1021 14678 1037 14742
rect 1101 14678 1117 14742
rect 1181 14678 1197 14742
rect 1261 14678 1277 14742
rect 1341 14678 1357 14742
rect 1421 14678 1437 14742
rect 1501 14678 1517 14742
rect 1581 14678 1597 14742
rect 1661 14678 1677 14742
rect 1741 14678 1757 14742
rect 1821 14678 1837 14742
rect 1901 14678 1917 14742
rect 1981 14678 1997 14742
rect 2061 14678 2077 14742
rect 2141 14678 2157 14742
rect 2221 14678 2237 14742
rect 2301 14678 2317 14742
rect 2381 14678 2397 14742
rect 2461 14678 2477 14742
rect 2541 14678 2557 14742
rect 2621 14678 2637 14742
rect 2701 14678 2717 14742
rect 2781 14678 2797 14742
rect 2861 14678 2877 14742
rect 2941 14678 2957 14742
rect 3021 14678 3037 14742
rect 3101 14678 3117 14742
rect 3181 14678 3197 14742
rect 3261 14678 3277 14742
rect 3341 14678 3357 14742
rect 3421 14678 3437 14742
rect 3501 14678 3517 14742
rect 3581 14678 3597 14742
rect 3661 14678 3677 14742
rect 3741 14678 3757 14742
rect 3821 14678 3837 14742
rect 3901 14678 3917 14742
rect 3981 14678 3997 14742
rect 4061 14678 4077 14742
rect 4141 14678 4157 14742
rect 4221 14678 4237 14742
rect 4301 14678 4317 14742
rect 4381 14678 4397 14742
rect 4461 14678 4477 14742
rect 4541 14678 4557 14742
rect 4621 14678 4637 14742
rect 4701 14678 4717 14742
rect 4781 14678 4797 14742
rect 4861 14678 14666 14742
rect 334 14661 14666 14678
rect 381 14597 397 14661
rect 461 14597 477 14661
rect 541 14597 557 14661
rect 621 14597 637 14661
rect 701 14597 717 14661
rect 781 14597 797 14661
rect 861 14597 877 14661
rect 941 14597 957 14661
rect 1021 14597 1037 14661
rect 1101 14597 1117 14661
rect 1181 14597 1197 14661
rect 1261 14597 1277 14661
rect 1341 14597 1357 14661
rect 1421 14597 1437 14661
rect 1501 14597 1517 14661
rect 1581 14597 1597 14661
rect 1661 14597 1677 14661
rect 1741 14597 1757 14661
rect 1821 14597 1837 14661
rect 1901 14597 1917 14661
rect 1981 14597 1997 14661
rect 2061 14597 2077 14661
rect 2141 14597 2157 14661
rect 2221 14597 2237 14661
rect 2301 14597 2317 14661
rect 2381 14597 2397 14661
rect 2461 14597 2477 14661
rect 2541 14597 2557 14661
rect 2621 14597 2637 14661
rect 2701 14597 2717 14661
rect 2781 14597 2797 14661
rect 2861 14597 2877 14661
rect 2941 14597 2957 14661
rect 3021 14597 3037 14661
rect 3101 14597 3117 14661
rect 3181 14597 3197 14661
rect 3261 14597 3277 14661
rect 3341 14597 3357 14661
rect 3421 14597 3437 14661
rect 3501 14597 3517 14661
rect 3581 14597 3597 14661
rect 3661 14597 3677 14661
rect 3741 14597 3757 14661
rect 3821 14597 3837 14661
rect 3901 14597 3917 14661
rect 3981 14597 3997 14661
rect 4061 14597 4077 14661
rect 4141 14597 4157 14661
rect 4221 14597 4237 14661
rect 4301 14597 4317 14661
rect 4381 14597 4397 14661
rect 4461 14597 4477 14661
rect 4541 14597 4557 14661
rect 4621 14597 4637 14661
rect 4701 14597 4717 14661
rect 4781 14597 4797 14661
rect 4861 14597 14666 14661
rect 334 14579 14666 14597
rect 381 14515 397 14579
rect 461 14515 477 14579
rect 541 14515 557 14579
rect 621 14515 637 14579
rect 701 14515 717 14579
rect 781 14515 797 14579
rect 861 14515 877 14579
rect 941 14515 957 14579
rect 1021 14515 1037 14579
rect 1101 14515 1117 14579
rect 1181 14515 1197 14579
rect 1261 14515 1277 14579
rect 1341 14515 1357 14579
rect 1421 14515 1437 14579
rect 1501 14515 1517 14579
rect 1581 14515 1597 14579
rect 1661 14515 1677 14579
rect 1741 14515 1757 14579
rect 1821 14515 1837 14579
rect 1901 14515 1917 14579
rect 1981 14515 1997 14579
rect 2061 14515 2077 14579
rect 2141 14515 2157 14579
rect 2221 14515 2237 14579
rect 2301 14515 2317 14579
rect 2381 14515 2397 14579
rect 2461 14515 2477 14579
rect 2541 14515 2557 14579
rect 2621 14515 2637 14579
rect 2701 14515 2717 14579
rect 2781 14515 2797 14579
rect 2861 14515 2877 14579
rect 2941 14515 2957 14579
rect 3021 14515 3037 14579
rect 3101 14515 3117 14579
rect 3181 14515 3197 14579
rect 3261 14515 3277 14579
rect 3341 14515 3357 14579
rect 3421 14515 3437 14579
rect 3501 14515 3517 14579
rect 3581 14515 3597 14579
rect 3661 14515 3677 14579
rect 3741 14515 3757 14579
rect 3821 14515 3837 14579
rect 3901 14515 3917 14579
rect 3981 14515 3997 14579
rect 4061 14515 4077 14579
rect 4141 14515 4157 14579
rect 4221 14515 4237 14579
rect 4301 14515 4317 14579
rect 4381 14515 4397 14579
rect 4461 14515 4477 14579
rect 4541 14515 4557 14579
rect 4621 14515 4637 14579
rect 4701 14515 4717 14579
rect 4781 14515 4797 14579
rect 4861 14515 14666 14579
rect 334 14497 14666 14515
rect 381 14433 397 14497
rect 461 14433 477 14497
rect 541 14433 557 14497
rect 621 14433 637 14497
rect 701 14433 717 14497
rect 781 14433 797 14497
rect 861 14433 877 14497
rect 941 14433 957 14497
rect 1021 14433 1037 14497
rect 1101 14433 1117 14497
rect 1181 14433 1197 14497
rect 1261 14433 1277 14497
rect 1341 14433 1357 14497
rect 1421 14433 1437 14497
rect 1501 14433 1517 14497
rect 1581 14433 1597 14497
rect 1661 14433 1677 14497
rect 1741 14433 1757 14497
rect 1821 14433 1837 14497
rect 1901 14433 1917 14497
rect 1981 14433 1997 14497
rect 2061 14433 2077 14497
rect 2141 14433 2157 14497
rect 2221 14433 2237 14497
rect 2301 14433 2317 14497
rect 2381 14433 2397 14497
rect 2461 14433 2477 14497
rect 2541 14433 2557 14497
rect 2621 14433 2637 14497
rect 2701 14433 2717 14497
rect 2781 14433 2797 14497
rect 2861 14433 2877 14497
rect 2941 14433 2957 14497
rect 3021 14433 3037 14497
rect 3101 14433 3117 14497
rect 3181 14433 3197 14497
rect 3261 14433 3277 14497
rect 3341 14433 3357 14497
rect 3421 14433 3437 14497
rect 3501 14433 3517 14497
rect 3581 14433 3597 14497
rect 3661 14433 3677 14497
rect 3741 14433 3757 14497
rect 3821 14433 3837 14497
rect 3901 14433 3917 14497
rect 3981 14433 3997 14497
rect 4061 14433 4077 14497
rect 4141 14433 4157 14497
rect 4221 14433 4237 14497
rect 4301 14433 4317 14497
rect 4381 14433 4397 14497
rect 4461 14433 4477 14497
rect 4541 14433 4557 14497
rect 4621 14433 4637 14497
rect 4701 14433 4717 14497
rect 4781 14433 4797 14497
rect 4861 14433 14666 14497
rect 334 14415 14666 14433
rect 381 14351 397 14415
rect 461 14351 477 14415
rect 541 14351 557 14415
rect 621 14351 637 14415
rect 701 14351 717 14415
rect 781 14351 797 14415
rect 861 14351 877 14415
rect 941 14351 957 14415
rect 1021 14351 1037 14415
rect 1101 14351 1117 14415
rect 1181 14351 1197 14415
rect 1261 14351 1277 14415
rect 1341 14351 1357 14415
rect 1421 14351 1437 14415
rect 1501 14351 1517 14415
rect 1581 14351 1597 14415
rect 1661 14351 1677 14415
rect 1741 14351 1757 14415
rect 1821 14351 1837 14415
rect 1901 14351 1917 14415
rect 1981 14351 1997 14415
rect 2061 14351 2077 14415
rect 2141 14351 2157 14415
rect 2221 14351 2237 14415
rect 2301 14351 2317 14415
rect 2381 14351 2397 14415
rect 2461 14351 2477 14415
rect 2541 14351 2557 14415
rect 2621 14351 2637 14415
rect 2701 14351 2717 14415
rect 2781 14351 2797 14415
rect 2861 14351 2877 14415
rect 2941 14351 2957 14415
rect 3021 14351 3037 14415
rect 3101 14351 3117 14415
rect 3181 14351 3197 14415
rect 3261 14351 3277 14415
rect 3341 14351 3357 14415
rect 3421 14351 3437 14415
rect 3501 14351 3517 14415
rect 3581 14351 3597 14415
rect 3661 14351 3677 14415
rect 3741 14351 3757 14415
rect 3821 14351 3837 14415
rect 3901 14351 3917 14415
rect 3981 14351 3997 14415
rect 4061 14351 4077 14415
rect 4141 14351 4157 14415
rect 4221 14351 4237 14415
rect 4301 14351 4317 14415
rect 4381 14351 4397 14415
rect 4461 14351 4477 14415
rect 4541 14351 4557 14415
rect 4621 14351 4637 14415
rect 4701 14351 4717 14415
rect 4781 14351 4797 14415
rect 4861 14351 14666 14415
rect 334 14333 14666 14351
rect 381 14269 397 14333
rect 461 14269 477 14333
rect 541 14269 557 14333
rect 621 14269 637 14333
rect 701 14269 717 14333
rect 781 14269 797 14333
rect 861 14269 877 14333
rect 941 14269 957 14333
rect 1021 14269 1037 14333
rect 1101 14269 1117 14333
rect 1181 14269 1197 14333
rect 1261 14269 1277 14333
rect 1341 14269 1357 14333
rect 1421 14269 1437 14333
rect 1501 14269 1517 14333
rect 1581 14269 1597 14333
rect 1661 14269 1677 14333
rect 1741 14269 1757 14333
rect 1821 14269 1837 14333
rect 1901 14269 1917 14333
rect 1981 14269 1997 14333
rect 2061 14269 2077 14333
rect 2141 14269 2157 14333
rect 2221 14269 2237 14333
rect 2301 14269 2317 14333
rect 2381 14269 2397 14333
rect 2461 14269 2477 14333
rect 2541 14269 2557 14333
rect 2621 14269 2637 14333
rect 2701 14269 2717 14333
rect 2781 14269 2797 14333
rect 2861 14269 2877 14333
rect 2941 14269 2957 14333
rect 3021 14269 3037 14333
rect 3101 14269 3117 14333
rect 3181 14269 3197 14333
rect 3261 14269 3277 14333
rect 3341 14269 3357 14333
rect 3421 14269 3437 14333
rect 3501 14269 3517 14333
rect 3581 14269 3597 14333
rect 3661 14269 3677 14333
rect 3741 14269 3757 14333
rect 3821 14269 3837 14333
rect 3901 14269 3917 14333
rect 3981 14269 3997 14333
rect 4061 14269 4077 14333
rect 4141 14269 4157 14333
rect 4221 14269 4237 14333
rect 4301 14269 4317 14333
rect 4381 14269 4397 14333
rect 4461 14269 4477 14333
rect 4541 14269 4557 14333
rect 4621 14269 4637 14333
rect 4701 14269 4717 14333
rect 4781 14269 4797 14333
rect 4861 14269 14666 14333
rect 334 14251 14666 14269
rect 381 14187 397 14251
rect 461 14187 477 14251
rect 541 14187 557 14251
rect 621 14187 637 14251
rect 701 14187 717 14251
rect 781 14187 797 14251
rect 861 14187 877 14251
rect 941 14187 957 14251
rect 1021 14187 1037 14251
rect 1101 14187 1117 14251
rect 1181 14187 1197 14251
rect 1261 14187 1277 14251
rect 1341 14187 1357 14251
rect 1421 14187 1437 14251
rect 1501 14187 1517 14251
rect 1581 14187 1597 14251
rect 1661 14187 1677 14251
rect 1741 14187 1757 14251
rect 1821 14187 1837 14251
rect 1901 14187 1917 14251
rect 1981 14187 1997 14251
rect 2061 14187 2077 14251
rect 2141 14187 2157 14251
rect 2221 14187 2237 14251
rect 2301 14187 2317 14251
rect 2381 14187 2397 14251
rect 2461 14187 2477 14251
rect 2541 14187 2557 14251
rect 2621 14187 2637 14251
rect 2701 14187 2717 14251
rect 2781 14187 2797 14251
rect 2861 14187 2877 14251
rect 2941 14187 2957 14251
rect 3021 14187 3037 14251
rect 3101 14187 3117 14251
rect 3181 14187 3197 14251
rect 3261 14187 3277 14251
rect 3341 14187 3357 14251
rect 3421 14187 3437 14251
rect 3501 14187 3517 14251
rect 3581 14187 3597 14251
rect 3661 14187 3677 14251
rect 3741 14187 3757 14251
rect 3821 14187 3837 14251
rect 3901 14187 3917 14251
rect 3981 14187 3997 14251
rect 4061 14187 4077 14251
rect 4141 14187 4157 14251
rect 4221 14187 4237 14251
rect 4301 14187 4317 14251
rect 4381 14187 4397 14251
rect 4461 14187 4477 14251
rect 4541 14187 4557 14251
rect 4621 14187 4637 14251
rect 4701 14187 4717 14251
rect 4781 14187 4797 14251
rect 4861 14187 14666 14251
rect 334 14169 14666 14187
rect 381 14105 397 14169
rect 461 14105 477 14169
rect 541 14105 557 14169
rect 621 14105 637 14169
rect 701 14105 717 14169
rect 781 14105 797 14169
rect 861 14105 877 14169
rect 941 14105 957 14169
rect 1021 14105 1037 14169
rect 1101 14105 1117 14169
rect 1181 14105 1197 14169
rect 1261 14105 1277 14169
rect 1341 14105 1357 14169
rect 1421 14105 1437 14169
rect 1501 14105 1517 14169
rect 1581 14105 1597 14169
rect 1661 14105 1677 14169
rect 1741 14105 1757 14169
rect 1821 14105 1837 14169
rect 1901 14105 1917 14169
rect 1981 14105 1997 14169
rect 2061 14105 2077 14169
rect 2141 14105 2157 14169
rect 2221 14105 2237 14169
rect 2301 14105 2317 14169
rect 2381 14105 2397 14169
rect 2461 14105 2477 14169
rect 2541 14105 2557 14169
rect 2621 14105 2637 14169
rect 2701 14105 2717 14169
rect 2781 14105 2797 14169
rect 2861 14105 2877 14169
rect 2941 14105 2957 14169
rect 3021 14105 3037 14169
rect 3101 14105 3117 14169
rect 3181 14105 3197 14169
rect 3261 14105 3277 14169
rect 3341 14105 3357 14169
rect 3421 14105 3437 14169
rect 3501 14105 3517 14169
rect 3581 14105 3597 14169
rect 3661 14105 3677 14169
rect 3741 14105 3757 14169
rect 3821 14105 3837 14169
rect 3901 14105 3917 14169
rect 3981 14105 3997 14169
rect 4061 14105 4077 14169
rect 4141 14105 4157 14169
rect 4221 14105 4237 14169
rect 4301 14105 4317 14169
rect 4381 14105 4397 14169
rect 4461 14105 4477 14169
rect 4541 14105 4557 14169
rect 4621 14105 4637 14169
rect 4701 14105 4717 14169
rect 4781 14105 4797 14169
rect 4861 14105 14666 14169
rect 334 14087 14666 14105
rect 381 14023 397 14087
rect 461 14023 477 14087
rect 541 14023 557 14087
rect 621 14023 637 14087
rect 701 14023 717 14087
rect 781 14023 797 14087
rect 861 14023 877 14087
rect 941 14023 957 14087
rect 1021 14023 1037 14087
rect 1101 14023 1117 14087
rect 1181 14023 1197 14087
rect 1261 14023 1277 14087
rect 1341 14023 1357 14087
rect 1421 14023 1437 14087
rect 1501 14023 1517 14087
rect 1581 14023 1597 14087
rect 1661 14023 1677 14087
rect 1741 14023 1757 14087
rect 1821 14023 1837 14087
rect 1901 14023 1917 14087
rect 1981 14023 1997 14087
rect 2061 14023 2077 14087
rect 2141 14023 2157 14087
rect 2221 14023 2237 14087
rect 2301 14023 2317 14087
rect 2381 14023 2397 14087
rect 2461 14023 2477 14087
rect 2541 14023 2557 14087
rect 2621 14023 2637 14087
rect 2701 14023 2717 14087
rect 2781 14023 2797 14087
rect 2861 14023 2877 14087
rect 2941 14023 2957 14087
rect 3021 14023 3037 14087
rect 3101 14023 3117 14087
rect 3181 14023 3197 14087
rect 3261 14023 3277 14087
rect 3341 14023 3357 14087
rect 3421 14023 3437 14087
rect 3501 14023 3517 14087
rect 3581 14023 3597 14087
rect 3661 14023 3677 14087
rect 3741 14023 3757 14087
rect 3821 14023 3837 14087
rect 3901 14023 3917 14087
rect 3981 14023 3997 14087
rect 4061 14023 4077 14087
rect 4141 14023 4157 14087
rect 4221 14023 4237 14087
rect 4301 14023 4317 14087
rect 4381 14023 4397 14087
rect 4461 14023 4477 14087
rect 4541 14023 4557 14087
rect 4621 14023 4637 14087
rect 4701 14023 4717 14087
rect 4781 14023 4797 14087
rect 4861 14023 14666 14087
rect 334 14005 14666 14023
rect 381 13941 397 14005
rect 461 13941 477 14005
rect 541 13941 557 14005
rect 621 13941 637 14005
rect 701 13941 717 14005
rect 781 13941 797 14005
rect 861 13941 877 14005
rect 941 13941 957 14005
rect 1021 13941 1037 14005
rect 1101 13941 1117 14005
rect 1181 13941 1197 14005
rect 1261 13941 1277 14005
rect 1341 13941 1357 14005
rect 1421 13941 1437 14005
rect 1501 13941 1517 14005
rect 1581 13941 1597 14005
rect 1661 13941 1677 14005
rect 1741 13941 1757 14005
rect 1821 13941 1837 14005
rect 1901 13941 1917 14005
rect 1981 13941 1997 14005
rect 2061 13941 2077 14005
rect 2141 13941 2157 14005
rect 2221 13941 2237 14005
rect 2301 13941 2317 14005
rect 2381 13941 2397 14005
rect 2461 13941 2477 14005
rect 2541 13941 2557 14005
rect 2621 13941 2637 14005
rect 2701 13941 2717 14005
rect 2781 13941 2797 14005
rect 2861 13941 2877 14005
rect 2941 13941 2957 14005
rect 3021 13941 3037 14005
rect 3101 13941 3117 14005
rect 3181 13941 3197 14005
rect 3261 13941 3277 14005
rect 3341 13941 3357 14005
rect 3421 13941 3437 14005
rect 3501 13941 3517 14005
rect 3581 13941 3597 14005
rect 3661 13941 3677 14005
rect 3741 13941 3757 14005
rect 3821 13941 3837 14005
rect 3901 13941 3917 14005
rect 3981 13941 3997 14005
rect 4061 13941 4077 14005
rect 4141 13941 4157 14005
rect 4221 13941 4237 14005
rect 4301 13941 4317 14005
rect 4381 13941 4397 14005
rect 4461 13941 4477 14005
rect 4541 13941 4557 14005
rect 4621 13941 4637 14005
rect 4701 13941 4717 14005
rect 4781 13941 4797 14005
rect 4861 13941 14666 14005
rect 334 13923 14666 13941
rect 381 13859 397 13923
rect 461 13859 477 13923
rect 541 13859 557 13923
rect 621 13859 637 13923
rect 701 13859 717 13923
rect 781 13859 797 13923
rect 861 13859 877 13923
rect 941 13859 957 13923
rect 1021 13859 1037 13923
rect 1101 13859 1117 13923
rect 1181 13859 1197 13923
rect 1261 13859 1277 13923
rect 1341 13859 1357 13923
rect 1421 13859 1437 13923
rect 1501 13859 1517 13923
rect 1581 13859 1597 13923
rect 1661 13859 1677 13923
rect 1741 13859 1757 13923
rect 1821 13859 1837 13923
rect 1901 13859 1917 13923
rect 1981 13859 1997 13923
rect 2061 13859 2077 13923
rect 2141 13859 2157 13923
rect 2221 13859 2237 13923
rect 2301 13859 2317 13923
rect 2381 13859 2397 13923
rect 2461 13859 2477 13923
rect 2541 13859 2557 13923
rect 2621 13859 2637 13923
rect 2701 13859 2717 13923
rect 2781 13859 2797 13923
rect 2861 13859 2877 13923
rect 2941 13859 2957 13923
rect 3021 13859 3037 13923
rect 3101 13859 3117 13923
rect 3181 13859 3197 13923
rect 3261 13859 3277 13923
rect 3341 13859 3357 13923
rect 3421 13859 3437 13923
rect 3501 13859 3517 13923
rect 3581 13859 3597 13923
rect 3661 13859 3677 13923
rect 3741 13859 3757 13923
rect 3821 13859 3837 13923
rect 3901 13859 3917 13923
rect 3981 13859 3997 13923
rect 4061 13859 4077 13923
rect 4141 13859 4157 13923
rect 4221 13859 4237 13923
rect 4301 13859 4317 13923
rect 4381 13859 4397 13923
rect 4461 13859 4477 13923
rect 4541 13859 4557 13923
rect 4621 13859 4637 13923
rect 4701 13859 4717 13923
rect 4781 13859 4797 13923
rect 4861 13859 14666 13923
rect 334 13841 14666 13859
rect 381 13777 397 13841
rect 461 13777 477 13841
rect 541 13777 557 13841
rect 621 13777 637 13841
rect 701 13777 717 13841
rect 781 13777 797 13841
rect 861 13777 877 13841
rect 941 13777 957 13841
rect 1021 13777 1037 13841
rect 1101 13777 1117 13841
rect 1181 13777 1197 13841
rect 1261 13777 1277 13841
rect 1341 13777 1357 13841
rect 1421 13777 1437 13841
rect 1501 13777 1517 13841
rect 1581 13777 1597 13841
rect 1661 13777 1677 13841
rect 1741 13777 1757 13841
rect 1821 13777 1837 13841
rect 1901 13777 1917 13841
rect 1981 13777 1997 13841
rect 2061 13777 2077 13841
rect 2141 13777 2157 13841
rect 2221 13777 2237 13841
rect 2301 13777 2317 13841
rect 2381 13777 2397 13841
rect 2461 13777 2477 13841
rect 2541 13777 2557 13841
rect 2621 13777 2637 13841
rect 2701 13777 2717 13841
rect 2781 13777 2797 13841
rect 2861 13777 2877 13841
rect 2941 13777 2957 13841
rect 3021 13777 3037 13841
rect 3101 13777 3117 13841
rect 3181 13777 3197 13841
rect 3261 13777 3277 13841
rect 3341 13777 3357 13841
rect 3421 13777 3437 13841
rect 3501 13777 3517 13841
rect 3581 13777 3597 13841
rect 3661 13777 3677 13841
rect 3741 13777 3757 13841
rect 3821 13777 3837 13841
rect 3901 13777 3917 13841
rect 3981 13777 3997 13841
rect 4061 13777 4077 13841
rect 4141 13777 4157 13841
rect 4221 13777 4237 13841
rect 4301 13777 4317 13841
rect 4381 13777 4397 13841
rect 4461 13777 4477 13841
rect 4541 13777 4557 13841
rect 4621 13777 4637 13841
rect 4701 13777 4717 13841
rect 4781 13777 4797 13841
rect 4861 13777 14666 13841
rect 334 13759 14666 13777
rect 381 13695 397 13759
rect 461 13695 477 13759
rect 541 13695 557 13759
rect 621 13695 637 13759
rect 701 13695 717 13759
rect 781 13695 797 13759
rect 861 13695 877 13759
rect 941 13695 957 13759
rect 1021 13695 1037 13759
rect 1101 13695 1117 13759
rect 1181 13695 1197 13759
rect 1261 13695 1277 13759
rect 1341 13695 1357 13759
rect 1421 13695 1437 13759
rect 1501 13695 1517 13759
rect 1581 13695 1597 13759
rect 1661 13695 1677 13759
rect 1741 13695 1757 13759
rect 1821 13695 1837 13759
rect 1901 13695 1917 13759
rect 1981 13695 1997 13759
rect 2061 13695 2077 13759
rect 2141 13695 2157 13759
rect 2221 13695 2237 13759
rect 2301 13695 2317 13759
rect 2381 13695 2397 13759
rect 2461 13695 2477 13759
rect 2541 13695 2557 13759
rect 2621 13695 2637 13759
rect 2701 13695 2717 13759
rect 2781 13695 2797 13759
rect 2861 13695 2877 13759
rect 2941 13695 2957 13759
rect 3021 13695 3037 13759
rect 3101 13695 3117 13759
rect 3181 13695 3197 13759
rect 3261 13695 3277 13759
rect 3341 13695 3357 13759
rect 3421 13695 3437 13759
rect 3501 13695 3517 13759
rect 3581 13695 3597 13759
rect 3661 13695 3677 13759
rect 3741 13695 3757 13759
rect 3821 13695 3837 13759
rect 3901 13695 3917 13759
rect 3981 13695 3997 13759
rect 4061 13695 4077 13759
rect 4141 13695 4157 13759
rect 4221 13695 4237 13759
rect 4301 13695 4317 13759
rect 4381 13695 4397 13759
rect 4461 13695 4477 13759
rect 4541 13695 4557 13759
rect 4621 13695 4637 13759
rect 4701 13695 4717 13759
rect 4781 13695 4797 13759
rect 4861 13695 14666 13759
rect 334 13677 14666 13695
rect 381 13613 397 13677
rect 461 13613 477 13677
rect 541 13613 557 13677
rect 621 13613 637 13677
rect 701 13613 717 13677
rect 781 13613 797 13677
rect 861 13613 877 13677
rect 941 13613 957 13677
rect 1021 13613 1037 13677
rect 1101 13613 1117 13677
rect 1181 13613 1197 13677
rect 1261 13613 1277 13677
rect 1341 13613 1357 13677
rect 1421 13613 1437 13677
rect 1501 13613 1517 13677
rect 1581 13613 1597 13677
rect 1661 13613 1677 13677
rect 1741 13613 1757 13677
rect 1821 13613 1837 13677
rect 1901 13613 1917 13677
rect 1981 13613 1997 13677
rect 2061 13613 2077 13677
rect 2141 13613 2157 13677
rect 2221 13613 2237 13677
rect 2301 13613 2317 13677
rect 2381 13613 2397 13677
rect 2461 13613 2477 13677
rect 2541 13613 2557 13677
rect 2621 13613 2637 13677
rect 2701 13613 2717 13677
rect 2781 13613 2797 13677
rect 2861 13613 2877 13677
rect 2941 13613 2957 13677
rect 3021 13613 3037 13677
rect 3101 13613 3117 13677
rect 3181 13613 3197 13677
rect 3261 13613 3277 13677
rect 3341 13613 3357 13677
rect 3421 13613 3437 13677
rect 3501 13613 3517 13677
rect 3581 13613 3597 13677
rect 3661 13613 3677 13677
rect 3741 13613 3757 13677
rect 3821 13613 3837 13677
rect 3901 13613 3917 13677
rect 3981 13613 3997 13677
rect 4061 13613 4077 13677
rect 4141 13613 4157 13677
rect 4221 13613 4237 13677
rect 4301 13613 4317 13677
rect 4381 13613 4397 13677
rect 4461 13613 4477 13677
rect 4541 13613 4557 13677
rect 4621 13613 4637 13677
rect 4701 13613 4717 13677
rect 4781 13613 4797 13677
rect 4861 13613 14666 13677
rect 334 13527 14666 13613
rect 193 13387 14807 13527
rect 334 13304 14666 13387
rect 352 13240 369 13304
rect 433 13240 450 13304
rect 514 13240 531 13304
rect 595 13240 612 13304
rect 676 13240 693 13304
rect 757 13240 774 13304
rect 838 13240 855 13304
rect 919 13240 936 13304
rect 1000 13240 1017 13304
rect 1081 13240 1098 13304
rect 1162 13240 1179 13304
rect 1243 13240 1260 13304
rect 1324 13240 1341 13304
rect 1405 13240 1422 13304
rect 1486 13240 1503 13304
rect 1567 13240 1584 13304
rect 1648 13240 1665 13304
rect 1729 13240 1746 13304
rect 1810 13240 1827 13304
rect 1891 13240 1908 13304
rect 1972 13240 1989 13304
rect 2053 13240 2070 13304
rect 2134 13240 2151 13304
rect 2215 13240 2232 13304
rect 2296 13240 2313 13304
rect 2377 13240 2394 13304
rect 2458 13240 2475 13304
rect 2539 13240 2556 13304
rect 2620 13240 2637 13304
rect 2701 13240 2718 13304
rect 2782 13240 2799 13304
rect 2863 13240 2880 13304
rect 2944 13240 2961 13304
rect 3025 13240 3042 13304
rect 3106 13240 3123 13304
rect 3187 13240 3204 13304
rect 3268 13240 3285 13304
rect 3349 13240 3366 13304
rect 3430 13240 3447 13304
rect 3511 13240 3528 13304
rect 3592 13240 3609 13304
rect 3673 13240 3690 13304
rect 3754 13240 3771 13304
rect 3835 13240 3852 13304
rect 3916 13240 3933 13304
rect 3997 13240 4014 13304
rect 4078 13240 4095 13304
rect 4159 13240 4176 13304
rect 4240 13240 4257 13304
rect 4321 13240 4338 13304
rect 4402 13240 4420 13304
rect 4484 13240 4502 13304
rect 4566 13240 4584 13304
rect 4648 13240 4666 13304
rect 4730 13240 4748 13304
rect 4812 13240 4830 13304
rect 4894 13240 14666 13304
rect 334 13222 14666 13240
rect 352 13158 369 13222
rect 433 13158 450 13222
rect 514 13158 531 13222
rect 595 13158 612 13222
rect 676 13158 693 13222
rect 757 13158 774 13222
rect 838 13158 855 13222
rect 919 13158 936 13222
rect 1000 13158 1017 13222
rect 1081 13158 1098 13222
rect 1162 13158 1179 13222
rect 1243 13158 1260 13222
rect 1324 13158 1341 13222
rect 1405 13158 1422 13222
rect 1486 13158 1503 13222
rect 1567 13158 1584 13222
rect 1648 13158 1665 13222
rect 1729 13158 1746 13222
rect 1810 13158 1827 13222
rect 1891 13158 1908 13222
rect 1972 13158 1989 13222
rect 2053 13158 2070 13222
rect 2134 13158 2151 13222
rect 2215 13158 2232 13222
rect 2296 13158 2313 13222
rect 2377 13158 2394 13222
rect 2458 13158 2475 13222
rect 2539 13158 2556 13222
rect 2620 13158 2637 13222
rect 2701 13158 2718 13222
rect 2782 13158 2799 13222
rect 2863 13158 2880 13222
rect 2944 13158 2961 13222
rect 3025 13158 3042 13222
rect 3106 13158 3123 13222
rect 3187 13158 3204 13222
rect 3268 13158 3285 13222
rect 3349 13158 3366 13222
rect 3430 13158 3447 13222
rect 3511 13158 3528 13222
rect 3592 13158 3609 13222
rect 3673 13158 3690 13222
rect 3754 13158 3771 13222
rect 3835 13158 3852 13222
rect 3916 13158 3933 13222
rect 3997 13158 4014 13222
rect 4078 13158 4095 13222
rect 4159 13158 4176 13222
rect 4240 13158 4257 13222
rect 4321 13158 4338 13222
rect 4402 13158 4420 13222
rect 4484 13158 4502 13222
rect 4566 13158 4584 13222
rect 4648 13158 4666 13222
rect 4730 13158 4748 13222
rect 4812 13158 4830 13222
rect 4894 13158 14666 13222
rect 334 13140 14666 13158
rect 352 13076 369 13140
rect 433 13076 450 13140
rect 514 13076 531 13140
rect 595 13076 612 13140
rect 676 13076 693 13140
rect 757 13076 774 13140
rect 838 13076 855 13140
rect 919 13076 936 13140
rect 1000 13076 1017 13140
rect 1081 13076 1098 13140
rect 1162 13076 1179 13140
rect 1243 13076 1260 13140
rect 1324 13076 1341 13140
rect 1405 13076 1422 13140
rect 1486 13076 1503 13140
rect 1567 13076 1584 13140
rect 1648 13076 1665 13140
rect 1729 13076 1746 13140
rect 1810 13076 1827 13140
rect 1891 13076 1908 13140
rect 1972 13076 1989 13140
rect 2053 13076 2070 13140
rect 2134 13076 2151 13140
rect 2215 13076 2232 13140
rect 2296 13076 2313 13140
rect 2377 13076 2394 13140
rect 2458 13076 2475 13140
rect 2539 13076 2556 13140
rect 2620 13076 2637 13140
rect 2701 13076 2718 13140
rect 2782 13076 2799 13140
rect 2863 13076 2880 13140
rect 2944 13076 2961 13140
rect 3025 13076 3042 13140
rect 3106 13076 3123 13140
rect 3187 13076 3204 13140
rect 3268 13076 3285 13140
rect 3349 13076 3366 13140
rect 3430 13076 3447 13140
rect 3511 13076 3528 13140
rect 3592 13076 3609 13140
rect 3673 13076 3690 13140
rect 3754 13076 3771 13140
rect 3835 13076 3852 13140
rect 3916 13076 3933 13140
rect 3997 13076 4014 13140
rect 4078 13076 4095 13140
rect 4159 13076 4176 13140
rect 4240 13076 4257 13140
rect 4321 13076 4338 13140
rect 4402 13076 4420 13140
rect 4484 13076 4502 13140
rect 4566 13076 4584 13140
rect 4648 13076 4666 13140
rect 4730 13076 4748 13140
rect 4812 13076 4830 13140
rect 4894 13076 14666 13140
rect 334 13058 14666 13076
rect 352 12994 369 13058
rect 433 12994 450 13058
rect 514 12994 531 13058
rect 595 12994 612 13058
rect 676 12994 693 13058
rect 757 12994 774 13058
rect 838 12994 855 13058
rect 919 12994 936 13058
rect 1000 12994 1017 13058
rect 1081 12994 1098 13058
rect 1162 12994 1179 13058
rect 1243 12994 1260 13058
rect 1324 12994 1341 13058
rect 1405 12994 1422 13058
rect 1486 12994 1503 13058
rect 1567 12994 1584 13058
rect 1648 12994 1665 13058
rect 1729 12994 1746 13058
rect 1810 12994 1827 13058
rect 1891 12994 1908 13058
rect 1972 12994 1989 13058
rect 2053 12994 2070 13058
rect 2134 12994 2151 13058
rect 2215 12994 2232 13058
rect 2296 12994 2313 13058
rect 2377 12994 2394 13058
rect 2458 12994 2475 13058
rect 2539 12994 2556 13058
rect 2620 12994 2637 13058
rect 2701 12994 2718 13058
rect 2782 12994 2799 13058
rect 2863 12994 2880 13058
rect 2944 12994 2961 13058
rect 3025 12994 3042 13058
rect 3106 12994 3123 13058
rect 3187 12994 3204 13058
rect 3268 12994 3285 13058
rect 3349 12994 3366 13058
rect 3430 12994 3447 13058
rect 3511 12994 3528 13058
rect 3592 12994 3609 13058
rect 3673 12994 3690 13058
rect 3754 12994 3771 13058
rect 3835 12994 3852 13058
rect 3916 12994 3933 13058
rect 3997 12994 4014 13058
rect 4078 12994 4095 13058
rect 4159 12994 4176 13058
rect 4240 12994 4257 13058
rect 4321 12994 4338 13058
rect 4402 12994 4420 13058
rect 4484 12994 4502 13058
rect 4566 12994 4584 13058
rect 4648 12994 4666 13058
rect 4730 12994 4748 13058
rect 4812 12994 4830 13058
rect 4894 12994 14666 13058
rect 334 12976 14666 12994
rect 352 12912 369 12976
rect 433 12912 450 12976
rect 514 12912 531 12976
rect 595 12912 612 12976
rect 676 12912 693 12976
rect 757 12912 774 12976
rect 838 12912 855 12976
rect 919 12912 936 12976
rect 1000 12912 1017 12976
rect 1081 12912 1098 12976
rect 1162 12912 1179 12976
rect 1243 12912 1260 12976
rect 1324 12912 1341 12976
rect 1405 12912 1422 12976
rect 1486 12912 1503 12976
rect 1567 12912 1584 12976
rect 1648 12912 1665 12976
rect 1729 12912 1746 12976
rect 1810 12912 1827 12976
rect 1891 12912 1908 12976
rect 1972 12912 1989 12976
rect 2053 12912 2070 12976
rect 2134 12912 2151 12976
rect 2215 12912 2232 12976
rect 2296 12912 2313 12976
rect 2377 12912 2394 12976
rect 2458 12912 2475 12976
rect 2539 12912 2556 12976
rect 2620 12912 2637 12976
rect 2701 12912 2718 12976
rect 2782 12912 2799 12976
rect 2863 12912 2880 12976
rect 2944 12912 2961 12976
rect 3025 12912 3042 12976
rect 3106 12912 3123 12976
rect 3187 12912 3204 12976
rect 3268 12912 3285 12976
rect 3349 12912 3366 12976
rect 3430 12912 3447 12976
rect 3511 12912 3528 12976
rect 3592 12912 3609 12976
rect 3673 12912 3690 12976
rect 3754 12912 3771 12976
rect 3835 12912 3852 12976
rect 3916 12912 3933 12976
rect 3997 12912 4014 12976
rect 4078 12912 4095 12976
rect 4159 12912 4176 12976
rect 4240 12912 4257 12976
rect 4321 12912 4338 12976
rect 4402 12912 4420 12976
rect 4484 12912 4502 12976
rect 4566 12912 4584 12976
rect 4648 12912 4666 12976
rect 4730 12912 4748 12976
rect 4812 12912 4830 12976
rect 4894 12912 14666 12976
rect 334 12894 14666 12912
rect 352 12830 369 12894
rect 433 12830 450 12894
rect 514 12830 531 12894
rect 595 12830 612 12894
rect 676 12830 693 12894
rect 757 12830 774 12894
rect 838 12830 855 12894
rect 919 12830 936 12894
rect 1000 12830 1017 12894
rect 1081 12830 1098 12894
rect 1162 12830 1179 12894
rect 1243 12830 1260 12894
rect 1324 12830 1341 12894
rect 1405 12830 1422 12894
rect 1486 12830 1503 12894
rect 1567 12830 1584 12894
rect 1648 12830 1665 12894
rect 1729 12830 1746 12894
rect 1810 12830 1827 12894
rect 1891 12830 1908 12894
rect 1972 12830 1989 12894
rect 2053 12830 2070 12894
rect 2134 12830 2151 12894
rect 2215 12830 2232 12894
rect 2296 12830 2313 12894
rect 2377 12830 2394 12894
rect 2458 12830 2475 12894
rect 2539 12830 2556 12894
rect 2620 12830 2637 12894
rect 2701 12830 2718 12894
rect 2782 12830 2799 12894
rect 2863 12830 2880 12894
rect 2944 12830 2961 12894
rect 3025 12830 3042 12894
rect 3106 12830 3123 12894
rect 3187 12830 3204 12894
rect 3268 12830 3285 12894
rect 3349 12830 3366 12894
rect 3430 12830 3447 12894
rect 3511 12830 3528 12894
rect 3592 12830 3609 12894
rect 3673 12830 3690 12894
rect 3754 12830 3771 12894
rect 3835 12830 3852 12894
rect 3916 12830 3933 12894
rect 3997 12830 4014 12894
rect 4078 12830 4095 12894
rect 4159 12830 4176 12894
rect 4240 12830 4257 12894
rect 4321 12830 4338 12894
rect 4402 12830 4420 12894
rect 4484 12830 4502 12894
rect 4566 12830 4584 12894
rect 4648 12830 4666 12894
rect 4730 12830 4748 12894
rect 4812 12830 4830 12894
rect 4894 12830 14666 12894
rect 334 12812 14666 12830
rect 352 12748 369 12812
rect 433 12748 450 12812
rect 514 12748 531 12812
rect 595 12748 612 12812
rect 676 12748 693 12812
rect 757 12748 774 12812
rect 838 12748 855 12812
rect 919 12748 936 12812
rect 1000 12748 1017 12812
rect 1081 12748 1098 12812
rect 1162 12748 1179 12812
rect 1243 12748 1260 12812
rect 1324 12748 1341 12812
rect 1405 12748 1422 12812
rect 1486 12748 1503 12812
rect 1567 12748 1584 12812
rect 1648 12748 1665 12812
rect 1729 12748 1746 12812
rect 1810 12748 1827 12812
rect 1891 12748 1908 12812
rect 1972 12748 1989 12812
rect 2053 12748 2070 12812
rect 2134 12748 2151 12812
rect 2215 12748 2232 12812
rect 2296 12748 2313 12812
rect 2377 12748 2394 12812
rect 2458 12748 2475 12812
rect 2539 12748 2556 12812
rect 2620 12748 2637 12812
rect 2701 12748 2718 12812
rect 2782 12748 2799 12812
rect 2863 12748 2880 12812
rect 2944 12748 2961 12812
rect 3025 12748 3042 12812
rect 3106 12748 3123 12812
rect 3187 12748 3204 12812
rect 3268 12748 3285 12812
rect 3349 12748 3366 12812
rect 3430 12748 3447 12812
rect 3511 12748 3528 12812
rect 3592 12748 3609 12812
rect 3673 12748 3690 12812
rect 3754 12748 3771 12812
rect 3835 12748 3852 12812
rect 3916 12748 3933 12812
rect 3997 12748 4014 12812
rect 4078 12748 4095 12812
rect 4159 12748 4176 12812
rect 4240 12748 4257 12812
rect 4321 12748 4338 12812
rect 4402 12748 4420 12812
rect 4484 12748 4502 12812
rect 4566 12748 4584 12812
rect 4648 12748 4666 12812
rect 4730 12748 4748 12812
rect 4812 12748 4830 12812
rect 4894 12748 14666 12812
rect 334 12730 14666 12748
rect 352 12666 369 12730
rect 433 12666 450 12730
rect 514 12666 531 12730
rect 595 12666 612 12730
rect 676 12666 693 12730
rect 757 12666 774 12730
rect 838 12666 855 12730
rect 919 12666 936 12730
rect 1000 12666 1017 12730
rect 1081 12666 1098 12730
rect 1162 12666 1179 12730
rect 1243 12666 1260 12730
rect 1324 12666 1341 12730
rect 1405 12666 1422 12730
rect 1486 12666 1503 12730
rect 1567 12666 1584 12730
rect 1648 12666 1665 12730
rect 1729 12666 1746 12730
rect 1810 12666 1827 12730
rect 1891 12666 1908 12730
rect 1972 12666 1989 12730
rect 2053 12666 2070 12730
rect 2134 12666 2151 12730
rect 2215 12666 2232 12730
rect 2296 12666 2313 12730
rect 2377 12666 2394 12730
rect 2458 12666 2475 12730
rect 2539 12666 2556 12730
rect 2620 12666 2637 12730
rect 2701 12666 2718 12730
rect 2782 12666 2799 12730
rect 2863 12666 2880 12730
rect 2944 12666 2961 12730
rect 3025 12666 3042 12730
rect 3106 12666 3123 12730
rect 3187 12666 3204 12730
rect 3268 12666 3285 12730
rect 3349 12666 3366 12730
rect 3430 12666 3447 12730
rect 3511 12666 3528 12730
rect 3592 12666 3609 12730
rect 3673 12666 3690 12730
rect 3754 12666 3771 12730
rect 3835 12666 3852 12730
rect 3916 12666 3933 12730
rect 3997 12666 4014 12730
rect 4078 12666 4095 12730
rect 4159 12666 4176 12730
rect 4240 12666 4257 12730
rect 4321 12666 4338 12730
rect 4402 12666 4420 12730
rect 4484 12666 4502 12730
rect 4566 12666 4584 12730
rect 4648 12666 4666 12730
rect 4730 12666 4748 12730
rect 4812 12666 4830 12730
rect 4894 12666 14666 12730
rect 334 12648 14666 12666
rect 352 12584 369 12648
rect 433 12584 450 12648
rect 514 12584 531 12648
rect 595 12584 612 12648
rect 676 12584 693 12648
rect 757 12584 774 12648
rect 838 12584 855 12648
rect 919 12584 936 12648
rect 1000 12584 1017 12648
rect 1081 12584 1098 12648
rect 1162 12584 1179 12648
rect 1243 12584 1260 12648
rect 1324 12584 1341 12648
rect 1405 12584 1422 12648
rect 1486 12584 1503 12648
rect 1567 12584 1584 12648
rect 1648 12584 1665 12648
rect 1729 12584 1746 12648
rect 1810 12584 1827 12648
rect 1891 12584 1908 12648
rect 1972 12584 1989 12648
rect 2053 12584 2070 12648
rect 2134 12584 2151 12648
rect 2215 12584 2232 12648
rect 2296 12584 2313 12648
rect 2377 12584 2394 12648
rect 2458 12584 2475 12648
rect 2539 12584 2556 12648
rect 2620 12584 2637 12648
rect 2701 12584 2718 12648
rect 2782 12584 2799 12648
rect 2863 12584 2880 12648
rect 2944 12584 2961 12648
rect 3025 12584 3042 12648
rect 3106 12584 3123 12648
rect 3187 12584 3204 12648
rect 3268 12584 3285 12648
rect 3349 12584 3366 12648
rect 3430 12584 3447 12648
rect 3511 12584 3528 12648
rect 3592 12584 3609 12648
rect 3673 12584 3690 12648
rect 3754 12584 3771 12648
rect 3835 12584 3852 12648
rect 3916 12584 3933 12648
rect 3997 12584 4014 12648
rect 4078 12584 4095 12648
rect 4159 12584 4176 12648
rect 4240 12584 4257 12648
rect 4321 12584 4338 12648
rect 4402 12584 4420 12648
rect 4484 12584 4502 12648
rect 4566 12584 4584 12648
rect 4648 12584 4666 12648
rect 4730 12584 4748 12648
rect 4812 12584 4830 12648
rect 4894 12584 14666 12648
rect 334 12566 14666 12584
rect 352 12502 369 12566
rect 433 12502 450 12566
rect 514 12502 531 12566
rect 595 12502 612 12566
rect 676 12502 693 12566
rect 757 12502 774 12566
rect 838 12502 855 12566
rect 919 12502 936 12566
rect 1000 12502 1017 12566
rect 1081 12502 1098 12566
rect 1162 12502 1179 12566
rect 1243 12502 1260 12566
rect 1324 12502 1341 12566
rect 1405 12502 1422 12566
rect 1486 12502 1503 12566
rect 1567 12502 1584 12566
rect 1648 12502 1665 12566
rect 1729 12502 1746 12566
rect 1810 12502 1827 12566
rect 1891 12502 1908 12566
rect 1972 12502 1989 12566
rect 2053 12502 2070 12566
rect 2134 12502 2151 12566
rect 2215 12502 2232 12566
rect 2296 12502 2313 12566
rect 2377 12502 2394 12566
rect 2458 12502 2475 12566
rect 2539 12502 2556 12566
rect 2620 12502 2637 12566
rect 2701 12502 2718 12566
rect 2782 12502 2799 12566
rect 2863 12502 2880 12566
rect 2944 12502 2961 12566
rect 3025 12502 3042 12566
rect 3106 12502 3123 12566
rect 3187 12502 3204 12566
rect 3268 12502 3285 12566
rect 3349 12502 3366 12566
rect 3430 12502 3447 12566
rect 3511 12502 3528 12566
rect 3592 12502 3609 12566
rect 3673 12502 3690 12566
rect 3754 12502 3771 12566
rect 3835 12502 3852 12566
rect 3916 12502 3933 12566
rect 3997 12502 4014 12566
rect 4078 12502 4095 12566
rect 4159 12502 4176 12566
rect 4240 12502 4257 12566
rect 4321 12502 4338 12566
rect 4402 12502 4420 12566
rect 4484 12502 4502 12566
rect 4566 12502 4584 12566
rect 4648 12502 4666 12566
rect 4730 12502 4748 12566
rect 4812 12502 4830 12566
rect 4894 12502 14666 12566
rect 334 12484 14666 12502
rect 352 12420 369 12484
rect 433 12420 450 12484
rect 514 12420 531 12484
rect 595 12420 612 12484
rect 676 12420 693 12484
rect 757 12420 774 12484
rect 838 12420 855 12484
rect 919 12420 936 12484
rect 1000 12420 1017 12484
rect 1081 12420 1098 12484
rect 1162 12420 1179 12484
rect 1243 12420 1260 12484
rect 1324 12420 1341 12484
rect 1405 12420 1422 12484
rect 1486 12420 1503 12484
rect 1567 12420 1584 12484
rect 1648 12420 1665 12484
rect 1729 12420 1746 12484
rect 1810 12420 1827 12484
rect 1891 12420 1908 12484
rect 1972 12420 1989 12484
rect 2053 12420 2070 12484
rect 2134 12420 2151 12484
rect 2215 12420 2232 12484
rect 2296 12420 2313 12484
rect 2377 12420 2394 12484
rect 2458 12420 2475 12484
rect 2539 12420 2556 12484
rect 2620 12420 2637 12484
rect 2701 12420 2718 12484
rect 2782 12420 2799 12484
rect 2863 12420 2880 12484
rect 2944 12420 2961 12484
rect 3025 12420 3042 12484
rect 3106 12420 3123 12484
rect 3187 12420 3204 12484
rect 3268 12420 3285 12484
rect 3349 12420 3366 12484
rect 3430 12420 3447 12484
rect 3511 12420 3528 12484
rect 3592 12420 3609 12484
rect 3673 12420 3690 12484
rect 3754 12420 3771 12484
rect 3835 12420 3852 12484
rect 3916 12420 3933 12484
rect 3997 12420 4014 12484
rect 4078 12420 4095 12484
rect 4159 12420 4176 12484
rect 4240 12420 4257 12484
rect 4321 12420 4338 12484
rect 4402 12420 4420 12484
rect 4484 12420 4502 12484
rect 4566 12420 4584 12484
rect 4648 12420 4666 12484
rect 4730 12420 4748 12484
rect 4812 12420 4830 12484
rect 4894 12420 14666 12484
rect 334 12337 14666 12420
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10151 12418 14931 13306 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13252 14913 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13170 14913 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13088 14913 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13006 14913 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12924 14913 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12842 14913 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12760 14913 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12678 14913 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12596 14913 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12514 14913 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12432 14913 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13252 14831 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13170 14831 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13088 14831 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13006 14831 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12924 14831 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12842 14831 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12760 14831 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12678 14831 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12596 14831 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12514 14831 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12432 14831 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13252 14749 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13170 14749 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13088 14749 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13006 14749 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12924 14749 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12842 14749 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12760 14749 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12678 14749 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12596 14749 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12514 14749 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12432 14749 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13252 14667 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13170 14667 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13088 14667 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13006 14667 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12924 14667 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12842 14667 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12760 14667 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12678 14667 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12596 14667 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12514 14667 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12432 14667 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13252 14585 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13170 14585 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13088 14585 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13006 14585 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12924 14585 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12842 14585 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12760 14585 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12678 14585 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12596 14585 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12514 14585 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12432 14585 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13252 14503 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13170 14503 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13088 14503 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13006 14503 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12924 14503 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12842 14503 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12760 14503 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12678 14503 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12596 14503 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12514 14503 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12432 14503 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13252 14421 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13170 14421 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13088 14421 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13006 14421 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12924 14421 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12842 14421 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12760 14421 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12678 14421 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12596 14421 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12514 14421 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12432 14421 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13252 14340 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13170 14340 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13088 14340 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13006 14340 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12924 14340 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12842 14340 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12760 14340 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12678 14340 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12596 14340 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12514 14340 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12432 14340 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13252 14259 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13170 14259 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13088 14259 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13006 14259 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12924 14259 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12842 14259 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12760 14259 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12678 14259 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12596 14259 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12514 14259 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12432 14259 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13252 14178 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13170 14178 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13088 14178 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13006 14178 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12924 14178 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12842 14178 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12760 14178 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12678 14178 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12596 14178 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12514 14178 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12432 14178 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13252 14097 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13170 14097 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13088 14097 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13006 14097 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12924 14097 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12842 14097 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12760 14097 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12678 14097 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12596 14097 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12514 14097 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12432 14097 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13252 14016 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13170 14016 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13088 14016 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13006 14016 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12924 14016 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12842 14016 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12760 14016 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12678 14016 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12596 14016 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12514 14016 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12432 14016 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13252 13935 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13170 13935 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13088 13935 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13006 13935 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12924 13935 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12842 13935 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12760 13935 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12678 13935 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12596 13935 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12514 13935 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12432 13935 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13252 13854 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13170 13854 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13088 13854 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13006 13854 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12924 13854 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12842 13854 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12760 13854 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12678 13854 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12596 13854 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12514 13854 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12432 13854 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13252 13773 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13170 13773 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13088 13773 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13006 13773 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12924 13773 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12842 13773 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12760 13773 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12678 13773 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12596 13773 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12514 13773 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12432 13773 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13252 13692 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13170 13692 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13088 13692 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13006 13692 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12924 13692 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12842 13692 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12760 13692 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12678 13692 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12596 13692 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12514 13692 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12432 13692 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13252 13611 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13170 13611 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13088 13611 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13006 13611 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12924 13611 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12842 13611 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12760 13611 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12678 13611 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12596 13611 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12514 13611 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12432 13611 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13252 13530 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13170 13530 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13088 13530 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13006 13530 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12924 13530 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12842 13530 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12760 13530 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12678 13530 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12596 13530 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12514 13530 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12432 13530 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13252 13449 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13170 13449 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13088 13449 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13006 13449 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12924 13449 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12842 13449 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12760 13449 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12678 13449 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12596 13449 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12514 13449 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12432 13449 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13252 13368 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13170 13368 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13088 13368 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13006 13368 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12924 13368 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12842 13368 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12760 13368 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12678 13368 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12596 13368 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12514 13368 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12432 13368 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13252 13287 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13170 13287 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13088 13287 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13006 13287 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12924 13287 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12842 13287 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12760 13287 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12678 13287 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12596 13287 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12514 13287 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12432 13287 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13252 13206 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13170 13206 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13088 13206 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13006 13206 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12924 13206 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12842 13206 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12760 13206 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12678 13206 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12596 13206 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12514 13206 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12432 13206 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13252 13125 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13170 13125 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13088 13125 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13006 13125 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12924 13125 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12842 13125 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12760 13125 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12678 13125 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12596 13125 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12514 13125 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12432 13125 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13252 13044 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13170 13044 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13088 13044 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13006 13044 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12924 13044 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12842 13044 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12760 13044 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12678 13044 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12596 13044 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12514 13044 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12432 13044 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13252 12963 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13170 12963 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13088 12963 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13006 12963 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12924 12963 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12842 12963 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12760 12963 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12678 12963 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12596 12963 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12514 12963 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12432 12963 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13252 12882 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13170 12882 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13088 12882 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13006 12882 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12924 12882 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12842 12882 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12760 12882 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12678 12882 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12596 12882 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12514 12882 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12432 12882 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13252 12801 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13170 12801 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13088 12801 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13006 12801 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12924 12801 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12842 12801 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12760 12801 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12678 12801 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12596 12801 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12514 12801 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12432 12801 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13252 12720 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13170 12720 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13088 12720 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13006 12720 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12924 12720 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12842 12720 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12760 12720 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12678 12720 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12596 12720 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12514 12720 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12432 12720 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13252 12639 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13170 12639 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13088 12639 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13006 12639 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12924 12639 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12842 12639 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12760 12639 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12678 12639 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12596 12639 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12514 12639 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12432 12639 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13252 12558 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13170 12558 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13088 12558 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13006 12558 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12924 12558 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12842 12558 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12760 12558 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12678 12558 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12596 12558 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12514 12558 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12432 12558 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13252 12477 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13170 12477 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13088 12477 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13006 12477 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12924 12477 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12842 12477 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12760 12477 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12678 12477 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12596 12477 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12514 12477 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12432 12477 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13252 12396 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13170 12396 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13088 12396 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13006 12396 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12924 12396 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12842 12396 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12760 12396 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12678 12396 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12596 12396 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12514 12396 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12432 12396 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13252 12315 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13170 12315 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13088 12315 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13006 12315 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12924 12315 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12842 12315 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12760 12315 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12678 12315 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12596 12315 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12514 12315 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12432 12315 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13252 12234 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13170 12234 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13088 12234 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13006 12234 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12924 12234 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12842 12234 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12760 12234 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12678 12234 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12596 12234 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12514 12234 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12432 12234 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13252 12153 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13170 12153 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13088 12153 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13006 12153 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12924 12153 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12842 12153 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12760 12153 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12678 12153 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12596 12153 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12514 12153 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12432 12153 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13252 12072 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13170 12072 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13088 12072 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13006 12072 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12924 12072 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12842 12072 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12760 12072 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12678 12072 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12596 12072 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12514 12072 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12432 12072 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13252 11991 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13170 11991 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13088 11991 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13006 11991 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12924 11991 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12842 11991 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12760 11991 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12678 11991 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12596 11991 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12514 11991 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12432 11991 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13252 11910 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13170 11910 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13088 11910 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13006 11910 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12924 11910 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12842 11910 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12760 11910 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12678 11910 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12596 11910 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12514 11910 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12432 11910 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13252 11829 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13170 11829 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13088 11829 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13006 11829 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12924 11829 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12842 11829 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12760 11829 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12678 11829 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12596 11829 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12514 11829 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12432 11829 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13252 11748 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13170 11748 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13088 11748 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13006 11748 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12924 11748 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12842 11748 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12760 11748 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12678 11748 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12596 11748 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12514 11748 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12432 11748 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13252 11667 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13170 11667 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13088 11667 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13006 11667 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12924 11667 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12842 11667 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12760 11667 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12678 11667 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12596 11667 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12514 11667 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12432 11667 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13252 11586 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13170 11586 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13088 11586 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13006 11586 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12924 11586 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12842 11586 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12760 11586 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12678 11586 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12596 11586 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12514 11586 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12432 11586 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13252 11505 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13170 11505 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13088 11505 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13006 11505 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12924 11505 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12842 11505 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12760 11505 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12678 11505 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12596 11505 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12514 11505 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12432 11505 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13252 11424 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13170 11424 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13088 11424 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13006 11424 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12924 11424 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12842 11424 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12760 11424 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12678 11424 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12596 11424 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12514 11424 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12432 11424 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13252 11343 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13170 11343 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13088 11343 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13006 11343 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12924 11343 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12842 11343 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12760 11343 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12678 11343 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12596 11343 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12514 11343 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12432 11343 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13252 11262 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13170 11262 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13088 11262 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13006 11262 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12924 11262 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12842 11262 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12760 11262 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12678 11262 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12596 11262 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12514 11262 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12432 11262 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13252 11181 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13170 11181 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13088 11181 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13006 11181 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12924 11181 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12842 11181 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12760 11181 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12678 11181 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12596 11181 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12514 11181 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12432 11181 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13252 11100 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13170 11100 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13088 11100 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13006 11100 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12924 11100 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12842 11100 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12760 11100 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12678 11100 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12596 11100 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12514 11100 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12432 11100 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13252 11019 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13170 11019 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13088 11019 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13006 11019 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12924 11019 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12842 11019 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12760 11019 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12678 11019 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12596 11019 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12514 11019 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12432 11019 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13252 10938 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13170 10938 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13088 10938 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13006 10938 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12924 10938 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12842 10938 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12760 10938 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12678 10938 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12596 10938 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12514 10938 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12432 10938 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13252 10857 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13170 10857 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13088 10857 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13006 10857 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12924 10857 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12842 10857 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12760 10857 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12678 10857 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12596 10857 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12514 10857 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12432 10857 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13252 10776 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13170 10776 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13088 10776 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13006 10776 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12924 10776 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12842 10776 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12760 10776 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12678 10776 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12596 10776 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12514 10776 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12432 10776 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13252 10695 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13170 10695 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13088 10695 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13006 10695 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12924 10695 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12842 10695 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12760 10695 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12678 10695 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12596 10695 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12514 10695 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12432 10695 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13252 10614 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13170 10614 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13088 10614 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13006 10614 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12924 10614 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12842 10614 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12760 10614 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12678 10614 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12596 10614 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12514 10614 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12432 10614 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13252 10533 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13170 10533 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13088 10533 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13006 10533 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12924 10533 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12842 10533 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12760 10533 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12678 10533 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12596 10533 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12514 10533 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12432 10533 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13252 10452 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13170 10452 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13088 10452 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13006 10452 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12924 10452 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12842 10452 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12760 10452 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12678 10452 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12596 10452 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12514 10452 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12432 10452 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13252 10371 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13170 10371 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13088 10371 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13006 10371 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12924 10371 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12842 10371 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12760 10371 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12678 10371 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12596 10371 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12514 10371 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12432 10371 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13252 10290 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13170 10290 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13088 10290 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13006 10290 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12924 10290 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12842 10290 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12760 10290 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12678 10290 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12596 10290 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12514 10290 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12432 10290 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13252 10209 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13170 10209 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13088 10209 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13006 10209 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12924 10209 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12842 10209 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12760 10209 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12678 10209 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12596 10209 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12514 10209 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12432 10209 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 13240 4894 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13240 4894 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 13158 4894 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13158 4894 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 13076 4894 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13076 4894 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12994 4894 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12994 4894 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12912 4894 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12912 4894 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12830 4894 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12830 4894 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12748 4894 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12748 4894 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12666 4894 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12666 4894 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12584 4894 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12584 4894 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12502 4894 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12502 4894 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4830 12420 4894 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12420 4894 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 13240 4812 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13240 4812 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 13158 4812 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13158 4812 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 13076 4812 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13076 4812 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12994 4812 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12994 4812 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12912 4812 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12912 4812 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12830 4812 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12830 4812 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12748 4812 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12748 4812 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12666 4812 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12666 4812 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12584 4812 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12584 4812 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12502 4812 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12502 4812 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4748 12420 4812 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12420 4812 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 13240 4730 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13240 4730 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 13158 4730 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13158 4730 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 13076 4730 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13076 4730 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12994 4730 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12994 4730 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12912 4730 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12912 4730 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12830 4730 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12830 4730 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12748 4730 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12748 4730 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12666 4730 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12666 4730 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12584 4730 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12584 4730 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12502 4730 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12502 4730 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4666 12420 4730 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12420 4730 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 13240 4648 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13240 4648 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 13158 4648 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13158 4648 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 13076 4648 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13076 4648 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12994 4648 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12994 4648 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12912 4648 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12912 4648 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12830 4648 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12830 4648 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12748 4648 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12748 4648 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12666 4648 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12666 4648 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12584 4648 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12584 4648 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12502 4648 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12502 4648 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4584 12420 4648 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12420 4648 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 13240 4566 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13240 4566 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 13158 4566 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13158 4566 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 13076 4566 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13076 4566 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12994 4566 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12994 4566 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12912 4566 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12912 4566 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12830 4566 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12830 4566 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12748 4566 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12748 4566 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12666 4566 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12666 4566 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12584 4566 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12584 4566 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12502 4566 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12502 4566 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4502 12420 4566 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12420 4566 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 13240 4484 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13240 4484 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 13158 4484 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13158 4484 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 13076 4484 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13076 4484 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12994 4484 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12994 4484 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12912 4484 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12912 4484 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12830 4484 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12830 4484 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12748 4484 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12748 4484 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12666 4484 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12666 4484 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12584 4484 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12584 4484 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12502 4484 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12502 4484 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4420 12420 4484 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12420 4484 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 13240 4402 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13240 4402 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 13158 4402 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13158 4402 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 13076 4402 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13076 4402 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12994 4402 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12994 4402 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12912 4402 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12912 4402 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12830 4402 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12830 4402 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12748 4402 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12748 4402 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12666 4402 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12666 4402 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12584 4402 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12584 4402 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12502 4402 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12502 4402 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4338 12420 4402 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12420 4402 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 13240 4321 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13240 4321 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 13158 4321 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13158 4321 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 13076 4321 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13076 4321 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12994 4321 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12994 4321 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12912 4321 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12912 4321 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12830 4321 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12830 4321 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12748 4321 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12748 4321 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12666 4321 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12666 4321 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12584 4321 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12584 4321 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12502 4321 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12502 4321 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4257 12420 4321 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12420 4321 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 13240 4240 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13240 4240 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 13158 4240 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13158 4240 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 13076 4240 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13076 4240 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12994 4240 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12994 4240 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12912 4240 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12912 4240 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12830 4240 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12830 4240 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12748 4240 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12748 4240 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12666 4240 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12666 4240 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12584 4240 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12584 4240 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12502 4240 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12502 4240 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4176 12420 4240 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12420 4240 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 13240 4159 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13240 4159 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 13158 4159 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13158 4159 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 13076 4159 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13076 4159 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12994 4159 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12994 4159 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12912 4159 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12912 4159 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12830 4159 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12830 4159 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12748 4159 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12748 4159 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12666 4159 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12666 4159 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12584 4159 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12584 4159 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12502 4159 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12502 4159 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4095 12420 4159 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12420 4159 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 13240 4078 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13240 4078 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 13158 4078 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13158 4078 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 13076 4078 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13076 4078 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12994 4078 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12994 4078 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12912 4078 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12912 4078 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12830 4078 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12830 4078 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12748 4078 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12748 4078 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12666 4078 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12666 4078 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12584 4078 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12584 4078 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12502 4078 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12502 4078 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 4014 12420 4078 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12420 4078 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 13240 3997 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13240 3997 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 13158 3997 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13158 3997 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 13076 3997 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13076 3997 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12994 3997 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12994 3997 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12912 3997 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12912 3997 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12830 3997 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12830 3997 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12748 3997 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12748 3997 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12666 3997 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12666 3997 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12584 3997 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12584 3997 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12502 3997 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12502 3997 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3933 12420 3997 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12420 3997 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 13240 3916 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13240 3916 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 13158 3916 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13158 3916 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 13076 3916 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13076 3916 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12994 3916 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12994 3916 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12912 3916 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12912 3916 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12830 3916 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12830 3916 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12748 3916 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12748 3916 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12666 3916 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12666 3916 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12584 3916 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12584 3916 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12502 3916 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12502 3916 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3852 12420 3916 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12420 3916 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 13240 3835 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13240 3835 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 13158 3835 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13158 3835 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 13076 3835 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13076 3835 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12994 3835 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12994 3835 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12912 3835 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12912 3835 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12830 3835 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12830 3835 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12748 3835 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12748 3835 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12666 3835 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12666 3835 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12584 3835 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12584 3835 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12502 3835 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12502 3835 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3771 12420 3835 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12420 3835 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 13240 3754 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13240 3754 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 13158 3754 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13158 3754 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 13076 3754 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13076 3754 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12994 3754 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12994 3754 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12912 3754 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12912 3754 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12830 3754 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12830 3754 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12748 3754 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12748 3754 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12666 3754 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12666 3754 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12584 3754 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12584 3754 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12502 3754 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12502 3754 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3690 12420 3754 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12420 3754 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 13240 3673 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13240 3673 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 13158 3673 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13158 3673 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 13076 3673 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13076 3673 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12994 3673 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12994 3673 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12912 3673 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12912 3673 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12830 3673 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12830 3673 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12748 3673 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12748 3673 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12666 3673 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12666 3673 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12584 3673 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12584 3673 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12502 3673 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12502 3673 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3609 12420 3673 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12420 3673 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 13240 3592 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13240 3592 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 13158 3592 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13158 3592 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 13076 3592 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13076 3592 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12994 3592 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12994 3592 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12912 3592 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12912 3592 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12830 3592 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12830 3592 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12748 3592 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12748 3592 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12666 3592 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12666 3592 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12584 3592 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12584 3592 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12502 3592 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12502 3592 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3528 12420 3592 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12420 3592 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 13240 3511 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13240 3511 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 13158 3511 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13158 3511 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 13076 3511 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13076 3511 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12994 3511 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12994 3511 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12912 3511 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12912 3511 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12830 3511 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12830 3511 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12748 3511 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12748 3511 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12666 3511 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12666 3511 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12584 3511 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12584 3511 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12502 3511 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12502 3511 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3447 12420 3511 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12420 3511 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 13240 3430 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13240 3430 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 13158 3430 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13158 3430 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 13076 3430 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13076 3430 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12994 3430 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12994 3430 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12912 3430 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12912 3430 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12830 3430 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12830 3430 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12748 3430 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12748 3430 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12666 3430 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12666 3430 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12584 3430 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12584 3430 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12502 3430 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12502 3430 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3366 12420 3430 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12420 3430 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 13240 3349 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13240 3349 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 13158 3349 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13158 3349 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 13076 3349 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13076 3349 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12994 3349 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12994 3349 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12912 3349 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12912 3349 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12830 3349 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12830 3349 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12748 3349 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12748 3349 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12666 3349 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12666 3349 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12584 3349 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12584 3349 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12502 3349 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12502 3349 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3285 12420 3349 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12420 3349 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 13240 3268 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13240 3268 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 13158 3268 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13158 3268 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 13076 3268 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13076 3268 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12994 3268 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12994 3268 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12912 3268 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12912 3268 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12830 3268 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12830 3268 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12748 3268 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12748 3268 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12666 3268 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12666 3268 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12584 3268 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12584 3268 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12502 3268 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12502 3268 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3204 12420 3268 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12420 3268 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 13240 3187 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13240 3187 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 13158 3187 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13158 3187 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 13076 3187 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13076 3187 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12994 3187 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12994 3187 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12912 3187 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12912 3187 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12830 3187 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12830 3187 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12748 3187 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12748 3187 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12666 3187 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12666 3187 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12584 3187 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12584 3187 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12502 3187 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12502 3187 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3123 12420 3187 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12420 3187 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 13240 3106 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13240 3106 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 13158 3106 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13158 3106 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 13076 3106 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13076 3106 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12994 3106 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12994 3106 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12912 3106 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12912 3106 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12830 3106 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12830 3106 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12748 3106 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12748 3106 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12666 3106 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12666 3106 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12584 3106 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12584 3106 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12502 3106 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12502 3106 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 3042 12420 3106 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12420 3106 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 13240 3025 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13240 3025 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 13158 3025 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13158 3025 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 13076 3025 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13076 3025 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12994 3025 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12994 3025 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12912 3025 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12912 3025 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12830 3025 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12830 3025 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12748 3025 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12748 3025 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12666 3025 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12666 3025 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12584 3025 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12584 3025 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12502 3025 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12502 3025 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2961 12420 3025 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12420 3025 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 13240 2944 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13240 2944 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 13158 2944 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13158 2944 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 13076 2944 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13076 2944 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12994 2944 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12994 2944 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12912 2944 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12912 2944 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12830 2944 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12830 2944 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12748 2944 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12748 2944 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12666 2944 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12666 2944 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12584 2944 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12584 2944 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12502 2944 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12502 2944 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2880 12420 2944 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12420 2944 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 13240 2863 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13240 2863 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 13158 2863 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13158 2863 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 13076 2863 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13076 2863 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12994 2863 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12994 2863 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12912 2863 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12912 2863 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12830 2863 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12830 2863 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12748 2863 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12748 2863 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12666 2863 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12666 2863 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12584 2863 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12584 2863 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12502 2863 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12502 2863 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2799 12420 2863 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12420 2863 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 13240 2782 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13240 2782 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 13158 2782 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13158 2782 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 13076 2782 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13076 2782 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12994 2782 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12994 2782 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12912 2782 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12912 2782 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12830 2782 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12830 2782 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12748 2782 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12748 2782 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12666 2782 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12666 2782 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12584 2782 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12584 2782 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12502 2782 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12502 2782 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2718 12420 2782 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12420 2782 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 13240 2701 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13240 2701 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 13158 2701 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13158 2701 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 13076 2701 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13076 2701 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12994 2701 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12994 2701 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12912 2701 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12912 2701 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12830 2701 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12830 2701 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12748 2701 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12748 2701 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12666 2701 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12666 2701 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12584 2701 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12584 2701 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12502 2701 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12502 2701 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2637 12420 2701 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12420 2701 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 13240 2620 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13240 2620 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 13158 2620 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13158 2620 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 13076 2620 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13076 2620 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12994 2620 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12994 2620 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12912 2620 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12912 2620 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12830 2620 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12830 2620 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12748 2620 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12748 2620 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12666 2620 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12666 2620 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12584 2620 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12584 2620 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12502 2620 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12502 2620 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2556 12420 2620 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12420 2620 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 13240 2539 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13240 2539 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 13158 2539 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13158 2539 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 13076 2539 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13076 2539 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12994 2539 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12994 2539 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12912 2539 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12912 2539 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12830 2539 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12830 2539 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12748 2539 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12748 2539 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12666 2539 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12666 2539 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12584 2539 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12584 2539 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12502 2539 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12502 2539 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2475 12420 2539 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12420 2539 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 13240 2458 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13240 2458 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 13158 2458 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13158 2458 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 13076 2458 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13076 2458 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12994 2458 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12994 2458 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12912 2458 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12912 2458 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12830 2458 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12830 2458 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12748 2458 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12748 2458 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12666 2458 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12666 2458 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12584 2458 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12584 2458 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12502 2458 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12502 2458 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2394 12420 2458 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12420 2458 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 13240 2377 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13240 2377 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 13158 2377 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13158 2377 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 13076 2377 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13076 2377 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12994 2377 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12994 2377 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12912 2377 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12912 2377 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12830 2377 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12830 2377 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12748 2377 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12748 2377 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12666 2377 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12666 2377 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12584 2377 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12584 2377 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12502 2377 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12502 2377 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2313 12420 2377 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12420 2377 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 13240 2296 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13240 2296 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 13158 2296 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13158 2296 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 13076 2296 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13076 2296 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12994 2296 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12994 2296 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12912 2296 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12912 2296 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12830 2296 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12830 2296 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12748 2296 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12748 2296 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12666 2296 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12666 2296 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12584 2296 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12584 2296 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12502 2296 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12502 2296 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2232 12420 2296 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12420 2296 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 13240 2215 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13240 2215 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 13158 2215 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13158 2215 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 13076 2215 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13076 2215 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12994 2215 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12994 2215 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12912 2215 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12912 2215 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12830 2215 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12830 2215 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12748 2215 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12748 2215 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12666 2215 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12666 2215 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12584 2215 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12584 2215 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12502 2215 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12502 2215 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2151 12420 2215 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12420 2215 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 13240 2134 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13240 2134 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 13158 2134 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13158 2134 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 13076 2134 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13076 2134 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12994 2134 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12994 2134 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12912 2134 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12912 2134 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12830 2134 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12830 2134 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12748 2134 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12748 2134 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12666 2134 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12666 2134 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12584 2134 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12584 2134 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12502 2134 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12502 2134 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 2070 12420 2134 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12420 2134 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 13240 2053 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13240 2053 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 13158 2053 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13158 2053 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 13076 2053 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13076 2053 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12994 2053 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12994 2053 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12912 2053 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12912 2053 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12830 2053 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12830 2053 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12748 2053 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12748 2053 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12666 2053 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12666 2053 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12584 2053 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12584 2053 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12502 2053 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12502 2053 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1989 12420 2053 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12420 2053 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 13240 1972 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13240 1972 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 13158 1972 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13158 1972 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 13076 1972 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13076 1972 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12994 1972 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12994 1972 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12912 1972 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12912 1972 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12830 1972 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12830 1972 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12748 1972 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12748 1972 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12666 1972 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12666 1972 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12584 1972 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12584 1972 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12502 1972 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12502 1972 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1908 12420 1972 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12420 1972 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 13240 1891 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13240 1891 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 13158 1891 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13158 1891 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 13076 1891 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13076 1891 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12994 1891 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12994 1891 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12912 1891 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12912 1891 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12830 1891 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12830 1891 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12748 1891 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12748 1891 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12666 1891 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12666 1891 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12584 1891 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12584 1891 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12502 1891 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12502 1891 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1827 12420 1891 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12420 1891 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 13240 1810 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13240 1810 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 13158 1810 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13158 1810 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 13076 1810 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13076 1810 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12994 1810 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12994 1810 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12912 1810 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12912 1810 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12830 1810 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12830 1810 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12748 1810 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12748 1810 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12666 1810 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12666 1810 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12584 1810 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12584 1810 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12502 1810 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12502 1810 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1746 12420 1810 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12420 1810 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 13240 1729 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13240 1729 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 13158 1729 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13158 1729 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 13076 1729 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13076 1729 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12994 1729 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12994 1729 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12912 1729 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12912 1729 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12830 1729 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12830 1729 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12748 1729 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12748 1729 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12666 1729 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12666 1729 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12584 1729 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12584 1729 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12502 1729 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12502 1729 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1665 12420 1729 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12420 1729 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 13240 1648 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13240 1648 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 13158 1648 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13158 1648 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 13076 1648 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13076 1648 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12994 1648 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12994 1648 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12912 1648 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12912 1648 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12830 1648 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12830 1648 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12748 1648 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12748 1648 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12666 1648 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12666 1648 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12584 1648 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12584 1648 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12502 1648 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12502 1648 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1584 12420 1648 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12420 1648 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 13240 1567 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13240 1567 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 13158 1567 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13158 1567 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 13076 1567 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13076 1567 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12994 1567 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12994 1567 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12912 1567 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12912 1567 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12830 1567 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12830 1567 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12748 1567 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12748 1567 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12666 1567 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12666 1567 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12584 1567 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12584 1567 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12502 1567 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12502 1567 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1503 12420 1567 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12420 1567 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 13240 1486 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13240 1486 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 13158 1486 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13158 1486 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 13076 1486 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13076 1486 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12994 1486 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12994 1486 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12912 1486 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12912 1486 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12830 1486 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12830 1486 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12748 1486 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12748 1486 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12666 1486 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12666 1486 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12584 1486 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12584 1486 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12502 1486 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12502 1486 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1422 12420 1486 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12420 1486 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 13240 1405 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13240 1405 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 13158 1405 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13158 1405 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 13076 1405 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13076 1405 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12994 1405 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12994 1405 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12912 1405 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12912 1405 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12830 1405 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12830 1405 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12748 1405 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12748 1405 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12666 1405 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12666 1405 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12584 1405 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12584 1405 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12502 1405 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12502 1405 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1341 12420 1405 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12420 1405 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 13240 1324 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13240 1324 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 13158 1324 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13158 1324 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 13076 1324 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13076 1324 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12994 1324 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12994 1324 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12912 1324 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12912 1324 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12830 1324 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12830 1324 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12748 1324 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12748 1324 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12666 1324 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12666 1324 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12584 1324 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12584 1324 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12502 1324 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12502 1324 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1260 12420 1324 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12420 1324 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 13240 1243 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13240 1243 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 13158 1243 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13158 1243 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 13076 1243 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13076 1243 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12994 1243 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12994 1243 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12912 1243 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12912 1243 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12830 1243 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12830 1243 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12748 1243 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12748 1243 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12666 1243 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12666 1243 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12584 1243 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12584 1243 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12502 1243 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12502 1243 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1179 12420 1243 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12420 1243 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 13240 1162 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13240 1162 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 13158 1162 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13158 1162 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 13076 1162 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13076 1162 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12994 1162 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12994 1162 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12912 1162 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12912 1162 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12830 1162 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12830 1162 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12748 1162 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12748 1162 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12666 1162 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12666 1162 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12584 1162 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12584 1162 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12502 1162 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12502 1162 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1098 12420 1162 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12420 1162 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 13240 1081 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13240 1081 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 13158 1081 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13158 1081 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 13076 1081 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13076 1081 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12994 1081 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12994 1081 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12912 1081 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12912 1081 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12830 1081 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12830 1081 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12748 1081 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12748 1081 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12666 1081 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12666 1081 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12584 1081 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12584 1081 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12502 1081 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12502 1081 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 1017 12420 1081 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12420 1081 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 13240 1000 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13240 1000 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 13158 1000 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13158 1000 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 13076 1000 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13076 1000 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12994 1000 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12994 1000 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12912 1000 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12912 1000 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12830 1000 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12830 1000 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12748 1000 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12748 1000 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12666 1000 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12666 1000 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12584 1000 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12584 1000 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12502 1000 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12502 1000 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 936 12420 1000 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12420 1000 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 13240 919 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13240 919 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 13158 919 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13158 919 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 13076 919 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13076 919 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12994 919 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12994 919 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12912 919 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12912 919 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12830 919 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12830 919 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12748 919 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12748 919 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12666 919 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12666 919 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12584 919 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12584 919 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12502 919 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12502 919 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 855 12420 919 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12420 919 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 13240 838 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13240 838 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 13158 838 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13158 838 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 13076 838 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13076 838 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12994 838 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12994 838 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12912 838 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12912 838 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12830 838 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12830 838 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12748 838 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12748 838 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12666 838 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12666 838 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12584 838 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12584 838 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12502 838 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12502 838 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 774 12420 838 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12420 838 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 13240 757 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13240 757 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 13158 757 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13158 757 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 13076 757 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13076 757 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12994 757 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12994 757 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12912 757 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12912 757 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12830 757 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12830 757 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12748 757 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12748 757 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12666 757 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12666 757 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12584 757 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12584 757 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12502 757 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12502 757 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 693 12420 757 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12420 757 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 13240 676 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13240 676 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 13158 676 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13158 676 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 13076 676 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13076 676 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12994 676 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12994 676 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12912 676 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12912 676 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12830 676 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12830 676 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12748 676 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12748 676 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12666 676 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12666 676 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12584 676 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12584 676 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12502 676 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12502 676 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 612 12420 676 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12420 676 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 13240 595 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13240 595 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 13158 595 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13158 595 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 13076 595 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13076 595 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12994 595 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12994 595 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12912 595 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12912 595 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12830 595 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12830 595 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12748 595 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12748 595 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12666 595 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12666 595 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12584 595 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12584 595 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12502 595 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12502 595 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 531 12420 595 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12420 595 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 13240 514 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13240 514 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 13158 514 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13158 514 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 13076 514 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13076 514 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12994 514 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12994 514 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12912 514 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12912 514 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12830 514 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12830 514 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12748 514 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12748 514 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12666 514 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12666 514 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12584 514 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12584 514 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12502 514 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12502 514 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 450 12420 514 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12420 514 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 13240 433 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13240 433 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 13158 433 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13158 433 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 13076 433 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13076 433 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12994 433 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12994 433 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12912 433 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12912 433 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12830 433 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12830 433 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12748 433 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12748 433 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12666 433 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12666 433 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12584 433 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12584 433 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12502 433 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12502 433 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 369 12420 433 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12420 433 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 13240 352 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13240 352 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 13158 352 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13158 352 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 13076 352 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13076 352 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12994 352 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12994 352 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12912 352 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12912 352 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12830 352 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12830 352 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12748 352 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12748 352 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12666 352 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12666 352 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12584 352 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12584 352 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12502 352 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12502 352 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 288 12420 352 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12420 352 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 13240 271 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13240 271 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 13158 271 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13158 271 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 13076 271 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13076 271 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12994 271 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12994 271 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12912 271 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12912 271 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12830 271 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12830 271 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12748 271 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12748 271 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12666 271 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12666 271 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12584 271 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12584 271 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12502 271 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12502 271 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 254 12420 271 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12420 271 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13240 190 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13158 190 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13076 190 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12994 190 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12912 190 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12830 190 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12748 190 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12666 190 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12584 190 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12502 190 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12420 190 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 2 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 4 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 120 3558 4900 4486 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10151 3558 14931 4486 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12211 18573 14932 18592 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11966 18347 12211 18592 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11788 18169 11966 18347 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11530 17911 11788 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11283 17664 11530 17911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11027 17408 11283 17664 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10742 17123 11027 17408 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 16862 10742 17123 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10152 16533 10481 16862 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10152 13607 14932 16533 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2851 18190 3073 18342 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2854 17669 3250 18164 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2875 16598 3771 17628 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3283 17673 3505 17906 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3799 17162 4013 17403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3834 16589 4290 17118 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4330 16571 4554 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10497 16571 10721 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10761 16589 11217 17118 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11038 17162 11252 17403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11280 16598 12176 17628 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11546 17673 11768 17906 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11801 17669 12197 18164 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11978 18190 12200 18342 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4432 14913 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4346 14913 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4260 14913 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4174 14913 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4088 14913 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4002 14913 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3916 14913 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3830 14913 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3744 14913 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3658 14913 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3572 14913 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18539 14904 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18445 14916 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18363 14916 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18281 14916 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18199 14916 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18117 14916 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 18035 14916 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17953 14916 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17871 14916 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17789 14916 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17707 14916 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17625 14916 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17543 14916 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17461 14916 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17379 14916 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17297 14916 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17215 14916 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17133 14916 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 17051 14916 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16969 14916 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16887 14916 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16805 14916 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16723 14916 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16641 14916 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14852 16559 14916 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16472 14882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16391 14882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16310 14882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16229 14882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16148 14882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16067 14882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15986 14882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15905 14882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15824 14882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15743 14882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15662 14882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15581 14882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15500 14882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15419 14882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15338 14882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15257 14882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15176 14882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15095 14882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15014 14882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14933 14882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14852 14882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14771 14882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14690 14882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14609 14882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14527 14882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14445 14882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14363 14882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14281 14882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14199 14882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14117 14882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14035 14882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13953 14882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13871 14882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13789 14882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13707 14882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13625 14882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4432 14831 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4346 14831 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4260 14831 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4174 14831 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4088 14831 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4002 14831 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3916 14831 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3830 14831 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3744 14831 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3658 14831 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3572 14831 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18539 14822 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18445 14834 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18363 14834 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18281 14834 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18199 14834 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18117 14834 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 18035 14834 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17953 14834 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17871 14834 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17789 14834 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17707 14834 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17625 14834 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17543 14834 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17461 14834 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17379 14834 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17297 14834 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17215 14834 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17133 14834 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 17051 14834 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16969 14834 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16887 14834 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16805 14834 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16723 14834 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16641 14834 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14770 16559 14834 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16472 14802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16391 14802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16310 14802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16229 14802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16148 14802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16067 14802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15986 14802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15905 14802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15824 14802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15743 14802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15662 14802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15581 14802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15500 14802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15419 14802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15338 14802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15257 14802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15176 14802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15095 14802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15014 14802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14933 14802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14852 14802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14771 14802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14690 14802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14609 14802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14527 14802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14445 14802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14363 14802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14281 14802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14199 14802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14117 14802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14035 14802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13953 14802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13871 14802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13789 14802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13707 14802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13625 14802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4432 14749 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4346 14749 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4260 14749 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4174 14749 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4088 14749 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4002 14749 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3916 14749 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3830 14749 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3744 14749 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3658 14749 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3572 14749 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18539 14740 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18445 14746 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18445 14752 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18363 14746 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18363 14752 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18281 14746 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18281 14752 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18199 14746 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18199 14752 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18117 14746 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18117 14752 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 18035 14746 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 18035 14752 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17953 14746 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17953 14752 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17871 14746 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17871 14752 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17789 14746 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17789 14752 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17707 14746 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17707 14752 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17625 14746 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17625 14752 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17543 14746 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17543 14752 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17461 14746 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17461 14752 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17379 14746 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17379 14752 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17297 14746 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17297 14752 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17215 14746 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17215 14752 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17133 14746 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17133 14752 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 17051 14746 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 17051 14752 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16969 14746 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16969 14752 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16887 14746 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16887 14752 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16805 14746 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16805 14752 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16723 14746 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16723 14752 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16641 14746 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16641 14752 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14688 16559 14746 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14688 16559 14752 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16472 14722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16391 14722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16310 14722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16229 14722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16148 14722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16067 14722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15986 14722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15905 14722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15824 14722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15743 14722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15662 14722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15581 14722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15500 14722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15419 14722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15338 14722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15257 14722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15176 14722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15095 14722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15014 14722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14933 14722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14852 14722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14771 14722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14690 14722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14609 14722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14527 14722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14445 14722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14363 14722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14281 14722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14199 14722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14117 14722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14035 14722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13953 14722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13871 14722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13789 14722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13707 14722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13625 14722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4432 14667 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4346 14667 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4260 14667 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4174 14667 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4088 14667 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4002 14667 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3916 14667 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3830 14667 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3744 14667 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3658 14667 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3572 14667 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18539 14658 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18445 14670 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18445 14670 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18363 14670 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18363 14670 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18281 14670 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18281 14670 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18199 14670 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18199 14670 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18117 14670 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18117 14670 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 18035 14670 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 18035 14670 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17953 14670 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17953 14670 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17871 14670 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17871 14670 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17789 14670 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17789 14670 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17707 14670 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17707 14670 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17625 14670 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17625 14670 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17543 14670 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17543 14670 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17461 14670 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17461 14670 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17379 14670 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17379 14670 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17297 14670 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17297 14670 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17215 14670 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17215 14670 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17133 14670 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17133 14670 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 17051 14670 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 17051 14670 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16969 14670 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16969 14670 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16887 14670 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16887 14670 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16805 14670 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16805 14670 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16723 14670 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16723 14670 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16641 14670 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16641 14670 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14606 16559 14670 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14606 16559 14670 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16472 14642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16391 14642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16310 14642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16229 14642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16148 14642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16067 14642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15986 14642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15905 14642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15824 14642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15743 14642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15662 14642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15581 14642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15500 14642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15419 14642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15338 14642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15257 14642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15176 14642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15095 14642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15014 14642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14933 14642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14852 14642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14771 14642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14690 14642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14609 14642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14527 14642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14445 14642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14363 14642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14281 14642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14199 14642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14117 14642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14035 14642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13953 14642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13871 14642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13789 14642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13707 14642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13625 14642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4432 14585 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4346 14585 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4260 14585 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4174 14585 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4088 14585 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4002 14585 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3916 14585 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3830 14585 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3744 14585 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3658 14585 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3572 14585 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18539 14576 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18445 14588 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18445 14588 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18363 14588 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18363 14588 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18281 14588 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18281 14588 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18199 14588 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18199 14588 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18117 14588 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18117 14588 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 18035 14588 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 18035 14588 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17953 14588 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17953 14588 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17871 14588 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17871 14588 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17789 14588 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17789 14588 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17707 14588 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17707 14588 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17625 14588 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17625 14588 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17543 14588 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17543 14588 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17461 14588 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17461 14588 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17379 14588 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17379 14588 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17297 14588 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17297 14588 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17215 14588 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17215 14588 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17133 14588 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17133 14588 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 17051 14588 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 17051 14588 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16969 14588 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16969 14588 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16887 14588 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16887 14588 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16805 14588 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16805 14588 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16723 14588 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16723 14588 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16641 14588 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16641 14588 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14524 16559 14588 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14524 16559 14588 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16472 14562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16391 14562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16310 14562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16229 14562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16148 14562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16067 14562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15986 14562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15905 14562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15824 14562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15743 14562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15662 14562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15581 14562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15500 14562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15419 14562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15338 14562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15257 14562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15176 14562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15095 14562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15014 14562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14933 14562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14852 14562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14771 14562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14690 14562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14609 14562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14527 14562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14445 14562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14363 14562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14281 14562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14199 14562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14117 14562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14035 14562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13953 14562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13871 14562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13789 14562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13707 14562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13625 14562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4432 14503 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4346 14503 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4260 14503 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4174 14503 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4088 14503 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4002 14503 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3916 14503 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3830 14503 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3744 14503 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3658 14503 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3572 14503 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18539 14494 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18445 14506 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18445 14506 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18363 14506 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18363 14506 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18281 14506 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18281 14506 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18199 14506 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18199 14506 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18117 14506 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18117 14506 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 18035 14506 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 18035 14506 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17953 14506 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17953 14506 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17871 14506 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17871 14506 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17789 14506 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17789 14506 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17707 14506 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17707 14506 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17625 14506 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17625 14506 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17543 14506 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17543 14506 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17461 14506 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17461 14506 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17379 14506 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17379 14506 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17297 14506 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17297 14506 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17215 14506 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17215 14506 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17133 14506 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17133 14506 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 17051 14506 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 17051 14506 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16969 14506 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16969 14506 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16887 14506 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16887 14506 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16805 14506 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16805 14506 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16723 14506 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16723 14506 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16641 14506 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16641 14506 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14442 16559 14506 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16559 14506 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16472 14482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16391 14482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16310 14482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16229 14482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16148 14482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16067 14482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15986 14482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15905 14482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15824 14482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15743 14482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15662 14482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15581 14482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15500 14482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15419 14482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15338 14482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15257 14482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15176 14482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15095 14482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15014 14482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14933 14482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14852 14482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14771 14482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14690 14482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14609 14482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14527 14482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14445 14482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14363 14482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14281 14482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14199 14482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14117 14482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14035 14482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13953 14482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13871 14482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13789 14482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13707 14482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13625 14482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4432 14421 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4346 14421 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4260 14421 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4174 14421 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4088 14421 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4002 14421 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3916 14421 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3830 14421 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3744 14421 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3658 14421 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3572 14421 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18539 14412 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18445 14424 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18445 14424 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18363 14424 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18363 14424 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18281 14424 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18281 14424 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18199 14424 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18199 14424 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18117 14424 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18117 14424 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 18035 14424 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 18035 14424 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17953 14424 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17953 14424 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17871 14424 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17871 14424 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17789 14424 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17789 14424 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17707 14424 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17707 14424 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17625 14424 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17625 14424 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17543 14424 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17543 14424 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17461 14424 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17461 14424 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17379 14424 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17379 14424 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17297 14424 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17297 14424 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17215 14424 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17215 14424 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17133 14424 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17133 14424 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 17051 14424 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 17051 14424 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16969 14424 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16969 14424 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16887 14424 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16887 14424 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16805 14424 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16805 14424 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16723 14424 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16723 14424 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16641 14424 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16641 14424 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14360 16559 14424 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14360 16559 14424 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16472 14402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16391 14402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16310 14402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16229 14402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16148 14402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16067 14402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15986 14402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15905 14402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15824 14402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15743 14402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15662 14402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15581 14402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15500 14402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15419 14402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15338 14402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15257 14402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15176 14402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15095 14402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15014 14402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14933 14402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14852 14402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14771 14402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14690 14402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14609 14402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14527 14402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14445 14402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14363 14402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14281 14402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14199 14402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14117 14402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14035 14402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13953 14402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13871 14402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13789 14402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13707 14402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13625 14402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4432 14340 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4346 14340 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4260 14340 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4174 14340 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4088 14340 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4002 14340 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3916 14340 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3830 14340 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3744 14340 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3658 14340 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3572 14340 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18539 14330 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18445 14342 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18445 14342 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18363 14342 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18363 14342 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18281 14342 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18281 14342 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18199 14342 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18199 14342 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18117 14342 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18117 14342 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 18035 14342 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 18035 14342 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17953 14342 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17953 14342 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17871 14342 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17871 14342 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17789 14342 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17789 14342 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17707 14342 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17707 14342 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17625 14342 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17625 14342 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17543 14342 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17543 14342 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17461 14342 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17461 14342 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17379 14342 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17379 14342 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17297 14342 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17297 14342 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17215 14342 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17215 14342 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17133 14342 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17133 14342 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 17051 14342 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 17051 14342 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16969 14342 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16969 14342 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16887 14342 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16887 14342 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16805 14342 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16805 14342 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16723 14342 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16723 14342 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16641 14342 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16641 14342 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14278 16559 14342 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14278 16559 14342 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16472 14322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16391 14322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16310 14322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16229 14322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16148 14322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16067 14322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15986 14322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15905 14322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15824 14322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15743 14322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15662 14322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15581 14322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15500 14322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15419 14322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15338 14322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15257 14322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15176 14322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15095 14322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15014 14322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14933 14322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14852 14322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14771 14322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14690 14322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14609 14322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14527 14322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14445 14322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14363 14322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14281 14322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14199 14322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14117 14322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14035 14322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13953 14322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13871 14322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13789 14322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13707 14322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13625 14322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4432 14259 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4346 14259 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4260 14259 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4174 14259 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4088 14259 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4002 14259 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3916 14259 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3830 14259 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3744 14259 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3658 14259 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3572 14259 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18539 14248 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18445 14260 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18445 14260 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18363 14260 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18363 14260 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18281 14260 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18281 14260 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18199 14260 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18199 14260 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18117 14260 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18117 14260 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 18035 14260 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 18035 14260 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17953 14260 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17953 14260 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17871 14260 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17871 14260 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17789 14260 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17789 14260 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17707 14260 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17707 14260 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17625 14260 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17625 14260 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17543 14260 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17543 14260 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17461 14260 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17461 14260 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17379 14260 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17379 14260 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17297 14260 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17297 14260 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17215 14260 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17215 14260 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17133 14260 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17133 14260 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 17051 14260 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 17051 14260 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16969 14260 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16969 14260 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16887 14260 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16887 14260 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16805 14260 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16805 14260 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16723 14260 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16723 14260 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16641 14260 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16641 14260 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14196 16559 14260 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14196 16559 14260 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16472 14242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16391 14242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16310 14242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16229 14242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16148 14242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16067 14242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15986 14242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15905 14242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15824 14242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15743 14242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15662 14242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15581 14242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15500 14242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15419 14242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15338 14242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15257 14242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15176 14242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15095 14242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15014 14242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14933 14242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14852 14242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14771 14242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14690 14242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14609 14242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14527 14242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14445 14242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14363 14242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14281 14242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14199 14242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14117 14242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14035 14242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13953 14242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13871 14242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13789 14242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13707 14242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13625 14242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4432 14178 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4346 14178 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4260 14178 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4174 14178 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4088 14178 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4002 14178 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3916 14178 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3830 14178 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3744 14178 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3658 14178 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3572 14178 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18539 14166 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18445 14178 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18445 14178 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18363 14178 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18363 14178 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18281 14178 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18281 14178 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18199 14178 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18199 14178 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18117 14178 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18117 14178 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 18035 14178 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 18035 14178 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17953 14178 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17953 14178 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17871 14178 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17871 14178 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17789 14178 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17789 14178 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17707 14178 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17707 14178 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17625 14178 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17625 14178 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17543 14178 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17543 14178 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17461 14178 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17461 14178 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17379 14178 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17379 14178 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17297 14178 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17297 14178 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17215 14178 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17215 14178 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17133 14178 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17133 14178 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 17051 14178 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 17051 14178 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16969 14178 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16969 14178 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16887 14178 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16887 14178 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16805 14178 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16805 14178 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16723 14178 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16723 14178 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16641 14178 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16641 14178 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14114 16559 14178 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14114 16559 14178 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16472 14162 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16391 14162 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16310 14162 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16229 14162 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16148 14162 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16067 14162 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15986 14162 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15905 14162 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15824 14162 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15743 14162 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15662 14162 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15581 14162 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15500 14162 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15419 14162 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15338 14162 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15257 14162 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15176 14162 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15095 14162 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15014 14162 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14933 14162 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14852 14162 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14771 14162 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14690 14162 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14609 14162 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14527 14162 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14445 14162 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14363 14162 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14281 14162 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14199 14162 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14117 14162 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14035 14162 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13953 14162 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13871 14162 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13789 14162 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13707 14162 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13625 14162 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4432 14097 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4346 14097 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4260 14097 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4174 14097 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4088 14097 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4002 14097 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3916 14097 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3830 14097 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3744 14097 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3658 14097 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3572 14097 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18539 14084 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18445 14096 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18445 14096 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18363 14096 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18363 14096 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18281 14096 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18281 14096 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18199 14096 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18199 14096 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18117 14096 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18117 14096 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 18035 14096 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 18035 14096 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17953 14096 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17953 14096 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17871 14096 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17871 14096 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17789 14096 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17789 14096 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17707 14096 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17707 14096 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17625 14096 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17625 14096 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17543 14096 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17543 14096 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17461 14096 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17461 14096 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17379 14096 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17379 14096 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17297 14096 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17297 14096 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17215 14096 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17215 14096 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17133 14096 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17133 14096 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 17051 14096 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 17051 14096 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16969 14096 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16969 14096 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16887 14096 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16887 14096 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16805 14096 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16805 14096 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16723 14096 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16723 14096 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16641 14096 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16641 14096 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14032 16559 14096 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14032 16559 14096 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16472 14082 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16391 14082 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16310 14082 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16229 14082 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16148 14082 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16067 14082 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15986 14082 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15905 14082 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15824 14082 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15743 14082 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15662 14082 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15581 14082 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15500 14082 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15419 14082 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15338 14082 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15257 14082 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15176 14082 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15095 14082 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15014 14082 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14933 14082 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14852 14082 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14771 14082 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14690 14082 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14609 14082 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14527 14082 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14445 14082 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14363 14082 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14281 14082 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14199 14082 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14117 14082 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14035 14082 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13953 14082 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13871 14082 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13789 14082 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13707 14082 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13625 14082 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4432 14016 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4346 14016 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4260 14016 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4174 14016 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4088 14016 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4002 14016 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3916 14016 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3830 14016 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3744 14016 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3658 14016 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3572 14016 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18539 14002 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18445 14014 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18445 14014 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18363 14014 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18363 14014 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18281 14014 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18281 14014 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18199 14014 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18199 14014 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18117 14014 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18117 14014 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 18035 14014 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 18035 14014 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17953 14014 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17953 14014 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17871 14014 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17871 14014 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17789 14014 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17789 14014 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17707 14014 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17707 14014 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17625 14014 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17625 14014 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17543 14014 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17543 14014 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17461 14014 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17461 14014 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17379 14014 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17379 14014 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17297 14014 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17297 14014 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17215 14014 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17215 14014 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17133 14014 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17133 14014 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 17051 14014 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 17051 14014 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16969 14014 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16969 14014 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16887 14014 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16887 14014 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16805 14014 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16805 14014 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16723 14014 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16723 14014 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16641 14014 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16641 14014 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13950 16559 14014 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13950 16559 14014 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16472 14002 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16391 14002 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16310 14002 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16229 14002 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16148 14002 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16067 14002 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15986 14002 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15905 14002 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15824 14002 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15743 14002 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15662 14002 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15581 14002 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15500 14002 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15419 14002 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15338 14002 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15257 14002 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15176 14002 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15095 14002 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15014 14002 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14933 14002 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14852 14002 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14771 14002 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14690 14002 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14609 14002 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14527 14002 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14445 14002 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14363 14002 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14281 14002 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14199 14002 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14117 14002 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14035 14002 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13953 14002 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13871 14002 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13789 14002 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13707 14002 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13625 14002 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4432 13935 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4346 13935 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4260 13935 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4174 13935 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4088 13935 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4002 13935 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3916 13935 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3830 13935 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3744 13935 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3658 13935 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3572 13935 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16472 13922 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16391 13922 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16310 13922 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16229 13922 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16148 13922 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16067 13922 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15986 13922 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15905 13922 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15824 13922 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15743 13922 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15662 13922 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15581 13922 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15500 13922 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15419 13922 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15338 13922 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15257 13922 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15176 13922 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15095 13922 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15014 13922 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14933 13922 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14852 13922 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14771 13922 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14690 13922 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14609 13922 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14527 13922 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14445 13922 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14363 13922 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14281 13922 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14199 13922 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14117 13922 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14035 13922 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13953 13922 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13871 13922 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13789 13922 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13707 13922 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13625 13922 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18539 13920 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18445 13932 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18445 13932 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18363 13932 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18363 13932 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18281 13932 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18281 13932 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18199 13932 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18199 13932 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18117 13932 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18117 13932 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 18035 13932 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 18035 13932 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17953 13932 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17953 13932 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17871 13932 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17871 13932 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17789 13932 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17789 13932 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17707 13932 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17707 13932 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17625 13932 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17625 13932 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17543 13932 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17543 13932 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17461 13932 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17461 13932 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17379 13932 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17379 13932 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17297 13932 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17297 13932 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17215 13932 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17215 13932 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17133 13932 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17133 13932 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 17051 13932 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 17051 13932 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16969 13932 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16969 13932 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16887 13932 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16887 13932 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16805 13932 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16805 13932 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16723 13932 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16723 13932 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16641 13932 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16641 13932 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13868 16559 13932 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13868 16559 13932 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4432 13854 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4346 13854 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4260 13854 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4174 13854 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4088 13854 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4002 13854 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3916 13854 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3830 13854 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3744 13854 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3658 13854 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3572 13854 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16472 13842 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16391 13842 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16310 13842 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16229 13842 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16148 13842 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16067 13842 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15986 13842 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15905 13842 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15824 13842 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15743 13842 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15662 13842 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15581 13842 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15500 13842 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15419 13842 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15338 13842 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15257 13842 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15176 13842 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15095 13842 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15014 13842 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14933 13842 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14852 13842 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14771 13842 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14690 13842 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14609 13842 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14527 13842 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14445 13842 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14363 13842 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14281 13842 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14199 13842 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14117 13842 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14035 13842 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13953 13842 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13871 13842 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13789 13842 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13707 13842 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13625 13842 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18539 13838 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18445 13850 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18445 13850 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18363 13850 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18363 13850 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18281 13850 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18281 13850 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18199 13850 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18199 13850 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18117 13850 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18117 13850 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 18035 13850 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 18035 13850 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17953 13850 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17953 13850 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17871 13850 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17871 13850 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17789 13850 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17789 13850 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17707 13850 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17707 13850 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17625 13850 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17625 13850 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17543 13850 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17543 13850 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17461 13850 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17461 13850 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17379 13850 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17379 13850 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17297 13850 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17297 13850 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17215 13850 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17215 13850 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17133 13850 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17133 13850 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 17051 13850 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 17051 13850 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16969 13850 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16969 13850 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16887 13850 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16887 13850 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16805 13850 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16805 13850 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16723 13850 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16723 13850 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16641 13850 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16641 13850 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13786 16559 13850 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13786 16559 13850 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4432 13773 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4346 13773 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4260 13773 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4174 13773 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4088 13773 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4002 13773 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3916 13773 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3830 13773 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3744 13773 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3658 13773 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3572 13773 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16472 13762 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16391 13762 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16310 13762 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16229 13762 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16148 13762 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16067 13762 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15986 13762 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15905 13762 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15824 13762 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15743 13762 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15662 13762 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15581 13762 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15500 13762 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15419 13762 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15338 13762 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15257 13762 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15176 13762 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15095 13762 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15014 13762 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14933 13762 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14852 13762 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14771 13762 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14690 13762 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14609 13762 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14527 13762 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14445 13762 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14363 13762 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14281 13762 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14199 13762 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14117 13762 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14035 13762 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13953 13762 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13871 13762 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13789 13762 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13707 13762 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13625 13762 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18539 13756 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18445 13768 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18445 13768 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18363 13768 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18363 13768 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18281 13768 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18281 13768 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18199 13768 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18199 13768 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18117 13768 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18117 13768 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 18035 13768 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 18035 13768 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17953 13768 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17953 13768 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17871 13768 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17871 13768 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17789 13768 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17789 13768 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17707 13768 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17707 13768 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17625 13768 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17625 13768 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17543 13768 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17543 13768 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17461 13768 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17461 13768 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17379 13768 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17379 13768 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17297 13768 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17297 13768 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17215 13768 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17215 13768 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17133 13768 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17133 13768 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 17051 13768 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 17051 13768 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16969 13768 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16969 13768 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16887 13768 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16887 13768 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16805 13768 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16805 13768 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16723 13768 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16723 13768 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16641 13768 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16641 13768 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13704 16559 13768 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13704 16559 13768 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4432 13692 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4346 13692 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4260 13692 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4174 13692 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4088 13692 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4002 13692 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3916 13692 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3830 13692 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3744 13692 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3658 13692 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3572 13692 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16472 13682 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16391 13682 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16310 13682 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16229 13682 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16148 13682 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16067 13682 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15986 13682 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15905 13682 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15824 13682 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15743 13682 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15662 13682 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15581 13682 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15500 13682 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15419 13682 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15338 13682 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15257 13682 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15176 13682 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15095 13682 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15014 13682 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14933 13682 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14852 13682 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14771 13682 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14690 13682 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14609 13682 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14527 13682 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14445 13682 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14363 13682 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14281 13682 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14199 13682 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14117 13682 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14035 13682 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13953 13682 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13871 13682 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13789 13682 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13707 13682 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13625 13682 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18539 13674 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18445 13686 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18445 13686 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18363 13686 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18363 13686 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18281 13686 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18281 13686 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18199 13686 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18199 13686 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18117 13686 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18117 13686 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 18035 13686 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 18035 13686 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17953 13686 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17953 13686 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17871 13686 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17871 13686 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17789 13686 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17789 13686 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17707 13686 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17707 13686 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17625 13686 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17625 13686 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17543 13686 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17543 13686 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17461 13686 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17461 13686 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17379 13686 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17379 13686 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17297 13686 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17297 13686 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17215 13686 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17215 13686 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17133 13686 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17133 13686 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 17051 13686 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 17051 13686 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16969 13686 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16969 13686 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16887 13686 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16887 13686 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16805 13686 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16805 13686 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16723 13686 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16723 13686 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16641 13686 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16641 13686 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13622 16559 13686 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13622 16559 13686 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4432 13611 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4346 13611 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4260 13611 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4174 13611 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4088 13611 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4002 13611 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3916 13611 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3830 13611 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3744 13611 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3658 13611 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3572 13611 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16472 13602 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16391 13602 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16310 13602 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16229 13602 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16148 13602 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16067 13602 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15986 13602 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15905 13602 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15824 13602 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15743 13602 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15662 13602 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15581 13602 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15500 13602 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15419 13602 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15338 13602 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15257 13602 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15176 13602 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15095 13602 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15014 13602 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14933 13602 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14852 13602 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14771 13602 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14690 13602 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14609 13602 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14527 13602 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14445 13602 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14363 13602 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14281 13602 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14199 13602 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14117 13602 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14035 13602 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13953 13602 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13871 13602 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13789 13602 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13707 13602 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13625 13602 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18539 13592 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18445 13604 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18445 13604 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18363 13604 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18363 13604 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18281 13604 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18281 13604 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18199 13604 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18199 13604 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18117 13604 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18117 13604 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 18035 13604 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 18035 13604 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17953 13604 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17953 13604 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17871 13604 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17871 13604 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17789 13604 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17789 13604 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17707 13604 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17707 13604 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17625 13604 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17625 13604 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17543 13604 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17543 13604 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17461 13604 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17461 13604 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17379 13604 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17379 13604 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17297 13604 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17297 13604 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17215 13604 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17215 13604 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17133 13604 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17133 13604 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 17051 13604 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 17051 13604 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16969 13604 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16969 13604 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16887 13604 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16887 13604 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16805 13604 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16805 13604 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16723 13604 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16723 13604 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16641 13604 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16641 13604 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13540 16559 13604 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13540 16559 13604 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4432 13530 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4346 13530 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4260 13530 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4174 13530 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4088 13530 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4002 13530 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3916 13530 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3830 13530 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3744 13530 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3658 13530 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3572 13530 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16472 13522 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16391 13522 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16310 13522 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16229 13522 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16148 13522 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16067 13522 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15986 13522 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15905 13522 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15824 13522 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15743 13522 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15662 13522 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15581 13522 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15500 13522 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15419 13522 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15338 13522 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15257 13522 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15176 13522 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15095 13522 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15014 13522 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14933 13522 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14852 13522 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14771 13522 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14690 13522 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14609 13522 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14527 13522 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14445 13522 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14363 13522 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14281 13522 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14199 13522 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14117 13522 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14035 13522 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13953 13522 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13871 13522 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13789 13522 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13707 13522 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13625 13522 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18539 13510 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18445 13522 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18445 13522 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18363 13522 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18363 13522 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18281 13522 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18281 13522 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18199 13522 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18199 13522 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18117 13522 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18117 13522 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 18035 13522 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 18035 13522 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17953 13522 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17953 13522 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17871 13522 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17871 13522 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17789 13522 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17789 13522 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17707 13522 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17707 13522 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17625 13522 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17625 13522 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17543 13522 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17543 13522 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17461 13522 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17461 13522 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17379 13522 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17379 13522 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17297 13522 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17297 13522 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17215 13522 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17215 13522 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17133 13522 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17133 13522 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 17051 13522 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 17051 13522 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16969 13522 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16969 13522 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16887 13522 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16887 13522 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16805 13522 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16805 13522 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16723 13522 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16723 13522 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16641 13522 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16641 13522 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13458 16559 13522 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13458 16559 13522 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4432 13449 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4346 13449 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4260 13449 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4174 13449 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4088 13449 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4002 13449 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3916 13449 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3830 13449 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3744 13449 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3658 13449 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3572 13449 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16472 13442 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16391 13442 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16310 13442 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16229 13442 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16148 13442 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16067 13442 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15986 13442 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15905 13442 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15824 13442 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15743 13442 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15662 13442 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15581 13442 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15500 13442 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15419 13442 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15338 13442 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15257 13442 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15176 13442 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15095 13442 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15014 13442 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14933 13442 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14852 13442 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14771 13442 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14690 13442 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14609 13442 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14527 13442 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14445 13442 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14363 13442 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14281 13442 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14199 13442 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14117 13442 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14035 13442 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13953 13442 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13871 13442 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13789 13442 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13707 13442 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13625 13442 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18539 13428 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18445 13440 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18445 13440 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18363 13440 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18363 13440 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18281 13440 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18281 13440 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18199 13440 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18199 13440 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18117 13440 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18117 13440 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 18035 13440 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 18035 13440 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17953 13440 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17953 13440 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17871 13440 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17871 13440 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17789 13440 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17789 13440 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17707 13440 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17707 13440 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17625 13440 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17625 13440 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17543 13440 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17543 13440 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17461 13440 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17461 13440 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17379 13440 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17379 13440 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17297 13440 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17297 13440 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17215 13440 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17215 13440 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17133 13440 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17133 13440 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 17051 13440 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 17051 13440 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16969 13440 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16969 13440 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16887 13440 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16887 13440 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16805 13440 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16805 13440 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16723 13440 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16723 13440 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16641 13440 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16641 13440 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13376 16559 13440 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13376 16559 13440 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4432 13368 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4346 13368 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4260 13368 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4174 13368 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4088 13368 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4002 13368 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3916 13368 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3830 13368 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3744 13368 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3658 13368 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3572 13368 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16472 13362 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16391 13362 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16310 13362 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16229 13362 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16148 13362 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16067 13362 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15986 13362 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15905 13362 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15824 13362 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15743 13362 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15662 13362 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15581 13362 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15500 13362 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15419 13362 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15338 13362 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15257 13362 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15176 13362 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15095 13362 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15014 13362 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14933 13362 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14852 13362 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14771 13362 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14690 13362 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14609 13362 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14527 13362 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14445 13362 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14363 13362 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14281 13362 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14199 13362 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14117 13362 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14035 13362 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13953 13362 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13871 13362 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13789 13362 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13707 13362 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13625 13362 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18539 13346 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18445 13358 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18445 13358 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18363 13358 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18363 13358 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18281 13358 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18281 13358 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18199 13358 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18199 13358 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18117 13358 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18117 13358 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 18035 13358 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 18035 13358 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17953 13358 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17953 13358 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17871 13358 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17871 13358 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17789 13358 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17789 13358 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17707 13358 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17707 13358 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17625 13358 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17625 13358 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17543 13358 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17543 13358 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17461 13358 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17461 13358 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17379 13358 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17379 13358 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17297 13358 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17297 13358 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17215 13358 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17215 13358 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17133 13358 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17133 13358 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 17051 13358 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 17051 13358 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16969 13358 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16969 13358 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16887 13358 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16887 13358 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16805 13358 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16805 13358 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16723 13358 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16723 13358 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16641 13358 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16641 13358 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13294 16559 13358 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13294 16559 13358 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4432 13287 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4346 13287 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4260 13287 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4174 13287 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4088 13287 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4002 13287 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3916 13287 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3830 13287 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3744 13287 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3658 13287 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3572 13287 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16472 13282 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16391 13282 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16310 13282 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16229 13282 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16148 13282 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16067 13282 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15986 13282 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15905 13282 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15824 13282 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15743 13282 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15662 13282 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15581 13282 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15500 13282 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15419 13282 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15338 13282 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15257 13282 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15176 13282 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15095 13282 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15014 13282 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14933 13282 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14852 13282 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14771 13282 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14690 13282 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14609 13282 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14527 13282 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14445 13282 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14363 13282 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14281 13282 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14199 13282 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14117 13282 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14035 13282 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13953 13282 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13871 13282 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13789 13282 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13707 13282 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13625 13282 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18539 13264 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18445 13276 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18445 13276 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18363 13276 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18363 13276 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18281 13276 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18281 13276 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18199 13276 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18199 13276 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18117 13276 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18117 13276 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 18035 13276 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 18035 13276 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17953 13276 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17953 13276 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17871 13276 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17871 13276 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17789 13276 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17789 13276 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17707 13276 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17707 13276 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17625 13276 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17625 13276 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17543 13276 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17543 13276 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17461 13276 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17461 13276 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17379 13276 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17379 13276 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17297 13276 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17297 13276 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17215 13276 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17215 13276 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17133 13276 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17133 13276 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 17051 13276 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 17051 13276 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16969 13276 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16969 13276 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16887 13276 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16887 13276 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16805 13276 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16805 13276 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16723 13276 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16723 13276 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16641 13276 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16641 13276 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13212 16559 13276 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13212 16559 13276 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4432 13206 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4346 13206 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4260 13206 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4174 13206 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4088 13206 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4002 13206 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3916 13206 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3830 13206 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3744 13206 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3658 13206 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3572 13206 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16472 13202 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16391 13202 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16310 13202 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16229 13202 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16148 13202 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16067 13202 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15986 13202 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15905 13202 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15824 13202 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15743 13202 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15662 13202 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15581 13202 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15500 13202 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15419 13202 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15338 13202 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15257 13202 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15176 13202 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15095 13202 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15014 13202 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14933 13202 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14852 13202 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14771 13202 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14690 13202 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14609 13202 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14527 13202 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14445 13202 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14363 13202 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14281 13202 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14199 13202 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14117 13202 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14035 13202 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13953 13202 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13871 13202 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13789 13202 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13707 13202 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13625 13202 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18539 13182 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18445 13194 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18445 13194 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18363 13194 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18363 13194 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18281 13194 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18281 13194 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18199 13194 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18199 13194 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18117 13194 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18117 13194 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 18035 13194 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 18035 13194 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17953 13194 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17953 13194 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17871 13194 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17871 13194 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17789 13194 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17789 13194 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17707 13194 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17707 13194 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17625 13194 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17625 13194 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17543 13194 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17543 13194 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17461 13194 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17461 13194 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17379 13194 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17379 13194 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17297 13194 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17297 13194 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17215 13194 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17215 13194 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17133 13194 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17133 13194 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 17051 13194 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 17051 13194 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16969 13194 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16969 13194 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16887 13194 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16887 13194 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16805 13194 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16805 13194 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16723 13194 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16723 13194 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16641 13194 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16641 13194 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13130 16559 13194 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13130 16559 13194 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4432 13125 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4346 13125 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4260 13125 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4174 13125 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4088 13125 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4002 13125 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3916 13125 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3830 13125 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3744 13125 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3658 13125 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3572 13125 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16472 13122 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16391 13122 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16310 13122 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16229 13122 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16148 13122 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16067 13122 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15986 13122 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15905 13122 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15824 13122 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15743 13122 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15662 13122 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15581 13122 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15500 13122 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15419 13122 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15338 13122 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15257 13122 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15176 13122 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15095 13122 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15014 13122 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14933 13122 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14852 13122 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14771 13122 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14690 13122 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14609 13122 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14527 13122 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14445 13122 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14363 13122 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14281 13122 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14199 13122 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14117 13122 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14035 13122 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13953 13122 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13871 13122 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13789 13122 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13707 13122 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13625 13122 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18539 13100 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18445 13112 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18445 13112 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18363 13112 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18363 13112 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18281 13112 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18281 13112 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18199 13112 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18199 13112 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18117 13112 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18117 13112 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 18035 13112 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 18035 13112 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17953 13112 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17953 13112 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17871 13112 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17871 13112 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17789 13112 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17789 13112 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17707 13112 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17707 13112 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17625 13112 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17625 13112 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17543 13112 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17543 13112 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17461 13112 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17461 13112 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17379 13112 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17379 13112 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17297 13112 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17297 13112 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17215 13112 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17215 13112 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17133 13112 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17133 13112 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 17051 13112 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 17051 13112 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16969 13112 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16969 13112 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16887 13112 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16887 13112 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16805 13112 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16805 13112 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16723 13112 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16723 13112 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16641 13112 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16641 13112 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 13048 16559 13112 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13048 16559 13112 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4432 13044 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4346 13044 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4260 13044 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4174 13044 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4088 13044 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4002 13044 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3916 13044 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3830 13044 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3744 13044 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3658 13044 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3572 13044 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16472 13042 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16391 13042 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16310 13042 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16229 13042 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16148 13042 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16067 13042 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15986 13042 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15905 13042 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15824 13042 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15743 13042 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15662 13042 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15581 13042 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15500 13042 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15419 13042 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15338 13042 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15257 13042 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15176 13042 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15095 13042 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15014 13042 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14933 13042 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14852 13042 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14771 13042 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14690 13042 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14609 13042 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14527 13042 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14445 13042 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14363 13042 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14281 13042 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14199 13042 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14117 13042 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14035 13042 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13953 13042 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13871 13042 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13789 13042 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13707 13042 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13625 13042 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18539 13018 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18445 13030 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18445 13030 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18363 13030 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18363 13030 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18281 13030 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18281 13030 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18199 13030 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18199 13030 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18117 13030 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18117 13030 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 18035 13030 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 18035 13030 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17953 13030 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17953 13030 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17871 13030 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17871 13030 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17789 13030 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17789 13030 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17707 13030 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17707 13030 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17625 13030 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17625 13030 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17543 13030 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17543 13030 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17461 13030 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17461 13030 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17379 13030 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17379 13030 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17297 13030 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17297 13030 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17215 13030 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17215 13030 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17133 13030 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17133 13030 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 17051 13030 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 17051 13030 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16969 13030 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16969 13030 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16887 13030 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16887 13030 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16805 13030 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16805 13030 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16723 13030 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16723 13030 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16641 13030 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16641 13030 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12966 16559 13030 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12966 16559 13030 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4432 12963 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4346 12963 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4260 12963 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4174 12963 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4088 12963 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4002 12963 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3916 12963 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3830 12963 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3744 12963 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3658 12963 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3572 12963 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16472 12962 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16391 12962 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16310 12962 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16229 12962 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16148 12962 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16067 12962 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15986 12962 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15905 12962 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15824 12962 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15743 12962 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15662 12962 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15581 12962 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15500 12962 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15419 12962 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15338 12962 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15257 12962 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15176 12962 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15095 12962 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15014 12962 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14933 12962 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14852 12962 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14771 12962 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14690 12962 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14609 12962 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14527 12962 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14445 12962 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14363 12962 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14281 12962 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14199 12962 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14117 12962 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14035 12962 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13953 12962 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13871 12962 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13789 12962 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13707 12962 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13625 12962 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18539 12936 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18445 12948 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18445 12948 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18363 12948 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18363 12948 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18281 12948 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18281 12948 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18199 12948 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18199 12948 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18117 12948 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18117 12948 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 18035 12948 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 18035 12948 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17953 12948 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17953 12948 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17871 12948 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17871 12948 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17789 12948 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17789 12948 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17707 12948 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17707 12948 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17625 12948 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17625 12948 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17543 12948 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17543 12948 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17461 12948 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17461 12948 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17379 12948 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17379 12948 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17297 12948 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17297 12948 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17215 12948 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17215 12948 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17133 12948 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17133 12948 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 17051 12948 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 17051 12948 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16969 12948 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16969 12948 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16887 12948 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16887 12948 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16805 12948 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16805 12948 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16723 12948 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16723 12948 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16641 12948 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16641 12948 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12884 16559 12948 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12884 16559 12948 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16472 12882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16391 12882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16310 12882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16229 12882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16148 12882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16067 12882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15986 12882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15905 12882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15824 12882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15743 12882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15662 12882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15581 12882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15500 12882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15419 12882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15338 12882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15257 12882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15176 12882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15095 12882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15014 12882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14933 12882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14852 12882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14771 12882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14690 12882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14609 12882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14527 12882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14445 12882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14363 12882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14281 12882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14199 12882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14117 12882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14035 12882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13953 12882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13871 12882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13789 12882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13707 12882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13625 12882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4432 12882 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4346 12882 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4260 12882 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4174 12882 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4088 12882 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4002 12882 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3916 12882 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3830 12882 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3744 12882 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3658 12882 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3572 12882 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18539 12854 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18445 12866 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18445 12866 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18363 12866 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18363 12866 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18281 12866 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18281 12866 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18199 12866 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18199 12866 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18117 12866 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18117 12866 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 18035 12866 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 18035 12866 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17953 12866 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17953 12866 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17871 12866 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17871 12866 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17789 12866 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17789 12866 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17707 12866 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17707 12866 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17625 12866 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17625 12866 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17543 12866 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17543 12866 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17461 12866 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17461 12866 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17379 12866 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17379 12866 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17297 12866 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17297 12866 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17215 12866 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17215 12866 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17133 12866 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17133 12866 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 17051 12866 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 17051 12866 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16969 12866 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16969 12866 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16887 12866 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16887 12866 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16805 12866 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16805 12866 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16723 12866 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16723 12866 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16641 12866 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16641 12866 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12802 16559 12866 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12802 16559 12866 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16472 12802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16391 12802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16310 12802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16229 12802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16148 12802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16067 12802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15986 12802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15905 12802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15824 12802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15743 12802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15662 12802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15581 12802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15500 12802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15419 12802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15338 12802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15257 12802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15176 12802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15095 12802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15014 12802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14933 12802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14852 12802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14771 12802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14690 12802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14609 12802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14527 12802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14445 12802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14363 12802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14281 12802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14199 12802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14117 12802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14035 12802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13953 12802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13871 12802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13789 12802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13707 12802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13625 12802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4432 12801 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4346 12801 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4260 12801 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4174 12801 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4088 12801 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4002 12801 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3916 12801 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3830 12801 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3744 12801 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3658 12801 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3572 12801 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18539 12772 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18445 12784 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18445 12784 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18363 12784 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18363 12784 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18281 12784 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18281 12784 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18199 12784 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18199 12784 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18117 12784 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18117 12784 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 18035 12784 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 18035 12784 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17953 12784 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17953 12784 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17871 12784 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17871 12784 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17789 12784 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17789 12784 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17707 12784 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17707 12784 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17625 12784 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17625 12784 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17543 12784 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17543 12784 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17461 12784 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17461 12784 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17379 12784 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17379 12784 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17297 12784 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17297 12784 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17215 12784 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17215 12784 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17133 12784 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17133 12784 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 17051 12784 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 17051 12784 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16969 12784 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16969 12784 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16887 12784 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16887 12784 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16805 12784 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16805 12784 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16723 12784 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16723 12784 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16641 12784 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16641 12784 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12720 16559 12784 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12720 16559 12784 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16472 12722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16391 12722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16310 12722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16229 12722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16148 12722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16067 12722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15986 12722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15905 12722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15824 12722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15743 12722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15662 12722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15581 12722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15500 12722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15419 12722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15338 12722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15257 12722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15176 12722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15095 12722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15014 12722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14933 12722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14852 12722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14771 12722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14690 12722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14609 12722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14527 12722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14445 12722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14363 12722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14281 12722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14199 12722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14117 12722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14035 12722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13953 12722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13871 12722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13789 12722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13707 12722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13625 12722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4432 12720 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4346 12720 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4260 12720 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4174 12720 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4088 12720 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4002 12720 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3916 12720 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3830 12720 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3744 12720 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3658 12720 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3572 12720 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18539 12690 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18445 12702 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18445 12702 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18363 12702 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18363 12702 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18281 12702 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18281 12702 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18199 12702 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18199 12702 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18117 12702 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18117 12702 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 18035 12702 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 18035 12702 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17953 12702 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17953 12702 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17871 12702 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17871 12702 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17789 12702 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17789 12702 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17707 12702 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17707 12702 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17625 12702 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17625 12702 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17543 12702 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17543 12702 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17461 12702 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17461 12702 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17379 12702 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17379 12702 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17297 12702 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17297 12702 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17215 12702 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17215 12702 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17133 12702 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17133 12702 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 17051 12702 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 17051 12702 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16969 12702 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16969 12702 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16887 12702 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16887 12702 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16805 12702 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16805 12702 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16723 12702 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16723 12702 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16641 12702 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16641 12702 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12638 16559 12702 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12638 16559 12702 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16472 12642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16391 12642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16310 12642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16229 12642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16148 12642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16067 12642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15986 12642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15905 12642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15824 12642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15743 12642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15662 12642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15581 12642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15500 12642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15419 12642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15338 12642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15257 12642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15176 12642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15095 12642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15014 12642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14933 12642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14852 12642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14771 12642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14690 12642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14609 12642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14527 12642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14445 12642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14363 12642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14281 12642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14199 12642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14117 12642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14035 12642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13953 12642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13871 12642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13789 12642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13707 12642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13625 12642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4432 12639 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4346 12639 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4260 12639 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4174 12639 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4088 12639 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4002 12639 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3916 12639 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3830 12639 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3744 12639 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3658 12639 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3572 12639 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18539 12608 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18445 12620 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18445 12620 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18363 12620 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18363 12620 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18281 12620 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18281 12620 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18199 12620 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18199 12620 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18117 12620 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18117 12620 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 18035 12620 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 18035 12620 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17953 12620 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17953 12620 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17871 12620 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17871 12620 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17789 12620 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17789 12620 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17707 12620 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17707 12620 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17625 12620 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17625 12620 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17543 12620 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17543 12620 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17461 12620 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17461 12620 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17379 12620 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17379 12620 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17297 12620 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17297 12620 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17215 12620 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17215 12620 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17133 12620 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17133 12620 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 17051 12620 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 17051 12620 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16969 12620 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16969 12620 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16887 12620 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16887 12620 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16805 12620 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16805 12620 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16723 12620 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16723 12620 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16641 12620 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16641 12620 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12556 16559 12620 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12556 16559 12620 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16472 12562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16391 12562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16310 12562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16229 12562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16148 12562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16067 12562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15986 12562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15905 12562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15824 12562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15743 12562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15662 12562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15581 12562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15500 12562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15419 12562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15338 12562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15257 12562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15176 12562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15095 12562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15014 12562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14933 12562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14852 12562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14771 12562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14690 12562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14609 12562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14527 12562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14445 12562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14363 12562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14281 12562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14199 12562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14117 12562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14035 12562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13953 12562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13871 12562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13789 12562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13707 12562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13625 12562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4432 12558 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4346 12558 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4260 12558 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4174 12558 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4088 12558 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4002 12558 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3916 12558 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3830 12558 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3744 12558 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3658 12558 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3572 12558 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18539 12526 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18445 12538 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18445 12538 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18363 12538 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18363 12538 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18281 12538 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18281 12538 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18199 12538 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18199 12538 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18117 12538 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18117 12538 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 18035 12538 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 18035 12538 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17953 12538 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17953 12538 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17871 12538 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17871 12538 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17789 12538 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17789 12538 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17707 12538 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17707 12538 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17625 12538 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17625 12538 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17543 12538 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17543 12538 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17461 12538 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17461 12538 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17379 12538 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17379 12538 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17297 12538 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17297 12538 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17215 12538 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17215 12538 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17133 12538 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17133 12538 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 17051 12538 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 17051 12538 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16969 12538 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16969 12538 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16887 12538 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16887 12538 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16805 12538 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16805 12538 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16723 12538 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16723 12538 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16641 12538 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16641 12538 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12474 16559 12538 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12474 16559 12538 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16472 12482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16391 12482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16310 12482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16229 12482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16148 12482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16067 12482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15986 12482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15905 12482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15824 12482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15743 12482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15662 12482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15581 12482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15500 12482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15419 12482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15338 12482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15257 12482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15176 12482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15095 12482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15014 12482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14933 12482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14852 12482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14771 12482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14690 12482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14609 12482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14527 12482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14445 12482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14363 12482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14281 12482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14199 12482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14117 12482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14035 12482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13953 12482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13871 12482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13789 12482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13707 12482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13625 12482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4432 12477 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4346 12477 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4260 12477 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4174 12477 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4088 12477 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4002 12477 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3916 12477 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3830 12477 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3744 12477 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3658 12477 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3572 12477 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18539 12445 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18445 12457 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18445 12457 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18363 12457 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18363 12457 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18281 12457 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18281 12457 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18199 12457 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18199 12457 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18117 12457 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18117 12457 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 18035 12457 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 18035 12457 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17953 12457 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17953 12457 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17871 12457 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17871 12457 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17789 12457 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17789 12457 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17707 12457 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17707 12457 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17625 12457 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17625 12457 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17543 12457 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17543 12457 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17461 12457 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17461 12457 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17379 12457 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17379 12457 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17297 12457 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17297 12457 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17215 12457 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17215 12457 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17133 12457 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17133 12457 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 17051 12457 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 17051 12457 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16969 12457 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16969 12457 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16887 12457 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16887 12457 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16805 12457 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16805 12457 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16723 12457 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16723 12457 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16641 12457 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16641 12457 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12393 16559 12457 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12393 16559 12457 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16472 12402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16391 12402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16310 12402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16229 12402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16148 12402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16067 12402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15986 12402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15905 12402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15824 12402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15743 12402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15662 12402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15581 12402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15500 12402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15419 12402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15338 12402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15257 12402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15176 12402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15095 12402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15014 12402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14933 12402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14852 12402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14771 12402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14690 12402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14609 12402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14527 12402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14445 12402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14363 12402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14281 12402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14199 12402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14117 12402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14035 12402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13953 12402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13871 12402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13789 12402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13707 12402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13625 12402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4432 12396 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4346 12396 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4260 12396 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4174 12396 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4088 12396 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4002 12396 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3916 12396 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3830 12396 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3744 12396 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3658 12396 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3572 12396 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18539 12364 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18445 12376 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18445 12376 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18363 12376 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18363 12376 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18281 12376 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18281 12376 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18199 12376 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18199 12376 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18117 12376 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18117 12376 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 18035 12376 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 18035 12376 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17953 12376 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17953 12376 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17871 12376 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17871 12376 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17789 12376 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17789 12376 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17707 12376 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17707 12376 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17625 12376 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17625 12376 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17543 12376 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17543 12376 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17461 12376 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17461 12376 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17379 12376 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17379 12376 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17297 12376 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17297 12376 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17215 12376 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17215 12376 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17133 12376 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17133 12376 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 17051 12376 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 17051 12376 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16969 12376 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16969 12376 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16887 12376 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16887 12376 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16805 12376 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16805 12376 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16723 12376 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16723 12376 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16641 12376 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16641 12376 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12312 16559 12376 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12312 16559 12376 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16472 12322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16391 12322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16310 12322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16229 12322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16148 12322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16067 12322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15986 12322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15905 12322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15824 12322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15743 12322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15662 12322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15581 12322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15500 12322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15419 12322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15338 12322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15257 12322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15176 12322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15095 12322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15014 12322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14933 12322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14852 12322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14771 12322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14690 12322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14609 12322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14527 12322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14445 12322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14363 12322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14281 12322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14199 12322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14117 12322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14035 12322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13953 12322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13871 12322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13789 12322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13707 12322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13625 12322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4432 12315 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4346 12315 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4260 12315 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4174 12315 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4088 12315 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4002 12315 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3916 12315 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3830 12315 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3744 12315 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3658 12315 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3572 12315 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18539 12283 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18445 12295 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18445 12295 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18363 12295 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18363 12295 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18281 12295 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18281 12295 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18199 12295 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18199 12295 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18117 12295 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18117 12295 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 18035 12295 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 18035 12295 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17953 12295 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17953 12295 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17871 12295 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17871 12295 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17789 12295 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17789 12295 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17707 12295 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17707 12295 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17625 12295 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17625 12295 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17543 12295 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17543 12295 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17461 12295 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17461 12295 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17379 12295 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17379 12295 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17297 12295 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17297 12295 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17215 12295 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17215 12295 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17133 12295 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17133 12295 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 17051 12295 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 17051 12295 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16969 12295 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16969 12295 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16887 12295 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16887 12295 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16805 12295 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16805 12295 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16723 12295 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16723 12295 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16641 12295 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16641 12295 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12231 16559 12295 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12231 16559 12295 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16472 12242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16391 12242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16310 12242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16229 12242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16148 12242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16067 12242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15986 12242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15905 12242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15824 12242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15743 12242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15662 12242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15581 12242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15500 12242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15419 12242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15338 12242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15257 12242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15176 12242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15095 12242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15014 12242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14933 12242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14852 12242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14771 12242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14690 12242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14609 12242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14527 12242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14445 12242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14363 12242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14281 12242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14199 12242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14117 12242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14035 12242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13953 12242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13871 12242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13789 12242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13707 12242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13625 12242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4432 12234 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4346 12234 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4260 12234 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4174 12234 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4088 12234 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4002 12234 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3916 12234 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3830 12234 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3744 12234 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3658 12234 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3572 12234 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12135 18277 12199 18341 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12135 18191 12199 18255 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 18099 12195 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 18013 12195 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17927 12195 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17841 12195 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17755 12195 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12131 17670 12195 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16472 12162 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16391 12162 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16310 12162 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16229 12162 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16148 12162 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16067 12162 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15986 12162 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15905 12162 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15824 12162 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15743 12162 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15662 12162 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15581 12162 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15500 12162 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15419 12162 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15338 12162 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15257 12162 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15176 12162 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15095 12162 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15014 12162 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14933 12162 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14852 12162 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14771 12162 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14690 12162 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14609 12162 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14527 12162 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14445 12162 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14363 12162 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14281 12162 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14199 12162 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14117 12162 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14035 12162 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13953 12162 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13871 12162 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13789 12162 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13707 12162 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13625 12162 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17563 12170 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17482 12170 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17401 12170 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17320 12170 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17239 12170 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17159 12170 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 17079 12170 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16999 12170 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16919 12170 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16839 12170 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16759 12170 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16679 12170 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12106 16599 12170 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4432 12153 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4346 12153 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4260 12153 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4174 12153 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4088 12153 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4002 12153 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3916 12153 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3830 12153 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3744 12153 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3658 12153 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3572 12153 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 18099 12113 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 18013 12113 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17927 12113 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17841 12113 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17755 12113 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12049 17670 12113 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16472 12082 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16391 12082 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16310 12082 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16229 12082 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16148 12082 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16067 12082 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15986 12082 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15905 12082 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15824 12082 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15743 12082 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15662 12082 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15581 12082 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15500 12082 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15419 12082 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15338 12082 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15257 12082 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15176 12082 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15095 12082 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15014 12082 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14933 12082 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14852 12082 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14771 12082 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14690 12082 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14609 12082 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14527 12082 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14445 12082 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14363 12082 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14281 12082 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14199 12082 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14117 12082 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14035 12082 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13953 12082 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13871 12082 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13789 12082 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13707 12082 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13625 12082 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17563 12088 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17482 12088 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17401 12088 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17320 12088 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17239 12088 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17159 12088 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 17079 12088 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16999 12088 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16919 12088 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16839 12088 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16759 12088 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16679 12088 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12024 16599 12088 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4432 12072 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4346 12072 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4260 12072 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4174 12072 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4088 12072 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4002 12072 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3916 12072 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3830 12072 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3744 12072 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3658 12072 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3572 12072 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18277 12043 18341 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18191 12043 18255 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 18099 12031 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 18013 12031 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17927 12031 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17841 12031 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17755 12031 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11967 17670 12031 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16472 12002 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16391 12002 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16310 12002 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16229 12002 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16148 12002 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16067 12002 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15986 12002 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15905 12002 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15824 12002 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15743 12002 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15662 12002 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15581 12002 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15500 12002 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15419 12002 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15338 12002 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15257 12002 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15176 12002 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15095 12002 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15014 12002 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14933 12002 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14852 12002 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14771 12002 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14690 12002 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14609 12002 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14527 12002 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14445 12002 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14363 12002 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14281 12002 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14199 12002 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14117 12002 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14035 12002 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13953 12002 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13871 12002 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13789 12002 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13707 12002 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13625 12002 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17563 12006 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17482 12006 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17401 12006 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17320 12006 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17239 12006 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17159 12006 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 17079 12006 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16999 12006 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16919 12006 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16839 12006 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16759 12006 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16679 12006 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11942 16599 12006 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4432 11991 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4346 11991 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4260 11991 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4174 11991 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4088 11991 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4002 11991 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3916 11991 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3830 11991 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3744 11991 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3658 11991 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3572 11991 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 18099 11949 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 18013 11949 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17927 11949 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17841 11949 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17755 11949 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11885 17670 11949 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16472 11922 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16391 11922 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16310 11922 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16229 11922 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16148 11922 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16067 11922 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15986 11922 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15905 11922 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15824 11922 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15743 11922 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15662 11922 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15581 11922 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15500 11922 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15419 11922 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15338 11922 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15257 11922 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15176 11922 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15095 11922 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15014 11922 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14933 11922 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14852 11922 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14771 11922 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14690 11922 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14609 11922 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14527 11922 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14445 11922 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14363 11922 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14281 11922 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14199 11922 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14117 11922 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14035 11922 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13953 11922 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13871 11922 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13789 11922 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13707 11922 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13625 11922 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17563 11924 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17482 11924 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17401 11924 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17320 11924 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17239 11924 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17159 11924 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 17079 11924 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16999 11924 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16919 11924 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16839 11924 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16759 11924 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16679 11924 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11860 16599 11924 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4432 11910 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4346 11910 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4260 11910 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4174 11910 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4088 11910 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4002 11910 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3916 11910 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3830 11910 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3744 11910 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3658 11910 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3572 11910 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 18099 11867 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 18013 11867 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17927 11867 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17841 11867 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17755 11867 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11803 17670 11867 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16472 11842 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16391 11842 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16310 11842 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16229 11842 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16148 11842 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16067 11842 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15986 11842 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15905 11842 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15824 11842 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15743 11842 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15662 11842 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15581 11842 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15500 11842 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15419 11842 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15338 11842 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15257 11842 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15176 11842 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15095 11842 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15014 11842 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14933 11842 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14852 11842 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14771 11842 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14690 11842 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14609 11842 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14527 11842 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14445 11842 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14363 11842 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14281 11842 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14199 11842 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14117 11842 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14035 11842 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13953 11842 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13871 11842 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13789 11842 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13707 11842 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13625 11842 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17563 11842 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17482 11842 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17401 11842 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17320 11842 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17239 11842 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17159 11842 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 17079 11842 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16999 11842 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16919 11842 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16839 11842 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16759 11842 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16679 11842 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11778 16599 11842 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4432 11829 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4346 11829 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4260 11829 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4174 11829 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4088 11829 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4002 11829 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3916 11829 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3830 11829 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3744 11829 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3658 11829 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3572 11829 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16472 11762 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16391 11762 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16310 11762 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16229 11762 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16148 11762 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16067 11762 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15986 11762 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15905 11762 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15824 11762 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15743 11762 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15662 11762 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15581 11762 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15500 11762 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15419 11762 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15338 11762 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15257 11762 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15176 11762 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15095 11762 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15014 11762 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14933 11762 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14852 11762 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14771 11762 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14690 11762 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14609 11762 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14527 11762 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14445 11762 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14363 11762 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14281 11762 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14199 11762 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14117 11762 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14035 11762 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13953 11762 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13871 11762 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13789 11762 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13707 11762 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13625 11762 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11703 17841 11767 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11703 17757 11767 17821 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11703 17674 11767 17738 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17563 11760 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17482 11760 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17401 11760 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17320 11760 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17239 11760 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17159 11760 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 17079 11760 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16999 11760 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16919 11760 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16839 11760 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16759 11760 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16679 11760 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11696 16599 11760 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4432 11748 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4346 11748 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4260 11748 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4174 11748 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4088 11748 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4002 11748 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3916 11748 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3830 11748 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3744 11748 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3658 11748 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3572 11748 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16472 11682 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16391 11682 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16310 11682 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16229 11682 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16148 11682 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16067 11682 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15986 11682 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15905 11682 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15824 11682 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15743 11682 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15662 11682 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15581 11682 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15500 11682 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15419 11682 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15338 11682 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15257 11682 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15176 11682 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15095 11682 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15014 11682 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14933 11682 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14852 11682 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14771 11682 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14690 11682 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14609 11682 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14527 11682 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14445 11682 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14363 11682 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14281 11682 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14199 11682 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14117 11682 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14035 11682 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13953 11682 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13871 11682 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13789 11682 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13707 11682 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13625 11682 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4432 11667 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4346 11667 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4260 11667 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4174 11667 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4088 11667 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4002 11667 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3916 11667 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3830 11667 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3744 11667 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3658 11667 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3572 11667 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17563 11678 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17482 11678 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17401 11678 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17320 11678 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17239 11678 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17159 11678 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 17079 11678 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16999 11678 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16919 11678 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16839 11678 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16759 11678 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16679 11678 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11614 16599 11678 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16472 11602 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16391 11602 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16310 11602 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16229 11602 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16148 11602 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16067 11602 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15986 11602 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15905 11602 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15824 11602 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15743 11602 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15662 11602 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15581 11602 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15500 11602 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15419 11602 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15338 11602 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15257 11602 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15176 11602 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15095 11602 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15014 11602 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14933 11602 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14852 11602 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14771 11602 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14690 11602 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14609 11602 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14527 11602 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14445 11602 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14363 11602 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14281 11602 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14199 11602 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14117 11602 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14035 11602 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13953 11602 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13871 11602 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13789 11602 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13707 11602 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13625 11602 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11547 17841 11611 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11547 17757 11611 17821 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11547 17674 11611 17738 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4432 11586 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4346 11586 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4260 11586 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4174 11586 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4088 11586 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4002 11586 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3916 11586 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3830 11586 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3744 11586 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3658 11586 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3572 11586 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17563 11596 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17482 11596 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17401 11596 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17320 11596 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17239 11596 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17159 11596 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17079 11596 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16999 11596 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16919 11596 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16839 11596 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16759 11596 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16679 11596 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 16599 11596 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16472 11522 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16391 11522 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16310 11522 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16229 11522 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16148 11522 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16067 11522 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15986 11522 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15905 11522 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15824 11522 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15743 11522 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15662 11522 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15581 11522 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15500 11522 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15419 11522 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15338 11522 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15257 11522 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15176 11522 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15095 11522 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15014 11522 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14933 11522 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14852 11522 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14771 11522 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14690 11522 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14609 11522 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14527 11522 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14445 11522 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14363 11522 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14281 11522 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14199 11522 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14117 11522 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14035 11522 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13953 11522 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13871 11522 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13789 11522 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13707 11522 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13625 11522 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4432 11505 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4346 11505 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4260 11505 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4174 11505 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4088 11505 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4002 11505 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3916 11505 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3830 11505 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3744 11505 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3658 11505 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3572 11505 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17563 11514 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17482 11514 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17401 11514 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17320 11514 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17239 11514 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17159 11514 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 17079 11514 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16999 11514 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16919 11514 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16839 11514 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16759 11514 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16679 11514 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11450 16599 11514 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16472 11442 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16391 11442 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16310 11442 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16229 11442 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16148 11442 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16067 11442 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15986 11442 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15905 11442 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15824 11442 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15743 11442 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15662 11442 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15581 11442 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15500 11442 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15419 11442 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15338 11442 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15257 11442 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15176 11442 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15095 11442 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15014 11442 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14933 11442 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14852 11442 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14771 11442 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14690 11442 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14609 11442 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14527 11442 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14445 11442 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14363 11442 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14281 11442 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14199 11442 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14117 11442 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14035 11442 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13953 11442 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13871 11442 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13789 11442 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13707 11442 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13625 11442 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4432 11424 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4346 11424 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4260 11424 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4174 11424 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4088 11424 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4002 11424 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3916 11424 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3830 11424 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3744 11424 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3658 11424 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3572 11424 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17563 11432 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17482 11432 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17401 11432 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17320 11432 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17239 11432 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17159 11432 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 17079 11432 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16999 11432 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16919 11432 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16839 11432 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16759 11432 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16679 11432 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11368 16599 11432 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16472 11362 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16391 11362 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16310 11362 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16229 11362 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16148 11362 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16067 11362 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15986 11362 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15905 11362 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15824 11362 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15743 11362 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15662 11362 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15581 11362 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15500 11362 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15419 11362 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15338 11362 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15257 11362 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15176 11362 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15095 11362 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15014 11362 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14933 11362 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14852 11362 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14771 11362 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14690 11362 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14609 11362 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14527 11362 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14445 11362 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14363 11362 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14281 11362 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14199 11362 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14117 11362 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14035 11362 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13953 11362 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13871 11362 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13789 11362 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13707 11362 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13625 11362 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4432 11343 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4346 11343 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4260 11343 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4174 11343 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4088 11343 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4002 11343 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3916 11343 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3830 11343 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3744 11343 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3658 11343 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3572 11343 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17563 11350 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17482 11350 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17401 11350 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17320 11350 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17239 11350 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17159 11350 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 17079 11350 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16999 11350 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16919 11350 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16839 11350 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16759 11350 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16679 11350 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11286 16599 11350 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16472 11282 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16391 11282 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16310 11282 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16229 11282 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16148 11282 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16067 11282 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15986 11282 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15905 11282 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15824 11282 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15743 11282 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15662 11282 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15581 11282 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15500 11282 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15419 11282 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15338 11282 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15257 11282 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15176 11282 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15095 11282 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15014 11282 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14933 11282 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14852 11282 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14771 11282 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14690 11282 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14609 11282 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14527 11282 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14445 11282 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14363 11282 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14281 11282 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14199 11282 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14117 11282 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14035 11282 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13953 11282 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13871 11282 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13789 11282 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13707 11282 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13625 11282 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4432 11262 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4346 11262 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4260 11262 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4174 11262 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4088 11262 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4002 11262 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3916 11262 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3830 11262 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3744 11262 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3658 11262 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3572 11262 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11187 17338 11251 17402 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11187 17250 11251 17314 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11187 17163 11251 17227 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16472 11202 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16391 11202 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16310 11202 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16229 11202 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16148 11202 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16067 11202 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15986 11202 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15905 11202 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15824 11202 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15743 11202 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15662 11202 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15581 11202 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15500 11202 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15419 11202 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15338 11202 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15257 11202 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15176 11202 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15095 11202 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15014 11202 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14933 11202 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14852 11202 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14771 11202 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14690 11202 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14609 11202 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14527 11202 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14445 11202 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14363 11202 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14281 11202 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14199 11202 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14117 11202 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14035 11202 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13953 11202 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13871 11202 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13789 11202 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13707 11202 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13625 11202 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 17053 11213 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16960 11213 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16867 11213 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16774 11213 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16682 11213 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11149 16590 11213 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4432 11181 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4346 11181 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4260 11181 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4174 11181 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4088 11181 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4002 11181 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3916 11181 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3830 11181 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3744 11181 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3658 11181 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3572 11181 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16472 11122 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16391 11122 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16310 11122 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16229 11122 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16148 11122 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16067 11122 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15986 11122 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15905 11122 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15824 11122 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15743 11122 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15662 11122 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15581 11122 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15500 11122 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15419 11122 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15338 11122 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15257 11122 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15176 11122 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15095 11122 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15014 11122 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14933 11122 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14852 11122 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14771 11122 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14690 11122 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14609 11122 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14527 11122 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14445 11122 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14363 11122 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14281 11122 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14199 11122 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14117 11122 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14035 11122 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13953 11122 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13871 11122 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13789 11122 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13707 11122 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13625 11122 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 17053 11117 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16960 11117 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16867 11117 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16774 11117 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16682 11117 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11053 16590 11117 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4432 11100 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4346 11100 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4260 11100 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4174 11100 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4088 11100 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4002 11100 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3916 11100 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3830 11100 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3744 11100 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3658 11100 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3572 11100 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11039 17338 11103 17402 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11039 17250 11103 17314 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11039 17163 11103 17227 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16472 11042 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16391 11042 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16310 11042 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16229 11042 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16148 11042 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16067 11042 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15986 11042 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15905 11042 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15824 11042 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15743 11042 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15662 11042 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15581 11042 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15500 11042 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15419 11042 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15338 11042 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15257 11042 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15176 11042 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15095 11042 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15014 11042 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14933 11042 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14852 11042 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14771 11042 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14690 11042 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14609 11042 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14527 11042 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14445 11042 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14363 11042 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14281 11042 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14199 11042 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14117 11042 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14035 11042 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13953 11042 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13871 11042 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13789 11042 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13707 11042 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13625 11042 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4432 11019 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4346 11019 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4260 11019 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4174 11019 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4088 11019 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4002 11019 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3916 11019 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3830 11019 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3744 11019 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3658 11019 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3572 11019 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 17053 11021 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16960 11021 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16867 11021 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16774 11021 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16682 11021 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10957 16590 11021 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16472 10962 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16391 10962 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16310 10962 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16229 10962 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16148 10962 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16067 10962 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15986 10962 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15905 10962 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15824 10962 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15743 10962 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15662 10962 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15581 10962 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15500 10962 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15419 10962 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15338 10962 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15257 10962 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15176 10962 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15095 10962 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15014 10962 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14933 10962 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14852 10962 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14771 10962 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14690 10962 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14609 10962 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14527 10962 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14445 10962 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14363 10962 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14281 10962 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14199 10962 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14117 10962 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14035 10962 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13953 10962 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13871 10962 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13789 10962 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13707 10962 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13625 10962 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4432 10938 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4346 10938 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4260 10938 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4174 10938 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4088 10938 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4002 10938 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3916 10938 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3830 10938 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3744 10938 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3658 10938 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3572 10938 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 17053 10925 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16960 10925 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16867 10925 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16774 10925 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16682 10925 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10861 16590 10925 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16472 10882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16391 10882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16310 10882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16229 10882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16148 10882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16067 10882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15986 10882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15905 10882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15824 10882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15743 10882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15662 10882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15581 10882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15500 10882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15419 10882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15338 10882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15257 10882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15176 10882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15095 10882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15014 10882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14933 10882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14852 10882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14771 10882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14690 10882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14609 10882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14527 10882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14445 10882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14363 10882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14281 10882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14199 10882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14117 10882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14035 10882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13953 10882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13871 10882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13789 10882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13707 10882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13625 10882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4432 10857 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4346 10857 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4260 10857 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4174 10857 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4088 10857 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4002 10857 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3916 10857 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3830 10857 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3744 10857 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3658 10857 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3572 10857 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 17053 10829 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16960 10829 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16867 10829 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16774 10829 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16682 10829 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10765 16590 10829 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16472 10802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16391 10802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16310 10802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16229 10802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16148 10802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16067 10802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15986 10802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15905 10802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15824 10802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15743 10802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15662 10802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15581 10802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15500 10802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15419 10802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15338 10802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15257 10802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15176 10802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15095 10802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15014 10802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14933 10802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14852 10802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14771 10802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14690 10802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14609 10802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14527 10802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14445 10802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14363 10802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14281 10802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14199 10802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14117 10802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14035 10802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13953 10802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13871 10802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13789 10802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13707 10802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13625 10802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4432 10776 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4346 10776 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4260 10776 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4174 10776 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4088 10776 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4002 10776 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3916 10776 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3830 10776 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3744 10776 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3658 10776 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3572 10776 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16472 10722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16391 10722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16310 10722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16229 10722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16148 10722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16067 10722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15986 10722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15905 10722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15824 10722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15743 10722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15662 10722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15581 10722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15500 10722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15419 10722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15338 10722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15257 10722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15176 10722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15095 10722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15014 10722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14933 10722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14852 10722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14771 10722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14690 10722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14609 10722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14527 10722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14445 10722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14363 10722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14281 10722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14199 10722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14117 10722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14035 10722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13953 10722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13871 10722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13789 10722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13707 10722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13625 10722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10656 16792 10720 16856 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10656 16682 10720 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10656 16572 10720 16636 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4432 10695 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4346 10695 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4260 10695 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4174 10695 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4088 10695 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4002 10695 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3916 10695 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3830 10695 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3744 10695 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3658 10695 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3572 10695 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16472 10642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16391 10642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16310 10642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16229 10642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16148 10642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16067 10642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15986 10642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15905 10642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15824 10642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15743 10642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15662 10642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15581 10642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15500 10642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15419 10642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15338 10642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15257 10642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15176 10642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15095 10642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15014 10642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14933 10642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14852 10642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14771 10642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14690 10642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14609 10642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14527 10642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14445 10642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14363 10642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14281 10642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14199 10642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14117 10642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14035 10642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13953 10642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13871 10642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13789 10642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13707 10642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13625 10642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4432 10614 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4346 10614 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4260 10614 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4174 10614 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4088 10614 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4002 10614 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3916 10614 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3830 10614 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3744 10614 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3658 10614 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3572 10614 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16472 10562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16391 10562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16310 10562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16229 10562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16148 10562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16067 10562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15986 10562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15905 10562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15824 10562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15743 10562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15662 10562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15581 10562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15500 10562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15419 10562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15338 10562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15257 10562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15176 10562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15095 10562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15014 10562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14933 10562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14852 10562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14771 10562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14690 10562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14609 10562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14527 10562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14445 10562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14363 10562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14281 10562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14199 10562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14117 10562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14035 10562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13953 10562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13871 10562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13789 10562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13707 10562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13625 10562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10498 16792 10562 16856 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10498 16682 10562 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10498 16572 10562 16636 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4432 10533 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4346 10533 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4260 10533 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4174 10533 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4088 10533 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4002 10533 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3916 10533 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3830 10533 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3744 10533 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3658 10533 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3572 10533 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16472 10482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16391 10482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16310 10482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16229 10482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16148 10482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16067 10482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15986 10482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15905 10482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15824 10482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15743 10482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15662 10482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15581 10482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15500 10482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15419 10482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15338 10482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15257 10482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15176 10482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15095 10482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15014 10482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14933 10482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14852 10482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14771 10482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14690 10482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14609 10482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14527 10482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14445 10482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14363 10482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14281 10482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14199 10482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14117 10482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14035 10482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13953 10482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13871 10482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13789 10482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13707 10482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13625 10482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4432 10452 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4346 10452 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4260 10452 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4174 10452 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4088 10452 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4002 10452 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3916 10452 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3830 10452 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3744 10452 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3658 10452 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3572 10452 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16472 10402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16391 10402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16310 10402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16229 10402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16148 10402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16067 10402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15986 10402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15905 10402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15824 10402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15743 10402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15662 10402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15581 10402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15500 10402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15419 10402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15338 10402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15257 10402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15176 10402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15095 10402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15014 10402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14933 10402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14852 10402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14771 10402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14690 10402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14609 10402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14527 10402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14445 10402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14363 10402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14281 10402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14199 10402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14117 10402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14035 10402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13953 10402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13871 10402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13789 10402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13707 10402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13625 10402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4432 10371 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4346 10371 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4260 10371 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4174 10371 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4088 10371 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4002 10371 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3916 10371 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3830 10371 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3744 10371 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3658 10371 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3572 10371 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16472 10322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16391 10322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16310 10322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16229 10322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16148 10322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16067 10322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15986 10322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15905 10322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15824 10322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15743 10322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15662 10322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15581 10322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15500 10322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15419 10322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15338 10322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15257 10322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15176 10322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15095 10322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15014 10322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14933 10322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14852 10322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14771 10322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14690 10322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14609 10322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14527 10322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14445 10322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14363 10322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14281 10322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14199 10322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14117 10322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14035 10322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13953 10322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13871 10322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13789 10322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13707 10322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13625 10322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4432 10290 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4346 10290 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4260 10290 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4174 10290 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4088 10290 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4002 10290 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3916 10290 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3830 10290 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3744 10290 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3658 10290 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3572 10290 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16472 10242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16391 10242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16310 10242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16229 10242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16148 10242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16067 10242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15986 10242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15905 10242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15824 10242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15743 10242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15662 10242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15581 10242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15500 10242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15419 10242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15338 10242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15257 10242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15176 10242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15095 10242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15014 10242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14933 10242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14852 10242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14771 10242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14690 10242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14609 10242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14527 10242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14445 10242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14363 10242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14281 10242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14199 10242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14117 10242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14035 10242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13953 10242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13871 10242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13789 10242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13707 10242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13625 10242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4432 10209 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4346 10209 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4260 10209 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4174 10209 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4088 10209 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4002 10209 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3916 10209 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3830 10209 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3744 10209 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3658 10209 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3572 10209 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4432 4882 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4346 4882 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4260 4882 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4174 4882 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4088 4882 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4002 4882 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3916 4882 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3830 4882 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3744 4882 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3658 4882 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3572 4882 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16460 4861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16460 4861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16379 4861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16379 4861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16298 4861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16298 4861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16217 4861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16217 4861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16136 4861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16136 4861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 16055 4861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16055 4861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15974 4861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15974 4861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15893 4861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15893 4861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15812 4861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15812 4861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15731 4861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15731 4861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15650 4861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15650 4861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15569 4861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15569 4861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15488 4861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15488 4861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15407 4861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15407 4861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15326 4861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15326 4861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15245 4861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15245 4861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15164 4861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15164 4861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15083 4861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15083 4861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 15002 4861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15002 4861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14921 4861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14921 4861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14840 4861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14840 4861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14759 4861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14759 4861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14678 4861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14678 4861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14597 4861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14597 4861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14515 4861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14515 4861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14433 4861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14433 4861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14351 4861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14351 4861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14269 4861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14269 4861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14187 4861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14187 4861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14105 4861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14105 4861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 14023 4861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14023 4861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13941 4861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13941 4861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13859 4861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13859 4861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13777 4861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13777 4861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13695 4861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13695 4861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4797 13613 4861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13613 4861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4432 4800 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4346 4800 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4260 4800 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4174 4800 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4088 4800 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4002 4800 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3916 4800 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3830 4800 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3744 4800 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3658 4800 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3572 4800 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16460 4781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16460 4781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16379 4781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16379 4781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16298 4781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16298 4781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16217 4781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16217 4781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16136 4781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16136 4781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 16055 4781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16055 4781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15974 4781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15974 4781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15893 4781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15893 4781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15812 4781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15812 4781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15731 4781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15731 4781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15650 4781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15650 4781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15569 4781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15569 4781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15488 4781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15488 4781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15407 4781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15407 4781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15326 4781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15326 4781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15245 4781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15245 4781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15164 4781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15164 4781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15083 4781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15083 4781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 15002 4781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15002 4781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14921 4781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14921 4781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14840 4781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14840 4781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14759 4781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14759 4781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14678 4781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14678 4781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14597 4781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14597 4781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14515 4781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14515 4781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14433 4781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14433 4781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14351 4781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14351 4781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14269 4781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14269 4781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14187 4781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14187 4781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14105 4781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14105 4781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 14023 4781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14023 4781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13941 4781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13941 4781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13859 4781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13859 4781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13777 4781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13777 4781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13695 4781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13695 4781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4717 13613 4781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13613 4781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4432 4718 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4346 4718 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4260 4718 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4174 4718 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4088 4718 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4002 4718 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3916 4718 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3830 4718 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3744 4718 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3658 4718 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3572 4718 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16460 4701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16460 4701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16379 4701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16379 4701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16298 4701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16298 4701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16217 4701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16217 4701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16136 4701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16136 4701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 16055 4701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16055 4701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15974 4701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15974 4701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15893 4701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15893 4701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15812 4701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15812 4701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15731 4701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15731 4701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15650 4701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15650 4701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15569 4701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15569 4701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15488 4701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15488 4701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15407 4701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15407 4701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15326 4701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15326 4701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15245 4701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15245 4701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15164 4701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15164 4701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15083 4701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15083 4701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 15002 4701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15002 4701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14921 4701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14921 4701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14840 4701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14840 4701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14759 4701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14759 4701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14678 4701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14678 4701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14597 4701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14597 4701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14515 4701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14515 4701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14433 4701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14433 4701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14351 4701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14351 4701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14269 4701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14269 4701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14187 4701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14187 4701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14105 4701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14105 4701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 14023 4701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14023 4701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13941 4701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13941 4701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13859 4701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13859 4701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13777 4701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13777 4701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13695 4701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13695 4701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4637 13613 4701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13613 4701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4432 4636 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4346 4636 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4260 4636 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4174 4636 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4088 4636 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4002 4636 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3916 4636 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3830 4636 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3744 4636 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3658 4636 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3572 4636 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16460 4621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16460 4621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16379 4621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16379 4621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16298 4621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16298 4621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16217 4621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16217 4621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16136 4621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16136 4621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 16055 4621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16055 4621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15974 4621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15974 4621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15893 4621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15893 4621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15812 4621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15812 4621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15731 4621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15731 4621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15650 4621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15650 4621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15569 4621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15569 4621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15488 4621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15488 4621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15407 4621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15407 4621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15326 4621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15326 4621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15245 4621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15245 4621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15164 4621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15164 4621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15083 4621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15083 4621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 15002 4621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15002 4621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14921 4621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14921 4621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14840 4621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14840 4621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14759 4621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14759 4621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14678 4621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14678 4621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14597 4621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14597 4621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14515 4621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14515 4621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14433 4621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14433 4621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14351 4621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14351 4621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14269 4621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14269 4621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14187 4621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14187 4621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14105 4621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14105 4621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 14023 4621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14023 4621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13941 4621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13941 4621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13859 4621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13859 4621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13777 4621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13777 4621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13695 4621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13695 4621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4557 13613 4621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13613 4621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4432 4554 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4346 4554 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4260 4554 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4174 4554 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4088 4554 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4002 4554 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3916 4554 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3830 4554 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3744 4554 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3658 4554 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3572 4554 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16792 4553 16856 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16682 4553 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16572 4553 16636 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16460 4541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16460 4541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16379 4541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16379 4541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16298 4541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16298 4541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16217 4541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16217 4541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16136 4541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16136 4541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 16055 4541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16055 4541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15974 4541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15974 4541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15893 4541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15893 4541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15812 4541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15812 4541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15731 4541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15731 4541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15650 4541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15650 4541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15569 4541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15569 4541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15488 4541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15488 4541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15407 4541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15407 4541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15326 4541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15326 4541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15245 4541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15245 4541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15164 4541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15164 4541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15083 4541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15083 4541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 15002 4541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15002 4541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14921 4541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14921 4541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14840 4541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14840 4541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14759 4541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14759 4541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14678 4541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14678 4541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14597 4541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14597 4541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14515 4541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14515 4541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14433 4541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14433 4541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14351 4541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14351 4541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14269 4541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14269 4541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14187 4541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14187 4541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14105 4541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14105 4541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 14023 4541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14023 4541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13941 4541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13941 4541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13859 4541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13859 4541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13777 4541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13777 4541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13695 4541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13695 4541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4477 13613 4541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13613 4541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4432 4472 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4346 4472 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4260 4472 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4174 4472 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4088 4472 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4002 4472 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3916 4472 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3830 4472 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3744 4472 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3658 4472 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3572 4472 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16460 4461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16460 4461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16379 4461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16379 4461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16298 4461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16298 4461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16217 4461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16217 4461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16136 4461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16136 4461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 16055 4461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16055 4461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15974 4461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15974 4461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15893 4461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15893 4461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15812 4461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15812 4461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15731 4461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15731 4461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15650 4461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15650 4461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15569 4461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15569 4461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15488 4461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15488 4461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15407 4461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15407 4461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15326 4461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15326 4461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15245 4461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15245 4461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15164 4461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15164 4461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15083 4461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15083 4461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 15002 4461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15002 4461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14921 4461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14921 4461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14840 4461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14840 4461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14759 4461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14759 4461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14678 4461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14678 4461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14597 4461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14597 4461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14515 4461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14515 4461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14433 4461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14433 4461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14351 4461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14351 4461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14269 4461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14269 4461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14187 4461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14187 4461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14105 4461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14105 4461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 14023 4461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14023 4461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13941 4461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13941 4461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13859 4461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13859 4461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13777 4461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13777 4461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13695 4461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13695 4461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4397 13613 4461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13613 4461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4432 4390 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4346 4390 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4260 4390 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4174 4390 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4088 4390 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4002 4390 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3916 4390 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3830 4390 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3744 4390 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3658 4390 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3572 4390 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16792 4395 16856 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16682 4395 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16572 4395 16636 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16460 4381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16460 4381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16379 4381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16379 4381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16298 4381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16298 4381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16217 4381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16217 4381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16136 4381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16136 4381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 16055 4381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16055 4381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15974 4381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15974 4381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15893 4381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15893 4381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15812 4381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15812 4381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15731 4381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15731 4381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15650 4381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15650 4381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15569 4381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15569 4381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15488 4381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15488 4381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15407 4381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15407 4381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15326 4381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15326 4381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15245 4381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15245 4381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15164 4381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15164 4381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15083 4381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15083 4381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 15002 4381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15002 4381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14921 4381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14921 4381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14840 4381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14840 4381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14759 4381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14759 4381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14678 4381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14678 4381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14597 4381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14597 4381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14515 4381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14515 4381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14433 4381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14433 4381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14351 4381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14351 4381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14269 4381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14269 4381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14187 4381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14187 4381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14105 4381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14105 4381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 14023 4381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14023 4381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13941 4381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13941 4381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13859 4381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13859 4381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13777 4381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13777 4381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13695 4381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13695 4381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4317 13613 4381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13613 4381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4432 4309 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4346 4309 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4260 4309 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4174 4309 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4088 4309 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4002 4309 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3916 4309 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3830 4309 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3744 4309 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3658 4309 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3572 4309 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16460 4301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16460 4301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16379 4301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16379 4301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16298 4301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16298 4301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16217 4301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16217 4301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16136 4301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16136 4301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 16055 4301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16055 4301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15974 4301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15974 4301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15893 4301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15893 4301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15812 4301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15812 4301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15731 4301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15731 4301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15650 4301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15650 4301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15569 4301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15569 4301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15488 4301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15488 4301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15407 4301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15407 4301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15326 4301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15326 4301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15245 4301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15245 4301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15164 4301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15164 4301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15083 4301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15083 4301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 15002 4301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15002 4301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14921 4301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14921 4301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14840 4301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14840 4301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14759 4301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14759 4301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14678 4301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14678 4301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14597 4301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14597 4301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14515 4301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14515 4301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14433 4301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14433 4301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14351 4301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14351 4301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14269 4301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14269 4301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14187 4301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14187 4301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14105 4301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14105 4301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 14023 4301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14023 4301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13941 4301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13941 4301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13859 4301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13859 4301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13777 4301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13777 4301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13695 4301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13695 4301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4237 13613 4301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13613 4301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 17053 4286 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16960 4286 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16867 4286 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16774 4286 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16682 4286 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16590 4286 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4432 4228 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4346 4228 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4260 4228 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4174 4228 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4088 4228 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4002 4228 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3916 4228 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3830 4228 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3744 4228 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3658 4228 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3572 4228 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16460 4221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16460 4221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16379 4221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16379 4221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16298 4221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16298 4221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16217 4221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16217 4221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16136 4221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16136 4221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 16055 4221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16055 4221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15974 4221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15974 4221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15893 4221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15893 4221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15812 4221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15812 4221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15731 4221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15731 4221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15650 4221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15650 4221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15569 4221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15569 4221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15488 4221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15488 4221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15407 4221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15407 4221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15326 4221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15326 4221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15245 4221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15245 4221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15164 4221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15164 4221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15083 4221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15083 4221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 15002 4221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15002 4221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14921 4221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14921 4221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14840 4221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14840 4221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14759 4221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14759 4221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14678 4221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14678 4221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14597 4221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14597 4221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14515 4221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14515 4221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14433 4221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14433 4221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14351 4221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14351 4221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14269 4221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14269 4221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14187 4221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14187 4221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14105 4221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14105 4221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 14023 4221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14023 4221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13941 4221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13941 4221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13859 4221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13859 4221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13777 4221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13777 4221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13695 4221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13695 4221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4157 13613 4221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13613 4221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 17053 4190 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16960 4190 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16867 4190 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16774 4190 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16682 4190 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16590 4190 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4432 4147 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4346 4147 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4260 4147 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4174 4147 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4088 4147 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4002 4147 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3916 4147 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3830 4147 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3744 4147 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3658 4147 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3572 4147 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16460 4141 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16460 4141 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16379 4141 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16379 4141 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16298 4141 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16298 4141 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16217 4141 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16217 4141 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16136 4141 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16136 4141 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 16055 4141 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16055 4141 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15974 4141 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15974 4141 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15893 4141 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15893 4141 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15812 4141 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15812 4141 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15731 4141 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15731 4141 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15650 4141 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15650 4141 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15569 4141 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15569 4141 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15488 4141 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15488 4141 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15407 4141 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15407 4141 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15326 4141 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15326 4141 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15245 4141 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15245 4141 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15164 4141 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15164 4141 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15083 4141 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15083 4141 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 15002 4141 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15002 4141 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14921 4141 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14921 4141 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14840 4141 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14840 4141 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14759 4141 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14759 4141 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14678 4141 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14678 4141 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14597 4141 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14597 4141 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14515 4141 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14515 4141 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14433 4141 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14433 4141 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14351 4141 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14351 4141 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14269 4141 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14269 4141 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14187 4141 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14187 4141 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14105 4141 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14105 4141 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 14023 4141 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14023 4141 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13941 4141 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13941 4141 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13859 4141 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13859 4141 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13777 4141 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13777 4141 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13695 4141 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13695 4141 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4077 13613 4141 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13613 4141 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 17053 4094 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16960 4094 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16867 4094 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16774 4094 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16682 4094 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16590 4094 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4432 4066 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4346 4066 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4260 4066 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4174 4066 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4088 4066 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4002 4066 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3916 4066 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3830 4066 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3744 4066 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3658 4066 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3572 4066 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16460 4061 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16460 4061 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16379 4061 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16379 4061 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16298 4061 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16298 4061 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16217 4061 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16217 4061 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16136 4061 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16136 4061 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 16055 4061 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16055 4061 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15974 4061 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15974 4061 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15893 4061 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15893 4061 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15812 4061 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15812 4061 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15731 4061 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15731 4061 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15650 4061 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15650 4061 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15569 4061 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15569 4061 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15488 4061 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15488 4061 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15407 4061 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15407 4061 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15326 4061 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15326 4061 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15245 4061 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15245 4061 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15164 4061 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15164 4061 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15083 4061 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15083 4061 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 15002 4061 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15002 4061 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14921 4061 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14921 4061 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14840 4061 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14840 4061 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14759 4061 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14759 4061 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14678 4061 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14678 4061 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14597 4061 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14597 4061 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14515 4061 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14515 4061 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14433 4061 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14433 4061 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14351 4061 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14351 4061 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14269 4061 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14269 4061 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14187 4061 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14187 4061 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14105 4061 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14105 4061 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 14023 4061 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14023 4061 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13941 4061 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13941 4061 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13859 4061 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13859 4061 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13777 4061 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13777 4061 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13695 4061 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13695 4061 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3997 13613 4061 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13613 4061 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17338 4012 17402 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17250 4012 17314 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17163 4012 17227 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 17053 3998 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16960 3998 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16867 3998 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16774 3998 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16682 3998 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16590 3998 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4432 3985 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4346 3985 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4260 3985 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4174 3985 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4088 3985 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4002 3985 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3916 3985 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3830 3985 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3744 3985 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3658 3985 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3572 3985 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16460 3981 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16460 3981 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16379 3981 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16379 3981 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16298 3981 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16298 3981 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16217 3981 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16217 3981 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16136 3981 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16136 3981 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 16055 3981 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16055 3981 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15974 3981 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15974 3981 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15893 3981 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15893 3981 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15812 3981 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15812 3981 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15731 3981 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15731 3981 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15650 3981 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15650 3981 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15569 3981 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15569 3981 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15488 3981 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15488 3981 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15407 3981 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15407 3981 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15326 3981 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15326 3981 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15245 3981 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15245 3981 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15164 3981 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15164 3981 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15083 3981 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15083 3981 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 15002 3981 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15002 3981 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14921 3981 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14921 3981 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14840 3981 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14840 3981 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14759 3981 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14759 3981 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14678 3981 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14678 3981 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14597 3981 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14597 3981 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14515 3981 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14515 3981 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14433 3981 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14433 3981 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14351 3981 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14351 3981 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14269 3981 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14269 3981 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14187 3981 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14187 3981 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14105 3981 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14105 3981 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 14023 3981 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14023 3981 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13941 3981 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13941 3981 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13859 3981 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13859 3981 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13777 3981 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13777 3981 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13695 3981 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13695 3981 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3917 13613 3981 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13613 3981 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4432 3904 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4346 3904 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4260 3904 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4174 3904 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4088 3904 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4002 3904 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3916 3904 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3830 3904 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3744 3904 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3658 3904 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3572 3904 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 17053 3902 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16960 3902 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16867 3902 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16774 3902 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16682 3902 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16590 3902 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16460 3901 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16460 3901 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16379 3901 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16379 3901 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16298 3901 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16298 3901 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16217 3901 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16217 3901 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16136 3901 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16136 3901 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 16055 3901 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16055 3901 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15974 3901 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15974 3901 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15893 3901 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15893 3901 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15812 3901 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15812 3901 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15731 3901 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15731 3901 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15650 3901 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15650 3901 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15569 3901 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15569 3901 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15488 3901 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15488 3901 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15407 3901 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15407 3901 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15326 3901 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15326 3901 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15245 3901 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15245 3901 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15164 3901 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15164 3901 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15083 3901 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15083 3901 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 15002 3901 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15002 3901 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14921 3901 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14921 3901 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14840 3901 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14840 3901 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14759 3901 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14759 3901 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14678 3901 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14678 3901 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14597 3901 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14597 3901 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14515 3901 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14515 3901 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14433 3901 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14433 3901 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14351 3901 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14351 3901 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14269 3901 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14269 3901 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14187 3901 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14187 3901 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14105 3901 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14105 3901 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 14023 3901 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14023 3901 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13941 3901 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13941 3901 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13859 3901 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13859 3901 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13777 3901 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13777 3901 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13695 3901 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13695 3901 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3837 13613 3901 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13613 3901 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17338 3864 17402 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17250 3864 17314 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17163 3864 17227 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4432 3823 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4346 3823 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4260 3823 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4174 3823 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4088 3823 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4002 3823 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3916 3823 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3830 3823 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3744 3823 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3658 3823 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3572 3823 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16460 3821 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16460 3821 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16379 3821 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16379 3821 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16298 3821 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16298 3821 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16217 3821 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16217 3821 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16136 3821 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16136 3821 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 16055 3821 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16055 3821 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15974 3821 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15974 3821 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15893 3821 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15893 3821 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15812 3821 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15812 3821 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15731 3821 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15731 3821 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15650 3821 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15650 3821 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15569 3821 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15569 3821 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15488 3821 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15488 3821 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15407 3821 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15407 3821 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15326 3821 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15326 3821 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15245 3821 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15245 3821 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15164 3821 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15164 3821 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15083 3821 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15083 3821 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 15002 3821 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15002 3821 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14921 3821 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14921 3821 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14840 3821 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14840 3821 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14759 3821 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14759 3821 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14678 3821 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14678 3821 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14597 3821 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14597 3821 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14515 3821 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14515 3821 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14433 3821 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14433 3821 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14351 3821 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14351 3821 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14269 3821 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14269 3821 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14187 3821 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14187 3821 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14105 3821 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14105 3821 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 14023 3821 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14023 3821 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13941 3821 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13941 3821 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13859 3821 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13859 3821 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13777 3821 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13777 3821 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13695 3821 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13695 3821 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3757 13613 3821 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13613 3821 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17563 3765 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17482 3765 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17401 3765 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17320 3765 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17239 3765 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17159 3765 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17079 3765 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16999 3765 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16919 3765 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16839 3765 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16759 3765 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16679 3765 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16599 3765 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4432 3742 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4346 3742 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4260 3742 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4174 3742 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4088 3742 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4002 3742 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3916 3742 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3830 3742 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3744 3742 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3658 3742 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3572 3742 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16460 3741 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16460 3741 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16379 3741 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16379 3741 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16298 3741 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16298 3741 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16217 3741 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16217 3741 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16136 3741 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16136 3741 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 16055 3741 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16055 3741 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15974 3741 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15974 3741 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15893 3741 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15893 3741 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15812 3741 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15812 3741 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15731 3741 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15731 3741 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15650 3741 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15650 3741 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15569 3741 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15569 3741 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15488 3741 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15488 3741 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15407 3741 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15407 3741 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15326 3741 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15326 3741 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15245 3741 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15245 3741 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15164 3741 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15164 3741 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15083 3741 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15083 3741 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 15002 3741 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15002 3741 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14921 3741 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14921 3741 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14840 3741 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14840 3741 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14759 3741 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14759 3741 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14678 3741 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14678 3741 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14597 3741 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14597 3741 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14515 3741 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14515 3741 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14433 3741 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14433 3741 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14351 3741 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14351 3741 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14269 3741 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14269 3741 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14187 3741 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14187 3741 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14105 3741 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14105 3741 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 14023 3741 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14023 3741 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13941 3741 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13941 3741 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13859 3741 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13859 3741 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13777 3741 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13777 3741 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13695 3741 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13695 3741 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3677 13613 3741 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13613 3741 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17563 3683 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17482 3683 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17401 3683 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17320 3683 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17239 3683 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17159 3683 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17079 3683 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16999 3683 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16919 3683 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16839 3683 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16759 3683 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16679 3683 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16599 3683 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4432 3661 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4346 3661 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4260 3661 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4174 3661 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4088 3661 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4002 3661 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3916 3661 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3830 3661 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3744 3661 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3658 3661 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3572 3661 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16460 3661 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16460 3661 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16379 3661 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16379 3661 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16298 3661 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16298 3661 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16217 3661 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16217 3661 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16136 3661 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16136 3661 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 16055 3661 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16055 3661 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15974 3661 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15974 3661 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15893 3661 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15893 3661 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15812 3661 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15812 3661 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15731 3661 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15731 3661 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15650 3661 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15650 3661 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15569 3661 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15569 3661 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15488 3661 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15488 3661 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15407 3661 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15407 3661 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15326 3661 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15326 3661 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15245 3661 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15245 3661 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15164 3661 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15164 3661 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15083 3661 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15083 3661 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 15002 3661 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15002 3661 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14921 3661 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14921 3661 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14840 3661 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14840 3661 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14759 3661 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14759 3661 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14678 3661 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14678 3661 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14597 3661 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14597 3661 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14515 3661 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14515 3661 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14433 3661 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14433 3661 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14351 3661 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14351 3661 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14269 3661 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14269 3661 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14187 3661 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14187 3661 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14105 3661 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14105 3661 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 14023 3661 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14023 3661 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13941 3661 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13941 3661 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13859 3661 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13859 3661 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13777 3661 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13777 3661 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13695 3661 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13695 3661 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3597 13613 3661 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13613 3661 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17563 3601 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17482 3601 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17401 3601 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17320 3601 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17239 3601 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17159 3601 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17079 3601 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16999 3601 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16919 3601 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16839 3601 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16759 3601 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16679 3601 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16599 3601 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4432 3580 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4346 3580 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4260 3580 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4174 3580 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4088 3580 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4002 3580 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3916 3580 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3830 3580 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3744 3580 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3658 3580 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3572 3580 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16460 3581 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16460 3581 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16379 3581 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16379 3581 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16298 3581 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16298 3581 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16217 3581 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16217 3581 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16136 3581 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16136 3581 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 16055 3581 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16055 3581 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15974 3581 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15974 3581 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15893 3581 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15893 3581 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15812 3581 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15812 3581 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15731 3581 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15731 3581 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15650 3581 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15650 3581 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15569 3581 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15569 3581 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15488 3581 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15488 3581 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15407 3581 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15407 3581 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15326 3581 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15326 3581 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15245 3581 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15245 3581 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15164 3581 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15164 3581 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15083 3581 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15083 3581 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 15002 3581 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15002 3581 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14921 3581 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14921 3581 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14840 3581 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14840 3581 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14759 3581 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14759 3581 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14678 3581 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14678 3581 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14597 3581 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14597 3581 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14515 3581 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14515 3581 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14433 3581 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14433 3581 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14351 3581 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14351 3581 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14269 3581 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14269 3581 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14187 3581 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14187 3581 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14105 3581 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14105 3581 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 14023 3581 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14023 3581 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13941 3581 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13941 3581 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13859 3581 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13859 3581 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13777 3581 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13777 3581 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13695 3581 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13695 3581 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3517 13613 3581 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13613 3581 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17563 3519 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17482 3519 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17401 3519 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17320 3519 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17239 3519 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17159 3519 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17079 3519 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16999 3519 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16919 3519 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16839 3519 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16759 3519 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16679 3519 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16599 3519 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4432 3499 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4346 3499 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4260 3499 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4174 3499 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4088 3499 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4002 3499 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3916 3499 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3830 3499 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3744 3499 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3658 3499 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3572 3499 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17841 3504 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17757 3504 17821 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17674 3504 17738 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16460 3501 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16460 3501 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16379 3501 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16379 3501 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16298 3501 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16298 3501 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16217 3501 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16217 3501 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16136 3501 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16136 3501 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 16055 3501 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16055 3501 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15974 3501 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15974 3501 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15893 3501 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15893 3501 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15812 3501 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15812 3501 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15731 3501 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15731 3501 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15650 3501 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15650 3501 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15569 3501 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15569 3501 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15488 3501 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15488 3501 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15407 3501 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15407 3501 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15326 3501 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15326 3501 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15245 3501 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15245 3501 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15164 3501 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15164 3501 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15083 3501 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15083 3501 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 15002 3501 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15002 3501 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14921 3501 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14921 3501 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14840 3501 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14840 3501 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14759 3501 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14759 3501 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14678 3501 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14678 3501 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14597 3501 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14597 3501 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14515 3501 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14515 3501 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14433 3501 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14433 3501 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14351 3501 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14351 3501 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14269 3501 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14269 3501 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14187 3501 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14187 3501 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14105 3501 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14105 3501 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 14023 3501 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14023 3501 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13941 3501 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13941 3501 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13859 3501 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13859 3501 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13777 3501 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13777 3501 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13695 3501 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13695 3501 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3437 13613 3501 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13613 3501 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17563 3437 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17482 3437 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17401 3437 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17320 3437 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17239 3437 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17159 3437 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17079 3437 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16999 3437 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16919 3437 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16839 3437 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16759 3437 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16679 3437 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16599 3437 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4432 3418 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4346 3418 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4260 3418 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4174 3418 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4088 3418 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4002 3418 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3916 3418 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3830 3418 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3744 3418 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3658 3418 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3572 3418 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16460 3421 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16460 3421 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16379 3421 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16379 3421 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16298 3421 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16298 3421 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16217 3421 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16217 3421 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16136 3421 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16136 3421 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 16055 3421 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16055 3421 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15974 3421 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15974 3421 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15893 3421 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15893 3421 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15812 3421 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15812 3421 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15731 3421 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15731 3421 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15650 3421 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15650 3421 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15569 3421 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15569 3421 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15488 3421 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15488 3421 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15407 3421 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15407 3421 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15326 3421 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15326 3421 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15245 3421 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15245 3421 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15164 3421 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15164 3421 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15083 3421 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15083 3421 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 15002 3421 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15002 3421 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14921 3421 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14921 3421 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14840 3421 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14840 3421 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14759 3421 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14759 3421 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14678 3421 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14678 3421 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14597 3421 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14597 3421 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14515 3421 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14515 3421 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14433 3421 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14433 3421 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14351 3421 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14351 3421 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14269 3421 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14269 3421 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14187 3421 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14187 3421 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14105 3421 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14105 3421 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 14023 3421 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14023 3421 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13941 3421 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13941 3421 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13859 3421 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13859 3421 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13777 3421 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13777 3421 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13695 3421 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13695 3421 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3357 13613 3421 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13613 3421 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17563 3355 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17482 3355 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17401 3355 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17320 3355 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17239 3355 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17159 3355 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17079 3355 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16999 3355 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16919 3355 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16839 3355 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16759 3355 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16679 3355 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16599 3355 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4432 3337 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4346 3337 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4260 3337 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4174 3337 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4088 3337 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4002 3337 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3916 3337 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3830 3337 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3744 3337 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3658 3337 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3572 3337 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17841 3348 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17757 3348 17821 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17674 3348 17738 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16460 3341 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16460 3341 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16379 3341 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16379 3341 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16298 3341 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16298 3341 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16217 3341 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16217 3341 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16136 3341 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16136 3341 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 16055 3341 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16055 3341 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15974 3341 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15974 3341 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15893 3341 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15893 3341 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15812 3341 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15812 3341 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15731 3341 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15731 3341 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15650 3341 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15650 3341 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15569 3341 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15569 3341 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15488 3341 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15488 3341 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15407 3341 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15407 3341 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15326 3341 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15326 3341 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15245 3341 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15245 3341 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15164 3341 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15164 3341 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15083 3341 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15083 3341 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 15002 3341 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15002 3341 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14921 3341 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14921 3341 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14840 3341 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14840 3341 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14759 3341 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14759 3341 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14678 3341 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14678 3341 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14597 3341 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14597 3341 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14515 3341 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14515 3341 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14433 3341 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14433 3341 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14351 3341 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14351 3341 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14269 3341 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14269 3341 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14187 3341 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14187 3341 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14105 3341 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14105 3341 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 14023 3341 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14023 3341 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13941 3341 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13941 3341 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13859 3341 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13859 3341 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13777 3341 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13777 3341 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13695 3341 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13695 3341 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3277 13613 3341 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13613 3341 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17563 3273 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17482 3273 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17401 3273 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17320 3273 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17239 3273 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17159 3273 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17079 3273 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16999 3273 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16919 3273 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16839 3273 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16759 3273 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16679 3273 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16599 3273 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4432 3256 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4346 3256 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4260 3256 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4174 3256 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4088 3256 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4002 3256 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3916 3256 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3830 3256 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3744 3256 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3658 3256 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3572 3256 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16460 3261 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16460 3261 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16379 3261 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16379 3261 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16298 3261 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16298 3261 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16217 3261 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16217 3261 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16136 3261 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16136 3261 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 16055 3261 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16055 3261 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15974 3261 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15974 3261 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15893 3261 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15893 3261 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15812 3261 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15812 3261 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15731 3261 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15731 3261 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15650 3261 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15650 3261 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15569 3261 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15569 3261 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15488 3261 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15488 3261 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15407 3261 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15407 3261 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15326 3261 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15326 3261 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15245 3261 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15245 3261 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15164 3261 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15164 3261 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15083 3261 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15083 3261 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 15002 3261 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15002 3261 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14921 3261 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14921 3261 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14840 3261 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14840 3261 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14759 3261 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14759 3261 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14678 3261 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14678 3261 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14597 3261 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14597 3261 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14515 3261 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14515 3261 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14433 3261 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14433 3261 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14351 3261 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14351 3261 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14269 3261 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14269 3261 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14187 3261 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14187 3261 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14105 3261 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14105 3261 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 14023 3261 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14023 3261 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13941 3261 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13941 3261 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13859 3261 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13859 3261 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13777 3261 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13777 3261 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13695 3261 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13695 3261 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3197 13613 3261 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13613 3261 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 18099 3248 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 18013 3248 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17927 3248 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17841 3248 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17755 3248 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17670 3248 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17563 3191 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17482 3191 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17401 3191 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17320 3191 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17239 3191 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17159 3191 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17079 3191 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16999 3191 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16919 3191 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16839 3191 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16759 3191 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16679 3191 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16599 3191 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4432 3175 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4346 3175 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4260 3175 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4174 3175 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4088 3175 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4002 3175 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3916 3175 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3830 3175 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3744 3175 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3658 3175 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3572 3175 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16460 3181 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16460 3181 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16379 3181 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16379 3181 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16298 3181 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16298 3181 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16217 3181 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16217 3181 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16136 3181 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16136 3181 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 16055 3181 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16055 3181 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15974 3181 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15974 3181 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15893 3181 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15893 3181 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15812 3181 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15812 3181 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15731 3181 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15731 3181 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15650 3181 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15650 3181 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15569 3181 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15569 3181 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15488 3181 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15488 3181 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15407 3181 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15407 3181 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15326 3181 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15326 3181 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15245 3181 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15245 3181 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15164 3181 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15164 3181 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15083 3181 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15083 3181 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 15002 3181 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15002 3181 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14921 3181 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14921 3181 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14840 3181 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14840 3181 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14759 3181 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14759 3181 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14678 3181 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14678 3181 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14597 3181 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14597 3181 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14515 3181 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14515 3181 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14433 3181 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14433 3181 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14351 3181 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14351 3181 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14269 3181 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14269 3181 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14187 3181 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14187 3181 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14105 3181 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14105 3181 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 14023 3181 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14023 3181 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13941 3181 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13941 3181 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13859 3181 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13859 3181 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13777 3181 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13777 3181 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13695 3181 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13695 3181 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3117 13613 3181 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13613 3181 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 18099 3166 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 18013 3166 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17927 3166 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17841 3166 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17755 3166 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17670 3166 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17563 3109 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17482 3109 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17401 3109 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17320 3109 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17239 3109 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17159 3109 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17079 3109 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16999 3109 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16919 3109 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16839 3109 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16759 3109 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16679 3109 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16599 3109 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4432 3094 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4346 3094 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4260 3094 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4174 3094 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4088 3094 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4002 3094 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3916 3094 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3830 3094 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3744 3094 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3658 3094 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3572 3094 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16460 3101 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16460 3101 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16379 3101 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16379 3101 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16298 3101 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16298 3101 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16217 3101 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16217 3101 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16136 3101 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16136 3101 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 16055 3101 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16055 3101 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15974 3101 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15974 3101 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15893 3101 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15893 3101 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15812 3101 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15812 3101 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15731 3101 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15731 3101 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15650 3101 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15650 3101 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15569 3101 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15569 3101 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15488 3101 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15488 3101 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15407 3101 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15407 3101 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15326 3101 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15326 3101 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15245 3101 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15245 3101 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15164 3101 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15164 3101 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15083 3101 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15083 3101 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 15002 3101 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15002 3101 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14921 3101 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14921 3101 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14840 3101 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14840 3101 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14759 3101 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14759 3101 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14678 3101 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14678 3101 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14597 3101 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14597 3101 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14515 3101 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14515 3101 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14433 3101 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14433 3101 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14351 3101 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14351 3101 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14269 3101 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14269 3101 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14187 3101 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14187 3101 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14105 3101 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14105 3101 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 14023 3101 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14023 3101 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13941 3101 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13941 3101 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13859 3101 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13859 3101 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13777 3101 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13777 3101 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13695 3101 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13695 3101 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3037 13613 3101 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13613 3101 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18099 3084 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18013 3084 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17927 3084 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17841 3084 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17755 3084 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17670 3084 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3008 18277 3072 18341 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3008 18191 3072 18255 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17563 3027 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17482 3027 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17401 3027 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17320 3027 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17239 3027 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17159 3027 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17079 3027 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16999 3027 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16919 3027 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16839 3027 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16759 3027 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16679 3027 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16599 3027 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4432 3013 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4346 3013 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4260 3013 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4174 3013 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4088 3013 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4002 3013 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3916 3013 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3830 3013 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3744 3013 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3658 3013 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3572 3013 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16460 3021 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16460 3021 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16379 3021 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16379 3021 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16298 3021 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16298 3021 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16217 3021 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16217 3021 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16136 3021 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16136 3021 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 16055 3021 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16055 3021 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15974 3021 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15974 3021 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15893 3021 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15893 3021 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15812 3021 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15812 3021 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15731 3021 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15731 3021 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15650 3021 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15650 3021 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15569 3021 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15569 3021 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15488 3021 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15488 3021 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15407 3021 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15407 3021 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15326 3021 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15326 3021 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15245 3021 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15245 3021 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15164 3021 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15164 3021 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15083 3021 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15083 3021 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 15002 3021 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15002 3021 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14921 3021 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14921 3021 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14840 3021 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14840 3021 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14759 3021 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14759 3021 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14678 3021 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14678 3021 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14597 3021 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14597 3021 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14515 3021 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14515 3021 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14433 3021 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14433 3021 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14351 3021 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14351 3021 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14269 3021 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14269 3021 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14187 3021 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14187 3021 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14105 3021 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14105 3021 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 14023 3021 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14023 3021 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13941 3021 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13941 3021 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13859 3021 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13859 3021 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13777 3021 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13777 3021 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13695 3021 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13695 3021 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2957 13613 3021 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13613 3021 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 18099 3002 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 18013 3002 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17927 3002 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17841 3002 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17755 3002 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17670 3002 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17563 2945 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17482 2945 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17401 2945 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17320 2945 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17239 2945 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17159 2945 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17079 2945 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16999 2945 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16919 2945 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16839 2945 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16759 2945 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16679 2945 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16599 2945 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4432 2932 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4346 2932 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4260 2932 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4174 2932 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4088 2932 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4002 2932 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3916 2932 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3830 2932 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3744 2932 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3658 2932 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3572 2932 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16460 2941 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16460 2941 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16379 2941 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16379 2941 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16298 2941 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16298 2941 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16217 2941 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16217 2941 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16136 2941 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16136 2941 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 16055 2941 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16055 2941 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15974 2941 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15974 2941 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15893 2941 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15893 2941 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15812 2941 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15812 2941 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15731 2941 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15731 2941 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15650 2941 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15650 2941 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15569 2941 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15569 2941 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15488 2941 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15488 2941 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15407 2941 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15407 2941 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15326 2941 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15326 2941 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15245 2941 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15245 2941 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15164 2941 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15164 2941 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15083 2941 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15083 2941 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 15002 2941 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15002 2941 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14921 2941 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14921 2941 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14840 2941 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14840 2941 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14759 2941 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14759 2941 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14678 2941 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14678 2941 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14597 2941 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14597 2941 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14515 2941 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14515 2941 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14433 2941 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14433 2941 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14351 2941 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14351 2941 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14269 2941 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14269 2941 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14187 2941 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14187 2941 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14105 2941 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14105 2941 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 14023 2941 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14023 2941 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13941 2941 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13941 2941 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13859 2941 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13859 2941 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13777 2941 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13777 2941 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13695 2941 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13695 2941 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2877 13613 2941 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13613 2941 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 18099 2920 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 18013 2920 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17927 2920 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17841 2920 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17755 2920 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17670 2920 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2852 18277 2916 18341 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2852 18191 2916 18255 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4432 2851 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4346 2851 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4260 2851 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4174 2851 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4088 2851 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4002 2851 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3916 2851 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3830 2851 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3744 2851 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3658 2851 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3572 2851 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16460 2861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16460 2861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16379 2861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16379 2861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16298 2861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16298 2861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16217 2861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16217 2861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16136 2861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16136 2861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 16055 2861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16055 2861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15974 2861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15974 2861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15893 2861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15893 2861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15812 2861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15812 2861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15731 2861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15731 2861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15650 2861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15650 2861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15569 2861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15569 2861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15488 2861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15488 2861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15407 2861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15407 2861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15326 2861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15326 2861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15245 2861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15245 2861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15164 2861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15164 2861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15083 2861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15083 2861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 15002 2861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15002 2861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14921 2861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14921 2861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14840 2861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14840 2861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14759 2861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14759 2861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14678 2861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14678 2861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14597 2861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14597 2861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14515 2861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14515 2861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14433 2861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14433 2861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14351 2861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14351 2861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14269 2861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14269 2861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14187 2861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14187 2861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14105 2861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14105 2861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 14023 2861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14023 2861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13941 2861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13941 2861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13859 2861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13859 2861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13777 2861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13777 2861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13695 2861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13695 2861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2797 13613 2861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13613 2861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18527 2820 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18527 2820 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18445 2820 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18445 2820 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18363 2820 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18363 2820 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18281 2820 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18281 2820 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18199 2820 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18199 2820 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18117 2820 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18117 2820 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 18035 2820 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18035 2820 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17953 2820 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17953 2820 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17871 2820 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17871 2820 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17789 2820 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17789 2820 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17707 2820 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17707 2820 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17625 2820 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17625 2820 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17543 2820 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17543 2820 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17461 2820 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17461 2820 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17379 2820 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17379 2820 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17297 2820 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17297 2820 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17215 2820 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17215 2820 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17133 2820 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17133 2820 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 17051 2820 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17051 2820 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16969 2820 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16969 2820 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16887 2820 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16887 2820 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16805 2820 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16805 2820 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16723 2820 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16723 2820 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16641 2820 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16641 2820 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2756 16559 2820 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16559 2820 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4432 2770 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4346 2770 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4260 2770 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4174 2770 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4088 2770 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4002 2770 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3916 2770 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3830 2770 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3744 2770 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3658 2770 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3572 2770 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16460 2781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16460 2781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16379 2781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16379 2781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16298 2781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16298 2781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16217 2781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16217 2781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16136 2781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16136 2781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 16055 2781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16055 2781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15974 2781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15974 2781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15893 2781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15893 2781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15812 2781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15812 2781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15731 2781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15731 2781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15650 2781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15650 2781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15569 2781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15569 2781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15488 2781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15488 2781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15407 2781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15407 2781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15326 2781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15326 2781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15245 2781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15245 2781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15164 2781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15164 2781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15083 2781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15083 2781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 15002 2781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15002 2781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14921 2781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14921 2781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14840 2781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14840 2781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14759 2781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14759 2781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14678 2781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14678 2781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14597 2781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14597 2781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14515 2781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14515 2781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14433 2781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14433 2781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14351 2781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14351 2781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14269 2781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14269 2781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14187 2781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14187 2781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14105 2781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14105 2781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 14023 2781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14023 2781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13941 2781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13941 2781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13859 2781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13859 2781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13777 2781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13777 2781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13695 2781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13695 2781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2717 13613 2781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13613 2781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18527 2739 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18527 2739 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18445 2739 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18445 2739 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18363 2739 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18363 2739 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18281 2739 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18281 2739 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18199 2739 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18199 2739 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18117 2739 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18117 2739 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 18035 2739 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18035 2739 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17953 2739 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17953 2739 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17871 2739 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17871 2739 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17789 2739 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17789 2739 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17707 2739 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17707 2739 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17625 2739 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17625 2739 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17543 2739 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17543 2739 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17461 2739 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17461 2739 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17379 2739 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17379 2739 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17297 2739 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17297 2739 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17215 2739 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17215 2739 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17133 2739 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17133 2739 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 17051 2739 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17051 2739 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16969 2739 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16969 2739 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16887 2739 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16887 2739 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16805 2739 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16805 2739 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16723 2739 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16723 2739 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16641 2739 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16641 2739 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2675 16559 2739 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16559 2739 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16460 2701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16460 2701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16379 2701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16379 2701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16298 2701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16298 2701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16217 2701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16217 2701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16136 2701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16136 2701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 16055 2701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16055 2701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15974 2701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15974 2701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15893 2701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15893 2701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15812 2701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15812 2701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15731 2701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15731 2701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15650 2701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15650 2701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15569 2701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15569 2701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15488 2701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15488 2701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15407 2701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15407 2701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15326 2701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15326 2701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15245 2701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15245 2701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15164 2701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15164 2701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15083 2701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15083 2701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 15002 2701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15002 2701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14921 2701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14921 2701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14840 2701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14840 2701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14759 2701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14759 2701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14678 2701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14678 2701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14597 2701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14597 2701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14515 2701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14515 2701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14433 2701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14433 2701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14351 2701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14351 2701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14269 2701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14269 2701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14187 2701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14187 2701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14105 2701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14105 2701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 14023 2701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14023 2701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13941 2701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13941 2701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13859 2701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13859 2701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13777 2701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13777 2701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13695 2701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13695 2701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2637 13613 2701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13613 2701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4432 2689 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4346 2689 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4260 2689 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4174 2689 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4088 2689 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4002 2689 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3916 2689 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3830 2689 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3744 2689 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3658 2689 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3572 2689 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18527 2658 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18527 2658 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18445 2658 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18445 2658 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18363 2658 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18363 2658 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18281 2658 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18281 2658 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18199 2658 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18199 2658 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18117 2658 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18117 2658 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 18035 2658 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18035 2658 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17953 2658 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17953 2658 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17871 2658 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17871 2658 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17789 2658 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17789 2658 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17707 2658 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17707 2658 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17625 2658 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17625 2658 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17543 2658 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17543 2658 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17461 2658 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17461 2658 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17379 2658 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17379 2658 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17297 2658 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17297 2658 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17215 2658 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17215 2658 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17133 2658 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17133 2658 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 17051 2658 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17051 2658 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16969 2658 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16969 2658 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16887 2658 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16887 2658 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16805 2658 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16805 2658 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16723 2658 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16723 2658 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16641 2658 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16641 2658 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2594 16559 2658 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16559 2658 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16460 2621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16460 2621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16379 2621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16379 2621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16298 2621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16298 2621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16217 2621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16217 2621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16136 2621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16136 2621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 16055 2621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16055 2621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15974 2621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15974 2621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15893 2621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15893 2621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15812 2621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15812 2621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15731 2621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15731 2621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15650 2621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15650 2621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15569 2621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15569 2621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15488 2621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15488 2621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15407 2621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15407 2621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15326 2621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15326 2621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15245 2621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15245 2621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15164 2621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15164 2621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15083 2621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15083 2621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 15002 2621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15002 2621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14921 2621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14921 2621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14840 2621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14840 2621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14759 2621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14759 2621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14678 2621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14678 2621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14597 2621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14597 2621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14515 2621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14515 2621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14433 2621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14433 2621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14351 2621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14351 2621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14269 2621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14269 2621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14187 2621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14187 2621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14105 2621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14105 2621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 14023 2621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14023 2621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13941 2621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13941 2621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13859 2621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13859 2621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13777 2621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13777 2621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13695 2621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13695 2621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2557 13613 2621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13613 2621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4432 2608 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4346 2608 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4260 2608 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4174 2608 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4088 2608 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4002 2608 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3916 2608 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3830 2608 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3744 2608 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3658 2608 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3572 2608 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18527 2577 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18527 2577 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18445 2577 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18445 2577 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18363 2577 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18363 2577 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18281 2577 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18281 2577 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18199 2577 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18199 2577 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18117 2577 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18117 2577 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 18035 2577 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18035 2577 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17953 2577 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17953 2577 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17871 2577 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17871 2577 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17789 2577 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17789 2577 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17707 2577 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17707 2577 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17625 2577 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17625 2577 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17543 2577 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17543 2577 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17461 2577 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17461 2577 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17379 2577 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17379 2577 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17297 2577 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17297 2577 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17215 2577 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17215 2577 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17133 2577 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17133 2577 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 17051 2577 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17051 2577 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16969 2577 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16969 2577 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16887 2577 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16887 2577 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16805 2577 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16805 2577 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16723 2577 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16723 2577 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16641 2577 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16641 2577 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2513 16559 2577 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16559 2577 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16460 2541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16460 2541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16379 2541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16379 2541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16298 2541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16298 2541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16217 2541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16217 2541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16136 2541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16136 2541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 16055 2541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16055 2541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15974 2541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15974 2541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15893 2541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15893 2541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15812 2541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15812 2541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15731 2541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15731 2541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15650 2541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15650 2541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15569 2541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15569 2541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15488 2541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15488 2541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15407 2541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15407 2541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15326 2541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15326 2541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15245 2541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15245 2541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15164 2541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15164 2541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15083 2541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15083 2541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 15002 2541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15002 2541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14921 2541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14921 2541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14840 2541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14840 2541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14759 2541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14759 2541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14678 2541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14678 2541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14597 2541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14597 2541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14515 2541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14515 2541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14433 2541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14433 2541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14351 2541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14351 2541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14269 2541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14269 2541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14187 2541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14187 2541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14105 2541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14105 2541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 14023 2541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14023 2541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13941 2541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13941 2541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13859 2541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13859 2541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13777 2541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13777 2541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13695 2541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13695 2541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2477 13613 2541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13613 2541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4432 2527 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4346 2527 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4260 2527 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4174 2527 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4088 2527 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4002 2527 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3916 2527 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3830 2527 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3744 2527 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3658 2527 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3572 2527 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18527 2495 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18527 2495 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18445 2495 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18445 2495 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18363 2495 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18363 2495 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18281 2495 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18281 2495 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18199 2495 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18199 2495 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18117 2495 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18117 2495 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 18035 2495 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18035 2495 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17953 2495 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17953 2495 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17871 2495 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17871 2495 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17789 2495 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17789 2495 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17707 2495 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17707 2495 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17625 2495 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17625 2495 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17543 2495 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17543 2495 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17461 2495 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17461 2495 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17379 2495 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17379 2495 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17297 2495 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17297 2495 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17215 2495 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17215 2495 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17133 2495 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17133 2495 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 17051 2495 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17051 2495 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16969 2495 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16969 2495 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16887 2495 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16887 2495 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16805 2495 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16805 2495 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16723 2495 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16723 2495 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16641 2495 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16641 2495 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2431 16559 2495 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16559 2495 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16460 2461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16460 2461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16379 2461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16379 2461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16298 2461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16298 2461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16217 2461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16217 2461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16136 2461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16136 2461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 16055 2461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16055 2461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15974 2461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15974 2461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15893 2461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15893 2461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15812 2461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15812 2461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15731 2461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15731 2461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15650 2461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15650 2461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15569 2461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15569 2461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15488 2461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15488 2461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15407 2461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15407 2461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15326 2461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15326 2461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15245 2461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15245 2461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15164 2461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15164 2461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15083 2461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15083 2461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 15002 2461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15002 2461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14921 2461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14921 2461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14840 2461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14840 2461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14759 2461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14759 2461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14678 2461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14678 2461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14597 2461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14597 2461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14515 2461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14515 2461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14433 2461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14433 2461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14351 2461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14351 2461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14269 2461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14269 2461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14187 2461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14187 2461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14105 2461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14105 2461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 14023 2461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14023 2461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13941 2461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13941 2461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13859 2461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13859 2461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13777 2461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13777 2461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13695 2461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13695 2461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2397 13613 2461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13613 2461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4432 2446 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4346 2446 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4260 2446 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4174 2446 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4088 2446 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4002 2446 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3916 2446 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3830 2446 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3744 2446 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3658 2446 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3572 2446 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18527 2413 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18527 2413 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18445 2413 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18445 2413 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18363 2413 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18363 2413 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18281 2413 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18281 2413 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18199 2413 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18199 2413 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18117 2413 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18117 2413 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 18035 2413 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18035 2413 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17953 2413 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17953 2413 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17871 2413 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17871 2413 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17789 2413 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17789 2413 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17707 2413 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17707 2413 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17625 2413 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17625 2413 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17543 2413 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17543 2413 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17461 2413 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17461 2413 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17379 2413 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17379 2413 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17297 2413 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17297 2413 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17215 2413 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17215 2413 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17133 2413 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17133 2413 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 17051 2413 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17051 2413 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16969 2413 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16969 2413 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16887 2413 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16887 2413 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16805 2413 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16805 2413 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16723 2413 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16723 2413 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16641 2413 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16641 2413 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2349 16559 2413 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16559 2413 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16460 2381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16460 2381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16379 2381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16379 2381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16298 2381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16298 2381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16217 2381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16217 2381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16136 2381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16136 2381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 16055 2381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16055 2381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15974 2381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15974 2381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15893 2381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15893 2381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15812 2381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15812 2381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15731 2381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15731 2381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15650 2381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15650 2381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15569 2381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15569 2381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15488 2381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15488 2381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15407 2381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15407 2381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15326 2381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15326 2381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15245 2381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15245 2381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15164 2381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15164 2381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15083 2381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15083 2381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 15002 2381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15002 2381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14921 2381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14921 2381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14840 2381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14840 2381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14759 2381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14759 2381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14678 2381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14678 2381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14597 2381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14597 2381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14515 2381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14515 2381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14433 2381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14433 2381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14351 2381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14351 2381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14269 2381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14269 2381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14187 2381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14187 2381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14105 2381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14105 2381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 14023 2381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14023 2381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13941 2381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13941 2381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13859 2381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13859 2381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13777 2381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13777 2381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13695 2381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13695 2381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2317 13613 2381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13613 2381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4432 2365 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4346 2365 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4260 2365 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4174 2365 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4088 2365 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4002 2365 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3916 2365 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3830 2365 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3744 2365 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3658 2365 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3572 2365 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18527 2331 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18527 2331 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18445 2331 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18445 2331 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18363 2331 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18363 2331 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18281 2331 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18281 2331 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18199 2331 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18199 2331 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18117 2331 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18117 2331 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 18035 2331 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18035 2331 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17953 2331 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17953 2331 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17871 2331 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17871 2331 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17789 2331 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17789 2331 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17707 2331 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17707 2331 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17625 2331 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17625 2331 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17543 2331 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17543 2331 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17461 2331 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17461 2331 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17379 2331 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17379 2331 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17297 2331 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17297 2331 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17215 2331 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17215 2331 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17133 2331 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17133 2331 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 17051 2331 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17051 2331 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16969 2331 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16969 2331 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16887 2331 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16887 2331 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16805 2331 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16805 2331 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16723 2331 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16723 2331 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16641 2331 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16641 2331 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2267 16559 2331 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16559 2331 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16460 2301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16460 2301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16379 2301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16379 2301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16298 2301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16298 2301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16217 2301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16217 2301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16136 2301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16136 2301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 16055 2301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16055 2301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15974 2301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15974 2301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15893 2301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15893 2301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15812 2301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15812 2301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15731 2301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15731 2301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15650 2301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15650 2301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15569 2301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15569 2301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15488 2301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15488 2301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15407 2301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15407 2301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15326 2301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15326 2301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15245 2301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15245 2301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15164 2301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15164 2301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15083 2301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15083 2301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 15002 2301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15002 2301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14921 2301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14921 2301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14840 2301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14840 2301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14759 2301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14759 2301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14678 2301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14678 2301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14597 2301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14597 2301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14515 2301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14515 2301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14433 2301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14433 2301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14351 2301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14351 2301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14269 2301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14269 2301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14187 2301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14187 2301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14105 2301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14105 2301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 14023 2301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14023 2301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13941 2301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13941 2301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13859 2301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13859 2301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13777 2301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13777 2301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13695 2301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13695 2301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2237 13613 2301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13613 2301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4432 2284 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4346 2284 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4260 2284 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4174 2284 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4088 2284 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4002 2284 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3916 2284 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3830 2284 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3744 2284 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3658 2284 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3572 2284 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18527 2249 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18527 2249 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18445 2249 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18445 2249 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18363 2249 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18363 2249 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18281 2249 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18281 2249 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18199 2249 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18199 2249 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18117 2249 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18117 2249 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 18035 2249 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18035 2249 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17953 2249 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17953 2249 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17871 2249 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17871 2249 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17789 2249 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17789 2249 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17707 2249 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17707 2249 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17625 2249 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17625 2249 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17543 2249 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17543 2249 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17461 2249 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17461 2249 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17379 2249 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17379 2249 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17297 2249 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17297 2249 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17215 2249 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17215 2249 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17133 2249 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17133 2249 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 17051 2249 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17051 2249 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16969 2249 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16969 2249 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16887 2249 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16887 2249 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16805 2249 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16805 2249 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16723 2249 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16723 2249 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16641 2249 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16641 2249 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2185 16559 2249 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16559 2249 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16460 2221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16460 2221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16379 2221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16379 2221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16298 2221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16298 2221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16217 2221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16217 2221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16136 2221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16136 2221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 16055 2221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16055 2221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15974 2221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15974 2221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15893 2221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15893 2221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15812 2221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15812 2221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15731 2221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15731 2221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15650 2221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15650 2221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15569 2221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15569 2221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15488 2221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15488 2221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15407 2221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15407 2221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15326 2221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15326 2221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15245 2221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15245 2221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15164 2221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15164 2221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15083 2221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15083 2221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 15002 2221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15002 2221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14921 2221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14921 2221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14840 2221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14840 2221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14759 2221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14759 2221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14678 2221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14678 2221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14597 2221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14597 2221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14515 2221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14515 2221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14433 2221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14433 2221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14351 2221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14351 2221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14269 2221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14269 2221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14187 2221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14187 2221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14105 2221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14105 2221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 14023 2221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14023 2221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13941 2221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13941 2221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13859 2221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13859 2221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13777 2221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13777 2221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13695 2221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13695 2221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2157 13613 2221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13613 2221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4432 2203 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4346 2203 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4260 2203 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4174 2203 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4088 2203 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4002 2203 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3916 2203 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3830 2203 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3744 2203 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3658 2203 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3572 2203 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18527 2167 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18527 2167 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18445 2167 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18445 2167 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18363 2167 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18363 2167 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18281 2167 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18281 2167 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18199 2167 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18199 2167 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18117 2167 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18117 2167 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 18035 2167 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18035 2167 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17953 2167 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17953 2167 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17871 2167 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17871 2167 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17789 2167 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17789 2167 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17707 2167 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17707 2167 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17625 2167 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17625 2167 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17543 2167 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17543 2167 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17461 2167 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17461 2167 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17379 2167 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17379 2167 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17297 2167 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17297 2167 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17215 2167 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17215 2167 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17133 2167 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17133 2167 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 17051 2167 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17051 2167 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16969 2167 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16969 2167 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16887 2167 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16887 2167 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16805 2167 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16805 2167 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16723 2167 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16723 2167 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16641 2167 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16641 2167 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2103 16559 2167 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16559 2167 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16460 2141 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16460 2141 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16379 2141 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16379 2141 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16298 2141 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16298 2141 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16217 2141 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16217 2141 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16136 2141 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16136 2141 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 16055 2141 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16055 2141 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15974 2141 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15974 2141 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15893 2141 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15893 2141 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15812 2141 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15812 2141 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15731 2141 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15731 2141 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15650 2141 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15650 2141 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15569 2141 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15569 2141 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15488 2141 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15488 2141 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15407 2141 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15407 2141 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15326 2141 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15326 2141 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15245 2141 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15245 2141 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15164 2141 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15164 2141 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15083 2141 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15083 2141 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 15002 2141 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15002 2141 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14921 2141 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14921 2141 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14840 2141 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14840 2141 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14759 2141 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14759 2141 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14678 2141 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14678 2141 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14597 2141 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14597 2141 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14515 2141 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14515 2141 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14433 2141 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14433 2141 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14351 2141 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14351 2141 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14269 2141 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14269 2141 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14187 2141 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14187 2141 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14105 2141 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14105 2141 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 14023 2141 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14023 2141 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13941 2141 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13941 2141 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13859 2141 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13859 2141 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13777 2141 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13777 2141 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13695 2141 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13695 2141 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2077 13613 2141 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13613 2141 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4432 2122 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4346 2122 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4260 2122 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4174 2122 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4088 2122 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4002 2122 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3916 2122 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3830 2122 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3744 2122 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3658 2122 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3572 2122 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18527 2085 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18527 2085 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18445 2085 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18445 2085 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18363 2085 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18363 2085 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18281 2085 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18281 2085 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18199 2085 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18199 2085 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18117 2085 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18117 2085 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 18035 2085 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18035 2085 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17953 2085 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17953 2085 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17871 2085 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17871 2085 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17789 2085 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17789 2085 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17707 2085 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17707 2085 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17625 2085 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17625 2085 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17543 2085 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17543 2085 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17461 2085 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17461 2085 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17379 2085 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17379 2085 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17297 2085 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17297 2085 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17215 2085 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17215 2085 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17133 2085 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17133 2085 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 17051 2085 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17051 2085 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16969 2085 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16969 2085 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16887 2085 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16887 2085 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16805 2085 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16805 2085 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16723 2085 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16723 2085 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16641 2085 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16641 2085 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2021 16559 2085 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16559 2085 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16460 2061 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16460 2061 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16379 2061 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16379 2061 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16298 2061 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16298 2061 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16217 2061 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16217 2061 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16136 2061 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16136 2061 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 16055 2061 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16055 2061 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15974 2061 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15974 2061 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15893 2061 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15893 2061 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15812 2061 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15812 2061 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15731 2061 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15731 2061 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15650 2061 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15650 2061 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15569 2061 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15569 2061 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15488 2061 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15488 2061 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15407 2061 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15407 2061 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15326 2061 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15326 2061 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15245 2061 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15245 2061 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15164 2061 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15164 2061 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15083 2061 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15083 2061 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 15002 2061 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15002 2061 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14921 2061 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14921 2061 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14840 2061 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14840 2061 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14759 2061 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14759 2061 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14678 2061 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14678 2061 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14597 2061 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14597 2061 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14515 2061 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14515 2061 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14433 2061 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14433 2061 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14351 2061 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14351 2061 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14269 2061 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14269 2061 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14187 2061 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14187 2061 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14105 2061 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14105 2061 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 14023 2061 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14023 2061 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13941 2061 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13941 2061 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13859 2061 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13859 2061 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13777 2061 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13777 2061 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13695 2061 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13695 2061 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1997 13613 2061 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13613 2061 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4432 2041 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4346 2041 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4260 2041 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4174 2041 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4088 2041 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4002 2041 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3916 2041 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3830 2041 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3744 2041 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3658 2041 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3572 2041 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18527 2003 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18527 2003 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18445 2003 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18445 2003 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18363 2003 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18363 2003 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18281 2003 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18281 2003 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18199 2003 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18199 2003 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18117 2003 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18117 2003 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 18035 2003 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18035 2003 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17953 2003 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17953 2003 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17871 2003 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17871 2003 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17789 2003 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17789 2003 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17707 2003 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17707 2003 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17625 2003 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17625 2003 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17543 2003 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17543 2003 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17461 2003 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17461 2003 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17379 2003 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17379 2003 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17297 2003 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17297 2003 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17215 2003 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17215 2003 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17133 2003 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17133 2003 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 17051 2003 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17051 2003 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16969 2003 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16969 2003 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16887 2003 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16887 2003 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16805 2003 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16805 2003 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16723 2003 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16723 2003 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16641 2003 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16641 2003 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1939 16559 2003 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16559 2003 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16460 1981 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16460 1981 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16379 1981 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16379 1981 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16298 1981 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16298 1981 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16217 1981 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16217 1981 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16136 1981 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16136 1981 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 16055 1981 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16055 1981 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15974 1981 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15974 1981 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15893 1981 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15893 1981 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15812 1981 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15812 1981 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15731 1981 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15731 1981 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15650 1981 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15650 1981 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15569 1981 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15569 1981 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15488 1981 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15488 1981 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15407 1981 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15407 1981 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15326 1981 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15326 1981 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15245 1981 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15245 1981 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15164 1981 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15164 1981 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15083 1981 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15083 1981 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 15002 1981 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15002 1981 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14921 1981 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14921 1981 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14840 1981 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14840 1981 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14759 1981 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14759 1981 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14678 1981 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14678 1981 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14597 1981 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14597 1981 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14515 1981 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14515 1981 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14433 1981 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14433 1981 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14351 1981 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14351 1981 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14269 1981 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14269 1981 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14187 1981 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14187 1981 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14105 1981 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14105 1981 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 14023 1981 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14023 1981 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13941 1981 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13941 1981 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13859 1981 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13859 1981 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13777 1981 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13777 1981 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13695 1981 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13695 1981 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1917 13613 1981 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13613 1981 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4432 1960 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4346 1960 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4260 1960 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4174 1960 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4088 1960 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4002 1960 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3916 1960 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3830 1960 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3744 1960 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3658 1960 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3572 1960 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18527 1921 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18527 1921 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18445 1921 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18445 1921 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18363 1921 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18363 1921 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18281 1921 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18281 1921 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18199 1921 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18199 1921 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18117 1921 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18117 1921 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 18035 1921 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18035 1921 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17953 1921 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17953 1921 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17871 1921 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17871 1921 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17789 1921 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17789 1921 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17707 1921 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17707 1921 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17625 1921 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17625 1921 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17543 1921 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17543 1921 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17461 1921 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17461 1921 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17379 1921 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17379 1921 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17297 1921 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17297 1921 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17215 1921 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17215 1921 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17133 1921 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17133 1921 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 17051 1921 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17051 1921 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16969 1921 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16969 1921 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16887 1921 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16887 1921 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16805 1921 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16805 1921 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16723 1921 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16723 1921 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16641 1921 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16641 1921 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1857 16559 1921 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16559 1921 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16460 1901 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16460 1901 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16379 1901 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16379 1901 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16298 1901 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16298 1901 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16217 1901 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16217 1901 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16136 1901 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16136 1901 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 16055 1901 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16055 1901 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15974 1901 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15974 1901 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15893 1901 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15893 1901 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15812 1901 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15812 1901 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15731 1901 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15731 1901 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15650 1901 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15650 1901 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15569 1901 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15569 1901 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15488 1901 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15488 1901 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15407 1901 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15407 1901 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15326 1901 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15326 1901 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15245 1901 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15245 1901 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15164 1901 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15164 1901 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15083 1901 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15083 1901 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 15002 1901 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15002 1901 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14921 1901 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14921 1901 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14840 1901 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14840 1901 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14759 1901 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14759 1901 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14678 1901 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14678 1901 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14597 1901 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14597 1901 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14515 1901 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14515 1901 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14433 1901 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14433 1901 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14351 1901 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14351 1901 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14269 1901 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14269 1901 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14187 1901 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14187 1901 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14105 1901 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14105 1901 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 14023 1901 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14023 1901 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13941 1901 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13941 1901 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13859 1901 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13859 1901 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13777 1901 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13777 1901 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13695 1901 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13695 1901 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1837 13613 1901 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13613 1901 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4432 1879 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4346 1879 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4260 1879 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4174 1879 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4088 1879 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4002 1879 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3916 1879 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3830 1879 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3744 1879 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3658 1879 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3572 1879 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18527 1839 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18527 1839 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18445 1839 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18445 1839 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18363 1839 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18363 1839 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18281 1839 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18281 1839 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18199 1839 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18199 1839 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18117 1839 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18117 1839 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 18035 1839 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18035 1839 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17953 1839 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17953 1839 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17871 1839 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17871 1839 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17789 1839 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17789 1839 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17707 1839 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17707 1839 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17625 1839 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17625 1839 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17543 1839 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17543 1839 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17461 1839 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17461 1839 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17379 1839 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17379 1839 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17297 1839 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17297 1839 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17215 1839 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17215 1839 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17133 1839 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17133 1839 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 17051 1839 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17051 1839 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16969 1839 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16969 1839 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16887 1839 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16887 1839 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16805 1839 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16805 1839 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16723 1839 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16723 1839 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16641 1839 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16641 1839 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1775 16559 1839 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16559 1839 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16460 1821 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16460 1821 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16379 1821 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16379 1821 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16298 1821 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16298 1821 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16217 1821 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16217 1821 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16136 1821 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16136 1821 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 16055 1821 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16055 1821 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15974 1821 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15974 1821 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15893 1821 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15893 1821 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15812 1821 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15812 1821 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15731 1821 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15731 1821 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15650 1821 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15650 1821 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15569 1821 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15569 1821 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15488 1821 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15488 1821 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15407 1821 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15407 1821 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15326 1821 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15326 1821 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15245 1821 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15245 1821 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15164 1821 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15164 1821 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15083 1821 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15083 1821 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 15002 1821 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15002 1821 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14921 1821 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14921 1821 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14840 1821 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14840 1821 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14759 1821 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14759 1821 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14678 1821 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14678 1821 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14597 1821 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14597 1821 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14515 1821 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14515 1821 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14433 1821 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14433 1821 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14351 1821 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14351 1821 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14269 1821 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14269 1821 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14187 1821 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14187 1821 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14105 1821 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14105 1821 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 14023 1821 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14023 1821 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13941 1821 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13941 1821 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13859 1821 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13859 1821 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13777 1821 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13777 1821 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13695 1821 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13695 1821 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1757 13613 1821 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13613 1821 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4432 1798 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4346 1798 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4260 1798 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4174 1798 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4088 1798 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4002 1798 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3916 1798 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3830 1798 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3744 1798 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3658 1798 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3572 1798 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18527 1757 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18527 1757 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18445 1757 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18445 1757 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18363 1757 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18363 1757 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18281 1757 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18281 1757 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18199 1757 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18199 1757 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18117 1757 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18117 1757 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 18035 1757 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18035 1757 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17953 1757 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17953 1757 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17871 1757 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17871 1757 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17789 1757 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17789 1757 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17707 1757 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17707 1757 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17625 1757 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17625 1757 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17543 1757 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17543 1757 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17461 1757 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17461 1757 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17379 1757 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17379 1757 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17297 1757 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17297 1757 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17215 1757 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17215 1757 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17133 1757 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17133 1757 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 17051 1757 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17051 1757 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16969 1757 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16969 1757 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16887 1757 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16887 1757 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16805 1757 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16805 1757 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16723 1757 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16723 1757 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16641 1757 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16641 1757 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1693 16559 1757 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16559 1757 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16460 1741 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16460 1741 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16379 1741 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16379 1741 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16298 1741 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16298 1741 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16217 1741 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16217 1741 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16136 1741 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16136 1741 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 16055 1741 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16055 1741 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15974 1741 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15974 1741 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15893 1741 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15893 1741 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15812 1741 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15812 1741 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15731 1741 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15731 1741 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15650 1741 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15650 1741 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15569 1741 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15569 1741 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15488 1741 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15488 1741 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15407 1741 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15407 1741 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15326 1741 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15326 1741 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15245 1741 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15245 1741 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15164 1741 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15164 1741 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15083 1741 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15083 1741 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 15002 1741 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15002 1741 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14921 1741 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14921 1741 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14840 1741 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14840 1741 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14759 1741 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14759 1741 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14678 1741 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14678 1741 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14597 1741 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14597 1741 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14515 1741 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14515 1741 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14433 1741 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14433 1741 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14351 1741 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14351 1741 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14269 1741 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14269 1741 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14187 1741 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14187 1741 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14105 1741 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14105 1741 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 14023 1741 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14023 1741 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13941 1741 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13941 1741 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13859 1741 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13859 1741 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13777 1741 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13777 1741 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13695 1741 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13695 1741 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1677 13613 1741 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13613 1741 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4432 1717 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4346 1717 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4260 1717 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4174 1717 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4088 1717 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4002 1717 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3916 1717 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3830 1717 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3744 1717 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3658 1717 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3572 1717 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18527 1675 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18527 1675 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18445 1675 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18445 1675 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18363 1675 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18363 1675 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18281 1675 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18281 1675 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18199 1675 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18199 1675 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18117 1675 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18117 1675 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 18035 1675 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18035 1675 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17953 1675 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17953 1675 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17871 1675 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17871 1675 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17789 1675 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17789 1675 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17707 1675 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17707 1675 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17625 1675 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17625 1675 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17543 1675 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17543 1675 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17461 1675 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17461 1675 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17379 1675 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17379 1675 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17297 1675 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17297 1675 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17215 1675 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17215 1675 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17133 1675 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17133 1675 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 17051 1675 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17051 1675 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16969 1675 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16969 1675 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16887 1675 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16887 1675 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16805 1675 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16805 1675 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16723 1675 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16723 1675 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16641 1675 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16641 1675 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1611 16559 1675 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16559 1675 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16460 1661 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16460 1661 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16379 1661 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16379 1661 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16298 1661 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16298 1661 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16217 1661 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16217 1661 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16136 1661 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16136 1661 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 16055 1661 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16055 1661 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15974 1661 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15974 1661 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15893 1661 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15893 1661 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15812 1661 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15812 1661 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15731 1661 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15731 1661 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15650 1661 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15650 1661 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15569 1661 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15569 1661 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15488 1661 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15488 1661 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15407 1661 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15407 1661 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15326 1661 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15326 1661 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15245 1661 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15245 1661 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15164 1661 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15164 1661 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15083 1661 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15083 1661 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 15002 1661 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15002 1661 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14921 1661 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14921 1661 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14840 1661 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14840 1661 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14759 1661 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14759 1661 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14678 1661 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14678 1661 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14597 1661 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14597 1661 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14515 1661 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14515 1661 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14433 1661 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14433 1661 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14351 1661 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14351 1661 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14269 1661 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14269 1661 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14187 1661 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14187 1661 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14105 1661 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14105 1661 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 14023 1661 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14023 1661 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13941 1661 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13941 1661 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13859 1661 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13859 1661 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13777 1661 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13777 1661 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13695 1661 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13695 1661 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1597 13613 1661 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13613 1661 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4432 1636 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4346 1636 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4260 1636 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4174 1636 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4088 1636 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4002 1636 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3916 1636 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3830 1636 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3744 1636 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3658 1636 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3572 1636 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18527 1593 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18527 1593 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18445 1593 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18445 1593 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18363 1593 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18363 1593 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18281 1593 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18281 1593 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18199 1593 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18199 1593 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18117 1593 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18117 1593 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 18035 1593 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18035 1593 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17953 1593 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17953 1593 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17871 1593 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17871 1593 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17789 1593 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17789 1593 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17707 1593 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17707 1593 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17625 1593 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17625 1593 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17543 1593 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17543 1593 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17461 1593 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17461 1593 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17379 1593 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17379 1593 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17297 1593 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17297 1593 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17215 1593 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17215 1593 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17133 1593 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17133 1593 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 17051 1593 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17051 1593 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16969 1593 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16969 1593 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16887 1593 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16887 1593 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16805 1593 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16805 1593 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16723 1593 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16723 1593 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16641 1593 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16641 1593 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1529 16559 1593 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16559 1593 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16460 1581 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16460 1581 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16379 1581 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16379 1581 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16298 1581 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16298 1581 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16217 1581 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16217 1581 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16136 1581 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16136 1581 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 16055 1581 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16055 1581 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15974 1581 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15974 1581 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15893 1581 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15893 1581 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15812 1581 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15812 1581 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15731 1581 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15731 1581 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15650 1581 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15650 1581 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15569 1581 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15569 1581 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15488 1581 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15488 1581 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15407 1581 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15407 1581 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15326 1581 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15326 1581 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15245 1581 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15245 1581 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15164 1581 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15164 1581 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15083 1581 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15083 1581 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 15002 1581 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15002 1581 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14921 1581 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14921 1581 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14840 1581 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14840 1581 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14759 1581 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14759 1581 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14678 1581 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14678 1581 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14597 1581 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14597 1581 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14515 1581 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14515 1581 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14433 1581 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14433 1581 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14351 1581 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14351 1581 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14269 1581 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14269 1581 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14187 1581 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14187 1581 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14105 1581 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14105 1581 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 14023 1581 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14023 1581 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13941 1581 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13941 1581 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13859 1581 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13859 1581 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13777 1581 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13777 1581 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13695 1581 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13695 1581 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1517 13613 1581 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13613 1581 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4432 1555 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4346 1555 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4260 1555 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4174 1555 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4088 1555 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4002 1555 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3916 1555 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3830 1555 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3744 1555 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3658 1555 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3572 1555 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18527 1511 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18527 1511 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18445 1511 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18445 1511 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18363 1511 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18363 1511 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18281 1511 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18281 1511 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18199 1511 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18199 1511 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18117 1511 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18117 1511 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 18035 1511 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18035 1511 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17953 1511 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17953 1511 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17871 1511 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17871 1511 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17789 1511 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17789 1511 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17707 1511 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17707 1511 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17625 1511 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17625 1511 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17543 1511 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17543 1511 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17461 1511 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17461 1511 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17379 1511 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17379 1511 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17297 1511 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17297 1511 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17215 1511 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17215 1511 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17133 1511 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17133 1511 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 17051 1511 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17051 1511 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16969 1511 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16969 1511 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16887 1511 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16887 1511 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16805 1511 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16805 1511 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16723 1511 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16723 1511 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16641 1511 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16641 1511 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1447 16559 1511 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16559 1511 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16460 1501 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16460 1501 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16379 1501 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16379 1501 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16298 1501 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16298 1501 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16217 1501 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16217 1501 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16136 1501 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16136 1501 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 16055 1501 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16055 1501 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15974 1501 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15974 1501 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15893 1501 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15893 1501 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15812 1501 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15812 1501 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15731 1501 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15731 1501 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15650 1501 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15650 1501 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15569 1501 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15569 1501 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15488 1501 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15488 1501 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15407 1501 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15407 1501 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15326 1501 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15326 1501 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15245 1501 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15245 1501 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15164 1501 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15164 1501 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15083 1501 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15083 1501 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 15002 1501 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15002 1501 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14921 1501 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14921 1501 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14840 1501 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14840 1501 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14759 1501 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14759 1501 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14678 1501 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14678 1501 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14597 1501 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14597 1501 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14515 1501 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14515 1501 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14433 1501 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14433 1501 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14351 1501 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14351 1501 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14269 1501 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14269 1501 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14187 1501 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14187 1501 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14105 1501 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14105 1501 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 14023 1501 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14023 1501 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13941 1501 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13941 1501 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13859 1501 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13859 1501 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13777 1501 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13777 1501 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13695 1501 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13695 1501 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1437 13613 1501 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13613 1501 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4432 1474 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4346 1474 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4260 1474 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4174 1474 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4088 1474 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4002 1474 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3916 1474 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3830 1474 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3744 1474 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3658 1474 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3572 1474 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18527 1429 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18527 1429 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18445 1429 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18445 1429 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18363 1429 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18363 1429 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18281 1429 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18281 1429 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18199 1429 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18199 1429 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18117 1429 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18117 1429 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 18035 1429 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18035 1429 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17953 1429 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17953 1429 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17871 1429 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17871 1429 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17789 1429 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17789 1429 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17707 1429 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17707 1429 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17625 1429 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17625 1429 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17543 1429 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17543 1429 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17461 1429 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17461 1429 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17379 1429 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17379 1429 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17297 1429 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17297 1429 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17215 1429 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17215 1429 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17133 1429 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17133 1429 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 17051 1429 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17051 1429 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16969 1429 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16969 1429 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16887 1429 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16887 1429 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16805 1429 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16805 1429 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16723 1429 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16723 1429 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16641 1429 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16641 1429 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1365 16559 1429 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16559 1429 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16460 1421 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16460 1421 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16379 1421 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16379 1421 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16298 1421 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16298 1421 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16217 1421 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16217 1421 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16136 1421 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16136 1421 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 16055 1421 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16055 1421 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15974 1421 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15974 1421 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15893 1421 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15893 1421 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15812 1421 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15812 1421 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15731 1421 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15731 1421 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15650 1421 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15650 1421 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15569 1421 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15569 1421 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15488 1421 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15488 1421 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15407 1421 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15407 1421 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15326 1421 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15326 1421 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15245 1421 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15245 1421 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15164 1421 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15164 1421 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15083 1421 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15083 1421 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 15002 1421 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15002 1421 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14921 1421 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14921 1421 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14840 1421 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14840 1421 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14759 1421 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14759 1421 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14678 1421 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14678 1421 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14597 1421 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14597 1421 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14515 1421 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14515 1421 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14433 1421 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14433 1421 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14351 1421 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14351 1421 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14269 1421 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14269 1421 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14187 1421 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14187 1421 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14105 1421 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14105 1421 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 14023 1421 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14023 1421 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13941 1421 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13941 1421 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13859 1421 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13859 1421 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13777 1421 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13777 1421 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13695 1421 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13695 1421 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1357 13613 1421 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13613 1421 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4432 1393 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4346 1393 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4260 1393 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4174 1393 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4088 1393 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4002 1393 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3916 1393 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3830 1393 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3744 1393 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3658 1393 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3572 1393 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18527 1347 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18527 1347 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18445 1347 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18445 1347 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18363 1347 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18363 1347 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18281 1347 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18281 1347 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18199 1347 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18199 1347 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18117 1347 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18117 1347 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 18035 1347 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18035 1347 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17953 1347 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17953 1347 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17871 1347 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17871 1347 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17789 1347 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17789 1347 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17707 1347 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17707 1347 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17625 1347 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17625 1347 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17543 1347 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17543 1347 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17461 1347 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17461 1347 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17379 1347 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17379 1347 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17297 1347 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17297 1347 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17215 1347 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17215 1347 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17133 1347 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17133 1347 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 17051 1347 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17051 1347 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16969 1347 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16969 1347 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16887 1347 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16887 1347 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16805 1347 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16805 1347 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16723 1347 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16723 1347 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16641 1347 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16641 1347 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1283 16559 1347 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16559 1347 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16460 1341 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16460 1341 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16379 1341 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16379 1341 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16298 1341 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16298 1341 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16217 1341 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16217 1341 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16136 1341 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16136 1341 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 16055 1341 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16055 1341 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15974 1341 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15974 1341 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15893 1341 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15893 1341 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15812 1341 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15812 1341 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15731 1341 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15731 1341 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15650 1341 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15650 1341 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15569 1341 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15569 1341 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15488 1341 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15488 1341 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15407 1341 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15407 1341 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15326 1341 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15326 1341 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15245 1341 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15245 1341 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15164 1341 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15164 1341 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15083 1341 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15083 1341 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 15002 1341 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15002 1341 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14921 1341 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14921 1341 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14840 1341 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14840 1341 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14759 1341 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14759 1341 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14678 1341 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14678 1341 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14597 1341 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14597 1341 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14515 1341 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14515 1341 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14433 1341 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14433 1341 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14351 1341 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14351 1341 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14269 1341 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14269 1341 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14187 1341 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14187 1341 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14105 1341 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14105 1341 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 14023 1341 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14023 1341 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13941 1341 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13941 1341 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13859 1341 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13859 1341 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13777 1341 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13777 1341 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13695 1341 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13695 1341 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1277 13613 1341 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13613 1341 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4432 1312 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4346 1312 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4260 1312 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4174 1312 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4088 1312 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4002 1312 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3916 1312 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3830 1312 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3744 1312 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3658 1312 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3572 1312 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18527 1265 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18527 1265 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18445 1265 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18445 1265 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18363 1265 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18363 1265 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18281 1265 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18281 1265 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18199 1265 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18199 1265 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18117 1265 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18117 1265 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 18035 1265 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18035 1265 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17953 1265 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17953 1265 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17871 1265 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17871 1265 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17789 1265 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17789 1265 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17707 1265 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17707 1265 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17625 1265 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17625 1265 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17543 1265 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17543 1265 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17461 1265 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17461 1265 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17379 1265 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17379 1265 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17297 1265 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17297 1265 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17215 1265 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17215 1265 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17133 1265 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17133 1265 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 17051 1265 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17051 1265 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16969 1265 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16969 1265 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16887 1265 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16887 1265 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16805 1265 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16805 1265 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16723 1265 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16723 1265 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16641 1265 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16641 1265 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1201 16559 1265 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16559 1265 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16460 1261 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16460 1261 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16379 1261 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16379 1261 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16298 1261 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16298 1261 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16217 1261 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16217 1261 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16136 1261 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16136 1261 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 16055 1261 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16055 1261 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15974 1261 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15974 1261 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15893 1261 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15893 1261 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15812 1261 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15812 1261 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15731 1261 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15731 1261 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15650 1261 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15650 1261 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15569 1261 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15569 1261 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15488 1261 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15488 1261 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15407 1261 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15407 1261 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15326 1261 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15326 1261 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15245 1261 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15245 1261 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15164 1261 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15164 1261 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15083 1261 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15083 1261 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 15002 1261 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15002 1261 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14921 1261 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14921 1261 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14840 1261 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14840 1261 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14759 1261 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14759 1261 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14678 1261 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14678 1261 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14597 1261 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14597 1261 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14515 1261 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14515 1261 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14433 1261 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14433 1261 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14351 1261 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14351 1261 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14269 1261 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14269 1261 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14187 1261 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14187 1261 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14105 1261 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14105 1261 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 14023 1261 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14023 1261 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13941 1261 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13941 1261 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13859 1261 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13859 1261 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13777 1261 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13777 1261 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13695 1261 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13695 1261 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1197 13613 1261 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13613 1261 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4432 1231 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4346 1231 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4260 1231 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4174 1231 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4088 1231 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4002 1231 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3916 1231 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3830 1231 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3744 1231 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3658 1231 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3572 1231 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18527 1183 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18527 1183 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18445 1183 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18445 1183 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18363 1183 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18363 1183 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18281 1183 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18281 1183 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18199 1183 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18199 1183 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18117 1183 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18117 1183 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 18035 1183 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18035 1183 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17953 1183 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17953 1183 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17871 1183 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17871 1183 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17789 1183 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17789 1183 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17707 1183 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17707 1183 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17625 1183 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17625 1183 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17543 1183 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17543 1183 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17461 1183 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17461 1183 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17379 1183 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17379 1183 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17297 1183 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17297 1183 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17215 1183 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17215 1183 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17133 1183 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17133 1183 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 17051 1183 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17051 1183 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16969 1183 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16969 1183 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16887 1183 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16887 1183 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16805 1183 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16805 1183 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16723 1183 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16723 1183 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16641 1183 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16641 1183 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1119 16559 1183 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16559 1183 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16460 1181 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16460 1181 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16379 1181 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16379 1181 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16298 1181 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16298 1181 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16217 1181 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16217 1181 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16136 1181 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16136 1181 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 16055 1181 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16055 1181 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15974 1181 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15974 1181 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15893 1181 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15893 1181 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15812 1181 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15812 1181 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15731 1181 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15731 1181 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15650 1181 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15650 1181 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15569 1181 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15569 1181 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15488 1181 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15488 1181 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15407 1181 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15407 1181 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15326 1181 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15326 1181 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15245 1181 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15245 1181 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15164 1181 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15164 1181 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15083 1181 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15083 1181 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 15002 1181 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15002 1181 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14921 1181 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14921 1181 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14840 1181 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14840 1181 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14759 1181 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14759 1181 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14678 1181 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14678 1181 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14597 1181 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14597 1181 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14515 1181 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14515 1181 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14433 1181 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14433 1181 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14351 1181 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14351 1181 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14269 1181 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14269 1181 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14187 1181 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14187 1181 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14105 1181 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14105 1181 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 14023 1181 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14023 1181 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13941 1181 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13941 1181 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13859 1181 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13859 1181 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13777 1181 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13777 1181 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13695 1181 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13695 1181 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1117 13613 1181 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13613 1181 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4432 1150 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4346 1150 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4260 1150 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4174 1150 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4088 1150 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4002 1150 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3916 1150 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3830 1150 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3744 1150 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3658 1150 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3572 1150 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18527 1101 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18527 1101 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18445 1101 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18445 1101 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18363 1101 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18363 1101 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18281 1101 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18281 1101 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18199 1101 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18199 1101 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18117 1101 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18117 1101 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 18035 1101 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18035 1101 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17953 1101 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17953 1101 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17871 1101 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17871 1101 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17789 1101 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17789 1101 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17707 1101 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17707 1101 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17625 1101 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17625 1101 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17543 1101 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17543 1101 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17461 1101 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17461 1101 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17379 1101 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17379 1101 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17297 1101 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17297 1101 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17215 1101 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17215 1101 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17133 1101 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17133 1101 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 17051 1101 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17051 1101 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16969 1101 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16969 1101 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16887 1101 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16887 1101 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16805 1101 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16805 1101 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16723 1101 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16723 1101 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16641 1101 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16641 1101 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16559 1101 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16559 1101 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16460 1101 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16460 1101 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16379 1101 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16379 1101 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16298 1101 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16298 1101 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16217 1101 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16217 1101 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16136 1101 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16136 1101 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 16055 1101 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16055 1101 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15974 1101 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15974 1101 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15893 1101 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15893 1101 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15812 1101 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15812 1101 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15731 1101 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15731 1101 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15650 1101 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15650 1101 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15569 1101 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15569 1101 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15488 1101 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15488 1101 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15407 1101 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15407 1101 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15326 1101 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15326 1101 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15245 1101 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15245 1101 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15164 1101 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15164 1101 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15083 1101 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15083 1101 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 15002 1101 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15002 1101 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14921 1101 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14921 1101 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14840 1101 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14840 1101 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14759 1101 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14759 1101 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14678 1101 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14678 1101 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14597 1101 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14597 1101 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14515 1101 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14515 1101 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14433 1101 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14433 1101 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14351 1101 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14351 1101 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14269 1101 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14269 1101 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14187 1101 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14187 1101 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14105 1101 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14105 1101 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 14023 1101 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14023 1101 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13941 1101 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13941 1101 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13859 1101 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13859 1101 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13777 1101 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13777 1101 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13695 1101 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13695 1101 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 1037 13613 1101 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13613 1101 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4432 1069 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4346 1069 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4260 1069 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4174 1069 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4088 1069 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4002 1069 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3916 1069 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3830 1069 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3744 1069 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3658 1069 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3572 1069 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16460 1021 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16460 1021 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16379 1021 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16379 1021 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16298 1021 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16298 1021 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16217 1021 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16217 1021 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16136 1021 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16136 1021 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 16055 1021 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16055 1021 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15974 1021 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15974 1021 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15893 1021 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15893 1021 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15812 1021 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15812 1021 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15731 1021 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15731 1021 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15650 1021 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15650 1021 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15569 1021 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15569 1021 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15488 1021 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15488 1021 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15407 1021 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15407 1021 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15326 1021 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15326 1021 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15245 1021 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15245 1021 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15164 1021 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15164 1021 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15083 1021 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15083 1021 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 15002 1021 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15002 1021 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14921 1021 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14921 1021 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14840 1021 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14840 1021 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14759 1021 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14759 1021 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14678 1021 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14678 1021 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14597 1021 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14597 1021 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14515 1021 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14515 1021 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14433 1021 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14433 1021 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14351 1021 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14351 1021 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14269 1021 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14269 1021 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14187 1021 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14187 1021 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14105 1021 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14105 1021 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 14023 1021 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14023 1021 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13941 1021 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13941 1021 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13859 1021 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13859 1021 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13777 1021 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13777 1021 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13695 1021 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13695 1021 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 957 13613 1021 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13613 1021 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18527 1019 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18527 1019 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18445 1019 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18445 1019 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18363 1019 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18363 1019 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18281 1019 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18281 1019 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18199 1019 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18199 1019 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18117 1019 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18117 1019 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 18035 1019 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18035 1019 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17953 1019 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17953 1019 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17871 1019 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17871 1019 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17789 1019 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17789 1019 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17707 1019 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17707 1019 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17625 1019 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17625 1019 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17543 1019 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17543 1019 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17461 1019 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17461 1019 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17379 1019 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17379 1019 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17297 1019 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17297 1019 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17215 1019 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17215 1019 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17133 1019 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17133 1019 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 17051 1019 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17051 1019 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16969 1019 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16969 1019 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16887 1019 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16887 1019 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16805 1019 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16805 1019 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16723 1019 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16723 1019 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16641 1019 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16641 1019 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 955 16559 1019 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16559 1019 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4432 988 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4346 988 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4260 988 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4174 988 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4088 988 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4002 988 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3916 988 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3830 988 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3744 988 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3658 988 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3572 988 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16460 941 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16460 941 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16379 941 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16379 941 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16298 941 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16298 941 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16217 941 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16217 941 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16136 941 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16136 941 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 16055 941 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16055 941 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15974 941 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15974 941 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15893 941 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15893 941 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15812 941 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15812 941 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15731 941 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15731 941 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15650 941 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15650 941 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15569 941 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15569 941 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15488 941 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15488 941 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15407 941 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15407 941 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15326 941 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15326 941 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15245 941 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15245 941 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15164 941 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15164 941 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15083 941 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15083 941 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 15002 941 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15002 941 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14921 941 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14921 941 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14840 941 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14840 941 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14759 941 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14759 941 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14678 941 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14678 941 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14597 941 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14597 941 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14515 941 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14515 941 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14433 941 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14433 941 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14351 941 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14351 941 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14269 941 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14269 941 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14187 941 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14187 941 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14105 941 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14105 941 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 14023 941 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14023 941 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13941 941 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13941 941 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13859 941 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13859 941 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13777 941 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13777 941 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13695 941 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13695 941 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 877 13613 941 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13613 941 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18527 937 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18527 937 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18445 937 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18445 937 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18363 937 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18363 937 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18281 937 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18281 937 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18199 937 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18199 937 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18117 937 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18117 937 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 18035 937 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18035 937 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17953 937 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17953 937 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17871 937 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17871 937 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17789 937 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17789 937 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17707 937 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17707 937 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17625 937 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17625 937 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17543 937 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17543 937 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17461 937 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17461 937 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17379 937 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17379 937 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17297 937 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17297 937 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17215 937 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17215 937 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17133 937 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17133 937 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 17051 937 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17051 937 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16969 937 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16969 937 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16887 937 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16887 937 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16805 937 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16805 937 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16723 937 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16723 937 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16641 937 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16641 937 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 873 16559 937 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16559 937 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4432 907 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4346 907 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4260 907 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4174 907 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4088 907 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4002 907 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3916 907 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3830 907 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3744 907 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3658 907 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3572 907 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16460 861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16460 861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16379 861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16379 861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16298 861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16298 861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16217 861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16217 861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16136 861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16136 861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 16055 861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16055 861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15974 861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15974 861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15893 861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15893 861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15812 861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15812 861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15731 861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15731 861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15650 861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15650 861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15569 861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15569 861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15488 861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15488 861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15407 861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15407 861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15326 861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15326 861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15245 861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15245 861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15164 861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15164 861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15083 861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15083 861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 15002 861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15002 861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14921 861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14921 861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14840 861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14840 861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14759 861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14759 861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14678 861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14678 861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14597 861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14597 861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14515 861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14515 861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14433 861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14433 861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14351 861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14351 861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14269 861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14269 861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14187 861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14187 861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14105 861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14105 861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 14023 861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14023 861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13941 861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13941 861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13859 861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13859 861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13777 861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13777 861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13695 861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13695 861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 797 13613 861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13613 861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18527 855 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18527 855 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18445 855 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18445 855 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18363 855 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18363 855 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18281 855 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18281 855 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18199 855 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18199 855 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18117 855 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18117 855 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 18035 855 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18035 855 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17953 855 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17953 855 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17871 855 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17871 855 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17789 855 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17789 855 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17707 855 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17707 855 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17625 855 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17625 855 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17543 855 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17543 855 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17461 855 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17461 855 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17379 855 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17379 855 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17297 855 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17297 855 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17215 855 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17215 855 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17133 855 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17133 855 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 17051 855 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17051 855 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16969 855 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16969 855 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16887 855 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16887 855 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16805 855 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16805 855 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16723 855 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16723 855 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16641 855 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16641 855 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 791 16559 855 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16559 855 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4432 826 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4346 826 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4260 826 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4174 826 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4088 826 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4002 826 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3916 826 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3830 826 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3744 826 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3658 826 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3572 826 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16460 781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16460 781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16379 781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16379 781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16298 781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16298 781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16217 781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16217 781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16136 781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16136 781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 16055 781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16055 781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15974 781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15974 781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15893 781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15893 781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15812 781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15812 781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15731 781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15731 781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15650 781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15650 781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15569 781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15569 781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15488 781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15488 781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15407 781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15407 781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15326 781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15326 781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15245 781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15245 781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15164 781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15164 781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15083 781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15083 781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 15002 781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15002 781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14921 781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14921 781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14840 781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14840 781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14759 781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14759 781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14678 781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14678 781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14597 781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14597 781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14515 781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14515 781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14433 781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14433 781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14351 781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14351 781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14269 781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14269 781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14187 781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14187 781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14105 781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14105 781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 14023 781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14023 781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13941 781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13941 781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13859 781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13859 781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13777 781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13777 781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13695 781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13695 781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 717 13613 781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13613 781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18527 773 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18527 773 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18445 773 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18445 773 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18363 773 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18363 773 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18281 773 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18281 773 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18199 773 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18199 773 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18117 773 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18117 773 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 18035 773 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18035 773 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17953 773 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17953 773 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17871 773 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17871 773 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17789 773 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17789 773 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17707 773 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17707 773 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17625 773 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17625 773 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17543 773 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17543 773 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17461 773 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17461 773 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17379 773 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17379 773 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17297 773 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17297 773 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17215 773 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17215 773 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17133 773 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17133 773 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 17051 773 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17051 773 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16969 773 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16969 773 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16887 773 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16887 773 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16805 773 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16805 773 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16723 773 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16723 773 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16641 773 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16641 773 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 709 16559 773 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16559 773 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4432 745 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4346 745 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4260 745 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4174 745 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4088 745 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4002 745 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3916 745 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3830 745 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3744 745 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3658 745 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3572 745 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16460 701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16460 701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16379 701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16379 701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16298 701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16298 701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16217 701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16217 701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16136 701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16136 701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 16055 701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16055 701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15974 701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15974 701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15893 701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15893 701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15812 701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15812 701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15731 701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15731 701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15650 701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15650 701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15569 701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15569 701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15488 701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15488 701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15407 701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15407 701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15326 701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15326 701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15245 701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15245 701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15164 701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15164 701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15083 701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15083 701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 15002 701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15002 701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14921 701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14921 701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14840 701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14840 701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14759 701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14759 701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14678 701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14678 701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14597 701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14597 701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14515 701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14515 701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14433 701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14433 701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14351 701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14351 701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14269 701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14269 701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14187 701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14187 701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14105 701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14105 701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 14023 701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14023 701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13941 701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13941 701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13859 701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13859 701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13777 701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13777 701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13695 701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13695 701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 637 13613 701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13613 701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18527 691 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18527 691 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18445 691 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18445 691 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18363 691 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18363 691 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18281 691 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18281 691 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18199 691 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18199 691 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18117 691 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18117 691 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 18035 691 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18035 691 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17953 691 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17953 691 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17871 691 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17871 691 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17789 691 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17789 691 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17707 691 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17707 691 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17625 691 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17625 691 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17543 691 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17543 691 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17461 691 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17461 691 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17379 691 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17379 691 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17297 691 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17297 691 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17215 691 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17215 691 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17133 691 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17133 691 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 17051 691 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17051 691 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16969 691 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16969 691 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16887 691 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16887 691 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16805 691 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16805 691 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16723 691 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16723 691 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16641 691 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16641 691 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 627 16559 691 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16559 691 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4432 664 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4346 664 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4260 664 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4174 664 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4088 664 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4002 664 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3916 664 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3830 664 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3744 664 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3658 664 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3572 664 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16460 621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16460 621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16379 621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16379 621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16298 621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16298 621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16217 621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16217 621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16136 621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16136 621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 16055 621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16055 621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15974 621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15974 621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15893 621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15893 621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15812 621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15812 621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15731 621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15731 621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15650 621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15650 621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15569 621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15569 621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15488 621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15488 621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15407 621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15407 621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15326 621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15326 621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15245 621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15245 621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15164 621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15164 621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15083 621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15083 621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 15002 621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15002 621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14921 621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14921 621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14840 621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14840 621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14759 621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14759 621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14678 621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14678 621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14597 621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14597 621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14515 621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14515 621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14433 621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14433 621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14351 621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14351 621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14269 621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14269 621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14187 621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14187 621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14105 621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14105 621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 14023 621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14023 621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13941 621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13941 621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13859 621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13859 621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13777 621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13777 621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13695 621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13695 621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 557 13613 621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13613 621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18527 609 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18527 609 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18445 609 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18445 609 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18363 609 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18363 609 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18281 609 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18281 609 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18199 609 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18199 609 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18117 609 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18117 609 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 18035 609 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18035 609 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17953 609 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17953 609 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17871 609 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17871 609 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17789 609 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17789 609 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17707 609 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17707 609 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17625 609 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17625 609 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17543 609 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17543 609 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17461 609 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17461 609 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17379 609 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17379 609 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17297 609 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17297 609 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17215 609 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17215 609 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17133 609 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17133 609 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 17051 609 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17051 609 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16969 609 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16969 609 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16887 609 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16887 609 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16805 609 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16805 609 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16723 609 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16723 609 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16641 609 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16641 609 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 545 16559 609 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16559 609 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4432 583 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4346 583 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4260 583 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4174 583 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4088 583 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4002 583 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3916 583 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3830 583 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3744 583 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3658 583 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3572 583 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16460 541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16460 541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16379 541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16379 541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16298 541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16298 541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16217 541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16217 541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16136 541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16136 541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 16055 541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16055 541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15974 541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15974 541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15893 541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15893 541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15812 541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15812 541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15731 541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15731 541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15650 541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15650 541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15569 541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15569 541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15488 541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15488 541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15407 541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15407 541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15326 541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15326 541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15245 541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15245 541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15164 541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15164 541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15083 541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15083 541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 15002 541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15002 541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14921 541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14921 541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14840 541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14840 541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14759 541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14759 541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14678 541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14678 541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14597 541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14597 541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14515 541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14515 541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14433 541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14433 541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14351 541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14351 541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14269 541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14269 541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14187 541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14187 541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14105 541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14105 541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 14023 541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14023 541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13941 541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13941 541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13859 541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13859 541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13777 541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13777 541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13695 541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13695 541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 477 13613 541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13613 541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18527 527 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18527 527 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18445 527 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18445 527 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18363 527 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18363 527 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18281 527 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18281 527 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18199 527 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18199 527 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18117 527 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18117 527 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 18035 527 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18035 527 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17953 527 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17953 527 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17871 527 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17871 527 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17789 527 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17789 527 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17707 527 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17707 527 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17625 527 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17625 527 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17543 527 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17543 527 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17461 527 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17461 527 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17379 527 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17379 527 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17297 527 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17297 527 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17215 527 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17215 527 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17133 527 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17133 527 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 17051 527 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17051 527 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16969 527 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16969 527 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16887 527 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16887 527 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16805 527 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16805 527 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16723 527 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16723 527 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16641 527 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16641 527 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 463 16559 527 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16559 527 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4432 502 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4346 502 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4260 502 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4174 502 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4088 502 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4002 502 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3916 502 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3830 502 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3744 502 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3658 502 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3572 502 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16460 461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16460 461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16379 461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16379 461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16298 461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16298 461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16217 461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16217 461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16136 461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16136 461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 16055 461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16055 461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15974 461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15974 461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15893 461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15893 461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15812 461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15812 461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15731 461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15731 461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15650 461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15650 461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15569 461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15569 461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15488 461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15488 461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15407 461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15407 461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15326 461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15326 461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15245 461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15245 461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15164 461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15164 461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15083 461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15083 461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 15002 461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15002 461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14921 461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14921 461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14840 461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14840 461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14759 461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14759 461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14678 461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14678 461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14597 461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14597 461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14515 461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14515 461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14433 461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14433 461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14351 461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14351 461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14269 461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14269 461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14187 461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14187 461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14105 461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14105 461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 14023 461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14023 461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13941 461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13941 461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13859 461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13859 461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13777 461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13777 461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13695 461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13695 461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 397 13613 461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13613 461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18527 445 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18527 445 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18445 445 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18445 445 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18363 445 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18363 445 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18281 445 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18281 445 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18199 445 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18199 445 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18117 445 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18117 445 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 18035 445 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18035 445 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17953 445 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17953 445 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17871 445 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17871 445 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17789 445 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17789 445 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17707 445 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17707 445 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17625 445 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17625 445 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17543 445 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17543 445 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17461 445 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17461 445 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17379 445 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17379 445 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17297 445 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17297 445 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17215 445 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17215 445 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17133 445 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17133 445 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 17051 445 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17051 445 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16969 445 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16969 445 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16887 445 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16887 445 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16805 445 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16805 445 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16723 445 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16723 445 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16641 445 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16641 445 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 381 16559 445 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16559 445 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4432 421 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4346 421 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4260 421 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4174 421 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4088 421 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4002 421 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3916 421 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3830 421 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3744 421 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3658 421 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3572 421 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16460 381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16460 381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16379 381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16379 381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16298 381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16298 381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16217 381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16217 381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16136 381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16136 381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 16055 381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16055 381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15974 381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15974 381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15893 381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15893 381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15812 381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15812 381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15731 381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15731 381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15650 381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15650 381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15569 381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15569 381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15488 381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15488 381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15407 381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15407 381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15326 381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15326 381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15245 381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15245 381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15164 381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15164 381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15083 381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15083 381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 15002 381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15002 381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14921 381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14921 381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14840 381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14840 381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14759 381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14759 381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14678 381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14678 381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14597 381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14597 381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14515 381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14515 381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14433 381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14433 381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14351 381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14351 381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14269 381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14269 381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14187 381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14187 381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14105 381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14105 381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 14023 381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14023 381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13941 381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13941 381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13859 381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13859 381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13777 381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13777 381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13695 381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13695 381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 317 13613 381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13613 381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18527 363 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18527 363 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18445 363 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18445 363 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18363 363 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18363 363 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18281 363 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18281 363 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18199 363 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18199 363 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18117 363 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18117 363 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 18035 363 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18035 363 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17953 363 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17953 363 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17871 363 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17871 363 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17789 363 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17789 363 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17707 363 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17707 363 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17625 363 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17625 363 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17543 363 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17543 363 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17461 363 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17461 363 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17379 363 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17379 363 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17297 363 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17297 363 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17215 363 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17215 363 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17133 363 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17133 363 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 17051 363 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17051 363 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16969 363 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16969 363 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16887 363 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16887 363 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16805 363 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16805 363 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16723 363 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16723 363 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16641 363 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16641 363 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 299 16559 363 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16559 363 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4432 340 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4346 340 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4260 340 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4174 340 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4088 340 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4002 340 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3916 340 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3830 340 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3744 340 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3658 340 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3572 340 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16460 301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16460 301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16379 301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16379 301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16298 301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16298 301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16217 301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16217 301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16136 301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16136 301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16055 301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16055 301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15974 301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15974 301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15893 301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15893 301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15812 301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15812 301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15731 301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15731 301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15650 301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15650 301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15569 301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15569 301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15488 301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15488 301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15407 301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15407 301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15326 301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15326 301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15245 301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15245 301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15164 301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15164 301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15083 301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15083 301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 15002 301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15002 301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14921 301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14921 301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14840 301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14840 301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14759 301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14759 301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14678 301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14678 301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14597 301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14597 301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14515 301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14515 301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14433 301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14433 301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14351 301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14351 301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14269 301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14269 301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14187 301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14187 301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14105 301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14105 301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 14023 301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14023 301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 13941 301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13941 301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 13859 301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13859 301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 13777 301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13777 301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 13695 301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13695 301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 13613 301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13613 301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 18527 281 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18527 281 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 18445 281 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18445 281 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 18363 281 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18363 281 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 18281 281 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18281 281 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 18199 281 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18199 281 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 18117 281 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18117 281 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 18035 281 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18035 281 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17953 281 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17953 281 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17871 281 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17871 281 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17789 281 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17789 281 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17707 281 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17707 281 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17625 281 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17625 281 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17543 281 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17543 281 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17461 281 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17461 281 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17379 281 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17379 281 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17297 281 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17297 281 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17215 281 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17215 281 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17133 281 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17133 281 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 17051 281 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17051 281 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16969 281 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16969 281 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16887 281 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16887 281 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16805 281 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16805 281 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16723 281 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16723 281 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16641 281 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16641 281 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 254 16559 281 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16559 281 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4432 259 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4346 259 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4260 259 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4174 259 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4088 259 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4002 259 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3916 259 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3830 259 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3744 259 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3658 259 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3572 259 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16460 221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16379 221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16298 221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16217 221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16136 221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16055 221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15974 221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15893 221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15812 221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15731 221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15650 221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15569 221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15488 221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15407 221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15326 221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15245 221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15164 221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15083 221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15002 221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14921 221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14840 221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14759 221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14678 221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14597 221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14515 221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14433 221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14351 221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14269 221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14187 221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14105 221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14023 221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13941 221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13859 221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13777 221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13695 221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13613 221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18527 199 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18445 199 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18363 199 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18281 199 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18199 199 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18117 199 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18035 199 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17953 199 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17871 199 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17789 199 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17707 199 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17625 199 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17543 199 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17461 199 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17379 199 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17297 199 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17215 199 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17133 199 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17051 199 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16969 199 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16887 199 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16805 199 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16723 199 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16641 199 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16559 199 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4432 178 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4346 178 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4260 178 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4174 178 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4088 178 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4002 178 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3916 178 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3830 178 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3744 178 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3658 178 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3572 178 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1884376
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 1300792
<< end >>
