magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 1 21 1217 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 97 163 177
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 165 247 177
rect 193 131 203 165
rect 237 131 247 165
rect 193 97 247 131
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 97 331 177
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 165 415 177
rect 361 131 371 165
rect 405 131 415 165
rect 361 47 415 131
rect 445 97 499 177
rect 445 63 455 97
rect 489 63 499 97
rect 445 47 499 63
rect 529 165 583 177
rect 529 131 539 165
rect 573 131 583 165
rect 529 47 583 131
rect 613 97 667 177
rect 613 63 623 97
rect 657 63 667 97
rect 613 47 667 63
rect 697 165 749 177
rect 697 131 707 165
rect 741 131 749 165
rect 697 47 749 131
rect 803 97 855 177
rect 803 63 811 97
rect 845 63 855 97
rect 803 47 855 63
rect 885 165 939 177
rect 885 131 895 165
rect 929 131 939 165
rect 885 47 939 131
rect 969 97 1023 177
rect 969 63 979 97
rect 1013 63 1023 97
rect 969 47 1023 63
rect 1053 165 1107 177
rect 1053 131 1063 165
rect 1097 131 1107 165
rect 1053 47 1107 131
rect 1137 97 1191 177
rect 1137 63 1147 97
rect 1181 63 1191 97
rect 1137 47 1191 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 349 331 383
rect 277 315 287 349
rect 321 315 331 349
rect 277 297 331 315
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 485 499 497
rect 445 451 455 485
rect 489 451 499 485
rect 445 417 499 451
rect 445 383 455 417
rect 489 383 499 417
rect 445 349 499 383
rect 445 315 455 349
rect 489 315 499 349
rect 445 297 499 315
rect 529 485 583 497
rect 529 451 539 485
rect 573 451 583 485
rect 529 417 583 451
rect 529 383 539 417
rect 573 383 583 417
rect 529 297 583 383
rect 613 485 667 497
rect 613 451 623 485
rect 657 451 667 485
rect 613 417 667 451
rect 613 383 623 417
rect 657 383 667 417
rect 613 349 667 383
rect 613 315 623 349
rect 657 315 667 349
rect 613 297 667 315
rect 697 485 749 497
rect 697 451 707 485
rect 741 451 749 485
rect 697 417 749 451
rect 697 383 707 417
rect 741 383 749 417
rect 697 297 749 383
rect 803 485 855 497
rect 803 451 811 485
rect 845 451 855 485
rect 803 417 855 451
rect 803 383 811 417
rect 845 383 855 417
rect 803 297 855 383
rect 885 485 939 497
rect 885 451 895 485
rect 929 451 939 485
rect 885 417 939 451
rect 885 383 895 417
rect 929 383 939 417
rect 885 349 939 383
rect 885 315 895 349
rect 929 315 939 349
rect 885 297 939 315
rect 969 485 1023 497
rect 969 451 979 485
rect 1013 451 1023 485
rect 969 417 1023 451
rect 969 383 979 417
rect 1013 383 1023 417
rect 969 297 1023 383
rect 1053 485 1107 497
rect 1053 451 1063 485
rect 1097 451 1107 485
rect 1053 417 1107 451
rect 1053 383 1063 417
rect 1097 383 1107 417
rect 1053 349 1107 383
rect 1053 315 1063 349
rect 1097 315 1107 349
rect 1053 297 1107 315
rect 1137 485 1191 497
rect 1137 451 1147 485
rect 1181 451 1191 485
rect 1137 417 1191 451
rect 1137 383 1147 417
rect 1181 383 1191 417
rect 1137 297 1191 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 63 153 97
rect 203 131 237 165
rect 203 63 237 97
rect 287 63 321 97
rect 371 131 405 165
rect 455 63 489 97
rect 539 131 573 165
rect 623 63 657 97
rect 707 131 741 165
rect 811 63 845 97
rect 895 131 929 165
rect 979 63 1013 97
rect 1063 131 1097 165
rect 1147 63 1181 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 287 451 321 485
rect 287 383 321 417
rect 287 315 321 349
rect 371 451 405 485
rect 371 383 405 417
rect 455 451 489 485
rect 455 383 489 417
rect 455 315 489 349
rect 539 451 573 485
rect 539 383 573 417
rect 623 451 657 485
rect 623 383 657 417
rect 623 315 657 349
rect 707 451 741 485
rect 707 383 741 417
rect 811 451 845 485
rect 811 383 845 417
rect 895 451 929 485
rect 895 383 929 417
rect 895 315 929 349
rect 979 451 1013 485
rect 979 383 1013 417
rect 1063 451 1097 485
rect 1063 383 1097 417
rect 1063 315 1097 349
rect 1147 451 1181 485
rect 1147 383 1181 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 79 261 109 297
rect 22 259 109 261
rect 163 259 193 297
rect 247 259 277 297
rect 331 259 361 297
rect 22 249 361 259
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 361 249
rect 22 205 361 215
rect 22 203 109 205
rect 79 177 109 203
rect 163 177 193 205
rect 247 177 277 205
rect 331 177 361 205
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 259 697 297
rect 855 259 885 297
rect 939 259 969 297
rect 1023 259 1053 297
rect 1107 259 1137 297
rect 415 249 697 259
rect 415 215 455 249
rect 489 215 539 249
rect 573 215 623 249
rect 657 215 697 249
rect 415 205 697 215
rect 789 249 1137 259
rect 789 215 805 249
rect 839 215 894 249
rect 928 215 979 249
rect 1013 215 1063 249
rect 1097 215 1137 249
rect 789 205 1137 215
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 667 177 697 205
rect 855 177 885 205
rect 939 177 969 205
rect 1023 177 1053 205
rect 1107 177 1137 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
<< polycont >>
rect 38 215 72 249
rect 119 215 153 249
rect 203 215 237 249
rect 287 215 321 249
rect 455 215 489 249
rect 539 215 573 249
rect 623 215 657 249
rect 805 215 839 249
rect 894 215 928 249
rect 979 215 1013 249
rect 1063 215 1097 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 289 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 271 485 337 493
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 103 315 119 349
rect 153 333 169 349
rect 271 349 337 383
rect 371 485 405 527
rect 371 417 405 451
rect 371 367 405 383
rect 439 485 505 493
rect 439 451 455 485
rect 489 451 505 485
rect 439 417 505 451
rect 439 383 455 417
rect 489 383 505 417
rect 271 333 287 349
rect 153 315 287 333
rect 321 333 337 349
rect 439 349 505 383
rect 539 485 573 527
rect 539 417 573 451
rect 539 367 573 383
rect 607 485 673 493
rect 607 451 623 485
rect 657 451 673 485
rect 607 417 673 451
rect 607 383 623 417
rect 657 383 673 417
rect 439 333 455 349
rect 321 315 455 333
rect 489 333 505 349
rect 607 349 673 383
rect 707 485 845 527
rect 741 451 811 485
rect 707 417 845 451
rect 741 383 811 417
rect 707 367 845 383
rect 879 485 945 493
rect 879 451 895 485
rect 929 451 945 485
rect 879 417 945 451
rect 879 383 895 417
rect 929 383 945 417
rect 607 333 623 349
rect 489 315 623 333
rect 657 333 673 349
rect 879 349 945 383
rect 979 485 1013 527
rect 979 417 1013 451
rect 979 367 1013 383
rect 1047 485 1113 493
rect 1047 451 1063 485
rect 1097 451 1113 485
rect 1047 417 1113 451
rect 1047 383 1063 417
rect 1097 383 1113 417
rect 879 333 895 349
rect 657 315 895 333
rect 929 333 945 349
rect 1047 349 1113 383
rect 1147 485 1200 527
rect 1181 451 1200 485
rect 1147 417 1200 451
rect 1181 383 1200 417
rect 1147 367 1200 383
rect 1047 333 1063 349
rect 929 315 1063 333
rect 1097 333 1113 349
rect 1097 315 1271 333
rect 103 289 1271 315
rect 22 249 340 255
rect 22 215 38 249
rect 72 215 119 249
rect 153 215 203 249
rect 237 215 287 249
rect 321 215 340 249
rect 398 249 708 255
rect 398 215 455 249
rect 489 215 539 249
rect 573 215 623 249
rect 657 215 708 249
rect 770 249 1113 255
rect 770 215 805 249
rect 839 215 894 249
rect 928 215 979 249
rect 1013 215 1063 249
rect 1097 215 1113 249
rect 1225 181 1271 289
rect 18 165 757 181
rect 18 131 35 165
rect 69 147 203 165
rect 69 131 85 147
rect 18 97 85 131
rect 187 131 203 147
rect 237 147 371 165
rect 237 131 253 147
rect 355 131 371 147
rect 405 147 539 165
rect 405 131 421 147
rect 523 131 539 147
rect 573 147 707 165
rect 573 131 589 147
rect 691 131 707 147
rect 741 131 757 165
rect 879 165 1271 181
rect 879 131 895 165
rect 929 131 1063 165
rect 1097 131 1271 165
rect 18 63 35 97
rect 69 63 85 97
rect 18 51 85 63
rect 119 97 153 113
rect 119 17 153 63
rect 187 97 253 131
rect 187 63 203 97
rect 237 63 253 97
rect 187 51 253 63
rect 287 97 321 113
rect 287 17 321 63
rect 439 63 455 97
rect 489 63 623 97
rect 657 63 811 97
rect 845 63 979 97
rect 1013 63 1147 97
rect 1181 63 1200 97
rect 439 51 1200 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel locali s 1225 153 1259 187 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 1225 289 1259 323 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 1046 221 1080 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand3_4
rlabel metal1 s 0 -48 1288 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 1852526
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1841390
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 32.200 0.000 
<< end >>
