/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/sky130_fd_pr__model__diode_pw2nd_11v0.model.spice