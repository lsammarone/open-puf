magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 475 936 813 998
rect -91 821 813 936
rect 2735 954 3201 1626
rect -91 189 953 821
rect 175 120 953 189
<< pwell >>
rect 1232 2195 2455 2228
rect 1232 2050 2563 2195
rect 639 1582 2563 2050
rect 639 1451 725 1582
rect 4 1116 464 1308
rect 1232 1275 2563 1582
rect 747 1083 2563 1275
rect 1225 880 2563 1083
rect 1053 798 2563 880
rect 1053 546 3126 798
rect 1053 102 2563 546
rect 1053 66 1187 102
rect 2477 82 2563 102
<< nmos >>
rect 2679 572 2729 772
rect 2785 572 2835 772
rect 2891 572 2941 772
rect 2997 572 3047 772
<< mvnmos >>
rect 829 1884 949 2024
rect 1005 1884 1125 2024
rect 829 1608 949 1748
rect 1005 1608 1125 1748
rect 86 1142 206 1282
rect 262 1142 382 1282
rect 826 1109 946 1249
rect 1002 1109 1122 1249
rect 1311 1202 1411 2202
rect 1620 1202 1720 2202
<< mvpmos >>
rect 28 670 128 870
rect 294 555 414 755
rect 594 732 694 932
rect 28 255 128 455
rect 594 459 694 659
rect 294 186 414 386
rect 594 186 694 386
<< mvnnmos >>
rect 1900 2002 2080 2202
rect 1900 1742 2080 1942
rect 1900 1482 2080 1682
rect 1900 1222 2080 1422
rect 1304 908 1484 1108
rect 1540 908 1720 1108
rect 1900 908 2080 1108
rect 1304 648 1484 848
rect 1540 648 1720 848
rect 1900 648 2080 848
rect 1304 388 1484 588
rect 1540 388 1720 588
rect 1900 388 2080 588
rect 1304 128 1484 328
rect 1540 128 1720 328
rect 1900 128 2080 328
<< pmoshvt >>
rect 2824 990 2874 1590
rect 2930 990 2980 1590
<< nmoslvt >>
rect 2260 2002 2290 2202
rect 2346 2002 2376 2202
rect 2260 1742 2290 1942
rect 2346 1742 2376 1942
rect 2260 1482 2290 1682
rect 2346 1482 2376 1682
rect 2260 1222 2290 1422
rect 2346 1222 2376 1422
rect 2260 908 2290 1108
rect 2346 908 2376 1108
rect 2260 648 2290 848
rect 2346 648 2376 848
rect 2260 388 2290 588
rect 2346 388 2376 588
rect 2260 128 2290 328
rect 2346 128 2376 328
<< ndiff >>
rect 2207 2184 2260 2202
rect 2207 2150 2215 2184
rect 2249 2150 2260 2184
rect 2207 2116 2260 2150
rect 2207 2082 2215 2116
rect 2249 2082 2260 2116
rect 2207 2048 2260 2082
rect 2207 2014 2215 2048
rect 2249 2014 2260 2048
rect 2207 2002 2260 2014
rect 2290 2184 2346 2202
rect 2290 2150 2301 2184
rect 2335 2150 2346 2184
rect 2290 2116 2346 2150
rect 2290 2082 2301 2116
rect 2335 2082 2346 2116
rect 2290 2048 2346 2082
rect 2290 2014 2301 2048
rect 2335 2014 2346 2048
rect 2290 2002 2346 2014
rect 2376 2184 2429 2202
rect 2376 2150 2387 2184
rect 2421 2150 2429 2184
rect 2376 2116 2429 2150
rect 2376 2082 2387 2116
rect 2421 2082 2429 2116
rect 2376 2048 2429 2082
rect 2376 2014 2387 2048
rect 2421 2014 2429 2048
rect 2376 2002 2429 2014
rect 2207 1924 2260 1942
rect 2207 1890 2215 1924
rect 2249 1890 2260 1924
rect 2207 1856 2260 1890
rect 2207 1822 2215 1856
rect 2249 1822 2260 1856
rect 2207 1788 2260 1822
rect 2207 1754 2215 1788
rect 2249 1754 2260 1788
rect 2207 1742 2260 1754
rect 2290 1924 2346 1942
rect 2290 1890 2301 1924
rect 2335 1890 2346 1924
rect 2290 1856 2346 1890
rect 2290 1822 2301 1856
rect 2335 1822 2346 1856
rect 2290 1788 2346 1822
rect 2290 1754 2301 1788
rect 2335 1754 2346 1788
rect 2290 1742 2346 1754
rect 2376 1924 2429 1942
rect 2376 1890 2387 1924
rect 2421 1890 2429 1924
rect 2376 1856 2429 1890
rect 2376 1822 2387 1856
rect 2421 1822 2429 1856
rect 2376 1788 2429 1822
rect 2376 1754 2387 1788
rect 2421 1754 2429 1788
rect 2376 1742 2429 1754
rect 2207 1664 2260 1682
rect 2207 1630 2215 1664
rect 2249 1630 2260 1664
rect 2207 1596 2260 1630
rect 2207 1562 2215 1596
rect 2249 1562 2260 1596
rect 2207 1528 2260 1562
rect 2207 1494 2215 1528
rect 2249 1494 2260 1528
rect 2207 1482 2260 1494
rect 2290 1664 2346 1682
rect 2290 1630 2301 1664
rect 2335 1630 2346 1664
rect 2290 1596 2346 1630
rect 2290 1562 2301 1596
rect 2335 1562 2346 1596
rect 2290 1528 2346 1562
rect 2290 1494 2301 1528
rect 2335 1494 2346 1528
rect 2290 1482 2346 1494
rect 2376 1664 2429 1682
rect 2376 1630 2387 1664
rect 2421 1630 2429 1664
rect 2376 1596 2429 1630
rect 2376 1562 2387 1596
rect 2421 1562 2429 1596
rect 2376 1528 2429 1562
rect 2376 1494 2387 1528
rect 2421 1494 2429 1528
rect 2376 1482 2429 1494
rect 2207 1404 2260 1422
rect 2207 1370 2215 1404
rect 2249 1370 2260 1404
rect 2207 1336 2260 1370
rect 2207 1302 2215 1336
rect 2249 1302 2260 1336
rect 2207 1268 2260 1302
rect 2207 1234 2215 1268
rect 2249 1234 2260 1268
rect 2207 1222 2260 1234
rect 2290 1404 2346 1422
rect 2290 1370 2301 1404
rect 2335 1370 2346 1404
rect 2290 1336 2346 1370
rect 2290 1302 2301 1336
rect 2335 1302 2346 1336
rect 2290 1268 2346 1302
rect 2290 1234 2301 1268
rect 2335 1234 2346 1268
rect 2290 1222 2346 1234
rect 2376 1404 2429 1422
rect 2376 1370 2387 1404
rect 2421 1370 2429 1404
rect 2376 1336 2429 1370
rect 2376 1302 2387 1336
rect 2421 1302 2429 1336
rect 2376 1268 2429 1302
rect 2376 1234 2387 1268
rect 2421 1234 2429 1268
rect 2376 1222 2429 1234
rect 2207 1090 2260 1108
rect 2207 1056 2215 1090
rect 2249 1056 2260 1090
rect 2207 1022 2260 1056
rect 2207 988 2215 1022
rect 2249 988 2260 1022
rect 2207 954 2260 988
rect 2207 920 2215 954
rect 2249 920 2260 954
rect 2207 908 2260 920
rect 2290 1090 2346 1108
rect 2290 1056 2301 1090
rect 2335 1056 2346 1090
rect 2290 1022 2346 1056
rect 2290 988 2301 1022
rect 2335 988 2346 1022
rect 2290 954 2346 988
rect 2290 920 2301 954
rect 2335 920 2346 954
rect 2290 908 2346 920
rect 2376 1090 2429 1108
rect 2376 1056 2387 1090
rect 2421 1056 2429 1090
rect 2376 1022 2429 1056
rect 2376 988 2387 1022
rect 2421 988 2429 1022
rect 2376 954 2429 988
rect 2376 920 2387 954
rect 2421 920 2429 954
rect 2376 908 2429 920
rect 2207 830 2260 848
rect 2207 796 2215 830
rect 2249 796 2260 830
rect 2207 762 2260 796
rect 2207 728 2215 762
rect 2249 728 2260 762
rect 2207 694 2260 728
rect 2207 660 2215 694
rect 2249 660 2260 694
rect 2207 648 2260 660
rect 2290 830 2346 848
rect 2290 796 2301 830
rect 2335 796 2346 830
rect 2290 762 2346 796
rect 2290 728 2301 762
rect 2335 728 2346 762
rect 2290 694 2346 728
rect 2290 660 2301 694
rect 2335 660 2346 694
rect 2290 648 2346 660
rect 2376 830 2429 848
rect 2376 796 2387 830
rect 2421 796 2429 830
rect 2376 762 2429 796
rect 2376 728 2387 762
rect 2421 728 2429 762
rect 2376 694 2429 728
rect 2376 660 2387 694
rect 2421 660 2429 694
rect 2376 648 2429 660
rect 2207 570 2260 588
rect 2207 536 2215 570
rect 2249 536 2260 570
rect 2207 502 2260 536
rect 2207 468 2215 502
rect 2249 468 2260 502
rect 2207 434 2260 468
rect 2207 400 2215 434
rect 2249 400 2260 434
rect 2207 388 2260 400
rect 2290 570 2346 588
rect 2290 536 2301 570
rect 2335 536 2346 570
rect 2290 502 2346 536
rect 2290 468 2301 502
rect 2335 468 2346 502
rect 2290 434 2346 468
rect 2290 400 2301 434
rect 2335 400 2346 434
rect 2290 388 2346 400
rect 2376 570 2429 588
rect 2376 536 2387 570
rect 2421 536 2429 570
rect 2376 502 2429 536
rect 2376 468 2387 502
rect 2421 468 2429 502
rect 2376 434 2429 468
rect 2376 400 2387 434
rect 2421 400 2429 434
rect 2376 388 2429 400
rect 2626 754 2679 772
rect 2626 720 2634 754
rect 2668 720 2679 754
rect 2626 686 2679 720
rect 2626 652 2634 686
rect 2668 652 2679 686
rect 2626 618 2679 652
rect 2626 584 2634 618
rect 2668 584 2679 618
rect 2626 572 2679 584
rect 2729 754 2785 772
rect 2729 720 2740 754
rect 2774 720 2785 754
rect 2729 686 2785 720
rect 2729 652 2740 686
rect 2774 652 2785 686
rect 2729 618 2785 652
rect 2729 584 2740 618
rect 2774 584 2785 618
rect 2729 572 2785 584
rect 2835 754 2891 772
rect 2835 720 2846 754
rect 2880 720 2891 754
rect 2835 686 2891 720
rect 2835 652 2846 686
rect 2880 652 2891 686
rect 2835 618 2891 652
rect 2835 584 2846 618
rect 2880 584 2891 618
rect 2835 572 2891 584
rect 2941 754 2997 772
rect 2941 720 2952 754
rect 2986 720 2997 754
rect 2941 686 2997 720
rect 2941 652 2952 686
rect 2986 652 2997 686
rect 2941 618 2997 652
rect 2941 584 2952 618
rect 2986 584 2997 618
rect 2941 572 2997 584
rect 3047 754 3100 772
rect 3047 720 3058 754
rect 3092 720 3100 754
rect 3047 686 3100 720
rect 3047 652 3058 686
rect 3092 652 3100 686
rect 3047 618 3100 652
rect 3047 584 3058 618
rect 3092 584 3100 618
rect 3047 572 3100 584
rect 2207 310 2260 328
rect 2207 276 2215 310
rect 2249 276 2260 310
rect 2207 242 2260 276
rect 2207 208 2215 242
rect 2249 208 2260 242
rect 2207 174 2260 208
rect 2207 140 2215 174
rect 2249 140 2260 174
rect 2207 128 2260 140
rect 2290 310 2346 328
rect 2290 276 2301 310
rect 2335 276 2346 310
rect 2290 242 2346 276
rect 2290 208 2301 242
rect 2335 208 2346 242
rect 2290 174 2346 208
rect 2290 140 2301 174
rect 2335 140 2346 174
rect 2290 128 2346 140
rect 2376 310 2429 328
rect 2376 276 2387 310
rect 2421 276 2429 310
rect 2376 242 2429 276
rect 2376 208 2387 242
rect 2421 208 2429 242
rect 2376 174 2429 208
rect 2376 140 2387 174
rect 2421 140 2429 174
rect 2376 128 2429 140
<< pdiff >>
rect 2771 1578 2824 1590
rect 2771 1544 2779 1578
rect 2813 1544 2824 1578
rect 2771 1510 2824 1544
rect 2771 1476 2779 1510
rect 2813 1476 2824 1510
rect 2771 1442 2824 1476
rect 2771 1408 2779 1442
rect 2813 1408 2824 1442
rect 2771 1374 2824 1408
rect 2771 1340 2779 1374
rect 2813 1340 2824 1374
rect 2771 1306 2824 1340
rect 2771 1272 2779 1306
rect 2813 1272 2824 1306
rect 2771 1238 2824 1272
rect 2771 1204 2779 1238
rect 2813 1204 2824 1238
rect 2771 1170 2824 1204
rect 2771 1136 2779 1170
rect 2813 1136 2824 1170
rect 2771 1102 2824 1136
rect 2771 1068 2779 1102
rect 2813 1068 2824 1102
rect 2771 990 2824 1068
rect 2874 1578 2930 1590
rect 2874 1544 2885 1578
rect 2919 1544 2930 1578
rect 2874 1510 2930 1544
rect 2874 1476 2885 1510
rect 2919 1476 2930 1510
rect 2874 1442 2930 1476
rect 2874 1408 2885 1442
rect 2919 1408 2930 1442
rect 2874 1374 2930 1408
rect 2874 1340 2885 1374
rect 2919 1340 2930 1374
rect 2874 1306 2930 1340
rect 2874 1272 2885 1306
rect 2919 1272 2930 1306
rect 2874 1238 2930 1272
rect 2874 1204 2885 1238
rect 2919 1204 2930 1238
rect 2874 1170 2930 1204
rect 2874 1136 2885 1170
rect 2919 1136 2930 1170
rect 2874 1102 2930 1136
rect 2874 1068 2885 1102
rect 2919 1068 2930 1102
rect 2874 990 2930 1068
rect 2980 1578 3033 1590
rect 2980 1544 2991 1578
rect 3025 1544 3033 1578
rect 2980 1510 3033 1544
rect 2980 1476 2991 1510
rect 3025 1476 3033 1510
rect 2980 1442 3033 1476
rect 2980 1408 2991 1442
rect 3025 1408 3033 1442
rect 2980 1374 3033 1408
rect 2980 1340 2991 1374
rect 3025 1340 3033 1374
rect 2980 1306 3033 1340
rect 2980 1272 2991 1306
rect 3025 1272 3033 1306
rect 2980 1238 3033 1272
rect 2980 1204 2991 1238
rect 3025 1204 3033 1238
rect 2980 1170 3033 1204
rect 2980 1136 2991 1170
rect 3025 1136 3033 1170
rect 2980 1102 3033 1136
rect 2980 1068 2991 1102
rect 3025 1068 3033 1102
rect 2980 990 3033 1068
<< mvndiff >>
rect 1258 2190 1311 2202
rect 1258 2156 1266 2190
rect 1300 2156 1311 2190
rect 1258 2122 1311 2156
rect 1258 2088 1266 2122
rect 1300 2088 1311 2122
rect 1258 2054 1311 2088
rect 773 1998 829 2024
rect 773 1964 784 1998
rect 818 1964 829 1998
rect 773 1930 829 1964
rect 773 1896 784 1930
rect 818 1896 829 1930
rect 773 1884 829 1896
rect 949 1998 1005 2024
rect 949 1964 960 1998
rect 994 1964 1005 1998
rect 949 1930 1005 1964
rect 949 1896 960 1930
rect 994 1896 1005 1930
rect 949 1884 1005 1896
rect 1125 1998 1181 2024
rect 1125 1964 1136 1998
rect 1170 1964 1181 1998
rect 1125 1930 1181 1964
rect 1125 1896 1136 1930
rect 1170 1896 1181 1930
rect 1125 1884 1181 1896
rect 1258 2020 1266 2054
rect 1300 2020 1311 2054
rect 1258 1986 1311 2020
rect 1258 1952 1266 1986
rect 1300 1952 1311 1986
rect 1258 1918 1311 1952
rect 1258 1884 1266 1918
rect 1300 1884 1311 1918
rect 1258 1850 1311 1884
rect 1258 1816 1266 1850
rect 1300 1816 1311 1850
rect 1258 1782 1311 1816
rect 1258 1748 1266 1782
rect 1300 1748 1311 1782
rect 773 1722 829 1748
rect 773 1688 784 1722
rect 818 1688 829 1722
rect 773 1654 829 1688
rect 773 1620 784 1654
rect 818 1620 829 1654
rect 773 1608 829 1620
rect 949 1722 1005 1748
rect 949 1688 960 1722
rect 994 1688 1005 1722
rect 949 1654 1005 1688
rect 949 1620 960 1654
rect 994 1620 1005 1654
rect 949 1608 1005 1620
rect 1125 1722 1181 1748
rect 1125 1688 1136 1722
rect 1170 1688 1181 1722
rect 1125 1654 1181 1688
rect 1125 1620 1136 1654
rect 1170 1620 1181 1654
rect 1125 1608 1181 1620
rect 1258 1714 1311 1748
rect 1258 1680 1266 1714
rect 1300 1680 1311 1714
rect 1258 1646 1311 1680
rect 1258 1612 1266 1646
rect 1300 1612 1311 1646
rect 1258 1578 1311 1612
rect 1258 1544 1266 1578
rect 1300 1544 1311 1578
rect 1258 1510 1311 1544
rect 1258 1476 1266 1510
rect 1300 1476 1311 1510
rect 1258 1442 1311 1476
rect 1258 1408 1266 1442
rect 1300 1408 1311 1442
rect 1258 1374 1311 1408
rect 1258 1340 1266 1374
rect 1300 1340 1311 1374
rect 1258 1306 1311 1340
rect 30 1270 86 1282
rect 30 1236 41 1270
rect 75 1236 86 1270
rect 30 1202 86 1236
rect 30 1168 41 1202
rect 75 1168 86 1202
rect 30 1142 86 1168
rect 206 1270 262 1282
rect 206 1236 217 1270
rect 251 1236 262 1270
rect 206 1202 262 1236
rect 206 1168 217 1202
rect 251 1168 262 1202
rect 206 1142 262 1168
rect 382 1270 438 1282
rect 382 1236 393 1270
rect 427 1236 438 1270
rect 1258 1272 1266 1306
rect 1300 1272 1311 1306
rect 382 1202 438 1236
rect 382 1168 393 1202
rect 427 1168 438 1202
rect 382 1142 438 1168
rect 773 1237 826 1249
rect 773 1203 781 1237
rect 815 1203 826 1237
rect 773 1169 826 1203
rect 773 1135 781 1169
rect 815 1135 826 1169
rect 773 1109 826 1135
rect 946 1237 1002 1249
rect 946 1203 957 1237
rect 991 1203 1002 1237
rect 946 1169 1002 1203
rect 946 1135 957 1169
rect 991 1135 1002 1169
rect 946 1109 1002 1135
rect 1122 1237 1175 1249
rect 1122 1203 1133 1237
rect 1167 1203 1175 1237
rect 1122 1169 1175 1203
rect 1258 1202 1311 1272
rect 1411 2190 1467 2202
rect 1411 2156 1422 2190
rect 1456 2156 1467 2190
rect 1411 2122 1467 2156
rect 1411 2088 1422 2122
rect 1456 2088 1467 2122
rect 1411 2054 1467 2088
rect 1411 2020 1422 2054
rect 1456 2020 1467 2054
rect 1411 1986 1467 2020
rect 1411 1952 1422 1986
rect 1456 1952 1467 1986
rect 1411 1918 1467 1952
rect 1411 1884 1422 1918
rect 1456 1884 1467 1918
rect 1411 1850 1467 1884
rect 1411 1816 1422 1850
rect 1456 1816 1467 1850
rect 1411 1782 1467 1816
rect 1411 1748 1422 1782
rect 1456 1748 1467 1782
rect 1411 1714 1467 1748
rect 1411 1680 1422 1714
rect 1456 1680 1467 1714
rect 1411 1646 1467 1680
rect 1411 1612 1422 1646
rect 1456 1612 1467 1646
rect 1411 1578 1467 1612
rect 1411 1544 1422 1578
rect 1456 1544 1467 1578
rect 1411 1510 1467 1544
rect 1411 1476 1422 1510
rect 1456 1476 1467 1510
rect 1411 1442 1467 1476
rect 1411 1408 1422 1442
rect 1456 1408 1467 1442
rect 1411 1374 1467 1408
rect 1411 1340 1422 1374
rect 1456 1340 1467 1374
rect 1411 1306 1467 1340
rect 1411 1272 1422 1306
rect 1456 1272 1467 1306
rect 1411 1202 1467 1272
rect 1567 2190 1620 2202
rect 1567 2156 1575 2190
rect 1609 2156 1620 2190
rect 1567 2122 1620 2156
rect 1567 2088 1575 2122
rect 1609 2088 1620 2122
rect 1567 2054 1620 2088
rect 1567 2020 1575 2054
rect 1609 2020 1620 2054
rect 1567 1986 1620 2020
rect 1567 1952 1575 1986
rect 1609 1952 1620 1986
rect 1567 1918 1620 1952
rect 1567 1884 1575 1918
rect 1609 1884 1620 1918
rect 1567 1850 1620 1884
rect 1567 1816 1575 1850
rect 1609 1816 1620 1850
rect 1567 1782 1620 1816
rect 1567 1748 1575 1782
rect 1609 1748 1620 1782
rect 1567 1714 1620 1748
rect 1567 1680 1575 1714
rect 1609 1680 1620 1714
rect 1567 1646 1620 1680
rect 1567 1612 1575 1646
rect 1609 1612 1620 1646
rect 1567 1578 1620 1612
rect 1567 1544 1575 1578
rect 1609 1544 1620 1578
rect 1567 1510 1620 1544
rect 1567 1476 1575 1510
rect 1609 1476 1620 1510
rect 1567 1442 1620 1476
rect 1567 1408 1575 1442
rect 1609 1408 1620 1442
rect 1567 1374 1620 1408
rect 1567 1340 1575 1374
rect 1609 1340 1620 1374
rect 1567 1306 1620 1340
rect 1567 1272 1575 1306
rect 1609 1272 1620 1306
rect 1567 1202 1620 1272
rect 1720 2190 1773 2202
rect 1720 2156 1731 2190
rect 1765 2156 1773 2190
rect 1720 2122 1773 2156
rect 1720 2088 1731 2122
rect 1765 2088 1773 2122
rect 1720 2054 1773 2088
rect 1720 2020 1731 2054
rect 1765 2020 1773 2054
rect 1720 1986 1773 2020
rect 1847 2184 1900 2202
rect 1847 2150 1855 2184
rect 1889 2150 1900 2184
rect 1847 2116 1900 2150
rect 1847 2082 1855 2116
rect 1889 2082 1900 2116
rect 1847 2048 1900 2082
rect 1847 2014 1855 2048
rect 1889 2014 1900 2048
rect 1847 2002 1900 2014
rect 2080 2184 2133 2202
rect 2080 2150 2091 2184
rect 2125 2150 2133 2184
rect 2080 2116 2133 2150
rect 2080 2082 2091 2116
rect 2125 2082 2133 2116
rect 2080 2048 2133 2082
rect 2080 2014 2091 2048
rect 2125 2014 2133 2048
rect 2080 2002 2133 2014
rect 1720 1952 1731 1986
rect 1765 1952 1773 1986
rect 1720 1918 1773 1952
rect 1720 1884 1731 1918
rect 1765 1884 1773 1918
rect 1720 1850 1773 1884
rect 1720 1816 1731 1850
rect 1765 1816 1773 1850
rect 1720 1782 1773 1816
rect 1720 1748 1731 1782
rect 1765 1748 1773 1782
rect 1720 1714 1773 1748
rect 1847 1924 1900 1942
rect 1847 1890 1855 1924
rect 1889 1890 1900 1924
rect 1847 1856 1900 1890
rect 1847 1822 1855 1856
rect 1889 1822 1900 1856
rect 1847 1788 1900 1822
rect 1847 1754 1855 1788
rect 1889 1754 1900 1788
rect 1847 1742 1900 1754
rect 2080 1924 2133 1942
rect 2080 1890 2091 1924
rect 2125 1890 2133 1924
rect 2080 1856 2133 1890
rect 2080 1822 2091 1856
rect 2125 1822 2133 1856
rect 2080 1788 2133 1822
rect 2080 1754 2091 1788
rect 2125 1754 2133 1788
rect 2080 1742 2133 1754
rect 1720 1680 1731 1714
rect 1765 1680 1773 1714
rect 1720 1646 1773 1680
rect 1720 1612 1731 1646
rect 1765 1612 1773 1646
rect 1720 1578 1773 1612
rect 1720 1544 1731 1578
rect 1765 1544 1773 1578
rect 1720 1510 1773 1544
rect 1720 1476 1731 1510
rect 1765 1476 1773 1510
rect 1847 1664 1900 1682
rect 1847 1630 1855 1664
rect 1889 1630 1900 1664
rect 1847 1596 1900 1630
rect 1847 1562 1855 1596
rect 1889 1562 1900 1596
rect 1847 1528 1900 1562
rect 1847 1494 1855 1528
rect 1889 1494 1900 1528
rect 1847 1482 1900 1494
rect 2080 1664 2133 1682
rect 2080 1630 2091 1664
rect 2125 1630 2133 1664
rect 2080 1596 2133 1630
rect 2080 1562 2091 1596
rect 2125 1562 2133 1596
rect 2080 1528 2133 1562
rect 2080 1494 2091 1528
rect 2125 1494 2133 1528
rect 2080 1482 2133 1494
rect 1720 1442 1773 1476
rect 1720 1408 1731 1442
rect 1765 1408 1773 1442
rect 1720 1374 1773 1408
rect 1720 1340 1731 1374
rect 1765 1340 1773 1374
rect 1720 1306 1773 1340
rect 1720 1272 1731 1306
rect 1765 1272 1773 1306
rect 1720 1202 1773 1272
rect 1847 1404 1900 1422
rect 1847 1370 1855 1404
rect 1889 1370 1900 1404
rect 1847 1336 1900 1370
rect 1847 1302 1855 1336
rect 1889 1302 1900 1336
rect 1847 1268 1900 1302
rect 1847 1234 1855 1268
rect 1889 1234 1900 1268
rect 1847 1222 1900 1234
rect 2080 1404 2133 1422
rect 2080 1370 2091 1404
rect 2125 1370 2133 1404
rect 2080 1336 2133 1370
rect 2080 1302 2091 1336
rect 2125 1302 2133 1336
rect 2080 1268 2133 1302
rect 2080 1234 2091 1268
rect 2125 1234 2133 1268
rect 2080 1222 2133 1234
rect 1122 1135 1133 1169
rect 1167 1135 1175 1169
rect 1122 1109 1175 1135
rect 1251 1090 1304 1108
rect 1251 1056 1259 1090
rect 1293 1056 1304 1090
rect 1251 1022 1304 1056
rect 1251 988 1259 1022
rect 1293 988 1304 1022
rect 1251 954 1304 988
rect 1251 920 1259 954
rect 1293 920 1304 954
rect 1251 908 1304 920
rect 1484 1090 1540 1108
rect 1484 1056 1495 1090
rect 1529 1056 1540 1090
rect 1484 1022 1540 1056
rect 1484 988 1495 1022
rect 1529 988 1540 1022
rect 1484 954 1540 988
rect 1484 920 1495 954
rect 1529 920 1540 954
rect 1484 908 1540 920
rect 1720 1090 1773 1108
rect 1720 1056 1731 1090
rect 1765 1056 1773 1090
rect 1720 1022 1773 1056
rect 1720 988 1731 1022
rect 1765 988 1773 1022
rect 1720 954 1773 988
rect 1720 920 1731 954
rect 1765 920 1773 954
rect 1720 908 1773 920
rect 1847 1090 1900 1108
rect 1847 1056 1855 1090
rect 1889 1056 1900 1090
rect 1847 1022 1900 1056
rect 1847 988 1855 1022
rect 1889 988 1900 1022
rect 1847 954 1900 988
rect 1847 920 1855 954
rect 1889 920 1900 954
rect 1847 908 1900 920
rect 2080 1090 2133 1108
rect 2080 1056 2091 1090
rect 2125 1056 2133 1090
rect 2080 1022 2133 1056
rect 2080 988 2091 1022
rect 2125 988 2133 1022
rect 2080 954 2133 988
rect 2080 920 2091 954
rect 2125 920 2133 954
rect 2080 908 2133 920
rect 1251 830 1304 848
rect 1251 796 1259 830
rect 1293 796 1304 830
rect 1251 762 1304 796
rect 1251 728 1259 762
rect 1293 728 1304 762
rect 1251 694 1304 728
rect 1251 660 1259 694
rect 1293 660 1304 694
rect 1251 648 1304 660
rect 1484 830 1540 848
rect 1484 796 1495 830
rect 1529 796 1540 830
rect 1484 762 1540 796
rect 1484 728 1495 762
rect 1529 728 1540 762
rect 1484 694 1540 728
rect 1484 660 1495 694
rect 1529 660 1540 694
rect 1484 648 1540 660
rect 1720 830 1773 848
rect 1720 796 1731 830
rect 1765 796 1773 830
rect 1720 762 1773 796
rect 1720 728 1731 762
rect 1765 728 1773 762
rect 1720 694 1773 728
rect 1720 660 1731 694
rect 1765 660 1773 694
rect 1720 648 1773 660
rect 1847 830 1900 848
rect 1847 796 1855 830
rect 1889 796 1900 830
rect 1847 762 1900 796
rect 1847 728 1855 762
rect 1889 728 1900 762
rect 1847 694 1900 728
rect 1847 660 1855 694
rect 1889 660 1900 694
rect 1847 648 1900 660
rect 2080 830 2133 848
rect 2080 796 2091 830
rect 2125 796 2133 830
rect 2080 762 2133 796
rect 2080 728 2091 762
rect 2125 728 2133 762
rect 2080 694 2133 728
rect 2080 660 2091 694
rect 2125 660 2133 694
rect 2080 648 2133 660
rect 1251 570 1304 588
rect 1251 536 1259 570
rect 1293 536 1304 570
rect 1251 502 1304 536
rect 1251 468 1259 502
rect 1293 468 1304 502
rect 1251 434 1304 468
rect 1251 400 1259 434
rect 1293 400 1304 434
rect 1251 388 1304 400
rect 1484 570 1540 588
rect 1484 536 1495 570
rect 1529 536 1540 570
rect 1484 502 1540 536
rect 1484 468 1495 502
rect 1529 468 1540 502
rect 1484 434 1540 468
rect 1484 400 1495 434
rect 1529 400 1540 434
rect 1484 388 1540 400
rect 1720 570 1773 588
rect 1720 536 1731 570
rect 1765 536 1773 570
rect 1720 502 1773 536
rect 1720 468 1731 502
rect 1765 468 1773 502
rect 1720 434 1773 468
rect 1720 400 1731 434
rect 1765 400 1773 434
rect 1720 388 1773 400
rect 1847 570 1900 588
rect 1847 536 1855 570
rect 1889 536 1900 570
rect 1847 502 1900 536
rect 1847 468 1855 502
rect 1889 468 1900 502
rect 1847 434 1900 468
rect 1847 400 1855 434
rect 1889 400 1900 434
rect 1847 388 1900 400
rect 2080 570 2133 588
rect 2080 536 2091 570
rect 2125 536 2133 570
rect 2080 502 2133 536
rect 2080 468 2091 502
rect 2125 468 2133 502
rect 2080 434 2133 468
rect 2080 400 2091 434
rect 2125 400 2133 434
rect 2080 388 2133 400
rect 1251 310 1304 328
rect 1251 276 1259 310
rect 1293 276 1304 310
rect 1251 242 1304 276
rect 1251 208 1259 242
rect 1293 208 1304 242
rect 1251 174 1304 208
rect 1251 140 1259 174
rect 1293 140 1304 174
rect 1251 128 1304 140
rect 1484 310 1540 328
rect 1484 276 1495 310
rect 1529 276 1540 310
rect 1484 242 1540 276
rect 1484 208 1495 242
rect 1529 208 1540 242
rect 1484 174 1540 208
rect 1484 140 1495 174
rect 1529 140 1540 174
rect 1484 128 1540 140
rect 1720 310 1773 328
rect 1720 276 1731 310
rect 1765 276 1773 310
rect 1720 242 1773 276
rect 1720 208 1731 242
rect 1765 208 1773 242
rect 1720 174 1773 208
rect 1720 140 1731 174
rect 1765 140 1773 174
rect 1720 128 1773 140
rect 1847 310 1900 328
rect 1847 276 1855 310
rect 1889 276 1900 310
rect 1847 242 1900 276
rect 1847 208 1855 242
rect 1889 208 1900 242
rect 1847 174 1900 208
rect 1847 140 1855 174
rect 1889 140 1900 174
rect 1847 128 1900 140
rect 2080 310 2133 328
rect 2080 276 2091 310
rect 2125 276 2133 310
rect 2080 242 2133 276
rect 2080 208 2091 242
rect 2125 208 2133 242
rect 2080 174 2133 208
rect 2080 140 2091 174
rect 2125 140 2133 174
rect 2080 128 2133 140
<< mvpdiff >>
rect -25 858 28 870
rect -25 824 -17 858
rect 17 824 28 858
rect -25 790 28 824
rect -25 756 -17 790
rect 17 756 28 790
rect -25 722 28 756
rect -25 688 -17 722
rect 17 688 28 722
rect -25 670 28 688
rect 128 858 181 870
rect 128 824 139 858
rect 173 824 181 858
rect 128 790 181 824
rect 128 756 139 790
rect 173 756 181 790
rect 128 722 181 756
rect 541 914 594 932
rect 541 880 549 914
rect 583 880 594 914
rect 541 846 594 880
rect 541 812 549 846
rect 583 812 594 846
rect 541 778 594 812
rect 128 688 139 722
rect 173 688 181 722
rect 128 670 181 688
rect 241 743 294 755
rect 241 709 249 743
rect 283 709 294 743
rect 241 675 294 709
rect 241 641 249 675
rect 283 641 294 675
rect 241 607 294 641
rect 241 573 249 607
rect 283 573 294 607
rect 241 555 294 573
rect 414 743 467 755
rect 414 709 425 743
rect 459 709 467 743
rect 541 744 549 778
rect 583 744 594 778
rect 541 732 594 744
rect 694 914 747 932
rect 694 880 705 914
rect 739 880 747 914
rect 694 846 747 880
rect 694 812 705 846
rect 739 812 747 846
rect 694 778 747 812
rect 694 744 705 778
rect 739 744 747 778
rect 694 732 747 744
rect 414 675 467 709
rect 414 641 425 675
rect 459 641 467 675
rect 414 607 467 641
rect 414 573 425 607
rect 459 573 467 607
rect 414 555 467 573
rect 541 641 594 659
rect 541 607 549 641
rect 583 607 594 641
rect 541 573 594 607
rect 541 539 549 573
rect 583 539 594 573
rect 541 505 594 539
rect -25 443 28 455
rect -25 409 -17 443
rect 17 409 28 443
rect -25 375 28 409
rect -25 341 -17 375
rect 17 341 28 375
rect -25 307 28 341
rect -25 273 -17 307
rect 17 273 28 307
rect -25 255 28 273
rect 128 443 181 455
rect 128 409 139 443
rect 173 409 181 443
rect 128 375 181 409
rect 541 471 549 505
rect 583 471 594 505
rect 541 459 594 471
rect 694 641 747 659
rect 694 607 705 641
rect 739 607 747 641
rect 694 573 747 607
rect 694 539 705 573
rect 739 539 747 573
rect 694 505 747 539
rect 694 471 705 505
rect 739 471 747 505
rect 694 459 747 471
rect 128 341 139 375
rect 173 341 181 375
rect 128 307 181 341
rect 128 273 139 307
rect 173 273 181 307
rect 128 255 181 273
rect 241 374 294 386
rect 241 340 249 374
rect 283 340 294 374
rect 241 306 294 340
rect 241 272 249 306
rect 283 272 294 306
rect 241 238 294 272
rect 241 204 249 238
rect 283 204 294 238
rect 241 186 294 204
rect 414 374 467 386
rect 414 340 425 374
rect 459 340 467 374
rect 414 306 467 340
rect 414 272 425 306
rect 459 272 467 306
rect 414 238 467 272
rect 414 204 425 238
rect 459 204 467 238
rect 414 186 467 204
rect 541 368 594 386
rect 541 334 549 368
rect 583 334 594 368
rect 541 300 594 334
rect 541 266 549 300
rect 583 266 594 300
rect 541 232 594 266
rect 541 198 549 232
rect 583 198 594 232
rect 541 186 594 198
rect 694 368 747 386
rect 694 334 705 368
rect 739 334 747 368
rect 694 300 747 334
rect 694 266 705 300
rect 739 266 747 300
rect 694 232 747 266
rect 694 198 705 232
rect 739 198 747 232
rect 694 186 747 198
<< ndiffc >>
rect 2215 2150 2249 2184
rect 2215 2082 2249 2116
rect 2215 2014 2249 2048
rect 2301 2150 2335 2184
rect 2301 2082 2335 2116
rect 2301 2014 2335 2048
rect 2387 2150 2421 2184
rect 2387 2082 2421 2116
rect 2387 2014 2421 2048
rect 2215 1890 2249 1924
rect 2215 1822 2249 1856
rect 2215 1754 2249 1788
rect 2301 1890 2335 1924
rect 2301 1822 2335 1856
rect 2301 1754 2335 1788
rect 2387 1890 2421 1924
rect 2387 1822 2421 1856
rect 2387 1754 2421 1788
rect 2215 1630 2249 1664
rect 2215 1562 2249 1596
rect 2215 1494 2249 1528
rect 2301 1630 2335 1664
rect 2301 1562 2335 1596
rect 2301 1494 2335 1528
rect 2387 1630 2421 1664
rect 2387 1562 2421 1596
rect 2387 1494 2421 1528
rect 2215 1370 2249 1404
rect 2215 1302 2249 1336
rect 2215 1234 2249 1268
rect 2301 1370 2335 1404
rect 2301 1302 2335 1336
rect 2301 1234 2335 1268
rect 2387 1370 2421 1404
rect 2387 1302 2421 1336
rect 2387 1234 2421 1268
rect 2215 1056 2249 1090
rect 2215 988 2249 1022
rect 2215 920 2249 954
rect 2301 1056 2335 1090
rect 2301 988 2335 1022
rect 2301 920 2335 954
rect 2387 1056 2421 1090
rect 2387 988 2421 1022
rect 2387 920 2421 954
rect 2215 796 2249 830
rect 2215 728 2249 762
rect 2215 660 2249 694
rect 2301 796 2335 830
rect 2301 728 2335 762
rect 2301 660 2335 694
rect 2387 796 2421 830
rect 2387 728 2421 762
rect 2387 660 2421 694
rect 2215 536 2249 570
rect 2215 468 2249 502
rect 2215 400 2249 434
rect 2301 536 2335 570
rect 2301 468 2335 502
rect 2301 400 2335 434
rect 2387 536 2421 570
rect 2387 468 2421 502
rect 2387 400 2421 434
rect 2634 720 2668 754
rect 2634 652 2668 686
rect 2634 584 2668 618
rect 2740 720 2774 754
rect 2740 652 2774 686
rect 2740 584 2774 618
rect 2846 720 2880 754
rect 2846 652 2880 686
rect 2846 584 2880 618
rect 2952 720 2986 754
rect 2952 652 2986 686
rect 2952 584 2986 618
rect 3058 720 3092 754
rect 3058 652 3092 686
rect 3058 584 3092 618
rect 2215 276 2249 310
rect 2215 208 2249 242
rect 2215 140 2249 174
rect 2301 276 2335 310
rect 2301 208 2335 242
rect 2301 140 2335 174
rect 2387 276 2421 310
rect 2387 208 2421 242
rect 2387 140 2421 174
<< pdiffc >>
rect 2779 1544 2813 1578
rect 2779 1476 2813 1510
rect 2779 1408 2813 1442
rect 2779 1340 2813 1374
rect 2779 1272 2813 1306
rect 2779 1204 2813 1238
rect 2779 1136 2813 1170
rect 2779 1068 2813 1102
rect 2885 1544 2919 1578
rect 2885 1476 2919 1510
rect 2885 1408 2919 1442
rect 2885 1340 2919 1374
rect 2885 1272 2919 1306
rect 2885 1204 2919 1238
rect 2885 1136 2919 1170
rect 2885 1068 2919 1102
rect 2991 1544 3025 1578
rect 2991 1476 3025 1510
rect 2991 1408 3025 1442
rect 2991 1340 3025 1374
rect 2991 1272 3025 1306
rect 2991 1204 3025 1238
rect 2991 1136 3025 1170
rect 2991 1068 3025 1102
<< mvndiffc >>
rect 1266 2156 1300 2190
rect 1266 2088 1300 2122
rect 784 1964 818 1998
rect 784 1896 818 1930
rect 960 1964 994 1998
rect 960 1896 994 1930
rect 1136 1964 1170 1998
rect 1136 1896 1170 1930
rect 1266 2020 1300 2054
rect 1266 1952 1300 1986
rect 1266 1884 1300 1918
rect 1266 1816 1300 1850
rect 1266 1748 1300 1782
rect 784 1688 818 1722
rect 784 1620 818 1654
rect 960 1688 994 1722
rect 960 1620 994 1654
rect 1136 1688 1170 1722
rect 1136 1620 1170 1654
rect 1266 1680 1300 1714
rect 1266 1612 1300 1646
rect 1266 1544 1300 1578
rect 1266 1476 1300 1510
rect 1266 1408 1300 1442
rect 1266 1340 1300 1374
rect 41 1236 75 1270
rect 41 1168 75 1202
rect 217 1236 251 1270
rect 217 1168 251 1202
rect 393 1236 427 1270
rect 1266 1272 1300 1306
rect 393 1168 427 1202
rect 781 1203 815 1237
rect 781 1135 815 1169
rect 957 1203 991 1237
rect 957 1135 991 1169
rect 1133 1203 1167 1237
rect 1422 2156 1456 2190
rect 1422 2088 1456 2122
rect 1422 2020 1456 2054
rect 1422 1952 1456 1986
rect 1422 1884 1456 1918
rect 1422 1816 1456 1850
rect 1422 1748 1456 1782
rect 1422 1680 1456 1714
rect 1422 1612 1456 1646
rect 1422 1544 1456 1578
rect 1422 1476 1456 1510
rect 1422 1408 1456 1442
rect 1422 1340 1456 1374
rect 1422 1272 1456 1306
rect 1575 2156 1609 2190
rect 1575 2088 1609 2122
rect 1575 2020 1609 2054
rect 1575 1952 1609 1986
rect 1575 1884 1609 1918
rect 1575 1816 1609 1850
rect 1575 1748 1609 1782
rect 1575 1680 1609 1714
rect 1575 1612 1609 1646
rect 1575 1544 1609 1578
rect 1575 1476 1609 1510
rect 1575 1408 1609 1442
rect 1575 1340 1609 1374
rect 1575 1272 1609 1306
rect 1731 2156 1765 2190
rect 1731 2088 1765 2122
rect 1731 2020 1765 2054
rect 1855 2150 1889 2184
rect 1855 2082 1889 2116
rect 1855 2014 1889 2048
rect 2091 2150 2125 2184
rect 2091 2082 2125 2116
rect 2091 2014 2125 2048
rect 1731 1952 1765 1986
rect 1731 1884 1765 1918
rect 1731 1816 1765 1850
rect 1731 1748 1765 1782
rect 1855 1890 1889 1924
rect 1855 1822 1889 1856
rect 1855 1754 1889 1788
rect 2091 1890 2125 1924
rect 2091 1822 2125 1856
rect 2091 1754 2125 1788
rect 1731 1680 1765 1714
rect 1731 1612 1765 1646
rect 1731 1544 1765 1578
rect 1731 1476 1765 1510
rect 1855 1630 1889 1664
rect 1855 1562 1889 1596
rect 1855 1494 1889 1528
rect 2091 1630 2125 1664
rect 2091 1562 2125 1596
rect 2091 1494 2125 1528
rect 1731 1408 1765 1442
rect 1731 1340 1765 1374
rect 1731 1272 1765 1306
rect 1855 1370 1889 1404
rect 1855 1302 1889 1336
rect 1855 1234 1889 1268
rect 2091 1370 2125 1404
rect 2091 1302 2125 1336
rect 2091 1234 2125 1268
rect 1133 1135 1167 1169
rect 1259 1056 1293 1090
rect 1259 988 1293 1022
rect 1259 920 1293 954
rect 1495 1056 1529 1090
rect 1495 988 1529 1022
rect 1495 920 1529 954
rect 1731 1056 1765 1090
rect 1731 988 1765 1022
rect 1731 920 1765 954
rect 1855 1056 1889 1090
rect 1855 988 1889 1022
rect 1855 920 1889 954
rect 2091 1056 2125 1090
rect 2091 988 2125 1022
rect 2091 920 2125 954
rect 1259 796 1293 830
rect 1259 728 1293 762
rect 1259 660 1293 694
rect 1495 796 1529 830
rect 1495 728 1529 762
rect 1495 660 1529 694
rect 1731 796 1765 830
rect 1731 728 1765 762
rect 1731 660 1765 694
rect 1855 796 1889 830
rect 1855 728 1889 762
rect 1855 660 1889 694
rect 2091 796 2125 830
rect 2091 728 2125 762
rect 2091 660 2125 694
rect 1259 536 1293 570
rect 1259 468 1293 502
rect 1259 400 1293 434
rect 1495 536 1529 570
rect 1495 468 1529 502
rect 1495 400 1529 434
rect 1731 536 1765 570
rect 1731 468 1765 502
rect 1731 400 1765 434
rect 1855 536 1889 570
rect 1855 468 1889 502
rect 1855 400 1889 434
rect 2091 536 2125 570
rect 2091 468 2125 502
rect 2091 400 2125 434
rect 1259 276 1293 310
rect 1259 208 1293 242
rect 1259 140 1293 174
rect 1495 276 1529 310
rect 1495 208 1529 242
rect 1495 140 1529 174
rect 1731 276 1765 310
rect 1731 208 1765 242
rect 1731 140 1765 174
rect 1855 276 1889 310
rect 1855 208 1889 242
rect 1855 140 1889 174
rect 2091 276 2125 310
rect 2091 208 2125 242
rect 2091 140 2125 174
<< mvpdiffc >>
rect -17 824 17 858
rect -17 756 17 790
rect -17 688 17 722
rect 139 824 173 858
rect 139 756 173 790
rect 549 880 583 914
rect 549 812 583 846
rect 139 688 173 722
rect 249 709 283 743
rect 249 641 283 675
rect 249 573 283 607
rect 425 709 459 743
rect 549 744 583 778
rect 705 880 739 914
rect 705 812 739 846
rect 705 744 739 778
rect 425 641 459 675
rect 425 573 459 607
rect 549 607 583 641
rect 549 539 583 573
rect -17 409 17 443
rect -17 341 17 375
rect -17 273 17 307
rect 139 409 173 443
rect 549 471 583 505
rect 705 607 739 641
rect 705 539 739 573
rect 705 471 739 505
rect 139 341 173 375
rect 139 273 173 307
rect 249 340 283 374
rect 249 272 283 306
rect 249 204 283 238
rect 425 340 459 374
rect 425 272 459 306
rect 425 204 459 238
rect 549 334 583 368
rect 549 266 583 300
rect 549 198 583 232
rect 705 334 739 368
rect 705 266 739 300
rect 705 198 739 232
<< psubdiff >>
rect 665 2000 699 2024
rect 665 1923 699 1966
rect 665 1846 699 1889
rect 665 1769 699 1812
rect 665 1691 699 1735
rect 665 1613 699 1657
rect 665 1535 699 1579
rect 665 1477 699 1501
rect 2503 2145 2537 2169
rect 2503 2076 2537 2111
rect 2503 2007 2537 2042
rect 2503 1938 2537 1973
rect 2503 1869 2537 1904
rect 2503 1800 2537 1835
rect 2503 1731 2537 1766
rect 2503 1662 2537 1697
rect 2503 1594 2537 1628
rect 2503 1526 2537 1560
rect 2503 1458 2537 1492
rect 2503 1390 2537 1424
rect 2503 1322 2537 1356
rect 2503 1254 2537 1288
rect 2503 1186 2537 1220
rect 2503 1118 2537 1152
rect 2503 1050 2537 1084
rect 2503 982 2537 1016
rect 2503 914 2537 948
rect 2503 846 2537 880
rect 2503 778 2537 812
rect 2503 710 2537 744
rect 2503 642 2537 676
rect 2503 574 2537 608
rect 2503 506 2537 540
rect 2503 438 2537 472
rect 2503 370 2537 404
rect 2503 302 2537 336
rect 2503 234 2537 268
rect 2503 166 2537 200
rect 2503 108 2537 132
<< mvpsubdiff >>
rect 1079 830 1161 854
rect 1079 796 1103 830
rect 1137 796 1161 830
rect 1079 762 1161 796
rect 1079 728 1103 762
rect 1137 728 1161 762
rect 1079 694 1161 728
rect 1079 660 1103 694
rect 1137 660 1161 694
rect 1079 626 1161 660
rect 1079 592 1103 626
rect 1137 592 1161 626
rect 1079 558 1161 592
rect 1079 524 1103 558
rect 1137 524 1161 558
rect 1079 490 1161 524
rect 1079 456 1103 490
rect 1137 456 1161 490
rect 1079 422 1161 456
rect 1079 388 1103 422
rect 1137 388 1161 422
rect 1079 354 1161 388
rect 1079 320 1103 354
rect 1137 320 1161 354
rect 1079 286 1161 320
rect 1079 252 1103 286
rect 1137 252 1161 286
rect 1079 218 1161 252
rect 1079 184 1103 218
rect 1137 184 1161 218
rect 1079 150 1161 184
rect 1079 116 1103 150
rect 1137 116 1161 150
rect 1079 92 1161 116
<< mvnsubdiff >>
rect 853 731 887 755
rect 853 662 887 697
rect 853 593 887 628
rect 853 524 887 559
rect 853 454 887 490
rect 853 384 887 420
rect 853 314 887 350
rect 853 244 887 280
rect 853 186 887 210
<< psubdiffcont >>
rect 665 1966 699 2000
rect 665 1889 699 1923
rect 665 1812 699 1846
rect 665 1735 699 1769
rect 665 1657 699 1691
rect 665 1579 699 1613
rect 665 1501 699 1535
rect 2503 2111 2537 2145
rect 2503 2042 2537 2076
rect 2503 1973 2537 2007
rect 2503 1904 2537 1938
rect 2503 1835 2537 1869
rect 2503 1766 2537 1800
rect 2503 1697 2537 1731
rect 2503 1628 2537 1662
rect 2503 1560 2537 1594
rect 2503 1492 2537 1526
rect 2503 1424 2537 1458
rect 2503 1356 2537 1390
rect 2503 1288 2537 1322
rect 2503 1220 2537 1254
rect 2503 1152 2537 1186
rect 2503 1084 2537 1118
rect 2503 1016 2537 1050
rect 2503 948 2537 982
rect 2503 880 2537 914
rect 2503 812 2537 846
rect 2503 744 2537 778
rect 2503 676 2537 710
rect 2503 608 2537 642
rect 2503 540 2537 574
rect 2503 472 2537 506
rect 2503 404 2537 438
rect 2503 336 2537 370
rect 2503 268 2537 302
rect 2503 200 2537 234
rect 2503 132 2537 166
<< mvpsubdiffcont >>
rect 1103 796 1137 830
rect 1103 728 1137 762
rect 1103 660 1137 694
rect 1103 592 1137 626
rect 1103 524 1137 558
rect 1103 456 1137 490
rect 1103 388 1137 422
rect 1103 320 1137 354
rect 1103 252 1137 286
rect 1103 184 1137 218
rect 1103 116 1137 150
<< mvnsubdiffcont >>
rect 853 697 887 731
rect 853 628 887 662
rect 853 559 887 593
rect 853 490 887 524
rect 853 420 887 454
rect 853 350 887 384
rect 853 280 887 314
rect 853 210 887 244
<< poly >>
rect 1311 2278 1720 2294
rect 1311 2244 1329 2278
rect 1363 2244 1397 2278
rect 1431 2244 1465 2278
rect 1499 2244 1533 2278
rect 1567 2244 1601 2278
rect 1635 2244 1669 2278
rect 1703 2244 1720 2278
rect 1311 2228 1720 2244
rect 1311 2202 1411 2228
rect 1620 2202 1720 2228
rect 1900 2278 2080 2294
rect 1900 2244 1939 2278
rect 1973 2244 2007 2278
rect 2041 2244 2080 2278
rect 1900 2202 2080 2244
rect 2251 2278 2385 2294
rect 2251 2244 2267 2278
rect 2301 2244 2335 2278
rect 2369 2244 2385 2278
rect 2251 2228 2385 2244
rect 2260 2202 2290 2228
rect 2346 2202 2376 2228
rect 822 2120 956 2136
rect 822 2086 838 2120
rect 872 2086 906 2120
rect 940 2086 956 2120
rect 822 2050 956 2086
rect 1005 2120 1139 2136
rect 1005 2086 1021 2120
rect 1055 2086 1089 2120
rect 1123 2086 1139 2120
rect 1005 2050 1139 2086
rect 829 2024 949 2050
rect 1005 2024 1125 2050
rect 829 1850 949 1884
rect 1005 1850 1125 1884
rect 820 1834 954 1850
rect 820 1800 836 1834
rect 870 1800 904 1834
rect 938 1800 954 1834
rect 820 1784 954 1800
rect 1001 1834 1135 1850
rect 1001 1800 1017 1834
rect 1051 1800 1085 1834
rect 1119 1800 1135 1834
rect 1001 1784 1135 1800
rect 829 1748 949 1784
rect 1005 1748 1125 1784
rect 829 1582 949 1608
rect 1005 1582 1125 1608
rect 86 1282 206 1308
rect 262 1282 382 1308
rect 826 1249 946 1275
rect 1002 1249 1122 1275
rect 86 1116 206 1142
rect 262 1116 382 1142
rect 86 1050 414 1116
rect 1900 1942 2080 2002
rect 2260 1942 2290 2002
rect 2346 1942 2376 2002
rect 1900 1682 2080 1742
rect 2260 1682 2290 1742
rect 2346 1682 2376 1742
rect 2824 1590 2874 1622
rect 2930 1590 2980 1622
rect 1900 1422 2080 1482
rect 2260 1422 2290 1482
rect 2346 1422 2376 1482
rect 1311 1176 1411 1202
rect 1620 1176 1720 1202
rect 1900 1182 2080 1222
rect 2260 1196 2290 1222
rect 2346 1196 2376 1222
rect 1900 1148 1939 1182
rect 1973 1148 2007 1182
rect 2041 1148 2080 1182
rect 262 1034 414 1050
rect 28 967 206 983
rect 28 933 67 967
rect 101 933 135 967
rect 169 933 206 967
rect 28 885 206 933
rect 262 932 278 1034
rect 380 932 414 1034
rect 594 1092 694 1108
rect 594 1058 640 1092
rect 674 1058 694 1092
rect 594 1024 694 1058
rect 594 990 640 1024
rect 674 990 694 1024
rect 594 932 694 990
rect 826 1060 946 1109
rect 826 1026 896 1060
rect 930 1026 946 1060
rect 826 992 946 1026
rect 826 958 896 992
rect 930 958 946 992
rect 28 870 128 885
rect 262 781 414 932
rect 294 755 414 781
rect 28 644 128 670
rect 826 922 946 958
rect 1002 1040 1122 1109
rect 1304 1108 1484 1134
rect 1540 1108 1720 1134
rect 1900 1108 2080 1148
rect 2260 1108 2290 1134
rect 2346 1108 2376 1134
rect 1002 1006 1018 1040
rect 1052 1006 1122 1040
rect 1002 972 1122 1006
rect 1002 938 1018 972
rect 1052 938 1122 972
rect 1002 922 1122 938
rect 2824 958 2874 990
rect 1304 848 1484 908
rect 1540 848 1720 908
rect 1900 848 2080 908
rect 2260 848 2290 908
rect 2346 848 2376 908
rect 594 659 694 732
rect 294 503 414 555
rect 294 487 431 503
rect 28 455 128 481
rect 294 453 313 487
rect 347 453 381 487
rect 415 453 431 487
rect 294 437 431 453
rect 294 386 414 437
rect 594 386 694 459
rect 28 129 128 255
rect 2740 942 2874 958
rect 2740 908 2756 942
rect 2790 908 2824 942
rect 2858 908 2874 942
rect 2740 892 2874 908
rect 2930 958 2980 990
rect 2930 942 3064 958
rect 2930 908 2946 942
rect 2980 908 3014 942
rect 3048 908 3064 942
rect 2930 892 3064 908
rect 2740 867 2835 892
rect 2930 867 3049 892
rect 2679 851 2835 867
rect 2908 852 3049 867
rect 2679 817 2695 851
rect 2729 817 2785 851
rect 2819 817 2835 851
rect 2679 801 2835 817
rect 2679 772 2729 801
rect 2785 772 2835 801
rect 2891 851 3049 852
rect 2891 817 2924 851
rect 2958 817 2999 851
rect 3033 817 3049 851
rect 2891 801 3049 817
rect 2891 772 2941 801
rect 2997 772 3047 801
rect 1304 588 1484 648
rect 1540 588 1720 648
rect 1900 588 2080 648
rect 2260 588 2290 648
rect 2346 588 2376 648
rect 2679 546 2729 572
rect 2785 546 2835 572
rect 2891 546 2941 572
rect 2997 546 3047 572
rect 1304 328 1484 388
rect 1540 328 1720 388
rect 1900 328 2080 388
rect 2260 328 2290 388
rect 2346 328 2376 388
rect 294 160 414 186
rect 594 153 694 186
rect 28 87 189 129
rect 28 53 67 87
rect 101 53 135 87
rect 169 53 189 87
rect 594 121 728 153
rect 594 87 610 121
rect 644 87 678 121
rect 712 87 728 121
rect 1304 103 1484 128
rect 1540 103 1720 128
rect 1900 103 2080 128
rect 2260 103 2290 128
rect 2346 103 2376 128
rect 594 71 728 87
rect 1304 87 2080 103
rect 28 37 189 53
rect 1304 53 1328 87
rect 1362 53 1396 87
rect 1430 53 1464 87
rect 1498 53 1532 87
rect 1566 53 1600 87
rect 1634 53 1668 87
rect 1702 53 1736 87
rect 1770 53 1804 87
rect 1838 53 1872 87
rect 1906 53 1940 87
rect 1974 53 2008 87
rect 2042 53 2080 87
rect 1304 37 2080 53
rect 2251 87 2385 103
rect 2251 53 2267 87
rect 2301 53 2335 87
rect 2369 53 2385 87
rect 2251 37 2385 53
<< polycont >>
rect 1329 2244 1363 2278
rect 1397 2244 1431 2278
rect 1465 2244 1499 2278
rect 1533 2244 1567 2278
rect 1601 2244 1635 2278
rect 1669 2244 1703 2278
rect 1939 2244 1973 2278
rect 2007 2244 2041 2278
rect 2267 2244 2301 2278
rect 2335 2244 2369 2278
rect 838 2086 872 2120
rect 906 2086 940 2120
rect 1021 2086 1055 2120
rect 1089 2086 1123 2120
rect 836 1800 870 1834
rect 904 1800 938 1834
rect 1017 1800 1051 1834
rect 1085 1800 1119 1834
rect 1939 1148 1973 1182
rect 2007 1148 2041 1182
rect 67 933 101 967
rect 135 933 169 967
rect 278 932 380 1034
rect 640 1058 674 1092
rect 640 990 674 1024
rect 896 1026 930 1060
rect 896 958 930 992
rect 1018 1006 1052 1040
rect 1018 938 1052 972
rect 313 453 347 487
rect 381 453 415 487
rect 2756 908 2790 942
rect 2824 908 2858 942
rect 2946 908 2980 942
rect 3014 908 3048 942
rect 2695 817 2729 851
rect 2785 817 2819 851
rect 2924 817 2958 851
rect 2999 817 3033 851
rect 67 53 101 87
rect 135 53 169 87
rect 610 87 644 121
rect 678 87 712 121
rect 1328 53 1362 87
rect 1396 53 1430 87
rect 1464 53 1498 87
rect 1532 53 1566 87
rect 1600 53 1634 87
rect 1668 53 1702 87
rect 1736 53 1770 87
rect 1804 53 1838 87
rect 1872 53 1906 87
rect 1940 53 1974 87
rect 2008 53 2042 87
rect 2267 53 2301 87
rect 2335 53 2369 87
<< locali >>
rect 2251 2317 2385 2323
rect 2251 2283 2279 2317
rect 2313 2283 2351 2317
rect 2251 2278 2385 2283
rect 1313 2244 1329 2278
rect 1363 2244 1397 2278
rect 1431 2244 1465 2278
rect 1499 2244 1533 2278
rect 1567 2244 1601 2278
rect 1635 2244 1669 2278
rect 1703 2244 1719 2278
rect 1923 2244 1939 2278
rect 1973 2244 2007 2278
rect 2041 2244 2057 2278
rect 2251 2244 2267 2278
rect 2301 2244 2335 2278
rect 2369 2244 2385 2278
rect 822 2120 1153 2198
rect 1266 2190 1300 2206
rect 1266 2122 1300 2156
rect 822 2086 838 2120
rect 872 2086 906 2120
rect 940 2086 956 2120
rect 1005 2086 1021 2120
rect 1055 2086 1089 2120
rect 1123 2086 1139 2120
rect 665 2000 699 2024
rect 665 1923 699 1966
rect 665 1849 699 1889
rect 665 1777 699 1812
rect 665 1705 699 1735
rect 665 1633 699 1657
rect 736 1998 818 2014
rect 736 1964 784 1998
rect 736 1930 818 1964
rect 736 1896 784 1930
rect 960 1998 994 2014
rect 960 1930 994 1964
rect 736 1880 818 1896
rect 922 1880 960 1914
rect 736 1758 785 1880
rect 1028 1842 1102 2086
rect 1266 2054 1300 2088
rect 1266 2014 1300 2020
rect 1136 1998 1300 2014
rect 1170 1986 1300 1998
rect 1170 1964 1266 1986
rect 1136 1952 1266 1964
rect 1136 1930 1300 1952
rect 1170 1918 1300 1930
rect 1170 1896 1266 1918
rect 1136 1884 1266 1896
rect 1136 1880 1300 1884
rect 1169 1850 1300 1880
rect 820 1834 1135 1842
rect 820 1800 836 1834
rect 870 1800 904 1834
rect 938 1800 1017 1834
rect 1051 1800 1085 1834
rect 1119 1800 1135 1834
rect 820 1798 1135 1800
rect 1169 1816 1266 1850
rect 1169 1782 1300 1816
rect 736 1724 781 1758
rect 815 1724 818 1738
rect 736 1722 818 1724
rect 736 1688 784 1722
rect 922 1718 960 1752
rect 1169 1751 1266 1782
rect 736 1686 818 1688
rect 736 1652 781 1686
rect 815 1654 818 1686
rect 736 1620 784 1652
rect 736 1604 818 1620
rect 960 1654 994 1688
rect 960 1604 994 1620
rect 1103 1722 1142 1751
rect 1176 1748 1266 1751
rect 1103 1688 1136 1722
rect 1176 1717 1300 1748
rect 1170 1714 1300 1717
rect 1170 1688 1266 1714
rect 1103 1680 1266 1688
rect 1103 1679 1300 1680
rect 1103 1654 1142 1679
rect 1103 1620 1136 1654
rect 1176 1646 1300 1679
rect 1176 1645 1266 1646
rect 1170 1620 1266 1645
rect 1103 1612 1266 1620
rect 665 1561 699 1579
rect 1103 1578 1300 1612
rect 1103 1544 1266 1578
rect 665 1477 699 1501
rect 806 1489 844 1523
rect 1103 1510 1300 1544
rect 41 1270 95 1286
rect 75 1236 95 1270
rect 41 1202 95 1236
rect 75 1168 95 1202
rect 41 1118 95 1168
rect 323 1403 641 1443
rect 323 1369 409 1403
rect 443 1369 481 1403
rect 515 1369 641 1403
rect 323 1331 641 1369
rect 323 1320 494 1331
rect 482 1297 494 1320
rect 528 1297 566 1331
rect 600 1297 641 1331
rect 393 1270 448 1286
rect 217 1202 251 1236
rect 217 1152 251 1168
rect 427 1236 448 1270
rect 482 1265 641 1297
rect 393 1202 448 1236
rect 427 1200 448 1202
rect 781 1237 815 1489
rect 427 1168 487 1200
rect 393 1118 487 1168
rect 41 1084 487 1118
rect 781 1169 815 1203
rect 278 1034 380 1050
rect 51 933 67 967
rect 122 933 135 967
rect -17 858 17 874
rect -17 790 17 824
rect -17 722 17 756
rect -17 443 17 688
rect 51 481 105 933
rect 308 910 346 932
rect 274 899 380 910
rect 139 862 380 899
rect 139 858 173 862
rect 139 790 173 824
rect 249 756 283 759
rect 139 722 173 756
rect 139 672 173 688
rect 233 743 283 756
rect 233 709 249 743
rect 233 675 283 709
rect 233 641 249 675
rect 233 607 283 641
rect 233 573 249 607
rect 233 557 283 573
rect 51 447 173 481
rect -17 375 17 409
rect -17 307 17 341
rect -17 222 17 260
rect 139 443 173 447
rect 139 375 173 409
rect 139 307 173 341
rect 139 257 173 273
rect 233 390 273 557
rect 341 503 380 862
rect 414 791 487 1084
rect 640 1092 674 1108
rect 640 1024 674 1058
rect 425 743 487 791
rect 459 709 487 743
rect 425 675 487 709
rect 459 641 487 675
rect 425 607 487 641
rect 459 573 487 607
rect 425 557 487 573
rect 313 487 415 503
rect 347 453 381 487
rect 313 437 415 453
rect 233 374 283 390
rect 233 340 249 374
rect 233 306 283 340
rect 233 272 249 306
rect 233 260 269 272
rect 233 238 303 260
rect 233 204 249 238
rect 283 222 303 238
rect 233 188 269 204
rect -17 150 17 188
rect 337 87 391 437
rect 453 390 487 557
rect 425 374 487 390
rect 459 340 487 374
rect 425 306 487 340
rect 459 272 487 306
rect 425 238 487 272
rect 459 204 487 238
rect 425 188 487 204
rect 546 938 583 990
rect 640 974 674 990
rect 580 914 583 938
rect 781 938 815 1135
rect 957 1443 991 1486
rect 957 1371 991 1409
rect 957 1299 991 1337
rect 957 1237 991 1265
rect 957 1169 991 1203
rect 957 1119 991 1135
rect 1103 1476 1266 1510
rect 1103 1442 1300 1476
rect 1103 1408 1266 1442
rect 1103 1374 1300 1408
rect 1103 1340 1266 1374
rect 1103 1306 1300 1340
rect 1103 1272 1266 1306
rect 1103 1256 1300 1272
rect 1422 2190 1456 2206
rect 1422 2122 1456 2156
rect 1422 2054 1456 2088
rect 1422 1986 1456 2020
rect 1422 1918 1456 1952
rect 1422 1850 1456 1884
rect 1422 1782 1456 1816
rect 1422 1714 1456 1748
rect 1422 1646 1456 1680
rect 1422 1578 1456 1612
rect 1422 1510 1456 1544
rect 1575 2190 1609 2206
rect 1575 2122 1609 2156
rect 1575 2054 1609 2088
rect 1575 1986 1609 2020
rect 1575 1918 1609 1952
rect 1575 1850 1609 1884
rect 1575 1782 1609 1816
rect 1575 1714 1609 1748
rect 1575 1646 1609 1680
rect 1575 1578 1609 1612
rect 1575 1523 1609 1544
rect 1731 2190 1889 2206
rect 1765 2184 1889 2190
rect 1765 2156 1855 2184
rect 1731 2150 1855 2156
rect 1731 2122 1889 2150
rect 1765 2116 1889 2122
rect 1765 2088 1855 2116
rect 1731 2082 1855 2088
rect 1731 2054 1889 2082
rect 1765 2048 1889 2054
rect 1765 2020 1855 2048
rect 1731 2014 1855 2020
rect 1731 1986 1889 2014
rect 1765 1952 1889 1986
rect 1731 1924 1889 1952
rect 1731 1918 1855 1924
rect 1765 1890 1855 1918
rect 1765 1884 1889 1890
rect 1731 1856 1889 1884
rect 1731 1850 1855 1856
rect 1765 1822 1855 1850
rect 1765 1816 1889 1822
rect 1731 1788 1889 1816
rect 1731 1782 1855 1788
rect 1765 1754 1855 1782
rect 1765 1748 1889 1754
rect 1731 1714 1889 1748
rect 1765 1680 1889 1714
rect 1731 1664 1889 1680
rect 1731 1646 1855 1664
rect 1765 1630 1855 1646
rect 1765 1612 1889 1630
rect 1731 1596 1889 1612
rect 1731 1578 1855 1596
rect 1765 1562 1855 1578
rect 1765 1544 1889 1562
rect 1731 1528 1889 1544
rect 1553 1510 1591 1523
rect 1553 1489 1575 1510
rect 1731 1510 1855 1528
rect 1422 1442 1456 1476
rect 1422 1374 1456 1408
rect 1422 1306 1456 1340
rect 1103 1237 1209 1256
rect 1103 1203 1133 1237
rect 1167 1203 1209 1237
rect 1103 1169 1209 1203
rect 1422 1180 1456 1272
rect 1575 1442 1609 1476
rect 1575 1374 1609 1408
rect 1575 1306 1609 1340
rect 1575 1256 1609 1272
rect 1765 1494 1855 1510
rect 1765 1476 1889 1494
rect 1731 1442 1889 1476
rect 1765 1408 1889 1442
rect 1731 1404 1889 1408
rect 1731 1374 1855 1404
rect 1765 1370 1855 1374
rect 1765 1340 1889 1370
rect 1731 1336 1889 1340
rect 1731 1306 1855 1336
rect 1765 1302 1855 1306
rect 1765 1272 1889 1302
rect 1731 1268 1889 1272
rect 1731 1256 1855 1268
rect 1103 1135 1133 1169
rect 1167 1135 1209 1169
rect 896 1060 930 1076
rect 896 1018 930 1026
rect 887 992 925 1018
rect 887 984 896 992
rect 1002 1006 1018 1040
rect 1052 1006 1068 1040
rect 896 942 930 958
rect 1002 972 1068 1006
rect 1103 1018 1209 1135
rect 1137 984 1175 1018
rect 1259 1140 1765 1180
rect 1259 1090 1293 1140
rect 1259 1022 1293 1056
rect 1002 944 1018 972
rect 1052 944 1068 972
rect 1259 954 1293 988
rect 546 880 549 904
rect 546 866 583 880
rect 580 846 583 866
rect 546 812 549 832
rect 546 778 583 812
rect 546 744 549 778
rect 546 641 583 744
rect 546 607 549 641
rect 546 573 583 607
rect 546 539 549 573
rect 546 505 583 539
rect 546 471 549 505
rect 546 368 583 471
rect 546 334 549 368
rect 546 300 583 334
rect 546 266 549 300
rect 546 232 583 266
rect 546 198 549 232
rect 546 182 583 198
rect 705 914 739 930
rect 705 846 739 880
rect 1052 938 1074 944
rect 1036 910 1074 938
rect 781 866 815 904
rect 705 778 739 812
rect 1103 830 1137 846
rect 1103 762 1137 796
rect 705 641 739 744
rect 705 573 739 607
rect 705 505 739 539
rect 705 368 739 471
rect 705 300 739 334
rect 705 232 739 260
rect 705 182 739 188
rect 853 731 887 755
rect 853 662 887 697
rect 853 593 887 628
rect 853 524 887 559
rect 853 454 887 490
rect 1103 694 1137 728
rect 1103 626 1137 660
rect 1103 558 1137 592
rect 1103 490 1137 524
rect 1103 452 1137 456
rect 853 384 887 420
rect 853 314 887 350
rect 853 244 887 260
rect 853 150 887 188
rect 594 87 610 121
rect 644 87 678 121
rect 712 87 728 121
rect 1103 286 1137 320
rect 1103 218 1137 252
rect 1103 150 1137 184
rect 1259 830 1293 920
rect 1259 762 1293 796
rect 1259 694 1293 728
rect 1259 570 1293 660
rect 1259 502 1293 536
rect 1259 434 1293 468
rect 1259 310 1293 400
rect 1259 242 1293 276
rect 1259 174 1293 208
rect 1259 124 1293 140
rect 1495 1090 1529 1106
rect 1495 1022 1529 1056
rect 1495 954 1529 988
rect 1495 830 1529 916
rect 1495 762 1529 796
rect 1495 694 1529 728
rect 1495 570 1529 660
rect 1495 502 1529 536
rect 1495 434 1529 468
rect 1495 310 1529 400
rect 1495 242 1529 276
rect 1495 174 1529 208
rect 1495 124 1529 140
rect 1731 1090 1765 1140
rect 1731 1022 1765 1056
rect 1731 954 1765 988
rect 1731 830 1765 920
rect 1731 762 1765 796
rect 1731 694 1765 728
rect 1731 570 1765 660
rect 1731 502 1765 536
rect 1731 434 1765 468
rect 1731 310 1765 400
rect 1731 242 1765 276
rect 1731 174 1765 208
rect 1731 124 1765 140
rect 1855 1090 1889 1234
rect 1855 1022 1889 1056
rect 1855 954 1889 988
rect 1855 830 1889 920
rect 1855 762 1889 796
rect 1855 694 1889 728
rect 1855 570 1889 660
rect 1855 502 1889 536
rect 1855 434 1889 468
rect 1855 310 1889 400
rect 1855 242 1889 276
rect 1855 174 1889 208
rect 1855 124 1889 140
rect 1923 2090 2057 2244
rect 1923 1912 1937 2090
rect 2043 1912 2057 2090
rect 1923 1182 2057 1912
rect 1923 1148 1939 1182
rect 1973 1148 2007 1182
rect 2041 1148 2057 1182
rect 1103 100 1137 116
rect 1923 90 2057 1148
rect 2091 2184 2125 2200
rect 2091 2116 2125 2150
rect 2091 2048 2125 2082
rect 2091 1924 2125 2014
rect 2091 1856 2125 1890
rect 2091 1788 2125 1810
rect 2091 1664 2125 1738
rect 2091 1596 2125 1630
rect 2091 1528 2125 1562
rect 2091 1404 2125 1494
rect 2091 1336 2125 1370
rect 2091 1268 2125 1302
rect 2091 1090 2125 1234
rect 2091 1022 2125 1056
rect 2091 954 2125 988
rect 2091 830 2125 920
rect 2091 762 2125 796
rect 2091 694 2125 728
rect 2091 570 2125 660
rect 2091 502 2125 536
rect 2091 434 2125 468
rect 2091 310 2125 400
rect 2091 242 2125 276
rect 2091 174 2125 208
rect 2091 124 2125 140
rect 2159 2184 2267 2200
rect 2159 2150 2215 2184
rect 2249 2150 2267 2184
rect 2159 2116 2267 2150
rect 2159 2082 2215 2116
rect 2249 2082 2267 2116
rect 2159 2048 2267 2082
rect 2159 2014 2215 2048
rect 2249 2014 2267 2048
rect 2159 1924 2267 2014
rect 2159 1890 2215 1924
rect 2249 1890 2267 1924
rect 2159 1856 2267 1890
rect 2159 1822 2215 1856
rect 2249 1822 2267 1856
rect 2159 1788 2267 1822
rect 2159 1754 2215 1788
rect 2249 1754 2267 1788
rect 2159 1664 2267 1754
rect 2159 1630 2215 1664
rect 2249 1630 2267 1664
rect 2159 1596 2267 1630
rect 2159 1562 2215 1596
rect 2249 1562 2267 1596
rect 2159 1528 2267 1562
rect 2159 1494 2215 1528
rect 2249 1494 2267 1528
rect 2159 1443 2267 1494
rect 2159 1409 2202 1443
rect 2236 1409 2267 1443
rect 2159 1404 2267 1409
rect 2159 1371 2215 1404
rect 2159 1337 2202 1371
rect 2249 1370 2267 1404
rect 2236 1337 2267 1370
rect 2159 1336 2267 1337
rect 2159 1302 2215 1336
rect 2249 1302 2267 1336
rect 2159 1299 2267 1302
rect 2159 1265 2202 1299
rect 2236 1268 2267 1299
rect 2159 1234 2215 1265
rect 2249 1234 2267 1268
rect 2159 1090 2267 1234
rect 2301 2184 2335 2200
rect 2301 2116 2335 2150
rect 2301 2048 2335 2082
rect 2301 1924 2335 2014
rect 2301 1856 2335 1890
rect 2301 1788 2335 1810
rect 2301 1664 2335 1738
rect 2301 1596 2335 1630
rect 2301 1528 2335 1562
rect 2301 1404 2335 1494
rect 2301 1336 2335 1370
rect 2301 1268 2335 1302
rect 2301 1218 2335 1234
rect 2369 2184 2537 2200
rect 2369 2150 2387 2184
rect 2421 2150 2537 2184
rect 2369 2145 2537 2150
rect 2369 2116 2503 2145
rect 2369 2082 2387 2116
rect 2421 2111 2503 2116
rect 2421 2082 2537 2111
rect 2369 2076 2537 2082
rect 2369 2048 2503 2076
rect 2369 2014 2387 2048
rect 2421 2042 2503 2048
rect 2421 2014 2537 2042
rect 2369 2007 2537 2014
rect 2369 1973 2503 2007
rect 2369 1938 2537 1973
rect 2369 1924 2503 1938
rect 2369 1890 2387 1924
rect 2421 1904 2503 1924
rect 2421 1890 2537 1904
rect 2369 1869 2537 1890
rect 2369 1856 2503 1869
rect 2369 1822 2387 1856
rect 2421 1835 2503 1856
rect 2421 1822 2537 1835
rect 2369 1800 2537 1822
rect 2369 1788 2503 1800
rect 2369 1754 2387 1788
rect 2421 1766 2503 1788
rect 2421 1754 2537 1766
rect 2369 1731 2537 1754
rect 2369 1697 2503 1731
rect 2369 1664 2537 1697
rect 2848 1705 2956 1734
rect 2369 1630 2387 1664
rect 2421 1662 2537 1664
rect 2421 1630 2503 1662
rect 2369 1628 2503 1630
rect 2369 1596 2537 1628
rect 2369 1562 2387 1596
rect 2421 1594 2537 1596
rect 2421 1562 2503 1594
rect 2369 1560 2503 1562
rect 2805 1662 2813 1696
rect 2771 1624 2813 1662
rect 2805 1590 2813 1624
rect 2369 1528 2537 1560
rect 2779 1578 2813 1590
rect 2369 1494 2387 1528
rect 2421 1526 2537 1528
rect 2421 1494 2503 1526
rect 2369 1492 2503 1494
rect 2369 1458 2537 1492
rect 2369 1443 2503 1458
rect 2369 1409 2387 1443
rect 2421 1409 2503 1443
rect 2369 1404 2537 1409
rect 2369 1337 2387 1404
rect 2421 1390 2537 1404
rect 2421 1337 2503 1390
rect 2369 1336 2537 1337
rect 2369 1302 2387 1336
rect 2421 1322 2537 1336
rect 2421 1302 2503 1322
rect 2369 1299 2503 1302
rect 2369 1234 2387 1299
rect 2421 1265 2503 1299
rect 2421 1254 2537 1265
rect 2421 1234 2503 1254
rect 2369 1220 2503 1234
rect 2369 1186 2537 1220
rect 2369 1152 2503 1186
rect 2369 1118 2537 1152
rect 2159 1056 2215 1090
rect 2249 1056 2267 1090
rect 2159 1022 2267 1056
rect 2159 988 2215 1022
rect 2249 988 2267 1022
rect 2159 954 2267 988
rect 2159 920 2215 954
rect 2249 920 2267 954
rect 2159 830 2267 920
rect 2159 796 2215 830
rect 2249 796 2267 830
rect 2159 762 2267 796
rect 2159 728 2215 762
rect 2249 728 2267 762
rect 2159 694 2267 728
rect 2159 660 2215 694
rect 2249 660 2267 694
rect 2159 570 2267 660
rect 2159 536 2215 570
rect 2249 536 2267 570
rect 2159 502 2267 536
rect 2159 468 2215 502
rect 2249 468 2267 502
rect 2159 452 2267 468
rect 2159 418 2203 452
rect 2237 434 2267 452
rect 2159 400 2215 418
rect 2249 400 2267 434
rect 2159 380 2267 400
rect 2159 346 2203 380
rect 2237 346 2267 380
rect 2159 310 2267 346
rect 2159 276 2215 310
rect 2249 276 2267 310
rect 2159 242 2267 276
rect 2159 208 2215 242
rect 2249 208 2267 242
rect 2159 174 2267 208
rect 2159 140 2215 174
rect 2249 140 2267 174
rect 2159 124 2267 140
rect 2301 1090 2335 1106
rect 2301 1022 2335 1056
rect 2301 954 2335 988
rect 2301 830 2335 916
rect 2301 762 2335 796
rect 2301 694 2335 728
rect 2301 570 2335 660
rect 2301 502 2335 536
rect 2301 434 2335 468
rect 2301 310 2335 400
rect 2301 242 2335 276
rect 2301 174 2335 208
rect 2301 124 2335 140
rect 2369 1090 2503 1118
rect 2369 1056 2387 1090
rect 2421 1084 2503 1090
rect 2421 1056 2537 1084
rect 2369 1050 2537 1056
rect 2369 1022 2503 1050
rect 2369 988 2387 1022
rect 2421 1016 2503 1022
rect 2421 988 2537 1016
rect 2369 982 2537 988
rect 2369 954 2503 982
rect 2369 920 2387 954
rect 2421 948 2503 954
rect 2421 920 2537 948
rect 2369 914 2537 920
rect 2369 880 2503 914
rect 2369 846 2537 880
rect 2369 830 2503 846
rect 2369 796 2387 830
rect 2421 812 2503 830
rect 2600 1542 2745 1549
rect 2600 1508 2612 1542
rect 2646 1508 2699 1542
rect 2733 1508 2745 1542
rect 2600 942 2745 1508
rect 2779 1510 2813 1544
rect 2779 1442 2813 1476
rect 2779 1374 2813 1408
rect 2779 1306 2813 1340
rect 2779 1238 2813 1272
rect 2779 1170 2813 1204
rect 2779 1102 2813 1136
rect 2779 1052 2813 1068
rect 2848 1671 2849 1705
rect 2883 1671 2922 1705
rect 2848 1633 2956 1671
rect 2848 1599 2849 1633
rect 2883 1599 2922 1633
rect 2848 1578 2956 1599
rect 2848 1544 2885 1578
rect 2919 1544 2956 1578
rect 2848 1510 2956 1544
rect 2848 1476 2885 1510
rect 2919 1476 2956 1510
rect 2848 1442 2956 1476
rect 2848 1408 2885 1442
rect 2919 1408 2956 1442
rect 2848 1374 2956 1408
rect 2848 1340 2885 1374
rect 2919 1340 2956 1374
rect 2848 1306 2956 1340
rect 2848 1272 2885 1306
rect 2919 1272 2956 1306
rect 2848 1238 2956 1272
rect 2848 1204 2885 1238
rect 2919 1204 2956 1238
rect 2848 1170 2956 1204
rect 2848 1136 2885 1170
rect 2919 1136 2956 1170
rect 2848 1102 2956 1136
rect 2848 1068 2885 1102
rect 2919 1068 2956 1102
rect 2848 1053 2956 1068
rect 2991 1620 3034 1625
rect 2991 1586 3000 1620
rect 2991 1578 3034 1586
rect 3025 1548 3034 1578
rect 2991 1514 3000 1544
rect 2991 1510 3034 1514
rect 3025 1476 3034 1510
rect 2991 1472 3034 1476
rect 2991 1442 3025 1472
rect 2991 1374 3025 1408
rect 2991 1306 3025 1340
rect 2991 1238 3025 1272
rect 2991 1170 3025 1204
rect 2991 1102 3025 1136
rect 2885 1052 2919 1053
rect 2991 1052 3025 1068
rect 2971 942 3009 944
rect 2600 908 2756 942
rect 2790 908 2824 942
rect 2858 908 2874 942
rect 2930 910 2937 942
rect 2980 910 3009 942
rect 2930 908 2946 910
rect 2980 908 3014 910
rect 3048 908 3064 942
rect 2600 851 2835 908
rect 2930 851 3049 908
rect 2600 817 2695 851
rect 2729 817 2785 851
rect 2819 817 2835 851
rect 2908 817 2924 851
rect 2958 817 2999 851
rect 3033 817 3049 851
rect 2421 796 2537 812
rect 2369 778 2537 796
rect 2369 762 2503 778
rect 2369 728 2387 762
rect 2421 744 2503 762
rect 2421 728 2537 744
rect 2369 710 2537 728
rect 2369 694 2503 710
rect 2369 660 2387 694
rect 2421 676 2503 694
rect 2421 660 2537 676
rect 2369 642 2537 660
rect 2369 608 2503 642
rect 2369 574 2537 608
rect 2369 570 2503 574
rect 2369 536 2387 570
rect 2421 540 2503 570
rect 2634 754 2668 770
rect 2740 754 2778 783
rect 2634 703 2668 720
rect 2634 631 2668 652
rect 2634 568 2668 584
rect 2774 749 2778 754
rect 2846 754 2880 770
rect 2740 686 2774 720
rect 2740 618 2774 652
rect 2740 568 2774 584
rect 2950 754 2988 783
rect 2950 749 2952 754
rect 2846 703 2880 720
rect 2846 631 2880 652
rect 2846 568 2880 584
rect 2986 749 2988 754
rect 3058 754 3092 770
rect 2952 686 2986 720
rect 2952 618 2986 652
rect 2952 568 2986 584
rect 3058 703 3092 720
rect 3058 631 3092 652
rect 3058 568 3092 584
rect 2421 536 2537 540
rect 2369 506 2537 536
rect 2369 502 2503 506
rect 2369 468 2387 502
rect 2421 472 2503 502
rect 2421 468 2537 472
rect 2369 452 2537 468
rect 2369 400 2387 452
rect 2421 404 2503 452
rect 2421 400 2537 404
rect 2369 380 2537 400
rect 2369 346 2387 380
rect 2421 346 2503 380
rect 2369 336 2503 346
rect 2369 310 2537 336
rect 2369 276 2387 310
rect 2421 302 2537 310
rect 2421 276 2503 302
rect 2369 268 2503 276
rect 2369 242 2537 268
rect 2369 208 2387 242
rect 2421 234 2537 242
rect 2421 208 2503 234
rect 2369 200 2503 208
rect 2369 174 2537 200
rect 2369 140 2387 174
rect 2421 166 2537 174
rect 2421 140 2503 166
rect 2369 132 2503 140
rect 2369 124 2537 132
rect 2503 108 2537 124
rect 1312 87 2058 90
rect 51 53 67 87
rect 101 53 135 87
rect 169 53 391 87
rect 1312 53 1328 87
rect 1362 53 1396 87
rect 1430 53 1464 87
rect 1498 53 1532 87
rect 1566 53 1600 87
rect 1634 53 1668 87
rect 1702 53 1736 87
rect 1770 53 1804 87
rect 1838 53 1872 87
rect 1906 53 1940 87
rect 1974 53 2008 87
rect 2042 53 2058 87
rect 1312 26 2058 53
rect 2251 66 2267 87
rect 2301 66 2335 87
rect 2251 40 2262 66
rect 2301 53 2334 66
rect 2369 53 2385 87
rect 2296 32 2334 53
rect 2368 40 2385 53
<< viali >>
rect 2279 2283 2313 2317
rect 2351 2283 2385 2317
rect 665 1846 699 1849
rect 665 1815 699 1846
rect 665 1769 699 1777
rect 665 1743 699 1769
rect 665 1691 699 1705
rect 665 1671 699 1691
rect 665 1613 699 1633
rect 665 1599 699 1613
rect 888 1880 922 1914
rect 960 1896 994 1914
rect 960 1880 994 1896
rect 781 1724 815 1758
rect 888 1718 922 1752
rect 960 1722 994 1752
rect 960 1718 994 1722
rect 781 1654 815 1686
rect 781 1652 784 1654
rect 784 1652 815 1654
rect 1142 1722 1176 1751
rect 1142 1717 1170 1722
rect 1170 1717 1176 1722
rect 1142 1654 1176 1679
rect 1142 1645 1170 1654
rect 1170 1645 1176 1654
rect 665 1535 699 1561
rect 665 1527 699 1535
rect 772 1489 806 1523
rect 844 1489 878 1523
rect 217 1270 323 1443
rect 409 1369 443 1403
rect 481 1369 515 1403
rect 494 1297 528 1331
rect 566 1297 600 1331
rect 217 1265 251 1270
rect 251 1265 323 1270
rect 641 1265 747 1443
rect 88 933 101 967
rect 101 933 122 967
rect 160 933 169 967
rect 169 933 194 967
rect 274 932 278 944
rect 278 932 308 944
rect 346 932 380 944
rect 274 910 308 932
rect 346 910 380 932
rect -17 273 17 294
rect -17 260 17 273
rect 269 272 283 294
rect 283 272 303 294
rect 269 260 303 272
rect -17 188 17 222
rect 269 204 283 222
rect 283 204 303 222
rect 269 188 303 204
rect -17 116 17 150
rect 546 914 580 938
rect 957 1409 991 1443
rect 957 1337 991 1371
rect 957 1265 991 1299
rect 1519 1489 1553 1523
rect 1591 1510 1625 1523
rect 1591 1489 1609 1510
rect 1609 1489 1625 1510
rect 853 984 887 1018
rect 925 992 959 1018
rect 925 984 930 992
rect 930 984 959 992
rect 1103 984 1137 1018
rect 1175 984 1209 1018
rect 546 904 549 914
rect 549 904 580 914
rect 546 846 580 866
rect 546 832 549 846
rect 549 832 580 846
rect 781 904 815 938
rect 1002 938 1018 944
rect 1018 938 1036 944
rect 1002 910 1036 938
rect 1074 910 1108 944
rect 781 832 815 866
rect 705 266 739 294
rect 705 260 739 266
rect 705 198 739 222
rect 705 188 739 198
rect 959 422 1137 452
rect 959 388 1103 422
rect 1103 388 1137 422
rect 959 354 1137 388
rect 959 346 1103 354
rect 1103 346 1137 354
rect 853 280 887 294
rect 853 260 887 280
rect 853 210 887 222
rect 853 188 887 210
rect 853 116 887 150
rect 1495 988 1529 1022
rect 1495 920 1529 950
rect 1495 916 1529 920
rect 1937 1912 2043 2090
rect 2091 1822 2125 1844
rect 2091 1810 2125 1822
rect 2091 1754 2125 1772
rect 2091 1738 2125 1754
rect 2202 1409 2236 1443
rect 2202 1370 2215 1371
rect 2215 1370 2236 1371
rect 2202 1337 2236 1370
rect 2202 1268 2236 1299
rect 2202 1265 2215 1268
rect 2215 1265 2236 1268
rect 2301 1822 2335 1844
rect 2301 1810 2335 1822
rect 2301 1754 2335 1772
rect 2301 1738 2335 1754
rect 2771 1662 2805 1696
rect 2771 1590 2805 1624
rect 2387 1409 2421 1443
rect 2503 1424 2537 1443
rect 2503 1409 2537 1424
rect 2387 1370 2421 1371
rect 2387 1337 2421 1370
rect 2503 1356 2537 1371
rect 2503 1337 2537 1356
rect 2387 1268 2421 1299
rect 2387 1265 2421 1268
rect 2503 1288 2537 1299
rect 2503 1265 2537 1288
rect 2203 434 2237 452
rect 2203 418 2215 434
rect 2215 418 2237 434
rect 2203 346 2237 380
rect 2301 988 2335 1022
rect 2301 920 2335 950
rect 2301 916 2335 920
rect 2612 1508 2646 1542
rect 2699 1508 2733 1542
rect 2849 1671 2883 1705
rect 2922 1671 2956 1705
rect 2849 1599 2883 1633
rect 2922 1599 2956 1633
rect 3000 1586 3034 1620
rect 3000 1544 3025 1548
rect 3025 1544 3034 1548
rect 3000 1514 3034 1544
rect 2937 942 2971 944
rect 3009 942 3043 944
rect 2937 910 2946 942
rect 2946 910 2971 942
rect 3009 910 3014 942
rect 3014 910 3043 942
rect 2706 749 2740 783
rect 2634 686 2668 703
rect 2634 669 2668 686
rect 2634 618 2668 631
rect 2634 597 2668 618
rect 2778 749 2812 783
rect 2916 749 2950 783
rect 2846 686 2880 703
rect 2846 669 2880 686
rect 2846 618 2880 631
rect 2846 597 2880 618
rect 2988 749 3022 783
rect 3058 686 3092 703
rect 3058 669 3092 686
rect 3058 618 3092 631
rect 3058 597 3092 618
rect 2387 434 2421 452
rect 2387 418 2421 434
rect 2503 438 2537 452
rect 2503 418 2537 438
rect 2387 346 2421 380
rect 2503 370 2537 380
rect 2503 346 2537 370
rect 2262 53 2267 66
rect 2267 53 2296 66
rect 2334 53 2335 66
rect 2335 53 2368 66
rect 2262 32 2296 53
rect 2334 32 2368 53
<< metal1 >>
rect 2755 2323 2761 2329
rect 2267 2317 2761 2323
rect 2267 2283 2279 2317
rect 2313 2283 2351 2317
rect 2385 2283 2761 2317
rect 2267 2277 2761 2283
rect 2813 2277 2825 2329
rect 2877 2277 2883 2329
rect 738 2090 3312 2246
rect 738 1995 1937 2090
rect 876 1914 1006 1920
rect 876 1880 888 1914
rect 922 1880 960 1914
rect 994 1880 1006 1914
rect 1925 1912 1937 1995
rect 2043 1995 3312 2090
rect 2043 1912 2055 1995
tri 2431 1920 2506 1995 ne
rect 2506 1920 3312 1995
rect 1925 1906 2055 1912
tri 2506 1906 2520 1920 ne
rect 2520 1906 3312 1920
rect 876 1861 1006 1880
rect 659 1849 1006 1861
tri 2520 1850 2576 1906 ne
rect 2576 1850 3312 1906
rect 659 1815 665 1849
rect 699 1815 1006 1849
rect 659 1801 1006 1815
rect 659 1777 711 1801
rect 659 1743 665 1777
rect 699 1772 711 1777
tri 711 1772 740 1801 nw
rect 699 1743 705 1772
tri 705 1766 711 1772 nw
rect 659 1705 705 1743
rect 659 1671 665 1705
rect 699 1671 705 1705
rect 659 1633 705 1671
rect 775 1758 821 1770
rect 775 1724 781 1758
rect 815 1724 821 1758
rect 775 1686 821 1724
rect 876 1752 1006 1801
rect 2079 1844 2347 1850
rect 2079 1810 2091 1844
rect 2125 1810 2301 1844
rect 2335 1810 2347 1844
tri 2576 1839 2587 1850 ne
rect 2587 1839 3312 1850
rect 2079 1772 2347 1810
rect 876 1718 888 1752
rect 922 1718 960 1752
rect 994 1718 1006 1752
rect 876 1712 1006 1718
rect 1136 1751 1182 1763
rect 1136 1717 1142 1751
rect 1176 1717 1182 1751
rect 2079 1738 2091 1772
rect 2125 1738 2301 1772
rect 2335 1738 2347 1772
tri 2752 1748 2843 1839 ne
rect 2079 1732 2347 1738
rect 775 1652 781 1686
rect 815 1680 821 1686
rect 1136 1680 1182 1717
rect 815 1679 1182 1680
rect 815 1652 1142 1679
rect 775 1645 1142 1652
rect 1176 1645 1182 1679
rect 775 1640 1182 1645
rect 1136 1633 1182 1640
rect 2762 1702 2814 1708
rect 2762 1636 2814 1650
rect 659 1599 665 1633
rect 699 1599 705 1633
rect 659 1561 705 1599
rect 2843 1705 2962 1839
tri 2962 1768 3033 1839 nw
rect 2843 1671 2849 1705
rect 2883 1671 2922 1705
rect 2956 1671 2962 1705
rect 2843 1633 2962 1671
rect 2843 1599 2849 1633
rect 2883 1599 2922 1633
rect 2956 1599 2962 1633
rect 2843 1587 2962 1599
rect 2994 1626 3046 1632
rect 2762 1578 2814 1584
rect 659 1527 665 1561
rect 699 1527 705 1561
rect 2994 1560 3046 1574
rect 2600 1542 2994 1549
tri 630 1455 659 1484 se
rect 659 1483 705 1527
rect 760 1523 1637 1529
rect 760 1489 772 1523
rect 806 1489 844 1523
rect 878 1489 1519 1523
rect 1553 1489 1591 1523
rect 1625 1489 1637 1523
rect 2600 1508 2612 1542
rect 2646 1508 2699 1542
rect 2733 1508 2994 1542
rect 2600 1502 3046 1508
tri 705 1483 708 1486 sw
rect 760 1483 1637 1489
rect 659 1455 708 1483
tri 708 1455 736 1483 sw
rect -96 1443 3312 1455
rect -96 1265 217 1443
rect 323 1403 641 1443
rect 323 1369 409 1403
rect 443 1369 481 1403
rect 515 1369 641 1403
rect 323 1331 641 1369
rect 323 1297 494 1331
rect 528 1297 566 1331
rect 600 1297 641 1331
rect 323 1265 641 1297
rect 747 1409 957 1443
rect 991 1409 2202 1443
rect 2236 1409 2387 1443
rect 2421 1409 2503 1443
rect 2537 1409 3312 1443
rect 747 1371 3312 1409
rect 747 1337 957 1371
rect 991 1337 2202 1371
rect 2236 1337 2387 1371
rect 2421 1337 2503 1371
rect 2537 1337 3312 1371
rect 747 1299 3312 1337
rect 747 1265 957 1299
rect 991 1265 2202 1299
rect 2236 1265 2387 1299
rect 2421 1265 2503 1299
rect 2537 1265 3312 1299
rect -96 1253 3312 1265
tri 186 1022 188 1024 se
rect 188 1022 1221 1024
tri 182 1018 186 1022 se
rect 186 1018 1221 1022
tri 148 984 182 1018 se
rect 182 984 853 1018
rect 887 984 925 1018
rect 959 984 1103 1018
rect 1137 984 1175 1018
rect 1209 984 1221 1018
tri 143 979 148 984 se
rect 148 979 1221 984
rect 76 978 1221 979
rect 1489 1022 2347 1034
rect 1489 988 1495 1022
rect 1529 988 2301 1022
rect 2335 988 2347 1022
rect 76 969 218 978
tri 218 969 227 978 nw
rect 76 967 206 969
rect 76 933 88 967
rect 122 933 160 967
rect 194 933 206 967
tri 206 957 218 969 nw
rect 1489 950 2347 988
rect 76 927 206 933
rect 262 944 1120 950
rect 262 910 274 944
rect 308 910 346 944
rect 380 938 1002 944
rect 380 910 546 938
rect 262 904 546 910
rect 580 904 781 938
rect 815 910 1002 938
rect 1036 910 1074 944
rect 1108 910 1120 944
rect 815 904 1120 910
rect 1489 916 1495 950
rect 1529 916 2301 950
rect 2335 916 2347 950
rect 1489 904 2347 916
rect 2843 963 2895 969
tri 2895 950 2914 969 sw
rect 2895 944 3055 950
rect 2895 911 2937 944
rect 2843 910 2937 911
rect 2971 910 3009 944
rect 3043 910 3055 944
rect 2843 904 3055 910
rect 540 866 586 904
rect 540 832 546 866
rect 580 832 586 866
rect 540 820 586 832
rect 775 866 821 904
rect 2843 901 2918 904
tri 2918 901 2921 904 nw
rect 2843 899 2895 901
rect 775 832 781 866
rect 815 832 821 866
rect 775 820 821 832
rect 2731 867 2783 873
tri 2726 820 2731 825 se
tri 2695 789 2726 820 se
rect 2726 815 2731 820
tri 2895 878 2918 901 nw
rect 2843 841 2895 847
rect 2943 867 2995 873
tri 2940 825 2943 828 se
rect 2726 801 2783 815
rect 2726 789 2731 801
rect 2694 783 2731 789
tri 2783 789 2819 825 sw
tri 2904 789 2940 825 se
rect 2940 815 2943 825
rect 2940 801 2995 815
rect 2940 789 2943 801
rect 2783 783 2824 789
rect 2694 749 2706 783
rect 2812 749 2824 783
rect 2694 743 2824 749
rect 2904 783 2943 789
tri 2995 789 3034 828 sw
rect 2995 783 3034 789
rect 2904 749 2916 783
rect 3022 749 3034 783
rect 2904 743 3034 749
rect 2628 709 3148 715
rect 2628 703 2885 709
rect 2628 669 2634 703
rect 2668 669 2846 703
rect 2880 669 2885 703
rect 2628 657 2885 669
rect 2937 657 2993 709
rect 3045 703 3148 709
rect 3045 669 3058 703
rect 3092 669 3148 703
rect 3045 657 3148 669
rect 2628 637 3148 657
rect 2628 631 2885 637
rect 2628 597 2634 631
rect 2668 597 2846 631
rect 2880 597 2885 631
rect 2628 585 2885 597
rect 2937 585 2993 637
rect 3045 631 3148 637
rect 3045 597 3058 631
rect 3092 597 3148 631
rect 3045 585 3148 597
rect -179 452 2885 464
rect -179 346 959 452
rect 1137 418 2203 452
rect 2237 418 2387 452
rect 2421 418 2503 452
rect 2537 418 2885 452
rect 1137 412 2885 418
rect 2937 412 2993 464
rect 3045 412 3312 464
rect 1137 386 3312 412
rect 1137 380 2885 386
rect 1137 346 2203 380
rect 2237 346 2387 380
rect 2421 346 2503 380
rect 2537 346 2885 380
rect -179 334 2885 346
rect 2937 334 2993 386
rect 3045 334 3312 386
rect -179 294 3312 306
rect -179 260 -17 294
rect 17 260 269 294
rect 303 260 705 294
rect 739 260 853 294
rect 887 260 3312 294
rect -179 222 3312 260
rect -179 188 -17 222
rect 17 188 269 222
rect 303 188 705 222
rect 739 188 853 222
rect 887 188 3312 222
rect -179 150 3312 188
rect -179 116 -17 150
rect 17 116 853 150
rect 887 116 3312 150
rect -179 104 3312 116
tri 2680 72 2683 75 se
rect 2683 72 2689 75
rect 2250 66 2689 72
rect 2250 32 2262 66
rect 2296 32 2334 66
rect 2368 32 2689 66
rect 2250 26 2689 32
tri 2680 23 2683 26 ne
rect 2683 23 2689 26
rect 2741 23 2755 75
rect 2807 23 2813 75
<< via1 >>
rect 2761 2277 2813 2329
rect 2825 2277 2877 2329
rect 2762 1696 2814 1702
rect 2762 1662 2771 1696
rect 2771 1662 2805 1696
rect 2805 1662 2814 1696
rect 2762 1650 2814 1662
rect 2762 1624 2814 1636
rect 2762 1590 2771 1624
rect 2771 1590 2805 1624
rect 2805 1590 2814 1624
rect 2762 1584 2814 1590
rect 2994 1620 3046 1626
rect 2994 1586 3000 1620
rect 3000 1586 3034 1620
rect 3034 1586 3046 1620
rect 2994 1574 3046 1586
rect 2994 1548 3046 1560
rect 2994 1514 3000 1548
rect 3000 1514 3034 1548
rect 3034 1514 3046 1548
rect 2994 1508 3046 1514
rect 2843 911 2895 963
rect 2731 815 2783 867
rect 2843 847 2895 899
rect 2731 783 2783 801
rect 2943 815 2995 867
rect 2731 749 2740 783
rect 2740 749 2778 783
rect 2778 749 2783 783
rect 2943 783 2995 801
rect 2943 749 2950 783
rect 2950 749 2988 783
rect 2988 749 2995 783
rect 2885 657 2937 709
rect 2993 657 3045 709
rect 2885 585 2937 637
rect 2993 585 3045 637
rect 2885 412 2937 464
rect 2993 412 3045 464
rect 2885 334 2937 386
rect 2993 334 3045 386
rect 2689 23 2741 75
rect 2755 23 2807 75
<< metal2 >>
rect 3004 2405 3060 2414
rect 3004 2329 3060 2349
rect 2755 2277 2761 2329
rect 2813 2277 2825 2329
rect 2877 2325 3060 2329
rect 2877 2277 3004 2325
rect 3004 2260 3060 2269
rect 2762 1702 2814 1708
rect 2762 1636 2814 1650
tri 2731 1106 2762 1137 se
rect 2762 1123 2814 1584
rect 2762 1106 2797 1123
tri 2797 1106 2814 1123 nw
rect 2982 1635 3060 1644
rect 2982 1626 3004 1635
rect 2982 1574 2994 1626
rect 3046 1574 3060 1579
rect 2982 1560 3060 1574
rect 2982 1508 2994 1560
rect 3046 1555 3060 1560
rect 2982 1499 3004 1508
rect 2982 1490 3060 1499
rect 2731 867 2783 1106
tri 2783 1092 2797 1106 nw
tri 2964 1000 2982 1018 se
rect 2982 1004 3034 1490
tri 3034 1464 3060 1490 nw
rect 2982 1000 3009 1004
rect 2843 963 2895 1000
rect 2843 899 2895 911
rect 2843 841 2895 847
tri 2943 979 2964 1000 se
rect 2964 979 3009 1000
tri 3009 979 3034 1004 nw
rect 2943 867 2995 979
tri 2995 965 3009 979 nw
rect 2731 801 2783 815
tri 2727 105 2731 109 se
rect 2731 105 2783 749
rect 2943 801 2995 815
rect 2943 743 2995 749
rect 2879 657 2885 709
rect 2937 657 2993 709
rect 3045 657 3051 709
rect 2879 637 3051 657
rect 2879 585 2885 637
rect 2937 585 2993 637
rect 3045 585 3051 637
rect 2879 464 3051 585
rect 2879 412 2885 464
rect 2937 412 2993 464
rect 3045 412 3051 464
rect 2879 386 3051 412
rect 2879 334 2885 386
rect 2937 334 2993 386
rect 3045 334 3051 386
tri 2697 75 2727 105 se
rect 2727 75 2783 105
tri 2783 75 2813 105 sw
rect 2683 23 2689 75
rect 2741 23 2755 75
rect 2807 23 2813 75
<< via2 >>
rect 3004 2349 3060 2405
rect 3004 2269 3060 2325
rect 3004 1626 3060 1635
rect 3004 1579 3046 1626
rect 3046 1579 3060 1626
rect 3004 1508 3046 1555
rect 3046 1508 3060 1555
rect 3004 1499 3060 1508
<< metal3 >>
rect 2999 2405 3065 2410
rect 2999 2349 3004 2405
rect 3060 2349 3065 2405
rect 2999 2325 3065 2349
rect 2999 2269 3004 2325
rect 3060 2269 3065 2325
rect 2999 1635 3065 2269
rect 2999 1579 3004 1635
rect 3060 1579 3065 1635
rect 2999 1555 3065 1579
rect 2999 1499 3004 1555
rect 3060 1499 3065 1555
rect 2999 1494 3065 1499
use sky130_fd_pr__nfet_01v8__example_55959141808375  sky130_fd_pr__nfet_01v8__example_55959141808375_0
timestamp 1648127584
transform 1 0 2679 0 1 572
box -28 0 396 97
use sky130_fd_pr__nfet_01v8__example_55959141808376  sky130_fd_pr__nfet_01v8__example_55959141808376_0
timestamp 1648127584
transform 1 0 1620 0 -1 2202
box -28 0 128 471
use sky130_fd_pr__nfet_01v8__example_55959141808377  sky130_fd_pr__nfet_01v8__example_55959141808377_0
timestamp 1648127584
transform -1 0 1411 0 -1 2202
box -28 0 128 471
use sky130_fd_pr__nfet_01v8__example_55959141808381  sky130_fd_pr__nfet_01v8__example_55959141808381_0
timestamp 1648127584
transform -1 0 946 0 -1 1249
box -28 0 148 63
use sky130_fd_pr__nfet_01v8__example_55959141808384  sky130_fd_pr__nfet_01v8__example_55959141808384_0
timestamp 1648127584
transform 1 0 1002 0 -1 1249
box -28 0 148 63
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_0
timestamp 1648127584
transform 1 0 1304 0 1 648
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_1
timestamp 1648127584
transform 1 0 1304 0 1 128
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_2
timestamp 1648127584
transform 1 0 1304 0 1 388
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808386  sky130_fd_pr__nfet_01v8__example_55959141808386_3
timestamp 1648127584
transform 1 0 1304 0 1 908
box -28 0 444 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_0
timestamp 1648127584
transform 1 0 1900 0 1 2002
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_1
timestamp 1648127584
transform 1 0 1900 0 1 1222
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_2
timestamp 1648127584
transform 1 0 1900 0 1 1742
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_3
timestamp 1648127584
transform 1 0 1900 0 1 388
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_4
timestamp 1648127584
transform 1 0 1900 0 1 1482
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_5
timestamp 1648127584
transform 1 0 1900 0 1 128
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_6
timestamp 1648127584
transform 1 0 1900 0 1 648
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808387  sky130_fd_pr__nfet_01v8__example_55959141808387_7
timestamp 1648127584
transform 1 0 1900 0 1 908
box -28 0 208 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_0
timestamp 1648127584
transform 1 0 2260 0 1 908
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_1
timestamp 1648127584
transform 1 0 2260 0 1 648
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_2
timestamp 1648127584
transform 1 0 2260 0 1 1482
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_3
timestamp 1648127584
transform 1 0 2260 0 1 1222
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_4
timestamp 1648127584
transform 1 0 2260 0 1 2002
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_5
timestamp 1648127584
transform 1 0 2260 0 1 1742
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_6
timestamp 1648127584
transform 1 0 2260 0 1 128
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808388  sky130_fd_pr__nfet_01v8__example_55959141808388_7
timestamp 1648127584
transform 1 0 2260 0 1 388
box -28 0 144 97
use sky130_fd_pr__nfet_01v8__example_55959141808412  sky130_fd_pr__nfet_01v8__example_55959141808412_0
timestamp 1648127584
transform 1 0 86 0 -1 1282
box -28 0 324 63
use sky130_fd_pr__nfet_01v8__example_55959141808413  sky130_fd_pr__nfet_01v8__example_55959141808413_0
timestamp 1648127584
transform 1 0 829 0 1 1608
box -28 0 324 63
use sky130_fd_pr__nfet_01v8__example_55959141808413  sky130_fd_pr__nfet_01v8__example_55959141808413_1
timestamp 1648127584
transform 1 0 829 0 1 1884
box -28 0 324 63
use sky130_fd_pr__pfet_01v8__example_55959141808389  sky130_fd_pr__pfet_01v8__example_55959141808389_0
timestamp 1648127584
transform 1 0 2824 0 -1 1590
box -28 0 184 267
use sky130_fd_pr__pfet_01v8__example_55959141808390  sky130_fd_pr__pfet_01v8__example_55959141808390_0
timestamp 1648127584
transform 1 0 28 0 -1 455
box -28 0 128 97
use sky130_fd_pr__pfet_01v8__example_55959141808391  sky130_fd_pr__pfet_01v8__example_55959141808391_0
timestamp 1648127584
transform 1 0 28 0 -1 870
box -28 0 128 97
use sky130_fd_pr__pfet_01v8__example_55959141808414  sky130_fd_pr__pfet_01v8__example_55959141808414_0
timestamp 1648127584
transform -1 0 414 0 -1 755
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_55959141808414  sky130_fd_pr__pfet_01v8__example_55959141808414_1
timestamp 1648127584
transform -1 0 414 0 -1 386
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_55959141808415  sky130_fd_pr__pfet_01v8__example_55959141808415_0
timestamp 1648127584
transform 1 0 594 0 1 459
box -28 0 128 97
use sky130_fd_pr__pfet_01v8__example_55959141808415  sky130_fd_pr__pfet_01v8__example_55959141808415_1
timestamp 1648127584
transform 1 0 594 0 1 732
box -28 0 128 97
use sky130_fd_pr__pfet_01v8__example_55959141808415  sky130_fd_pr__pfet_01v8__example_55959141808415_2
timestamp 1648127584
transform 1 0 594 0 1 186
box -28 0 128 97
use sky130_fd_pr__tpl1__example_55959141808411  sky130_fd_pr__tpl1__example_55959141808411_0
timestamp 1648127584
transform -1 0 1161 0 1 92
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1648127584
transform 0 1 781 -1 0 1758
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1648127584
transform 0 -1 2335 -1 0 1022
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1648127584
transform 0 -1 1529 -1 0 1022
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1648127584
transform 1 0 1103 0 1 984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1648127584
transform 0 -1 815 -1 0 938
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1648127584
transform 0 1 2203 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1648127584
transform 0 1 2503 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1648127584
transform -1 0 1108 0 1 910
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1648127584
transform 0 -1 2537 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1648127584
transform 1 0 888 0 1 1718
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1648127584
transform -1 0 959 0 1 984
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1648127584
transform 0 1 2387 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1648127584
transform -1 0 600 0 1 1297
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1648127584
transform 0 -1 303 1 0 188
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1648127584
transform -1 0 380 0 1 910
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1648127584
transform -1 0 515 0 -1 1403
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1648127584
transform 0 1 1142 -1 0 1751
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1648127584
transform 1 0 888 0 1 1880
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1648127584
transform 1 0 1519 0 1 1489
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_19
timestamp 1648127584
transform 1 0 772 0 1 1489
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_20
timestamp 1648127584
transform -1 0 194 0 1 933
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_21
timestamp 1648127584
transform 0 -1 739 1 0 188
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_22
timestamp 1648127584
transform 1 0 2279 0 1 2283
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180857  sky130_fd_pr__via_l1m1__example_5595914180857_0
timestamp 1648127584
transform 0 -1 747 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180857  sky130_fd_pr__via_l1m1__example_5595914180857_1
timestamp 1648127584
transform 0 1 217 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1648127584
transform 1 0 2091 0 -1 1844
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1648127584
transform 1 0 2301 0 -1 1844
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1648127584
transform 0 -1 2236 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1648127584
transform 0 -1 2421 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1648127584
transform 0 -1 887 1 0 116
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1648127584
transform 0 1 2503 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1648127584
transform 0 -1 17 1 0 116
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1648127584
transform 0 -1 991 -1 0 1443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_0
timestamp 1648127584
transform -1 0 2043 0 -1 2090
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808264  sky130_fd_pr__via_l1m1__example_55959141808264_1
timestamp 1648127584
transform 0 1 959 -1 0 452
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_0
timestamp 1648127584
transform 0 1 665 -1 0 1849
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1648127584
transform 0 1 1002 1 0 922
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1648127584
transform 1 0 297 0 -1 503
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1648127584
transform 0 1 1923 1 0 2228
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1648127584
transform 0 1 2251 1 0 37
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1648127584
transform 0 1 2251 1 0 2228
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1648127584
transform -1 0 690 0 1 974
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1648127584
transform 0 1 1005 -1 0 2136
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1648127584
transform 0 1 822 -1 0 2136
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_6
timestamp 1648127584
transform 0 1 594 1 0 71
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_7
timestamp 1648127584
transform 0 1 51 1 0 37
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_8
timestamp 1648127584
transform -1 0 946 0 1 942
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_9
timestamp 1648127584
transform 0 1 1923 1 0 1132
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_10
timestamp 1648127584
transform 0 1 51 -1 0 983
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808272  sky130_fd_pr__via_pol1__example_55959141808272_0
timestamp 1648127584
transform 0 -1 1719 -1 0 2294
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1648127584
transform 0 1 1312 1 0 37
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808373  sky130_fd_pr__via_pol1__example_55959141808373_0
timestamp 1648127584
transform 1 0 262 0 -1 1050
box 0 0 1 1
<< labels >>
flabel locali s 642 87 682 121 3 FreeSans 300 180 0 0 SET_H_N
port 1 nsew
flabel locali s 413 1105 448 1151 7 FreeSans 300 180 0 0 OUT_H_N
port 2 nsew
flabel locali s 1074 2136 1114 2182 7 FreeSans 300 180 0 0 SET_H
port 3 nsew
flabel locali s 1496 2245 1536 2277 0 FreeSans 200 0 0 0 HLD_H_N
port 4 nsew
flabel metal1 s 3277 104 3312 306 7 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s -179 334 -144 464 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s -179 104 -144 306 3 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel metal1 s 3277 334 3312 464 7 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 3277 1253 3312 1455 7 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel metal1 s 3277 1898 3312 2246 7 FreeSans 300 0 0 0 VPWR_KA
port 7 nsew
flabel metal1 s 738 1995 773 2246 3 FreeSans 300 180 0 0 VPWR_KA
port 7 nsew
flabel metal1 s -96 1253 -56 1455 3 FreeSans 300 180 0 0 VGND
port 6 nsew
flabel comment s 870 1048 870 1048 0 FreeSans 300 0 0 0 FBK_N
flabel comment s 1065 1048 1065 1048 0 FreeSans 300 0 0 0 FBK
flabel comment s 766 836 766 836 0 FreeSans 300 180 0 0 IN_I
flabel comment s 1516 2251 1516 2251 0 FreeSans 200 180 0 0 HLD_H_N
flabel comment s 1405 1655 1405 1655 0 FreeSans 300 0 0 0 IN_I_N
flabel comment s 1512 1295 1512 1295 0 FreeSans 200 0 0 0 TO HVNATIVES
flabel comment s 1274 1338 1274 1338 0 FreeSans 300 90 0 0 FBK_N
flabel comment s 812 1318 812 1318 0 FreeSans 300 270 0 0 FBK
flabel comment s 388 727 388 727 0 FreeSans 200 0 0 0 OUT_H_N
flabel comment s 1197 1497 1197 1497 0 FreeSans 300 180 0 0 FBK
flabel comment s 2578 63 2578 63 0 FreeSans 400 0 0 0 IN_I
flabel comment s 1272 1831 1272 1831 0 FreeSans 300 270 0 0 FBK_N
<< properties >>
string GDS_END 36706652
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36675236
<< end >>
