magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 0 415 886 1116
<< pwell >>
rect 216 118 670 310
<< mvnmos >>
rect 295 144 415 284
rect 471 144 591 284
<< mvpmos >>
rect 119 750 239 950
rect 295 750 415 950
rect 471 750 591 950
rect 647 750 767 950
rect 119 482 239 682
rect 295 482 415 682
rect 471 482 591 682
rect 647 482 767 682
<< mvndiff >>
rect 242 272 295 284
rect 242 238 250 272
rect 284 238 295 272
rect 242 204 295 238
rect 242 170 250 204
rect 284 170 295 204
rect 242 144 295 170
rect 415 144 471 284
rect 591 272 644 284
rect 591 238 602 272
rect 636 238 644 272
rect 591 204 644 238
rect 591 170 602 204
rect 636 170 644 204
rect 591 144 644 170
<< mvpdiff >>
rect 66 932 119 950
rect 66 898 74 932
rect 108 898 119 932
rect 66 864 119 898
rect 66 830 74 864
rect 108 830 119 864
rect 66 796 119 830
rect 66 762 74 796
rect 108 762 119 796
rect 66 750 119 762
rect 239 932 295 950
rect 239 898 250 932
rect 284 898 295 932
rect 239 864 295 898
rect 239 830 250 864
rect 284 830 295 864
rect 239 796 295 830
rect 239 762 250 796
rect 284 762 295 796
rect 239 750 295 762
rect 415 932 471 950
rect 415 898 426 932
rect 460 898 471 932
rect 415 864 471 898
rect 415 830 426 864
rect 460 830 471 864
rect 415 796 471 830
rect 415 762 426 796
rect 460 762 471 796
rect 415 750 471 762
rect 591 932 647 950
rect 591 898 602 932
rect 636 898 647 932
rect 591 864 647 898
rect 591 830 602 864
rect 636 830 647 864
rect 591 796 647 830
rect 591 762 602 796
rect 636 762 647 796
rect 591 750 647 762
rect 767 932 820 950
rect 767 898 778 932
rect 812 898 820 932
rect 767 864 820 898
rect 767 830 778 864
rect 812 830 820 864
rect 767 796 820 830
rect 767 762 778 796
rect 812 762 820 796
rect 767 750 820 762
rect 66 670 119 682
rect 66 636 74 670
rect 108 636 119 670
rect 66 602 119 636
rect 66 568 74 602
rect 108 568 119 602
rect 66 534 119 568
rect 66 500 74 534
rect 108 500 119 534
rect 66 482 119 500
rect 239 670 295 682
rect 239 636 250 670
rect 284 636 295 670
rect 239 602 295 636
rect 239 568 250 602
rect 284 568 295 602
rect 239 534 295 568
rect 239 500 250 534
rect 284 500 295 534
rect 239 482 295 500
rect 415 670 471 682
rect 415 636 426 670
rect 460 636 471 670
rect 415 602 471 636
rect 415 568 426 602
rect 460 568 471 602
rect 415 534 471 568
rect 415 500 426 534
rect 460 500 471 534
rect 415 482 471 500
rect 591 670 647 682
rect 591 636 602 670
rect 636 636 647 670
rect 591 602 647 636
rect 591 568 602 602
rect 636 568 647 602
rect 591 534 647 568
rect 591 500 602 534
rect 636 500 647 534
rect 591 482 647 500
rect 767 670 820 682
rect 767 636 778 670
rect 812 636 820 670
rect 767 602 820 636
rect 767 568 778 602
rect 812 568 820 602
rect 767 534 820 568
rect 767 500 778 534
rect 812 500 820 534
rect 767 482 820 500
<< mvndiffc >>
rect 250 238 284 272
rect 250 170 284 204
rect 602 238 636 272
rect 602 170 636 204
<< mvpdiffc >>
rect 74 898 108 932
rect 74 830 108 864
rect 74 762 108 796
rect 250 898 284 932
rect 250 830 284 864
rect 250 762 284 796
rect 426 898 460 932
rect 426 830 460 864
rect 426 762 460 796
rect 602 898 636 932
rect 602 830 636 864
rect 602 762 636 796
rect 778 898 812 932
rect 778 830 812 864
rect 778 762 812 796
rect 74 636 108 670
rect 74 568 108 602
rect 74 500 108 534
rect 250 636 284 670
rect 250 568 284 602
rect 250 500 284 534
rect 426 636 460 670
rect 426 568 460 602
rect 426 500 460 534
rect 602 636 636 670
rect 602 568 636 602
rect 602 500 636 534
rect 778 636 812 670
rect 778 568 812 602
rect 778 500 812 534
<< poly >>
rect 119 950 239 976
rect 295 950 415 976
rect 471 950 591 976
rect 647 950 767 976
rect 119 682 239 750
rect 295 682 415 750
rect 471 682 591 750
rect 647 682 767 750
rect 119 456 239 482
rect 295 456 415 482
rect 119 365 415 456
rect 119 331 156 365
rect 190 331 241 365
rect 275 331 325 365
rect 359 331 415 365
rect 119 306 415 331
rect 295 284 415 306
rect 471 456 591 482
rect 647 456 767 482
rect 471 365 767 456
rect 471 331 515 365
rect 549 331 600 365
rect 634 331 684 365
rect 718 331 767 365
rect 471 310 767 331
rect 471 284 591 310
rect 295 118 415 144
rect 471 118 591 144
<< polycont >>
rect 156 331 190 365
rect 241 331 275 365
rect 325 331 359 365
rect 515 331 549 365
rect 600 331 634 365
rect 684 331 718 365
<< locali >>
rect 74 932 108 944
rect 74 864 108 872
rect 74 796 108 830
rect 74 670 108 762
rect 74 602 108 636
rect 74 534 108 568
rect 74 484 108 500
rect 250 932 284 948
rect 250 864 284 898
rect 250 796 284 830
rect 250 670 284 762
rect 250 602 284 636
rect 250 534 284 568
rect 250 440 284 500
rect 426 932 460 944
rect 426 864 460 872
rect 426 796 460 830
rect 426 670 460 762
rect 426 602 460 636
rect 426 534 460 568
rect 426 475 460 500
rect 602 932 636 978
rect 602 864 636 898
rect 602 796 636 830
rect 602 670 636 762
rect 602 602 636 636
rect 602 534 636 568
rect 602 440 636 500
rect 778 932 812 944
rect 778 864 812 872
rect 778 796 812 830
rect 778 670 812 762
rect 778 602 812 636
rect 778 534 812 568
rect 778 484 812 500
rect 250 410 636 440
rect 250 406 459 410
rect 134 365 378 372
rect 134 331 156 365
rect 190 331 241 365
rect 275 331 325 365
rect 359 331 378 365
rect 134 323 378 331
rect 413 288 459 406
rect 493 365 737 372
rect 493 331 515 365
rect 549 331 600 365
rect 634 331 684 365
rect 718 331 737 365
rect 493 323 737 331
rect 250 272 284 288
rect 250 227 284 238
rect 413 272 636 288
rect 413 238 602 272
rect 413 225 636 238
rect 250 155 284 170
rect 602 204 636 225
rect 602 154 636 170
<< viali >>
rect 74 944 108 978
rect 74 898 108 906
rect 74 872 108 898
rect 426 944 460 978
rect 426 898 460 906
rect 426 872 460 898
rect 778 944 812 978
rect 778 898 812 906
rect 778 872 812 898
rect 250 204 284 227
rect 250 193 284 204
rect 250 121 284 155
<< metal1 >>
rect 25 978 820 1062
rect 25 944 74 978
rect 108 944 426 978
rect 460 944 778 978
rect 812 944 820 978
rect 25 906 820 944
rect 25 872 74 906
rect 108 872 426 906
rect 460 872 778 906
rect 812 872 820 906
rect 25 859 820 872
rect 25 227 820 239
rect 25 193 250 227
rect 284 193 820 227
rect 25 155 820 193
rect 25 121 250 155
rect 284 121 820 155
rect 25 24 820 121
use sky130_fd_pr__nfet_01v8__example_559591418087  sky130_fd_pr__nfet_01v8__example_559591418087_0
timestamp 1648127584
transform 1 0 471 0 -1 284
box -25 0 148 70
use sky130_fd_pr__nfet_01v8__example_559591418089  sky130_fd_pr__nfet_01v8__example_559591418089_0
timestamp 1648127584
transform 1 0 295 0 -1 284
box -28 0 145 70
use sky130_fd_pr__pfet_01v8__example_55959141808441  sky130_fd_pr__pfet_01v8__example_55959141808441_0
timestamp 1648127584
transform 1 0 119 0 1 750
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808441  sky130_fd_pr__pfet_01v8__example_55959141808441_1
timestamp 1648127584
transform 1 0 471 0 1 750
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808441  sky130_fd_pr__pfet_01v8__example_55959141808441_2
timestamp 1648127584
transform 1 0 119 0 -1 682
box -28 0 324 97
use sky130_fd_pr__pfet_01v8__example_55959141808441  sky130_fd_pr__pfet_01v8__example_55959141808441_3
timestamp 1648127584
transform 1 0 471 0 -1 682
box -28 0 324 97
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1648127584
transform 0 -1 812 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1648127584
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1648127584
transform 0 -1 460 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1648127584
transform 0 -1 284 -1 0 227
box 0 0 1 1
<< labels >>
flabel metal1 s 200 24 283 238 0 FreeSans 320 0 0 0 VGND
port 1 nsew
flabel metal1 s 737 859 820 1062 0 FreeSans 320 0 0 0 VPWR
port 2 nsew
flabel locali s 297 331 348 372 0 FreeSans 400 0 0 0 IN0
port 3 nsew
<< properties >>
string GDS_END 35747260
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35743836
<< end >>
