magic
tech sky130A
magscale 1 2
timestamp 1652832150
<< nwell >>
rect -396 700 772 1034
rect 258 -422 630 -22
<< poly >>
rect 194 218 224 220
rect 194 188 328 218
rect 298 20 328 188
rect 24 -10 506 20
rect 24 -168 54 -10
rect 474 -92 506 -10
rect 24 -198 110 -168
rect 80 -272 110 -198
<< locali >>
rect -459 970 -336 1004
rect -80 998 68 1003
rect 180 1002 458 1004
rect 346 998 460 1002
rect -459 -65 -425 970
rect -109 969 78 998
rect 342 969 487 998
rect 256 690 476 692
rect 224 658 544 690
rect -356 425 -330 458
rect -356 214 -322 425
rect -100 122 -66 460
rect 240 240 622 280
rect -100 118 0 122
rect -100 88 10 118
rect 442 80 488 82
rect 270 76 442 78
rect 10 44 46 62
rect 242 46 442 76
rect 484 46 488 80
rect 242 44 488 46
rect 442 38 488 44
rect 588 -118 622 240
rect -100 -162 106 -118
rect 306 -162 494 -118
rect 546 -158 622 -118
rect -78 -324 -64 -294
rect -74 -326 -64 -324
rect 636 -350 726 -348
rect 636 -362 768 -350
rect 488 -368 554 -366
rect 636 -368 792 -362
rect 488 -372 792 -368
rect 530 -382 792 -372
rect 530 -402 674 -382
rect 726 -388 792 -382
rect 222 -484 502 -450
rect -332 -526 -48 -494
rect -378 -530 128 -526
rect -378 -554 -318 -530
rect -84 -562 128 -530
rect 454 -572 502 -484
rect 454 -606 460 -572
rect 498 -606 502 -572
rect 454 -618 502 -606
rect 575 -629 719 -587
rect 575 -936 617 -629
rect 214 -978 617 -936
<< viali >>
rect -322 666 -286 700
rect -150 662 -112 696
rect 664 664 700 698
rect -240 544 -204 582
rect 578 540 614 576
rect -356 180 -322 214
rect 442 46 484 80
rect -456 -388 -420 -352
rect 822 -490 856 -456
rect 460 -606 498 -572
<< metal1 >>
rect -566 938 -200 1034
rect -116 938 520 1034
rect 724 938 976 1034
rect 102 922 146 938
rect -336 746 30 778
rect -336 708 -308 746
rect -336 700 -270 708
rect -336 666 -322 700
rect -286 666 -270 700
rect -336 654 -270 666
rect -164 704 -96 710
rect -164 652 -154 704
rect -102 652 -96 704
rect -164 646 -96 652
rect 652 706 716 712
rect 652 654 658 706
rect 710 654 716 706
rect 652 648 716 654
rect -254 592 -186 598
rect -254 540 -246 592
rect -194 540 -186 592
rect -254 530 -186 540
rect 564 590 628 596
rect 564 538 570 590
rect 622 538 628 590
rect 564 532 628 538
rect -374 358 -310 364
rect -374 324 -368 358
rect -316 324 -310 358
rect -198 358 -134 364
rect -198 324 -192 358
rect -316 304 -192 324
rect -140 304 -134 358
rect -368 296 -134 304
rect -218 244 -14 258
rect -218 230 36 244
rect -374 224 -308 230
rect -374 172 -366 224
rect -314 172 -308 224
rect -374 166 -308 172
rect -218 -120 -190 230
rect 368 -10 402 232
rect 430 90 458 422
rect 430 80 498 90
rect 430 46 442 80
rect 484 46 498 80
rect 430 32 498 46
rect -158 -38 402 -10
rect -158 -84 -92 -38
rect -218 -122 -146 -120
rect -218 -124 -190 -122
rect -218 -148 -192 -124
rect -102 -148 -36 -142
rect -102 -200 -96 -148
rect -44 -200 -36 -148
rect -102 -208 -36 -200
rect 368 -212 402 -38
rect 488 -86 554 -30
rect 446 -128 512 -122
rect 446 -180 454 -128
rect 506 -180 512 -128
rect 446 -186 512 -180
rect -524 -334 -450 -326
rect -524 -386 -506 -334
rect -454 -342 -450 -334
rect -454 -352 -408 -342
rect -524 -388 -456 -386
rect -420 -388 -408 -352
rect -524 -398 -408 -388
rect -158 -416 -92 -358
rect 488 -412 554 -356
rect 810 -456 868 -442
rect 810 -476 822 -456
rect 386 -490 822 -476
rect 856 -490 868 -456
rect 386 -510 868 -490
rect -36 -542 28 -536
rect -36 -596 -30 -542
rect 22 -596 28 -542
rect -36 -602 28 -596
rect 446 -560 522 -554
rect 446 -612 454 -560
rect 506 -612 522 -560
rect 446 -618 522 -612
rect -296 -654 -89 -620
rect -123 -930 -89 -654
rect -566 -1012 976 -930
<< via1 >>
rect -154 696 -102 704
rect -154 662 -150 696
rect -150 662 -112 696
rect -112 662 -102 696
rect -154 652 -102 662
rect 658 698 710 706
rect 658 664 664 698
rect 664 664 700 698
rect 700 664 710 698
rect 658 654 710 664
rect -246 582 -194 592
rect -246 544 -240 582
rect -240 544 -204 582
rect -204 544 -194 582
rect -246 540 -194 544
rect 570 576 622 590
rect 570 540 578 576
rect 578 540 614 576
rect 614 540 622 576
rect 570 538 622 540
rect -368 304 -316 358
rect -192 304 -140 358
rect -366 214 -314 224
rect -366 180 -356 214
rect -356 180 -322 214
rect -322 180 -314 214
rect -366 172 -314 180
rect -342 -86 -290 -34
rect 4 52 64 112
rect -96 -200 -44 -148
rect 692 -94 744 -38
rect 454 -180 506 -128
rect -506 -352 -454 -334
rect -506 -386 -456 -352
rect -456 -386 -454 -352
rect -414 -640 -356 -576
rect -30 -596 22 -542
rect 454 -572 506 -560
rect 454 -606 460 -572
rect 460 -606 498 -572
rect 498 -606 506 -572
rect 454 -612 506 -606
<< metal2 >>
rect -484 816 866 844
rect -124 710 -96 816
rect -164 704 -96 710
rect -164 652 -154 704
rect -102 652 -96 704
rect 650 712 678 816
rect 650 706 716 712
rect 650 692 658 706
rect -164 646 -96 652
rect 652 654 658 692
rect 710 654 716 706
rect 652 648 716 654
rect -254 592 -186 598
rect -254 540 -246 592
rect -194 540 -186 592
rect 564 590 628 596
rect 564 560 570 590
rect -254 530 -186 540
rect 354 538 570 560
rect 622 538 628 590
rect 354 532 628 538
rect -374 358 -310 364
rect -374 326 -368 358
rect -566 304 -368 326
rect -316 304 -310 358
rect -566 298 -310 304
rect -566 296 -368 298
rect -566 290 -374 296
rect -374 224 -308 230
rect -374 172 -366 224
rect -314 172 -308 224
rect -374 166 -308 172
rect -374 44 -346 166
rect -414 16 -346 44
rect -524 -334 -450 -326
rect -524 -386 -506 -334
rect -454 -386 -450 -334
rect -524 -398 -450 -386
rect -524 -1012 -496 -398
rect -414 -568 -386 16
rect -352 -34 -290 -28
rect -352 -86 -342 -34
rect -254 -42 -226 530
rect 136 462 168 504
rect -198 358 -134 364
rect -198 304 -192 358
rect -140 324 -134 358
rect -140 304 180 324
rect -198 296 180 304
rect -2 112 70 120
rect -2 52 4 112
rect 64 52 70 112
rect -2 44 70 52
rect 34 42 70 44
rect -254 -70 34 -42
rect -352 -92 -290 -86
rect -318 -138 -290 -92
rect -318 -142 -74 -138
rect -318 -148 -36 -142
rect -318 -166 -96 -148
rect -102 -200 -96 -166
rect -44 -200 -36 -148
rect -102 -208 -36 -200
rect 6 -536 34 -70
rect -36 -542 34 -536
rect -414 -576 -350 -568
rect -356 -640 -350 -576
rect -36 -596 -30 -542
rect 22 -596 34 -542
rect 138 -572 166 -536
rect -36 -602 34 -596
rect 354 -586 382 532
rect 786 290 976 326
rect 686 -38 750 -32
rect 686 -94 692 -38
rect 744 -94 750 -38
rect 686 -100 750 -94
rect 446 -128 512 -122
rect 446 -180 454 -128
rect 506 -158 512 -128
rect 686 -158 714 -100
rect 506 -180 714 -158
rect 446 -186 714 -180
rect 446 -560 522 -554
rect 446 -586 454 -560
rect 354 -612 454 -586
rect 506 -612 522 -560
rect 354 -614 522 -612
rect 446 -618 522 -614
rect -414 -650 -350 -640
rect 786 -776 814 290
rect 162 -804 814 -776
use sky130_fd_pr__pfet_01v8_hvt_UUWA33  1
timestamp 1652659832
transform 1 0 -125 0 1 -222
box -109 -200 109 200
use sky130_fd_pr__pfet_01v8_hvt_UUWA33  2
timestamp 1652659832
transform 1 0 521 0 1 -222
box -109 -200 109 200
use demux  demux_0
timestamp 1652676461
transform 1 0 36 0 1 156
box -54 -136 366 878
use mux  mux_0
timestamp 1652660405
transform 1 0 34 0 1 -900
box -54 -136 366 878
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 662 0 1 -604
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1650294714
transform 1 0 -528 0 1 -606
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 -356 0 1 442
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1650294714
transform 1 0 458 0 1 442
box -38 -48 314 592
<< labels >>
flabel metal2 136 462 168 504 1 FreeSans 160 0 0 0 IN
port 1 n
flabel viali -452 -386 -420 -354 1 FreeSans 160 0 0 0 C
port 2 n
flabel metal2 -150 660 -104 692 1 FreeSans 160 0 0 0 RESET
port 3 n
flabel metal1 102 922 146 966 1 FreeSans 160 0 0 0 VDD
port 5 n
flabel metal1 8 -998 48 -960 1 FreeSans 160 0 0 0 VSS
port 4 n
flabel metal2 138 -572 166 -536 1 FreeSans 160 0 0 0 OUT
port 6 n
<< end >>
