magic
tech sky130B
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__hvdftpl1s__example_55959141808646  sky130_fd_pr__hvdftpl1s__example_55959141808646_0
timestamp 1648127584
transform -1 0 -77 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 145 500 145 500 0 FreeSans 300 0 0 0 D
flabel comment s -139 477 -139 477 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 3742796
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3741938
<< end >>
