.subckt BR128 VDD VSS OUT
+ C[127] C[126] C[125] C[124] C[123] C[122] C[121] C[120] C[119] C[118] C[117] C[116] C[115] C[114] C[113] C[112] C[111] C[110] C[109] C[108] C[107] C[106] C[105] C[104] C[103] C[102] C[101] C[100] C[99] C[98] C[97] C[96] C[95] C[94] C[93] C[92] C[91] C[90] C[89] C[88] C[87] C[86] C[85] C[84] C[83] C[82] C[81] C[80] C[79] C[78] C[77] C[76] C[75] C[74] C[73] C[72] C[71] C[70] C[69] C[68] C[67] C[66] C[65] C[64] C[63] C[62] C[61] C[60] C[59] C[58] C[57] C[56] C[55] C[54] C[53] C[52] C[51] C[50] C[49] C[48] C[47] C[46] C[45] C[44] C[43] C[42] C[41] C[40] C[39] C[38] C[37] C[36] C[35] C[34] C[33] C[32] C[31] C[30] C[29] C[28] C[27] C[26] C[25] C[24] C[23] C[22] C[21] C[20] C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12] C[11] C[10] C[9] C[8] C[7] C[6] C[5] C[4] C[3] C[2] C[1] C[0] RESET
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin
*+ C[127],C[126],C[125],C[124],C[123],C[122],C[121],C[120],C[119],C[118],C[117],C[116],C[115],C[114],C[113],C[112],C[111],C[110],C[109],C[108],C[107],C[106],C[105],C[104],C[103],C[102],C[101],C[100],C[99],C[98],C[97],C[96],C[95],C[94],C[93],C[92],C[91],C[90],C[89],C[88],C[87],C[86],C[85],C[84],C[83],C[82],C[81],C[80],C[79],C[78],C[77],C[76],C[75],C[74],C[73],C[72],C[71],C[70],C[69],C[68],C[67],C[66],C[65],C[64],C[63],C[62],C[61],C[60],C[59],C[58],C[57],C[56],C[55],C[54],C[53],C[52],C[51],C[50],C[49],C[48],C[47],C[46],C[45],C[44],C[43],C[42],C[41],C[40],C[39],C[38],C[37],C[36],C[35],C[34],C[33],C[32],C[31],C[30],C[29],C[28],C[27],C[26],C[25],C[24],C[23],C[22],C[21],C[20],C[19],C[18],C[17],C[16],C[15],C[14],C[13],C[12],C[11],C[10],C[9],C[8],C[7],C[6],C[5],C[4],C[3],C[2],C[1],C[0]
*.ipin RESET
x47 net1 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x48 net1 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x4 net1 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x5 net1 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x6 net1 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x7 net1 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x8 net1 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x10 net1 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x11 net2 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_16
x12 net2 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_16
x13 net3 VSS VSS VDD VDD r6 sky130_fd_sc_hd__inv_16
x14 net3 VSS VSS VDD VDD r5 sky130_fd_sc_hd__inv_16
x15 net3 VSS VSS VDD VDD r5 sky130_fd_sc_hd__inv_16
x16 net3 VSS VSS VDD VDD r6 sky130_fd_sc_hd__inv_16
x17 net3 VSS VSS VDD VDD r8 sky130_fd_sc_hd__inv_16
x18 net3 VSS VSS VDD VDD r7 sky130_fd_sc_hd__inv_16
x19 net3 VSS VSS VDD VDD r7 sky130_fd_sc_hd__inv_16
x20 net3 VSS VSS VDD VDD r8 sky130_fd_sc_hd__inv_16
x21 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_16
x22 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_16
x23 net21 VSS VSS VDD VDD net2 sky130_fd_sc_hd__inv_16
x3[7] r1 VDD VSS out[8] out[7] net4[7] C[7] singlestage
x3[6] r1 VDD VSS out[7] out[6] net4[6] C[6] singlestage
x3[5] r1 VDD VSS out[6] out[5] net4[5] C[5] singlestage
x3[4] r1 VDD VSS out[5] out[4] net4[4] C[4] singlestage
x3[3] r1 VDD VSS out[4] out[3] net4[3] C[3] singlestage
x3[2] r1 VDD VSS out[3] out[2] net4[2] C[2] singlestage
x3[1] r1 VDD VSS out[2] out[1] net4[1] C[1] singlestage
x3[0] r1 VDD VSS out[1] out[0] net4[0] C[0] singlestage
x1[15] r2 VDD VSS out[16] out[15] net5[7] C[15] singlestage
x1[14] r2 VDD VSS out[15] out[14] net5[6] C[14] singlestage
x1[13] r2 VDD VSS out[14] out[13] net5[5] C[13] singlestage
x1[12] r2 VDD VSS out[13] out[12] net5[4] C[12] singlestage
x1[11] r2 VDD VSS out[12] out[11] net5[3] C[11] singlestage
x1[10] r2 VDD VSS out[11] out[10] net5[2] C[10] singlestage
x1[9] r2 VDD VSS out[10] out[9] net5[1] C[9] singlestage
x1[8] r2 VDD VSS out[9] out[8] net5[0] C[8] singlestage
x2[23] r5 VDD VSS out[24] out[23] net6[7] C[23] singlestage
x2[22] r5 VDD VSS out[23] out[22] net6[6] C[22] singlestage
x2[21] r5 VDD VSS out[22] out[21] net6[5] C[21] singlestage
x2[20] r5 VDD VSS out[21] out[20] net6[4] C[20] singlestage
x2[19] r5 VDD VSS out[20] out[19] net6[3] C[19] singlestage
x2[18] r5 VDD VSS out[19] out[18] net6[2] C[18] singlestage
x2[17] r5 VDD VSS out[18] out[17] net6[1] C[17] singlestage
x2[16] r5 VDD VSS out[17] out[16] net6[0] C[16] singlestage
x4[31] r6 VDD VSS out[32] out[31] net7[7] C[31] singlestage
x4[30] r6 VDD VSS out[31] out[30] net7[6] C[30] singlestage
x4[29] r6 VDD VSS out[30] out[29] net7[5] C[29] singlestage
x4[28] r6 VDD VSS out[29] out[28] net7[4] C[28] singlestage
x4[27] r6 VDD VSS out[28] out[27] net7[3] C[27] singlestage
x4[26] r6 VDD VSS out[27] out[26] net7[2] C[26] singlestage
x4[25] r6 VDD VSS out[26] out[25] net7[1] C[25] singlestage
x4[24] r6 VDD VSS out[25] out[24] net7[0] C[24] singlestage
x5[63] r13 VDD VSS out[64] out[63] net8[7] C[63] singlestage
x5[62] r13 VDD VSS out[63] out[62] net8[6] C[62] singlestage
x5[61] r13 VDD VSS out[62] out[61] net8[5] C[61] singlestage
x5[60] r13 VDD VSS out[61] out[60] net8[4] C[60] singlestage
x5[59] r13 VDD VSS out[60] out[59] net8[3] C[59] singlestage
x5[58] r13 VDD VSS out[59] out[58] net8[2] C[58] singlestage
x5[57] r13 VDD VSS out[58] out[57] net8[1] C[57] singlestage
x5[56] r13 VDD VSS out[57] out[56] net8[0] C[56] singlestage
x6[55] r14 VDD VSS out[56] out[55] net9[7] C[55] singlestage
x6[54] r14 VDD VSS out[55] out[54] net9[6] C[54] singlestage
x6[53] r14 VDD VSS out[54] out[53] net9[5] C[53] singlestage
x6[52] r14 VDD VSS out[53] out[52] net9[4] C[52] singlestage
x6[51] r14 VDD VSS out[52] out[51] net9[3] C[51] singlestage
x6[50] r14 VDD VSS out[51] out[50] net9[2] C[50] singlestage
x6[49] r14 VDD VSS out[50] out[49] net9[1] C[49] singlestage
x6[48] r14 VDD VSS out[49] out[48] net9[0] C[48] singlestage
x7[47] r9 VDD VSS out[48] out[47] net10[7] C[47] singlestage
x7[46] r9 VDD VSS out[47] out[46] net10[6] C[46] singlestage
x7[45] r9 VDD VSS out[46] out[45] net10[5] C[45] singlestage
x7[44] r9 VDD VSS out[45] out[44] net10[4] C[44] singlestage
x7[43] r9 VDD VSS out[44] out[43] net10[3] C[43] singlestage
x7[42] r9 VDD VSS out[43] out[42] net10[2] C[42] singlestage
x7[41] r9 VDD VSS out[42] out[41] net10[1] C[41] singlestage
x7[40] r9 VDD VSS out[41] out[40] net10[0] C[40] singlestage
x8[39] r10 VDD VSS out[40] out[39] net11[7] C[39] singlestage
x8[38] r10 VDD VSS out[39] out[38] net11[6] C[38] singlestage
x8[37] r10 VDD VSS out[38] out[37] net11[5] C[37] singlestage
x8[36] r10 VDD VSS out[37] out[36] net11[4] C[36] singlestage
x8[35] r10 VDD VSS out[36] out[35] net11[3] C[35] singlestage
x8[34] r10 VDD VSS out[35] out[34] net11[2] C[34] singlestage
x8[33] r10 VDD VSS out[34] out[33] net11[1] C[33] singlestage
x8[32] r10 VDD VSS out[33] out[32] net11[0] C[32] singlestage
x1 net21 VSS VSS VDD VDD net2 sky130_fd_sc_hd__inv_16
x2 net12 VSS VSS VDD VDD r10 sky130_fd_sc_hd__inv_16
x3 net12 VSS VSS VDD VDD r9 sky130_fd_sc_hd__inv_16
x9 net12 VSS VSS VDD VDD r9 sky130_fd_sc_hd__inv_16
x24 net12 VSS VSS VDD VDD r10 sky130_fd_sc_hd__inv_16
x25 net12 VSS VSS VDD VDD r12 sky130_fd_sc_hd__inv_16
x26 net12 VSS VSS VDD VDD r11 sky130_fd_sc_hd__inv_16
x27 net12 VSS VSS VDD VDD r11 sky130_fd_sc_hd__inv_16
x28 net12 VSS VSS VDD VDD r12 sky130_fd_sc_hd__inv_16
x29 net2 VSS VSS VDD VDD net12 sky130_fd_sc_hd__inv_16
x30 net2 VSS VSS VDD VDD net12 sky130_fd_sc_hd__inv_16
x31 net13 VSS VSS VDD VDD r14 sky130_fd_sc_hd__inv_16
x32 net13 VSS VSS VDD VDD r13 sky130_fd_sc_hd__inv_16
x33 net13 VSS VSS VDD VDD r13 sky130_fd_sc_hd__inv_16
x34 net13 VSS VSS VDD VDD r14 sky130_fd_sc_hd__inv_16
x35 net13 VSS VSS VDD VDD r16 sky130_fd_sc_hd__inv_16
x36 net13 VSS VSS VDD VDD r15 sky130_fd_sc_hd__inv_16
x37 net13 VSS VSS VDD VDD r15 sky130_fd_sc_hd__inv_16
x38 net13 VSS VSS VDD VDD r16 sky130_fd_sc_hd__inv_16
x39 net2 VSS VSS VDD VDD net13 sky130_fd_sc_hd__inv_16
x40 net2 VSS VSS VDD VDD net13 sky130_fd_sc_hd__inv_16
x6[71] r16 VDD VSS out[72] out[71] net14[7] C[71] singlestage
x6[70] r16 VDD VSS out[71] out[70] net14[6] C[70] singlestage
x6[69] r16 VDD VSS out[70] out[69] net14[5] C[69] singlestage
x6[68] r16 VDD VSS out[69] out[68] net14[4] C[68] singlestage
x6[67] r16 VDD VSS out[68] out[67] net14[3] C[67] singlestage
x6[66] r16 VDD VSS out[67] out[66] net14[2] C[66] singlestage
x6[65] r16 VDD VSS out[66] out[65] net14[1] C[65] singlestage
x6[64] r16 VDD VSS out[65] out[64] net14[0] C[64] singlestage
x7[79] r15 VDD VSS out[80] out[79] net15[7] C[79] singlestage
x7[78] r15 VDD VSS out[79] out[78] net15[6] C[78] singlestage
x7[77] r15 VDD VSS out[78] out[77] net15[5] C[77] singlestage
x7[76] r15 VDD VSS out[77] out[76] net15[4] C[76] singlestage
x7[75] r15 VDD VSS out[76] out[75] net15[3] C[75] singlestage
x7[74] r15 VDD VSS out[75] out[74] net15[2] C[74] singlestage
x7[73] r15 VDD VSS out[74] out[73] net15[1] C[73] singlestage
x7[72] r15 VDD VSS out[73] out[72] net15[0] C[72] singlestage
x8[87] r12 VDD VSS out[88] out[87] net16[7] C[87] singlestage
x8[86] r12 VDD VSS out[87] out[86] net16[6] C[86] singlestage
x8[85] r12 VDD VSS out[86] out[85] net16[5] C[85] singlestage
x8[84] r12 VDD VSS out[85] out[84] net16[4] C[84] singlestage
x8[83] r12 VDD VSS out[84] out[83] net16[3] C[83] singlestage
x8[82] r12 VDD VSS out[83] out[82] net16[2] C[82] singlestage
x8[81] r12 VDD VSS out[82] out[81] net16[1] C[81] singlestage
x8[80] r12 VDD VSS out[81] out[80] net16[0] C[80] singlestage
x9[95] r11 VDD VSS out[96] out[95] net17[7] C[95] singlestage
x9[94] r11 VDD VSS out[95] out[94] net17[6] C[94] singlestage
x9[93] r11 VDD VSS out[94] out[93] net17[5] C[93] singlestage
x9[92] r11 VDD VSS out[93] out[92] net17[4] C[92] singlestage
x9[91] r11 VDD VSS out[92] out[91] net17[3] C[91] singlestage
x9[90] r11 VDD VSS out[91] out[90] net17[2] C[90] singlestage
x9[89] r11 VDD VSS out[90] out[89] net17[1] C[89] singlestage
x9[88] r11 VDD VSS out[89] out[88] net17[0] C[88] singlestage
x1[127] r3 VDD VSS out[0] out[127] OUT C[127] singlestage
x1[126] r3 VDD VSS out[127] out[126] buf_out[6] C[126] singlestage
x1[125] r3 VDD VSS out[126] out[125] buf_out[5] C[125] singlestage
x1[124] r3 VDD VSS out[125] out[124] buf_out[4] C[124] singlestage
x1[123] r3 VDD VSS out[124] out[123] buf_out[3] C[123] singlestage
x1[122] r3 VDD VSS out[123] out[122] buf_out[2] C[122] singlestage
x1[121] r3 VDD VSS out[122] out[121] buf_out[1] C[121] singlestage
x1[120] r3 VDD VSS out[121] out[120] buf_out[0] C[120] singlestage
x2[119] r4 VDD VSS out[120] out[119] net18[7] C[119] singlestage
x2[118] r4 VDD VSS out[119] out[118] net18[6] C[118] singlestage
x2[117] r4 VDD VSS out[118] out[117] net18[5] C[117] singlestage
x2[116] r4 VDD VSS out[117] out[116] net18[4] C[116] singlestage
x2[115] r4 VDD VSS out[116] out[115] net18[3] C[115] singlestage
x2[114] r4 VDD VSS out[115] out[114] net18[2] C[114] singlestage
x2[113] r4 VDD VSS out[114] out[113] net18[1] C[113] singlestage
x2[112] r4 VDD VSS out[113] out[112] net18[0] C[112] singlestage
x3[111] r8 VDD VSS out[112] out[111] net19[7] C[111] singlestage
x3[110] r8 VDD VSS out[111] out[110] net19[6] C[110] singlestage
x3[109] r8 VDD VSS out[110] out[109] net19[5] C[109] singlestage
x3[108] r8 VDD VSS out[109] out[108] net19[4] C[108] singlestage
x3[107] r8 VDD VSS out[108] out[107] net19[3] C[107] singlestage
x3[106] r8 VDD VSS out[107] out[106] net19[2] C[106] singlestage
x3[105] r8 VDD VSS out[106] out[105] net19[1] C[105] singlestage
x3[104] r8 VDD VSS out[105] out[104] net19[0] C[104] singlestage
x4[103] r7 VDD VSS out[104] out[103] net20[7] C[103] singlestage
x4[102] r7 VDD VSS out[103] out[102] net20[6] C[102] singlestage
x4[101] r7 VDD VSS out[102] out[101] net20[5] C[101] singlestage
x4[100] r7 VDD VSS out[101] out[100] net20[4] C[100] singlestage
x4[99] r7 VDD VSS out[100] out[99] net20[3] C[99] singlestage
x4[98] r7 VDD VSS out[99] out[98] net20[2] C[98] singlestage
x4[97] r7 VDD VSS out[98] out[97] net20[1] C[97] singlestage
x4[96] r7 VDD VSS out[97] out[96] net20[0] C[96] singlestage
x41 RESET VSS VSS VDD VDD net22 sky130_fd_sc_hd__buf_2
x42 net22 VSS VSS VDD VDD net21 sky130_fd_sc_hd__inv_8
.ends

* expanding   symbol:  singlestage.sym # of pins=7
* sym_path: /home/users/lsammaro/open-puf/design/singlestage.sym
* sch_path: /home/users/lsammaro/open-puf/design/singlestage.sch
.subckt singlestage  RESET VDD VSS OUT IN buf_out C
*.ipin IN
*.ipin C
*.ipin RESET
*.iopin VSS
*.iopin VDD
*.opin OUT
*.opin buf_out
x1 RESET net1 VSS VSS VDD VDD net3 sky130_fd_sc_hd__nor2_1
x2 RESET net2 VSS VSS VDD VDD net4 sky130_fd_sc_hd__nor2_1
x3 net6 VSS net1 VDD IN net5 net2 demux2-1
x4 net6 VSS net3 VDD OUT net5 net4 mux2-1
x5 net5 VSS VSS VDD VDD net6 sky130_fd_sc_hd__inv_1
XM1 net1 net6 VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net2 net5 VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x6 C VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_1
x7 OUT VSS VSS VDD VDD buf_out sky130_fd_sc_hd__buf_1
.ends


* expanding   symbol:  demux2-1.sym # of pins=7
* sym_path: /home/users/lsammaro/open-puf/design/demux2-1.sym
* sch_path: /home/users/lsammaro/open-puf/design/demux2-1.sch
.subckt demux2-1  S VSS OUT1 VDD IN Sbar OUT2
*.ipin Sbar
*.ipin S
*.iopin VSS
*.iopin VDD
*.opin OUT1
*.opin OUT2
*.ipin IN
XM2 IN S OUT1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 IN Sbar OUT2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 IN Sbar OUT1 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 IN S OUT2 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  mux2-1.sym # of pins=7
* sym_path: /home/users/lsammaro/open-puf/design/mux2-1.sym
* sch_path: /home/users/lsammaro/open-puf/design/mux2-1.sch
.subckt mux2-1  S VSS IN1 VDD OUT Sbar IN2
*.ipin IN1
*.ipin IN2
*.ipin Sbar
*.ipin S
*.opin OUT
*.iopin VSS
*.iopin VDD
XM2 IN1 S OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 IN2 Sbar OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 IN1 Sbar OUT VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 IN2 S OUT VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='1 * W/nf * 0.29' as='3/2 * W/nf * 0.29'
+ pd='2*1 * (W/nf + 0.29)' ps='2*3/2 * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes

.subckt BR32 VDD VSS RESET OUT
+ C[31] C[30] C[29] C[28] C[27] C[26] C[25] C[24] C[23] C[22] C[21] C[20] C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12] C[11] C[10] C[9] C[8] C[7] C[6] C[5] C[4] C[3] C[2] C[1] C[0]
*.iopin VDD
*.iopin VSS
*.ipin RESET
*.opin OUT
*.ipin
*+ C[31],C[30],C[29],C[28],C[27],C[26],C[25],C[24],C[23],C[22],C[21],C[20],C[19],C[18],C[17],C[16],C[15],C[14],C[13],C[12],C[11],C[10],C[9],C[8],C[7],C[6],C[5],C[4],C[3],C[2],C[1],C[0]
x47 net3 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x48 net3 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x50 net4 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x51 net4 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x9 net3 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x10 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_16
x11 net2 VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_16
x12 net3 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x29 net4 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x30 net4 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x31 RESET VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_2
x32 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__inv_8
x41[6] r1 VDD VSS int_out[6] int_out[5] buf_out[6] C[6] singlestage
x41[5] r1 VDD VSS int_out[5] int_out[4] buf_out[5] C[5] singlestage
x41[4] r1 VDD VSS int_out[4] int_out[3] buf_out[4] C[4] singlestage
x41[3] r1 VDD VSS int_out[3] int_out[2] buf_out[3] C[3] singlestage
x41[2] r1 VDD VSS int_out[2] int_out[1] buf_out[2] C[2] singlestage
x41[1] r1 VDD VSS int_out[1] int_out[0] buf_out[1] C[1] singlestage
x41[0] r1 VDD VSS int_out[0] int_out[31] buf_out[0] C[0] singlestage
x1[7] r4 VDD VSS int_out[14] int_out[13] buf_out[14] C[14] singlestage
x1[6] r4 VDD VSS int_out[13] int_out[12] buf_out[13] C[13] singlestage
x1[5] r4 VDD VSS int_out[12] int_out[11] buf_out[12] C[12] singlestage
x1[4] r4 VDD VSS int_out[11] int_out[10] buf_out[11] C[11] singlestage
x1[3] r4 VDD VSS int_out[10] int_out[9] buf_out[10] C[10] singlestage
x1[2] r4 VDD VSS int_out[9] int_out[8] buf_out[9] C[9] singlestage
x1[1] r4 VDD VSS int_out[8] int_out[7] buf_out[8] C[8] singlestage
x1[0] r4 VDD VSS int_out[7] int_out[6] buf_out[7] C[7] singlestage
x2[8] r3 VDD VSS int_out[23] int_out[22] buf_out[23] C[23] singlestage
x2[7] r3 VDD VSS int_out[22] int_out[21] buf_out[22] C[22] singlestage
x2[6] r3 VDD VSS int_out[21] int_out[20] buf_out[21] C[21] singlestage
x2[5] r3 VDD VSS int_out[20] int_out[19] buf_out[20] C[20] singlestage
x2[4] r3 VDD VSS int_out[19] int_out[18] buf_out[19] C[19] singlestage
x2[3] r3 VDD VSS int_out[18] int_out[17] buf_out[18] C[18] singlestage
x2[2] r3 VDD VSS int_out[17] int_out[16] buf_out[17] C[17] singlestage
x2[1] r3 VDD VSS int_out[16] int_out[15] buf_out[16] C[16] singlestage
x2[0] r3 VDD VSS int_out[15] int_out[14] buf_out[15] C[15] singlestage
x3[7] r2 VDD VSS int_out[31] int_out[30] OUT C[31] singlestage
x3[6] r2 VDD VSS int_out[30] int_out[29] buf_out[30] C[30] singlestage
x3[5] r2 VDD VSS int_out[29] int_out[28] buf_out[29] C[29] singlestage
x3[4] r2 VDD VSS int_out[28] int_out[27] buf_out[28] C[28] singlestage
x3[3] r2 VDD VSS int_out[27] int_out[26] buf_out[27] C[27] singlestage
x3[2] r2 VDD VSS int_out[26] int_out[25] buf_out[26] C[26] singlestage
x3[1] r2 VDD VSS int_out[25] int_out[24] buf_out[25] C[25] singlestage
x3[0] r2 VDD VSS int_out[24] int_out[23] buf_out[24] C[24] singlestage
.ends









** flattened .save nodes

.subckt BR64 VDD VSS OUT
+ C[63] C[62] C[61] C[60] C[59] C[58] C[57] C[56] C[55] C[54] C[53] C[52] C[51] C[50] C[49] C[48] C[47] C[46] C[45] C[44] C[43] C[42] C[41] C[40] C[39] C[38] C[37] C[36] C[35] C[34] C[33] C[32] C[31] C[30] C[29] C[28] C[27] C[26] C[25] C[24] C[23] C[22] C[21] C[20] C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12] C[11] C[10] C[9] C[8] C[7] C[6] C[5] C[4] C[3] C[2] C[1] C[0] RESET
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin
*+ C[63],C[62],C[61],C[60],C[59],C[58],C[57],C[56],C[55],C[54],C[53],C[52],C[51],C[50],C[49],C[48],C[47],C[46],C[45],C[44],C[43],C[42],C[41],C[40],C[39],C[38],C[37],C[36],C[35],C[34],C[33],C[32],C[31],C[30],C[29],C[28],C[27],C[26],C[25],C[24],C[23],C[22],C[21],C[20],C[19],C[18],C[17],C[16],C[15],C[14],C[13],C[12],C[11],C[10],C[9],C[8],C[7],C[6],C[5],C[4],C[3],C[2],C[1],C[0]
*.ipin RESET
x43 RESET VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_4
x47 net1 VSS VSS VDD VDD r6 sky130_fd_sc_hd__inv_16
x48 net1 VSS VSS VDD VDD r5 sky130_fd_sc_hd__inv_16
x4 net1 VSS VSS VDD VDD r5 sky130_fd_sc_hd__inv_16
x5 net1 VSS VSS VDD VDD r6 sky130_fd_sc_hd__inv_16
x6 net1 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x7 net1 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x8 net1 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x10 net1 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x11 net2 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_16
x12 net2 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_16
x13 net3 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x14 net3 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x15 net3 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x16 net3 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x17 net3 VSS VSS VDD VDD r8 sky130_fd_sc_hd__inv_16
x18 net3 VSS VSS VDD VDD r7 sky130_fd_sc_hd__inv_16
x19 net3 VSS VSS VDD VDD r7 sky130_fd_sc_hd__inv_16
x20 net3 VSS VSS VDD VDD r8 sky130_fd_sc_hd__inv_16
x21 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_16
x22 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_16
x23 net4 VSS VSS VDD VDD net2 sky130_fd_sc_hd__inv_16
x3[7] r1 VDD VSS out[8] out[7] net5[7] C[7] singlestage
x3[6] r1 VDD VSS out[7] out[6] net5[6] C[6] singlestage
x3[5] r1 VDD VSS out[6] out[5] net5[5] C[5] singlestage
x3[4] r1 VDD VSS out[5] out[4] net5[4] C[4] singlestage
x3[3] r1 VDD VSS out[4] out[3] net5[3] C[3] singlestage
x3[2] r1 VDD VSS out[3] out[2] net5[2] C[2] singlestage
x3[1] r1 VDD VSS out[2] out[1] net5[1] C[1] singlestage
x3[0] r1 VDD VSS out[1] out[0] net5[0] C[0] singlestage
x1[15] r2 VDD VSS out[16] out[15] net6[7] C[15] singlestage
x1[14] r2 VDD VSS out[15] out[14] net6[6] C[14] singlestage
x1[13] r2 VDD VSS out[14] out[13] net6[5] C[13] singlestage
x1[12] r2 VDD VSS out[13] out[12] net6[4] C[12] singlestage
x1[11] r2 VDD VSS out[12] out[11] net6[3] C[11] singlestage
x1[10] r2 VDD VSS out[11] out[10] net6[2] C[10] singlestage
x1[9] r2 VDD VSS out[10] out[9] net6[1] C[9] singlestage
x1[8] r2 VDD VSS out[9] out[8] net6[0] C[8] singlestage
x2[23] r3 VDD VSS out[24] out[23] net7[7] C[23] singlestage
x2[22] r3 VDD VSS out[23] out[22] net7[6] C[22] singlestage
x2[21] r3 VDD VSS out[22] out[21] net7[5] C[21] singlestage
x2[20] r3 VDD VSS out[21] out[20] net7[4] C[20] singlestage
x2[19] r3 VDD VSS out[20] out[19] net7[3] C[19] singlestage
x2[18] r3 VDD VSS out[19] out[18] net7[2] C[18] singlestage
x2[17] r3 VDD VSS out[18] out[17] net7[1] C[17] singlestage
x2[16] r3 VDD VSS out[17] out[16] net7[0] C[16] singlestage
x4[31] r4 VDD VSS out[32] out[31] net8[7] C[31] singlestage
x4[30] r4 VDD VSS out[31] out[30] net8[6] C[30] singlestage
x4[29] r4 VDD VSS out[30] out[29] net8[5] C[29] singlestage
x4[28] r4 VDD VSS out[29] out[28] net8[4] C[28] singlestage
x4[27] r4 VDD VSS out[28] out[27] net8[3] C[27] singlestage
x4[26] r4 VDD VSS out[27] out[26] net8[2] C[26] singlestage
x4[25] r4 VDD VSS out[26] out[25] net8[1] C[25] singlestage
x4[24] r4 VDD VSS out[25] out[24] net8[0] C[24] singlestage
x5[63] r8 VDD VSS out[0] out[63] OUT C[63] singlestage
x5[62] r8 VDD VSS out[63] out[62] buf_out[6] C[62] singlestage
x5[61] r8 VDD VSS out[62] out[61] buf_out[5] C[61] singlestage
x5[60] r8 VDD VSS out[61] out[60] buf_out[4] C[60] singlestage
x5[59] r8 VDD VSS out[60] out[59] buf_out[3] C[59] singlestage
x5[58] r8 VDD VSS out[59] out[58] buf_out[2] C[58] singlestage
x5[57] r8 VDD VSS out[58] out[57] buf_out[1] C[57] singlestage
x5[56] r8 VDD VSS out[57] out[56] buf_out[0] C[56] singlestage
x6[55] r7 VDD VSS out[56] out[55] net9[7] C[55] singlestage
x6[54] r7 VDD VSS out[55] out[54] net9[6] C[54] singlestage
x6[53] r7 VDD VSS out[54] out[53] net9[5] C[53] singlestage
x6[52] r7 VDD VSS out[53] out[52] net9[4] C[52] singlestage
x6[51] r7 VDD VSS out[52] out[51] net9[3] C[51] singlestage
x6[50] r7 VDD VSS out[51] out[50] net9[2] C[50] singlestage
x6[49] r7 VDD VSS out[50] out[49] net9[1] C[49] singlestage
x6[48] r7 VDD VSS out[49] out[48] net9[0] C[48] singlestage
x7[47] r6 VDD VSS out[48] out[47] net10[7] C[47] singlestage
x7[46] r6 VDD VSS out[47] out[46] net10[6] C[46] singlestage
x7[45] r6 VDD VSS out[46] out[45] net10[5] C[45] singlestage
x7[44] r6 VDD VSS out[45] out[44] net10[4] C[44] singlestage
x7[43] r6 VDD VSS out[44] out[43] net10[3] C[43] singlestage
x7[42] r6 VDD VSS out[43] out[42] net10[2] C[42] singlestage
x7[41] r6 VDD VSS out[42] out[41] net10[1] C[41] singlestage
x7[40] r6 VDD VSS out[41] out[40] net10[0] C[40] singlestage
x8[39] r5 VDD VSS out[40] out[39] net11[7] C[39] singlestage
x8[38] r5 VDD VSS out[39] out[38] net11[6] C[38] singlestage
x8[37] r5 VDD VSS out[38] out[37] net11[5] C[37] singlestage
x8[36] r5 VDD VSS out[37] out[36] net11[4] C[36] singlestage
x8[35] r5 VDD VSS out[36] out[35] net11[3] C[35] singlestage
x8[34] r5 VDD VSS out[35] out[34] net11[2] C[34] singlestage
x8[33] r5 VDD VSS out[34] out[33] net11[1] C[33] singlestage
x8[32] r5 VDD VSS out[33] out[32] net11[0] C[32] singlestage
.ends






** flattened .save nodes

