/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/parasitics/sky130_fd_pr__model__parasitic__res_po.model.spice