magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 443 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 417 177
rect 365 61 375 95
rect 409 61 417 95
rect 365 47 417 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 485 167 497
rect 113 451 123 485
rect 157 451 167 485
rect 113 417 167 451
rect 113 383 123 417
rect 157 383 167 417
rect 113 297 167 383
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 409 335 497
rect 281 375 291 409
rect 325 375 335 409
rect 281 341 335 375
rect 281 307 291 341
rect 325 307 335 341
rect 281 297 335 307
rect 365 485 417 497
rect 365 451 375 485
rect 409 451 417 485
rect 365 417 417 451
rect 365 383 375 417
rect 409 383 417 417
rect 365 297 417 383
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 451 157 485
rect 123 383 157 417
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 375 325 409
rect 291 307 325 341
rect 375 451 409 485
rect 375 383 409 417
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 83 265 113 297
rect 167 265 197 297
rect 83 249 197 265
rect 83 215 112 249
rect 146 215 197 249
rect 83 199 197 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 265 281 297
rect 335 265 365 297
rect 251 249 365 265
rect 251 215 291 249
rect 325 215 365 249
rect 251 199 365 215
rect 251 177 281 199
rect 335 177 365 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
<< polycont >>
rect 112 215 146 249
rect 291 215 325 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 18 477 73 493
rect 18 443 39 477
rect 18 409 73 443
rect 18 375 39 409
rect 18 341 73 375
rect 107 485 173 527
rect 107 451 123 485
rect 157 451 173 485
rect 107 417 173 451
rect 107 383 123 417
rect 157 383 173 417
rect 107 367 173 383
rect 207 485 435 493
rect 207 477 375 485
rect 241 459 375 477
rect 207 409 241 443
rect 409 451 435 485
rect 18 307 39 341
rect 207 341 241 375
rect 73 307 207 333
rect 18 291 241 307
rect 275 409 341 425
rect 275 375 291 409
rect 325 375 341 409
rect 275 341 341 375
rect 375 417 435 451
rect 409 383 435 417
rect 375 367 435 383
rect 275 307 291 341
rect 325 333 341 341
rect 325 307 427 333
rect 275 289 427 307
rect 18 249 162 255
rect 18 215 112 249
rect 146 215 162 249
rect 196 249 350 255
rect 196 215 291 249
rect 325 215 350 249
rect 384 181 427 289
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 427 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 147 427 163
rect 325 129 341 147
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 433 111
rect 409 61 433 95
rect 375 17 433 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 214 221 248 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 306 357 340 391 0 FreeSans 400 0 0 0 Y
port 7 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor2_2
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 1640654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1635912
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
