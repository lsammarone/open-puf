magic
tech sky130A
timestamp 1648127584
<< properties >>
string GDS_END 15511496
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15505796
<< end >>
