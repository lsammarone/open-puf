magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< labels >>
flabel comment s 36 5 36 5 2 FreeSans 50 0 0 0 EM1C
flabel comment s 62 15 62 15 0 FreeSans 50 0 0 0 A
flabel comment s 30 15 30 15 0 FreeSans 50 0 0 0 A
<< properties >>
string GDS_END 30709420
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30708716
<< end >>
