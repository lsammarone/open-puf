magic
tech sky130B
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_0
timestamp 1648127584
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180819  sky130_fd_pr__dfl1sd__example_5595914180819_1
timestamp 1648127584
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7397032
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7396110
<< end >>
