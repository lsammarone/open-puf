**.subckt demux2-1
**.ends
** flattened .save nodes
.end
