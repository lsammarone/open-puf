magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 81 43 699 294
rect -26 -43 794 43
<< mvnmos >>
rect 160 118 360 268
rect 416 118 616 268
<< mvpmos >>
rect 147 540 347 740
rect 403 540 603 740
<< mvndiff >>
rect 107 256 160 268
rect 107 222 115 256
rect 149 222 160 256
rect 107 178 160 222
rect 107 144 115 178
rect 149 144 160 178
rect 107 118 160 144
rect 360 256 416 268
rect 360 222 371 256
rect 405 222 416 256
rect 360 178 416 222
rect 360 144 371 178
rect 405 144 416 178
rect 360 118 416 144
rect 616 256 673 268
rect 616 222 627 256
rect 661 222 673 256
rect 616 178 673 222
rect 616 144 627 178
rect 661 144 673 178
rect 616 118 673 144
<< mvpdiff >>
rect 92 728 147 740
rect 92 694 100 728
rect 134 694 147 728
rect 92 657 147 694
rect 92 623 100 657
rect 134 623 147 657
rect 92 586 147 623
rect 92 552 100 586
rect 134 552 147 586
rect 92 540 147 552
rect 347 728 403 740
rect 347 694 358 728
rect 392 694 403 728
rect 347 657 403 694
rect 347 623 358 657
rect 392 623 403 657
rect 347 586 403 623
rect 347 552 358 586
rect 392 552 403 586
rect 347 540 403 552
rect 603 728 660 740
rect 603 694 614 728
rect 648 694 660 728
rect 603 657 660 694
rect 603 623 614 657
rect 648 623 660 657
rect 603 586 660 623
rect 603 552 614 586
rect 648 552 660 586
rect 603 540 660 552
<< mvndiffc >>
rect 115 222 149 256
rect 115 144 149 178
rect 371 222 405 256
rect 371 144 405 178
rect 627 222 661 256
rect 627 144 661 178
<< mvpdiffc >>
rect 100 694 134 728
rect 100 623 134 657
rect 100 552 134 586
rect 358 694 392 728
rect 358 623 392 657
rect 358 552 392 586
rect 614 694 648 728
rect 614 623 648 657
rect 614 552 648 586
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
<< poly >>
rect 147 740 347 766
rect 403 740 603 766
rect 147 514 347 540
rect 403 514 603 540
rect 147 389 213 514
rect 147 355 163 389
rect 197 355 213 389
rect 147 339 213 355
rect 294 389 360 405
rect 294 355 310 389
rect 344 355 360 389
rect 294 294 360 355
rect 403 389 469 514
rect 403 355 419 389
rect 453 355 469 389
rect 403 339 469 355
rect 550 389 616 405
rect 550 355 566 389
rect 600 355 616 389
rect 550 294 616 355
rect 160 268 360 294
rect 416 268 616 294
rect 160 80 360 118
rect 416 80 616 118
<< polycont >>
rect 163 355 197 389
rect 310 355 344 389
rect 419 355 453 389
rect 566 355 600 389
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 100 745 648 750
rect 100 728 141 745
rect 134 711 141 728
rect 175 711 229 745
rect 263 711 312 745
rect 346 728 397 745
rect 346 711 358 728
rect 134 694 358 711
rect 392 711 397 728
rect 431 711 485 745
rect 519 711 568 745
rect 602 728 648 745
rect 602 711 614 728
rect 392 694 614 711
rect 100 657 648 694
rect 134 623 358 657
rect 392 623 614 657
rect 100 586 648 623
rect 134 552 358 586
rect 392 552 614 586
rect 100 536 648 552
rect 147 389 213 405
rect 147 355 163 389
rect 197 355 213 389
rect 147 272 213 355
rect 294 389 360 536
rect 294 355 310 389
rect 344 355 360 389
rect 294 339 360 355
rect 403 389 469 405
rect 403 355 419 389
rect 453 355 469 389
rect 403 272 469 355
rect 550 389 616 536
rect 550 355 566 389
rect 600 355 616 389
rect 550 339 616 355
rect 115 256 661 272
rect 149 222 371 256
rect 405 222 627 256
rect 115 178 661 222
rect 149 144 371 178
rect 405 144 627 178
rect 115 112 661 144
rect 115 78 149 112
rect 183 78 237 112
rect 271 78 320 112
rect 354 78 405 112
rect 439 78 493 112
rect 527 78 576 112
rect 610 78 661 112
rect 115 72 661 78
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 141 711 175 745
rect 229 711 263 745
rect 312 711 346 745
rect 397 711 431 745
rect 485 711 519 745
rect 568 711 602 745
rect 149 78 183 112
rect 237 78 271 112
rect 320 78 354 112
rect 405 78 439 112
rect 493 78 527 112
rect 576 78 610 112
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 745 768 763
rect 0 711 141 745
rect 175 711 229 745
rect 263 711 312 745
rect 346 711 397 745
rect 431 711 485 745
rect 519 711 568 745
rect 602 711 768 745
rect 0 689 768 711
rect 0 112 768 125
rect 0 78 149 112
rect 183 78 237 112
rect 271 78 320 112
rect 354 78 405 112
rect 439 78 493 112
rect 527 78 576 112
rect 610 78 768 112
rect 0 51 768 78
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 decap_8
flabel metal1 s 0 0 768 23 0 FreeSans 340 0 0 0 VNB
port 2 nsew ground bidirectional
flabel metal1 s 0 51 768 125 0 FreeSans 340 0 0 0 VGND
port 1 nsew ground bidirectional
flabel metal1 s 384 11 384 11 0 FreeSans 340 0 0 0 VNB
port 2 nsew
flabel metal1 s 0 689 768 763 0 FreeSans 340 0 0 0 VPWR
port 4 nsew power bidirectional
flabel metal1 s 0 791 768 814 0 FreeSans 340 0 0 0 VPB
port 3 nsew power bidirectional
flabel metal1 s 384 802 384 802 0 FreeSans 340 0 0 0 VPB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 768 814
string GDS_END 955054
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 948224
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
