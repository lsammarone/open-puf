magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< pwell >>
rect 0 66 700 720
<< nmoslvt >>
rect 194 92 230 694
rect 286 92 322 694
rect 378 92 414 694
rect 470 92 506 694
<< ndiff >>
rect 138 682 194 694
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 230 682 286 694
rect 230 648 241 682
rect 275 648 286 682
rect 230 614 286 648
rect 230 580 241 614
rect 275 580 286 614
rect 230 546 286 580
rect 230 512 241 546
rect 275 512 286 546
rect 230 478 286 512
rect 230 444 241 478
rect 275 444 286 478
rect 230 410 286 444
rect 230 376 241 410
rect 275 376 286 410
rect 230 342 286 376
rect 230 308 241 342
rect 275 308 286 342
rect 230 274 286 308
rect 230 240 241 274
rect 275 240 286 274
rect 230 206 286 240
rect 230 172 241 206
rect 275 172 286 206
rect 230 138 286 172
rect 230 104 241 138
rect 275 104 286 138
rect 230 92 286 104
rect 322 682 378 694
rect 322 648 333 682
rect 367 648 378 682
rect 322 614 378 648
rect 322 580 333 614
rect 367 580 378 614
rect 322 546 378 580
rect 322 512 333 546
rect 367 512 378 546
rect 322 478 378 512
rect 322 444 333 478
rect 367 444 378 478
rect 322 410 378 444
rect 322 376 333 410
rect 367 376 378 410
rect 322 342 378 376
rect 322 308 333 342
rect 367 308 378 342
rect 322 274 378 308
rect 322 240 333 274
rect 367 240 378 274
rect 322 206 378 240
rect 322 172 333 206
rect 367 172 378 206
rect 322 138 378 172
rect 322 104 333 138
rect 367 104 378 138
rect 322 92 378 104
rect 414 682 470 694
rect 414 648 425 682
rect 459 648 470 682
rect 414 614 470 648
rect 414 580 425 614
rect 459 580 470 614
rect 414 546 470 580
rect 414 512 425 546
rect 459 512 470 546
rect 414 478 470 512
rect 414 444 425 478
rect 459 444 470 478
rect 414 410 470 444
rect 414 376 425 410
rect 459 376 470 410
rect 414 342 470 376
rect 414 308 425 342
rect 459 308 470 342
rect 414 274 470 308
rect 414 240 425 274
rect 459 240 470 274
rect 414 206 470 240
rect 414 172 425 206
rect 459 172 470 206
rect 414 138 470 172
rect 414 104 425 138
rect 459 104 470 138
rect 414 92 470 104
rect 506 682 562 694
rect 506 648 517 682
rect 551 648 562 682
rect 506 614 562 648
rect 506 580 517 614
rect 551 580 562 614
rect 506 546 562 580
rect 506 512 517 546
rect 551 512 562 546
rect 506 478 562 512
rect 506 444 517 478
rect 551 444 562 478
rect 506 410 562 444
rect 506 376 517 410
rect 551 376 562 410
rect 506 342 562 376
rect 506 308 517 342
rect 551 308 562 342
rect 506 274 562 308
rect 506 240 517 274
rect 551 240 562 274
rect 506 206 562 240
rect 506 172 517 206
rect 551 172 562 206
rect 506 138 562 172
rect 506 104 517 138
rect 551 104 562 138
rect 506 92 562 104
<< ndiffc >>
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 241 648 275 682
rect 241 580 275 614
rect 241 512 275 546
rect 241 444 275 478
rect 241 376 275 410
rect 241 308 275 342
rect 241 240 275 274
rect 241 172 275 206
rect 241 104 275 138
rect 333 648 367 682
rect 333 580 367 614
rect 333 512 367 546
rect 333 444 367 478
rect 333 376 367 410
rect 333 308 367 342
rect 333 240 367 274
rect 333 172 367 206
rect 333 104 367 138
rect 425 648 459 682
rect 425 580 459 614
rect 425 512 459 546
rect 425 444 459 478
rect 425 376 459 410
rect 425 308 459 342
rect 425 240 459 274
rect 425 172 459 206
rect 425 104 459 138
rect 517 648 551 682
rect 517 580 551 614
rect 517 512 551 546
rect 517 444 551 478
rect 517 376 551 410
rect 517 308 551 342
rect 517 240 551 274
rect 517 172 551 206
rect 517 104 551 138
<< psubdiff >>
rect 26 648 84 694
rect 26 614 38 648
rect 72 614 84 648
rect 26 580 84 614
rect 26 546 38 580
rect 72 546 84 580
rect 26 512 84 546
rect 26 478 38 512
rect 72 478 84 512
rect 26 444 84 478
rect 26 410 38 444
rect 72 410 84 444
rect 26 376 84 410
rect 26 342 38 376
rect 72 342 84 376
rect 26 308 84 342
rect 26 274 38 308
rect 72 274 84 308
rect 26 240 84 274
rect 26 206 38 240
rect 72 206 84 240
rect 26 172 84 206
rect 26 138 38 172
rect 72 138 84 172
rect 26 92 84 138
rect 616 648 674 694
rect 616 614 628 648
rect 662 614 674 648
rect 616 580 674 614
rect 616 546 628 580
rect 662 546 674 580
rect 616 512 674 546
rect 616 478 628 512
rect 662 478 674 512
rect 616 444 674 478
rect 616 410 628 444
rect 662 410 674 444
rect 616 376 674 410
rect 616 342 628 376
rect 662 342 674 376
rect 616 308 674 342
rect 616 274 628 308
rect 662 274 674 308
rect 616 240 674 274
rect 616 206 628 240
rect 662 206 674 240
rect 616 172 674 206
rect 616 138 628 172
rect 662 138 674 172
rect 616 92 674 138
<< psubdiffcont >>
rect 38 614 72 648
rect 38 546 72 580
rect 38 478 72 512
rect 38 410 72 444
rect 38 342 72 376
rect 38 274 72 308
rect 38 206 72 240
rect 38 138 72 172
rect 628 614 662 648
rect 628 546 662 580
rect 628 478 662 512
rect 628 410 662 444
rect 628 342 662 376
rect 628 274 662 308
rect 628 206 662 240
rect 628 138 662 172
<< poly >>
rect 181 766 519 786
rect 181 732 197 766
rect 231 732 265 766
rect 299 732 333 766
rect 367 732 401 766
rect 435 732 469 766
rect 503 732 519 766
rect 181 716 519 732
rect 194 694 230 716
rect 286 694 322 716
rect 378 694 414 716
rect 470 694 506 716
rect 194 70 230 92
rect 286 70 322 92
rect 378 70 414 92
rect 470 70 506 92
rect 181 54 519 70
rect 181 20 197 54
rect 231 20 265 54
rect 299 20 333 54
rect 367 20 401 54
rect 435 20 469 54
rect 503 20 519 54
rect 181 0 519 20
<< polycont >>
rect 197 732 231 766
rect 265 732 299 766
rect 333 732 367 766
rect 401 732 435 766
rect 469 732 503 766
rect 197 20 231 54
rect 265 20 299 54
rect 333 20 367 54
rect 401 20 435 54
rect 469 20 503 54
<< locali >>
rect 181 732 189 766
rect 231 732 261 766
rect 299 732 333 766
rect 367 732 401 766
rect 439 732 469 766
rect 511 732 519 766
rect 149 682 183 698
rect 38 662 72 664
rect 38 590 72 614
rect 38 518 72 546
rect 38 446 72 478
rect 38 376 72 410
rect 38 308 72 340
rect 38 240 72 268
rect 38 172 72 196
rect 38 122 72 124
rect 149 614 183 628
rect 149 546 183 556
rect 149 478 183 484
rect 149 410 183 412
rect 149 374 183 376
rect 149 302 183 308
rect 149 230 183 240
rect 149 158 183 172
rect 149 88 183 104
rect 241 682 275 698
rect 241 614 275 628
rect 241 546 275 556
rect 241 478 275 484
rect 241 410 275 412
rect 241 374 275 376
rect 241 302 275 308
rect 241 230 275 240
rect 241 158 275 172
rect 241 88 275 104
rect 333 682 367 698
rect 333 614 367 628
rect 333 546 367 556
rect 333 478 367 484
rect 333 410 367 412
rect 333 374 367 376
rect 333 302 367 308
rect 333 230 367 240
rect 333 158 367 172
rect 333 88 367 104
rect 425 682 459 698
rect 425 614 459 628
rect 425 546 459 556
rect 425 478 459 484
rect 425 410 459 412
rect 425 374 459 376
rect 425 302 459 308
rect 425 230 459 240
rect 425 158 459 172
rect 425 88 459 104
rect 517 682 551 698
rect 517 614 551 628
rect 517 546 551 556
rect 517 478 551 484
rect 517 410 551 412
rect 517 374 551 376
rect 517 302 551 308
rect 517 230 551 240
rect 517 158 551 172
rect 628 662 662 664
rect 628 590 662 614
rect 628 518 662 546
rect 628 446 662 478
rect 628 376 662 410
rect 628 308 662 340
rect 628 240 662 268
rect 628 172 662 196
rect 628 122 662 124
rect 517 88 551 104
rect 181 20 189 54
rect 231 20 261 54
rect 299 20 333 54
rect 367 20 401 54
rect 439 20 469 54
rect 511 20 519 54
<< viali >>
rect 189 732 197 766
rect 197 732 223 766
rect 261 732 265 766
rect 265 732 295 766
rect 333 732 367 766
rect 405 732 435 766
rect 435 732 439 766
rect 477 732 503 766
rect 503 732 511 766
rect 38 648 72 662
rect 38 628 72 648
rect 38 580 72 590
rect 38 556 72 580
rect 38 512 72 518
rect 38 484 72 512
rect 38 444 72 446
rect 38 412 72 444
rect 38 342 72 374
rect 38 340 72 342
rect 38 274 72 302
rect 38 268 72 274
rect 38 206 72 230
rect 38 196 72 206
rect 38 138 72 158
rect 38 124 72 138
rect 149 648 183 662
rect 149 628 183 648
rect 149 580 183 590
rect 149 556 183 580
rect 149 512 183 518
rect 149 484 183 512
rect 149 444 183 446
rect 149 412 183 444
rect 149 342 183 374
rect 149 340 183 342
rect 149 274 183 302
rect 149 268 183 274
rect 149 206 183 230
rect 149 196 183 206
rect 149 138 183 158
rect 149 124 183 138
rect 241 648 275 662
rect 241 628 275 648
rect 241 580 275 590
rect 241 556 275 580
rect 241 512 275 518
rect 241 484 275 512
rect 241 444 275 446
rect 241 412 275 444
rect 241 342 275 374
rect 241 340 275 342
rect 241 274 275 302
rect 241 268 275 274
rect 241 206 275 230
rect 241 196 275 206
rect 241 138 275 158
rect 241 124 275 138
rect 333 648 367 662
rect 333 628 367 648
rect 333 580 367 590
rect 333 556 367 580
rect 333 512 367 518
rect 333 484 367 512
rect 333 444 367 446
rect 333 412 367 444
rect 333 342 367 374
rect 333 340 367 342
rect 333 274 367 302
rect 333 268 367 274
rect 333 206 367 230
rect 333 196 367 206
rect 333 138 367 158
rect 333 124 367 138
rect 425 648 459 662
rect 425 628 459 648
rect 425 580 459 590
rect 425 556 459 580
rect 425 512 459 518
rect 425 484 459 512
rect 425 444 459 446
rect 425 412 459 444
rect 425 342 459 374
rect 425 340 459 342
rect 425 274 459 302
rect 425 268 459 274
rect 425 206 459 230
rect 425 196 459 206
rect 425 138 459 158
rect 425 124 459 138
rect 517 648 551 662
rect 517 628 551 648
rect 517 580 551 590
rect 517 556 551 580
rect 517 512 551 518
rect 517 484 551 512
rect 517 444 551 446
rect 517 412 551 444
rect 517 342 551 374
rect 517 340 551 342
rect 517 274 551 302
rect 517 268 551 274
rect 517 206 551 230
rect 517 196 551 206
rect 517 138 551 158
rect 517 124 551 138
rect 628 648 662 662
rect 628 628 662 648
rect 628 580 662 590
rect 628 556 662 580
rect 628 512 662 518
rect 628 484 662 512
rect 628 444 662 446
rect 628 412 662 444
rect 628 342 662 374
rect 628 340 662 342
rect 628 274 662 302
rect 628 268 662 274
rect 628 206 662 230
rect 628 196 662 206
rect 628 138 662 158
rect 628 124 662 138
rect 189 20 197 54
rect 197 20 223 54
rect 261 20 265 54
rect 265 20 295 54
rect 333 20 367 54
rect 405 20 435 54
rect 435 20 439 54
rect 477 20 503 54
rect 503 20 511 54
<< metal1 >>
rect 177 766 523 786
rect 177 732 189 766
rect 223 732 261 766
rect 295 732 333 766
rect 367 732 405 766
rect 439 732 477 766
rect 511 732 523 766
rect 177 720 523 732
rect 26 662 84 674
rect 26 628 38 662
rect 72 628 84 662
rect 26 590 84 628
rect 26 556 38 590
rect 72 556 84 590
rect 26 518 84 556
rect 26 484 38 518
rect 72 484 84 518
rect 26 446 84 484
rect 26 412 38 446
rect 72 412 84 446
rect 26 374 84 412
rect 26 340 38 374
rect 72 340 84 374
rect 26 302 84 340
rect 26 268 38 302
rect 72 268 84 302
rect 26 230 84 268
rect 26 196 38 230
rect 72 196 84 230
rect 26 158 84 196
rect 26 124 38 158
rect 72 124 84 158
rect 26 112 84 124
rect 140 662 192 674
rect 140 628 149 662
rect 183 628 192 662
rect 140 590 192 628
rect 140 556 149 590
rect 183 556 192 590
rect 140 518 192 556
rect 140 484 149 518
rect 183 484 192 518
rect 140 446 192 484
rect 140 412 149 446
rect 183 412 192 446
rect 140 374 192 412
rect 140 362 149 374
rect 183 362 192 374
rect 140 302 192 310
rect 140 298 149 302
rect 183 298 192 302
rect 140 234 192 246
rect 140 170 192 182
rect 140 112 192 118
rect 232 668 284 674
rect 232 604 284 616
rect 232 540 284 552
rect 232 484 241 488
rect 275 484 284 488
rect 232 476 284 484
rect 232 412 241 424
rect 275 412 284 424
rect 232 374 284 412
rect 232 340 241 374
rect 275 340 284 374
rect 232 302 284 340
rect 232 268 241 302
rect 275 268 284 302
rect 232 230 284 268
rect 232 196 241 230
rect 275 196 284 230
rect 232 158 284 196
rect 232 124 241 158
rect 275 124 284 158
rect 232 112 284 124
rect 324 662 376 674
rect 324 628 333 662
rect 367 628 376 662
rect 324 590 376 628
rect 324 556 333 590
rect 367 556 376 590
rect 324 518 376 556
rect 324 484 333 518
rect 367 484 376 518
rect 324 446 376 484
rect 324 412 333 446
rect 367 412 376 446
rect 324 374 376 412
rect 324 362 333 374
rect 367 362 376 374
rect 324 302 376 310
rect 324 298 333 302
rect 367 298 376 302
rect 324 234 376 246
rect 324 170 376 182
rect 324 112 376 118
rect 416 668 468 674
rect 416 604 468 616
rect 416 540 468 552
rect 416 484 425 488
rect 459 484 468 488
rect 416 476 468 484
rect 416 412 425 424
rect 459 412 468 424
rect 416 374 468 412
rect 416 340 425 374
rect 459 340 468 374
rect 416 302 468 340
rect 416 268 425 302
rect 459 268 468 302
rect 416 230 468 268
rect 416 196 425 230
rect 459 196 468 230
rect 416 158 468 196
rect 416 124 425 158
rect 459 124 468 158
rect 416 112 468 124
rect 508 662 560 674
rect 508 628 517 662
rect 551 628 560 662
rect 508 590 560 628
rect 508 556 517 590
rect 551 556 560 590
rect 508 518 560 556
rect 508 484 517 518
rect 551 484 560 518
rect 508 446 560 484
rect 508 412 517 446
rect 551 412 560 446
rect 508 374 560 412
rect 508 362 517 374
rect 551 362 560 374
rect 508 302 560 310
rect 508 298 517 302
rect 551 298 560 302
rect 508 234 560 246
rect 508 170 560 182
rect 508 112 560 118
rect 616 662 674 674
rect 616 628 628 662
rect 662 628 674 662
rect 616 590 674 628
rect 616 556 628 590
rect 662 556 674 590
rect 616 518 674 556
rect 616 484 628 518
rect 662 484 674 518
rect 616 446 674 484
rect 616 412 628 446
rect 662 412 674 446
rect 616 374 674 412
rect 616 340 628 374
rect 662 340 674 374
rect 616 302 674 340
rect 616 268 628 302
rect 662 268 674 302
rect 616 230 674 268
rect 616 196 628 230
rect 662 196 674 230
rect 616 158 674 196
rect 616 124 628 158
rect 662 124 674 158
rect 616 112 674 124
rect 177 54 523 66
rect 177 20 189 54
rect 223 20 261 54
rect 295 20 333 54
rect 367 20 405 54
rect 439 20 477 54
rect 511 20 523 54
rect 177 0 523 20
<< via1 >>
rect 140 340 149 362
rect 149 340 183 362
rect 183 340 192 362
rect 140 310 192 340
rect 140 268 149 298
rect 149 268 183 298
rect 183 268 192 298
rect 140 246 192 268
rect 140 230 192 234
rect 140 196 149 230
rect 149 196 183 230
rect 183 196 192 230
rect 140 182 192 196
rect 140 158 192 170
rect 140 124 149 158
rect 149 124 183 158
rect 183 124 192 158
rect 140 118 192 124
rect 232 662 284 668
rect 232 628 241 662
rect 241 628 275 662
rect 275 628 284 662
rect 232 616 284 628
rect 232 590 284 604
rect 232 556 241 590
rect 241 556 275 590
rect 275 556 284 590
rect 232 552 284 556
rect 232 518 284 540
rect 232 488 241 518
rect 241 488 275 518
rect 275 488 284 518
rect 232 446 284 476
rect 232 424 241 446
rect 241 424 275 446
rect 275 424 284 446
rect 324 340 333 362
rect 333 340 367 362
rect 367 340 376 362
rect 324 310 376 340
rect 324 268 333 298
rect 333 268 367 298
rect 367 268 376 298
rect 324 246 376 268
rect 324 230 376 234
rect 324 196 333 230
rect 333 196 367 230
rect 367 196 376 230
rect 324 182 376 196
rect 324 158 376 170
rect 324 124 333 158
rect 333 124 367 158
rect 367 124 376 158
rect 324 118 376 124
rect 416 662 468 668
rect 416 628 425 662
rect 425 628 459 662
rect 459 628 468 662
rect 416 616 468 628
rect 416 590 468 604
rect 416 556 425 590
rect 425 556 459 590
rect 459 556 468 590
rect 416 552 468 556
rect 416 518 468 540
rect 416 488 425 518
rect 425 488 459 518
rect 459 488 468 518
rect 416 446 468 476
rect 416 424 425 446
rect 425 424 459 446
rect 459 424 468 446
rect 508 340 517 362
rect 517 340 551 362
rect 551 340 560 362
rect 508 310 560 340
rect 508 268 517 298
rect 517 268 551 298
rect 551 268 560 298
rect 508 246 560 268
rect 508 230 560 234
rect 508 196 517 230
rect 517 196 551 230
rect 551 196 560 230
rect 508 182 560 196
rect 508 158 560 170
rect 508 124 517 158
rect 517 124 551 158
rect 551 124 560 158
rect 508 118 560 124
<< metal2 >>
rect 0 668 700 674
rect 0 616 232 668
rect 284 616 416 668
rect 468 616 700 668
rect 0 604 700 616
rect 0 552 232 604
rect 284 552 416 604
rect 468 552 700 604
rect 0 540 700 552
rect 0 488 232 540
rect 284 488 416 540
rect 468 488 700 540
rect 0 476 700 488
rect 0 424 232 476
rect 284 424 416 476
rect 468 424 700 476
rect 0 418 700 424
rect 0 362 700 368
rect 0 310 140 362
rect 192 310 324 362
rect 376 310 508 362
rect 560 310 700 362
rect 0 298 700 310
rect 0 246 140 298
rect 192 246 324 298
rect 376 246 508 298
rect 560 246 700 298
rect 0 234 700 246
rect 0 182 140 234
rect 192 182 324 234
rect 376 182 508 234
rect 560 182 700 234
rect 0 170 700 182
rect 0 118 140 170
rect 192 118 324 170
rect 376 118 508 170
rect 560 118 700 170
rect 0 112 700 118
<< labels >>
flabel comment s 166 393 166 393 0 FreeSans 300 0 0 0 S
flabel comment s 350 393 350 393 0 FreeSans 300 0 0 0 S
flabel comment s 258 393 258 393 0 FreeSans 300 0 0 0 D
flabel comment s 534 393 534 393 0 FreeSans 300 0 0 0 S
flabel comment s 166 393 166 393 0 FreeSans 300 0 0 0 S
flabel comment s 442 393 442 393 0 FreeSans 300 0 0 0 S
flabel comment s 350 393 350 393 0 FreeSans 300 0 0 0 S
flabel comment s 258 393 258 393 0 FreeSans 300 0 0 0 S
flabel comment s 442 393 442 393 0 FreeSans 300 0 0 0 D
flabel metal2 s 4 509 23 579 0 FreeSans 400 90 0 0 DRAIN
port 1 nsew
flabel metal2 s 3 195 24 259 0 FreeSans 400 90 0 0 SOURCE
port 3 nsew
flabel metal1 s 48 511 48 511 7 FreeSans 400 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 643 492 643 492 7 FreeSans 400 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 311 23 393 48 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel metal1 s 298 737 380 762 0 FreeSans 400 0 0 0 GATE
port 2 nsew
<< properties >>
string GDS_END 6163736
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6148110
<< end >>
