magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1887 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 751 47 781 177
rect 835 47 865 177
rect 919 47 949 177
rect 1003 47 1033 177
rect 1191 47 1221 177
rect 1275 47 1305 177
rect 1359 47 1389 177
rect 1443 47 1473 177
rect 1527 47 1557 177
rect 1611 47 1641 177
rect 1695 47 1725 177
rect 1779 47 1809 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
rect 1003 297 1033 497
rect 1191 297 1221 497
rect 1275 297 1305 497
rect 1359 297 1389 497
rect 1443 297 1473 497
rect 1527 297 1557 497
rect 1611 297 1641 497
rect 1695 297 1725 497
rect 1779 297 1809 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 95 163 129
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 95 247 177
rect 193 61 203 95
rect 237 61 247 95
rect 193 47 247 61
rect 277 163 331 177
rect 277 129 287 163
rect 321 129 331 163
rect 277 95 331 129
rect 277 61 287 95
rect 321 61 331 95
rect 277 47 331 61
rect 361 163 415 177
rect 361 129 371 163
rect 405 129 415 163
rect 361 47 415 129
rect 445 95 499 177
rect 445 61 455 95
rect 489 61 499 95
rect 445 47 499 61
rect 529 163 583 177
rect 529 129 539 163
rect 573 129 583 163
rect 529 47 583 129
rect 613 95 667 177
rect 613 61 623 95
rect 657 61 667 95
rect 613 47 667 61
rect 697 95 751 177
rect 697 61 707 95
rect 741 61 751 95
rect 697 47 751 61
rect 781 163 835 177
rect 781 129 791 163
rect 825 129 835 163
rect 781 95 835 129
rect 781 61 791 95
rect 825 61 835 95
rect 781 47 835 61
rect 865 95 919 177
rect 865 61 875 95
rect 909 61 919 95
rect 865 47 919 61
rect 949 163 1003 177
rect 949 129 959 163
rect 993 129 1003 163
rect 949 95 1003 129
rect 949 61 959 95
rect 993 61 1003 95
rect 949 47 1003 61
rect 1033 95 1191 177
rect 1033 61 1043 95
rect 1077 61 1147 95
rect 1181 61 1191 95
rect 1033 47 1191 61
rect 1221 163 1275 177
rect 1221 129 1231 163
rect 1265 129 1275 163
rect 1221 95 1275 129
rect 1221 61 1231 95
rect 1265 61 1275 95
rect 1221 47 1275 61
rect 1305 95 1359 177
rect 1305 61 1315 95
rect 1349 61 1359 95
rect 1305 47 1359 61
rect 1389 163 1443 177
rect 1389 129 1399 163
rect 1433 129 1443 163
rect 1389 95 1443 129
rect 1389 61 1399 95
rect 1433 61 1443 95
rect 1389 47 1443 61
rect 1473 95 1527 177
rect 1473 61 1483 95
rect 1517 61 1527 95
rect 1473 47 1527 61
rect 1557 163 1611 177
rect 1557 129 1567 163
rect 1601 129 1611 163
rect 1557 95 1611 129
rect 1557 61 1567 95
rect 1601 61 1611 95
rect 1557 47 1611 61
rect 1641 95 1695 177
rect 1641 61 1651 95
rect 1685 61 1695 95
rect 1641 47 1695 61
rect 1725 163 1779 177
rect 1725 129 1735 163
rect 1769 129 1779 163
rect 1725 95 1779 129
rect 1725 61 1735 95
rect 1769 61 1779 95
rect 1725 47 1779 61
rect 1809 95 1861 177
rect 1809 61 1819 95
rect 1853 61 1861 95
rect 1809 47 1861 61
<< pdiff >>
rect 27 483 79 497
rect 27 449 35 483
rect 69 449 79 483
rect 27 415 79 449
rect 27 381 35 415
rect 69 381 79 415
rect 27 347 79 381
rect 27 313 35 347
rect 69 313 79 347
rect 27 297 79 313
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 341 247 375
rect 193 307 203 341
rect 237 307 247 341
rect 193 297 247 307
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 297 331 443
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 477 499 497
rect 445 443 455 477
rect 489 443 499 477
rect 445 297 499 443
rect 529 477 583 497
rect 529 443 539 477
rect 573 443 583 477
rect 529 409 583 443
rect 529 375 539 409
rect 573 375 583 409
rect 529 297 583 375
rect 613 477 667 497
rect 613 443 623 477
rect 657 443 667 477
rect 613 297 667 443
rect 697 477 751 497
rect 697 443 707 477
rect 741 443 751 477
rect 697 409 751 443
rect 697 375 707 409
rect 741 375 751 409
rect 697 297 751 375
rect 781 409 835 497
rect 781 375 791 409
rect 825 375 835 409
rect 781 341 835 375
rect 781 307 791 341
rect 825 307 835 341
rect 781 297 835 307
rect 865 477 919 497
rect 865 443 875 477
rect 909 443 919 477
rect 865 409 919 443
rect 865 375 875 409
rect 909 375 919 409
rect 865 297 919 375
rect 949 409 1003 497
rect 949 375 959 409
rect 993 375 1003 409
rect 949 341 1003 375
rect 949 307 959 341
rect 993 307 1003 341
rect 949 297 1003 307
rect 1033 483 1085 497
rect 1033 449 1043 483
rect 1077 449 1085 483
rect 1033 415 1085 449
rect 1033 381 1043 415
rect 1077 381 1085 415
rect 1033 347 1085 381
rect 1033 313 1043 347
rect 1077 313 1085 347
rect 1033 297 1085 313
rect 1139 483 1191 497
rect 1139 449 1147 483
rect 1181 449 1191 483
rect 1139 415 1191 449
rect 1139 381 1147 415
rect 1181 381 1191 415
rect 1139 347 1191 381
rect 1139 313 1147 347
rect 1181 313 1191 347
rect 1139 297 1191 313
rect 1221 477 1275 497
rect 1221 443 1231 477
rect 1265 443 1275 477
rect 1221 409 1275 443
rect 1221 375 1231 409
rect 1265 375 1275 409
rect 1221 297 1275 375
rect 1305 477 1359 497
rect 1305 443 1315 477
rect 1349 443 1359 477
rect 1305 409 1359 443
rect 1305 375 1315 409
rect 1349 375 1359 409
rect 1305 341 1359 375
rect 1305 307 1315 341
rect 1349 307 1359 341
rect 1305 297 1359 307
rect 1389 477 1443 497
rect 1389 443 1399 477
rect 1433 443 1443 477
rect 1389 409 1443 443
rect 1389 375 1399 409
rect 1433 375 1443 409
rect 1389 297 1443 375
rect 1473 477 1527 497
rect 1473 443 1483 477
rect 1517 443 1527 477
rect 1473 409 1527 443
rect 1473 375 1483 409
rect 1517 375 1527 409
rect 1473 341 1527 375
rect 1473 307 1483 341
rect 1517 307 1527 341
rect 1473 297 1527 307
rect 1557 409 1611 497
rect 1557 375 1567 409
rect 1601 375 1611 409
rect 1557 341 1611 375
rect 1557 307 1567 341
rect 1601 307 1611 341
rect 1557 297 1611 307
rect 1641 477 1695 497
rect 1641 443 1651 477
rect 1685 443 1695 477
rect 1641 297 1695 443
rect 1725 409 1779 497
rect 1725 375 1735 409
rect 1769 375 1779 409
rect 1725 341 1779 375
rect 1725 307 1735 341
rect 1769 307 1779 341
rect 1725 297 1779 307
rect 1809 477 1865 497
rect 1809 443 1819 477
rect 1853 443 1865 477
rect 1809 409 1865 443
rect 1809 375 1819 409
rect 1853 375 1865 409
rect 1809 297 1865 375
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 119 129 153 163
rect 119 61 153 95
rect 203 61 237 95
rect 287 129 321 163
rect 287 61 321 95
rect 371 129 405 163
rect 455 61 489 95
rect 539 129 573 163
rect 623 61 657 95
rect 707 61 741 95
rect 791 129 825 163
rect 791 61 825 95
rect 875 61 909 95
rect 959 129 993 163
rect 959 61 993 95
rect 1043 61 1077 95
rect 1147 61 1181 95
rect 1231 129 1265 163
rect 1231 61 1265 95
rect 1315 61 1349 95
rect 1399 129 1433 163
rect 1399 61 1433 95
rect 1483 61 1517 95
rect 1567 129 1601 163
rect 1567 61 1601 95
rect 1651 61 1685 95
rect 1735 129 1769 163
rect 1735 61 1769 95
rect 1819 61 1853 95
<< pdiffc >>
rect 35 449 69 483
rect 35 381 69 415
rect 35 313 69 347
rect 119 443 153 477
rect 119 375 153 409
rect 203 443 237 477
rect 203 375 237 409
rect 203 307 237 341
rect 287 443 321 477
rect 371 443 405 477
rect 371 375 405 409
rect 455 443 489 477
rect 539 443 573 477
rect 539 375 573 409
rect 623 443 657 477
rect 707 443 741 477
rect 707 375 741 409
rect 791 375 825 409
rect 791 307 825 341
rect 875 443 909 477
rect 875 375 909 409
rect 959 375 993 409
rect 959 307 993 341
rect 1043 449 1077 483
rect 1043 381 1077 415
rect 1043 313 1077 347
rect 1147 449 1181 483
rect 1147 381 1181 415
rect 1147 313 1181 347
rect 1231 443 1265 477
rect 1231 375 1265 409
rect 1315 443 1349 477
rect 1315 375 1349 409
rect 1315 307 1349 341
rect 1399 443 1433 477
rect 1399 375 1433 409
rect 1483 443 1517 477
rect 1483 375 1517 409
rect 1483 307 1517 341
rect 1567 375 1601 409
rect 1567 307 1601 341
rect 1651 443 1685 477
rect 1735 375 1769 409
rect 1735 307 1769 341
rect 1819 443 1853 477
rect 1819 375 1853 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 1003 497 1033 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 1359 497 1389 523
rect 1443 497 1473 523
rect 1527 497 1557 523
rect 1611 497 1641 523
rect 1695 497 1725 523
rect 1779 497 1809 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 79 249 277 265
rect 79 215 94 249
rect 128 215 162 249
rect 196 215 230 249
rect 264 215 277 249
rect 79 199 277 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 265 361 297
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 751 265 781 297
rect 835 265 865 297
rect 919 265 949 297
rect 1003 265 1033 297
rect 331 249 613 265
rect 331 215 361 249
rect 395 215 429 249
rect 463 215 497 249
rect 531 215 565 249
rect 599 215 613 249
rect 331 199 613 215
rect 655 249 709 265
rect 655 215 665 249
rect 699 215 709 249
rect 655 199 709 215
rect 751 249 1033 265
rect 751 215 836 249
rect 870 215 904 249
rect 938 215 972 249
rect 1006 215 1033 249
rect 751 199 1033 215
rect 331 177 361 199
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 751 177 781 199
rect 835 177 865 199
rect 919 177 949 199
rect 1003 177 1033 199
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 1359 265 1389 297
rect 1443 265 1473 297
rect 1191 249 1473 265
rect 1191 215 1210 249
rect 1244 215 1278 249
rect 1312 215 1346 249
rect 1380 215 1414 249
rect 1448 215 1473 249
rect 1191 199 1473 215
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 1359 177 1389 199
rect 1443 177 1473 199
rect 1527 265 1557 297
rect 1611 265 1641 297
rect 1695 265 1725 297
rect 1779 265 1809 297
rect 1527 249 1809 265
rect 1527 215 1550 249
rect 1584 215 1618 249
rect 1652 215 1686 249
rect 1720 215 1754 249
rect 1788 215 1809 249
rect 1527 199 1809 215
rect 1527 177 1557 199
rect 1611 177 1641 199
rect 1695 177 1725 199
rect 1779 177 1809 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 751 21 781 47
rect 835 21 865 47
rect 919 21 949 47
rect 1003 21 1033 47
rect 1191 21 1221 47
rect 1275 21 1305 47
rect 1359 21 1389 47
rect 1443 21 1473 47
rect 1527 21 1557 47
rect 1611 21 1641 47
rect 1695 21 1725 47
rect 1779 21 1809 47
<< polycont >>
rect 94 215 128 249
rect 162 215 196 249
rect 230 215 264 249
rect 361 215 395 249
rect 429 215 463 249
rect 497 215 531 249
rect 565 215 599 249
rect 665 215 699 249
rect 836 215 870 249
rect 904 215 938 249
rect 972 215 1006 249
rect 1210 215 1244 249
rect 1278 215 1312 249
rect 1346 215 1380 249
rect 1414 215 1448 249
rect 1550 215 1584 249
rect 1618 215 1652 249
rect 1686 215 1720 249
rect 1754 215 1788 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 483 85 493
rect 17 449 35 483
rect 69 449 85 483
rect 17 415 85 449
rect 17 381 35 415
rect 69 381 85 415
rect 17 347 85 381
rect 119 477 161 527
rect 153 443 161 477
rect 119 409 161 443
rect 153 375 161 409
rect 119 359 161 375
rect 195 477 243 493
rect 195 443 203 477
rect 237 443 243 477
rect 195 409 243 443
rect 279 477 329 527
rect 279 443 287 477
rect 321 443 329 477
rect 279 427 329 443
rect 363 477 413 493
rect 363 443 371 477
rect 405 443 413 477
rect 195 375 203 409
rect 237 393 243 409
rect 363 409 413 443
rect 447 477 497 527
rect 447 443 455 477
rect 489 443 497 477
rect 447 427 497 443
rect 531 477 581 493
rect 531 443 539 477
rect 573 443 581 477
rect 363 393 371 409
rect 237 375 371 393
rect 405 393 413 409
rect 531 409 581 443
rect 615 477 665 527
rect 615 443 623 477
rect 657 443 665 477
rect 615 427 665 443
rect 699 483 1093 493
rect 699 477 1043 483
rect 699 443 707 477
rect 741 459 875 477
rect 741 443 749 459
rect 531 393 539 409
rect 405 375 539 393
rect 573 393 581 409
rect 699 409 749 443
rect 867 443 875 459
rect 909 459 1043 477
rect 909 443 915 459
rect 699 393 707 409
rect 573 375 707 393
rect 741 375 749 409
rect 195 359 749 375
rect 783 409 833 425
rect 783 375 791 409
rect 825 375 833 409
rect 17 313 35 347
rect 69 325 85 347
rect 195 341 243 359
rect 195 325 203 341
rect 69 313 203 325
rect 17 307 203 313
rect 237 307 243 341
rect 783 341 833 375
rect 867 409 915 443
rect 1027 449 1043 459
rect 1077 449 1093 483
rect 867 375 875 409
rect 909 375 915 409
rect 867 359 915 375
rect 949 409 993 425
rect 949 375 959 409
rect 783 323 791 341
rect 17 291 243 307
rect 277 289 715 323
rect 277 257 311 289
rect 20 249 311 257
rect 20 215 94 249
rect 128 215 162 249
rect 196 215 230 249
rect 264 215 311 249
rect 345 249 615 255
rect 345 215 361 249
rect 395 215 429 249
rect 463 215 497 249
rect 531 215 565 249
rect 599 215 615 249
rect 649 249 715 289
rect 649 215 665 249
rect 699 215 715 249
rect 749 307 791 323
rect 825 323 833 341
rect 949 341 993 375
rect 949 323 959 341
rect 825 307 959 323
rect 749 283 993 307
rect 1027 415 1093 449
rect 1027 381 1043 415
rect 1077 381 1093 415
rect 1027 347 1093 381
rect 1027 313 1043 347
rect 1077 313 1093 347
rect 1027 291 1093 313
rect 1131 483 1197 493
rect 1131 449 1147 483
rect 1181 449 1197 483
rect 1131 415 1197 449
rect 1131 381 1147 415
rect 1181 381 1197 415
rect 1131 347 1197 381
rect 1231 477 1273 527
rect 1265 443 1273 477
rect 1231 409 1273 443
rect 1265 375 1273 409
rect 1231 359 1273 375
rect 1308 477 1356 493
rect 1308 443 1315 477
rect 1349 443 1356 477
rect 1308 409 1356 443
rect 1308 375 1315 409
rect 1349 375 1356 409
rect 1131 313 1147 347
rect 1181 325 1197 347
rect 1308 341 1356 375
rect 1391 477 1441 527
rect 1391 443 1399 477
rect 1433 443 1441 477
rect 1391 409 1441 443
rect 1391 375 1399 409
rect 1433 375 1441 409
rect 1391 359 1441 375
rect 1475 477 1862 493
rect 1475 443 1483 477
rect 1517 459 1651 477
rect 1517 443 1525 459
rect 1475 409 1525 443
rect 1643 443 1651 459
rect 1685 459 1819 477
rect 1685 443 1693 459
rect 1475 375 1483 409
rect 1517 375 1525 409
rect 1308 325 1315 341
rect 1181 313 1315 325
rect 1131 307 1315 313
rect 1349 325 1356 341
rect 1475 341 1525 375
rect 1475 325 1483 341
rect 1349 307 1483 325
rect 1517 307 1525 341
rect 1131 291 1525 307
rect 1559 409 1609 425
rect 1559 375 1567 409
rect 1601 375 1609 409
rect 1559 341 1609 375
rect 1643 359 1693 443
rect 1812 443 1819 459
rect 1853 443 1862 477
rect 1727 409 1777 425
rect 1727 375 1735 409
rect 1769 375 1777 409
rect 1559 307 1567 341
rect 1601 325 1609 341
rect 1727 341 1777 375
rect 1812 409 1862 443
rect 1812 375 1819 409
rect 1853 375 1862 409
rect 1812 359 1862 375
rect 1727 325 1735 341
rect 1601 307 1735 325
rect 1769 325 1777 341
rect 1769 307 1915 325
rect 1559 291 1915 307
rect 749 181 783 283
rect 1189 249 1464 255
rect 817 215 836 249
rect 870 215 904 249
rect 938 215 972 249
rect 1006 215 1145 249
rect 1189 215 1210 249
rect 1244 215 1278 249
rect 1312 215 1346 249
rect 1380 215 1414 249
rect 1448 215 1464 249
rect 1519 249 1809 255
rect 1519 215 1550 249
rect 1584 215 1618 249
rect 1652 215 1686 249
rect 1720 215 1754 249
rect 1788 215 1809 249
rect 1111 181 1145 215
rect 1843 181 1915 291
rect 35 163 69 179
rect 35 95 69 129
rect 35 17 69 61
rect 103 163 321 181
rect 103 129 119 163
rect 153 145 287 163
rect 153 129 169 145
rect 103 95 169 129
rect 271 129 287 145
rect 355 163 1009 181
rect 355 129 371 163
rect 405 129 539 163
rect 573 145 791 163
rect 573 129 599 145
rect 775 129 791 145
rect 825 145 959 163
rect 825 129 841 145
rect 103 61 119 95
rect 153 61 169 95
rect 103 51 169 61
rect 203 95 237 111
rect 203 17 237 61
rect 271 95 321 129
rect 707 95 741 111
rect 271 61 287 95
rect 321 61 455 95
rect 489 61 623 95
rect 657 61 673 95
rect 271 51 673 61
rect 707 17 741 61
rect 775 95 841 129
rect 943 129 959 145
rect 993 129 1009 163
rect 1111 163 1915 181
rect 1111 147 1231 163
rect 775 61 791 95
rect 825 61 841 95
rect 775 55 841 61
rect 875 95 909 111
rect 875 17 909 61
rect 943 95 1009 129
rect 1215 129 1231 147
rect 1265 145 1399 163
rect 1265 129 1281 145
rect 943 61 959 95
rect 993 61 1009 95
rect 943 55 1009 61
rect 1043 95 1181 111
rect 1077 61 1147 95
rect 1043 17 1181 61
rect 1215 95 1281 129
rect 1383 129 1399 145
rect 1433 145 1567 163
rect 1433 129 1449 145
rect 1215 61 1231 95
rect 1265 61 1281 95
rect 1215 51 1281 61
rect 1315 95 1349 111
rect 1315 17 1349 61
rect 1383 95 1449 129
rect 1551 129 1567 145
rect 1601 145 1735 163
rect 1601 129 1617 145
rect 1383 61 1399 95
rect 1433 61 1449 95
rect 1383 51 1449 61
rect 1483 95 1517 111
rect 1483 17 1517 61
rect 1551 95 1617 129
rect 1719 129 1735 145
rect 1769 147 1915 163
rect 1769 129 1785 147
rect 1551 61 1567 95
rect 1601 61 1617 95
rect 1551 51 1617 61
rect 1651 95 1685 111
rect 1651 17 1685 61
rect 1719 95 1785 129
rect 1719 61 1735 95
rect 1769 61 1785 95
rect 1719 51 1785 61
rect 1819 95 1853 111
rect 1819 17 1853 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 950 289 984 323 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 1598 221 1632 255 0 FreeSans 400 180 0 0 A2_N
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 400 180 0 0 B2
port 4 nsew signal input
flabel locali s 1322 221 1356 255 0 FreeSans 400 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a2bb2oi_4
rlabel metal1 s 0 -48 1932 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 3976018
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3961776
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 48.300 0.000 
<< end >>
