/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/capacitors/sky130_fd_pr__model__cap_var.model.spice