magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 106 157 584 203
rect 1 21 735 157
rect 30 -17 64 21
<< scnmos >>
rect 81 47 111 131
rect 194 47 244 177
rect 408 47 458 177
rect 580 47 610 131
<< scpmoshvt >>
rect 81 297 111 497
rect 194 333 244 497
rect 408 333 458 497
rect 580 297 610 497
<< ndiff >>
rect 132 131 194 177
rect 27 101 81 131
rect 27 67 36 101
rect 70 67 81 101
rect 27 47 81 67
rect 111 97 194 131
rect 111 63 132 97
rect 166 63 194 97
rect 111 47 194 63
rect 244 97 297 177
rect 244 63 255 97
rect 289 63 297 97
rect 244 47 297 63
rect 355 101 408 177
rect 355 67 363 101
rect 397 67 408 101
rect 355 47 408 67
rect 458 131 558 177
rect 458 97 580 131
rect 458 63 519 97
rect 553 63 580 97
rect 458 47 580 63
rect 610 97 709 131
rect 610 63 621 97
rect 655 63 709 97
rect 610 47 709 63
<< pdiff >>
rect 27 484 81 497
rect 27 450 36 484
rect 70 450 81 484
rect 27 416 81 450
rect 27 382 36 416
rect 70 382 81 416
rect 27 297 81 382
rect 111 484 194 497
rect 111 450 135 484
rect 169 450 194 484
rect 111 416 194 450
rect 111 382 135 416
rect 169 382 194 416
rect 111 333 194 382
rect 244 484 297 497
rect 244 450 255 484
rect 289 450 297 484
rect 244 416 297 450
rect 244 382 255 416
rect 289 382 297 416
rect 244 333 297 382
rect 355 477 408 497
rect 355 443 363 477
rect 397 443 408 477
rect 355 409 408 443
rect 355 375 363 409
rect 397 375 408 409
rect 355 333 408 375
rect 458 484 580 497
rect 458 450 519 484
rect 553 450 580 484
rect 458 416 580 450
rect 458 382 519 416
rect 553 382 580 416
rect 458 333 580 382
rect 111 297 161 333
rect 530 297 580 333
rect 610 477 709 497
rect 610 443 621 477
rect 655 443 709 477
rect 610 409 709 443
rect 610 375 621 409
rect 655 375 709 409
rect 610 297 709 375
<< ndiffc >>
rect 36 67 70 101
rect 132 63 166 97
rect 255 63 289 97
rect 363 67 397 101
rect 519 63 553 97
rect 621 63 655 97
<< pdiffc >>
rect 36 450 70 484
rect 36 382 70 416
rect 135 450 169 484
rect 135 382 169 416
rect 255 450 289 484
rect 255 382 289 416
rect 363 443 397 477
rect 363 375 397 409
rect 519 450 553 484
rect 519 382 553 416
rect 621 443 655 477
rect 621 375 655 409
<< poly >>
rect 81 497 111 523
rect 194 497 244 523
rect 408 497 458 523
rect 580 497 610 523
rect 81 261 111 297
rect 31 249 111 261
rect 194 259 244 333
rect 408 259 458 333
rect 580 265 610 297
rect 31 215 47 249
rect 81 215 111 249
rect 31 203 111 215
rect 155 249 244 259
rect 155 215 171 249
rect 205 215 244 249
rect 155 205 244 215
rect 350 249 484 259
rect 350 215 366 249
rect 400 215 434 249
rect 468 215 484 249
rect 350 205 484 215
rect 556 249 610 265
rect 556 215 566 249
rect 600 215 610 249
rect 81 131 111 203
rect 194 177 244 205
rect 408 177 458 205
rect 556 199 610 215
rect 580 131 610 199
rect 81 21 111 47
rect 194 21 244 47
rect 408 21 458 47
rect 580 21 610 47
<< polycont >>
rect 47 215 81 249
rect 171 215 205 249
rect 366 215 400 249
rect 434 215 468 249
rect 566 215 600 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 484 86 493
rect 17 450 36 484
rect 70 450 86 484
rect 17 416 86 450
rect 17 382 36 416
rect 70 382 86 416
rect 17 332 86 382
rect 120 484 185 527
rect 120 450 135 484
rect 169 450 185 484
rect 120 416 185 450
rect 120 382 135 416
rect 169 382 185 416
rect 120 366 185 382
rect 239 484 329 493
rect 239 450 255 484
rect 289 450 329 484
rect 239 416 329 450
rect 239 382 255 416
rect 289 382 329 416
rect 239 358 329 382
rect 17 298 201 332
rect 17 249 97 264
rect 17 215 47 249
rect 81 215 97 249
rect 131 259 201 298
rect 131 249 221 259
rect 131 215 171 249
rect 205 215 221 249
rect 131 205 221 215
rect 294 250 329 358
rect 363 477 413 493
rect 397 443 413 477
rect 363 409 413 443
rect 397 375 413 409
rect 363 333 413 375
rect 447 484 569 527
rect 447 450 519 484
rect 553 450 569 484
rect 447 416 569 450
rect 447 382 519 416
rect 553 382 569 416
rect 447 367 569 382
rect 607 477 719 493
rect 607 443 621 477
rect 655 443 719 477
rect 607 409 719 443
rect 607 375 621 409
rect 655 375 719 409
rect 363 299 553 333
rect 607 313 719 375
rect 519 265 553 299
rect 294 249 484 250
rect 294 215 366 249
rect 400 215 434 249
rect 468 215 484 249
rect 519 249 610 265
rect 519 215 566 249
rect 600 215 610 249
rect 131 181 201 205
rect 17 147 201 181
rect 294 171 329 215
rect 519 198 610 215
rect 519 181 553 198
rect 17 101 82 147
rect 17 67 36 101
rect 70 67 82 101
rect 17 51 82 67
rect 116 97 182 113
rect 116 63 132 97
rect 166 63 182 97
rect 116 17 182 63
rect 235 97 329 171
rect 235 63 255 97
rect 289 63 329 97
rect 235 51 329 63
rect 363 147 553 181
rect 363 101 413 147
rect 646 128 719 313
rect 397 67 413 101
rect 363 51 413 67
rect 448 97 569 113
rect 448 63 519 97
rect 553 63 569 97
rect 448 17 569 63
rect 603 97 719 128
rect 603 63 621 97
rect 655 63 719 97
rect 603 51 719 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 672 425 706 459 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 672 357 706 391 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 672 289 706 323 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 672 221 706 255 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 672 153 706 187 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 672 85 706 119 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 clkdlybuf4s25_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3261692
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3255572
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
