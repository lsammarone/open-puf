magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< locali >>
rect 191 1160 195 1194
rect 229 1160 267 1194
rect 301 1160 339 1194
rect 373 1160 411 1194
rect 445 1160 483 1194
rect 517 1160 555 1194
rect 589 1160 627 1194
rect 661 1160 665 1194
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 774 1020 808 1058
rect 774 948 808 986
rect 774 876 808 914
rect 774 804 808 842
rect 774 732 808 770
rect 774 660 808 698
rect 774 588 808 626
rect 774 516 808 554
rect 774 444 808 482
rect 774 372 808 410
rect 774 300 808 338
rect 774 228 808 266
rect 774 122 808 194
rect 191 20 195 54
rect 229 20 267 54
rect 301 20 339 54
rect 373 20 411 54
rect 445 20 483 54
rect 517 20 555 54
rect 589 20 627 54
rect 661 20 665 54
<< viali >>
rect 195 1160 229 1194
rect 267 1160 301 1194
rect 339 1160 373 1194
rect 411 1160 445 1194
rect 483 1160 517 1194
rect 555 1160 589 1194
rect 627 1160 661 1194
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 774 1058 808 1092
rect 774 986 808 1020
rect 774 914 808 948
rect 774 842 808 876
rect 774 770 808 804
rect 774 698 808 732
rect 774 626 808 660
rect 774 554 808 588
rect 774 482 808 516
rect 774 410 808 444
rect 774 338 808 372
rect 774 266 808 300
rect 774 194 808 228
rect 195 20 229 54
rect 267 20 301 54
rect 339 20 373 54
rect 411 20 445 54
rect 483 20 517 54
rect 555 20 589 54
rect 627 20 661 54
<< obsli1 >>
rect 159 98 193 1116
rect 285 98 319 1116
rect 411 98 445 1116
rect 537 98 571 1116
rect 663 98 697 1116
<< metal1 >>
rect 183 1194 673 1214
rect 183 1160 195 1194
rect 229 1160 267 1194
rect 301 1160 339 1194
rect 373 1160 411 1194
rect 445 1160 483 1194
rect 517 1160 555 1194
rect 589 1160 627 1194
rect 661 1160 673 1194
rect 183 1148 673 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 762 1092 820 1104
rect 762 1058 774 1092
rect 808 1058 820 1092
rect 762 1020 820 1058
rect 762 986 774 1020
rect 808 986 820 1020
rect 762 948 820 986
rect 762 914 774 948
rect 808 914 820 948
rect 762 876 820 914
rect 762 842 774 876
rect 808 842 820 876
rect 762 804 820 842
rect 762 770 774 804
rect 808 770 820 804
rect 762 732 820 770
rect 762 698 774 732
rect 808 698 820 732
rect 762 660 820 698
rect 762 626 774 660
rect 808 626 820 660
rect 762 588 820 626
rect 762 554 774 588
rect 808 554 820 588
rect 762 516 820 554
rect 762 482 774 516
rect 808 482 820 516
rect 762 444 820 482
rect 762 410 774 444
rect 808 410 820 444
rect 762 372 820 410
rect 762 338 774 372
rect 808 338 820 372
rect 762 300 820 338
rect 762 266 774 300
rect 808 266 820 300
rect 762 228 820 266
rect 762 194 774 228
rect 808 194 820 228
rect 762 110 820 194
rect 183 54 673 66
rect 183 20 195 54
rect 229 20 267 54
rect 301 20 339 54
rect 373 20 411 54
rect 445 20 483 54
rect 517 20 555 54
rect 589 20 627 54
rect 661 20 673 54
rect 183 0 673 20
<< obsm1 >>
rect 150 110 202 1104
rect 276 110 328 1104
rect 402 110 454 1104
rect 528 110 580 1104
rect 654 110 706 1104
<< metal2 >>
rect 10 632 846 1104
rect 10 110 846 582
<< labels >>
rlabel viali s 774 1058 808 1092 6 BULK
port 1 nsew
rlabel viali s 774 986 808 1020 6 BULK
port 1 nsew
rlabel viali s 774 914 808 948 6 BULK
port 1 nsew
rlabel viali s 774 842 808 876 6 BULK
port 1 nsew
rlabel viali s 774 770 808 804 6 BULK
port 1 nsew
rlabel viali s 774 698 808 732 6 BULK
port 1 nsew
rlabel viali s 774 626 808 660 6 BULK
port 1 nsew
rlabel viali s 774 554 808 588 6 BULK
port 1 nsew
rlabel viali s 774 482 808 516 6 BULK
port 1 nsew
rlabel viali s 774 410 808 444 6 BULK
port 1 nsew
rlabel viali s 774 338 808 372 6 BULK
port 1 nsew
rlabel viali s 774 266 808 300 6 BULK
port 1 nsew
rlabel viali s 774 194 808 228 6 BULK
port 1 nsew
rlabel viali s 48 1058 82 1092 6 BULK
port 1 nsew
rlabel viali s 48 986 82 1020 6 BULK
port 1 nsew
rlabel viali s 48 914 82 948 6 BULK
port 1 nsew
rlabel viali s 48 842 82 876 6 BULK
port 1 nsew
rlabel viali s 48 770 82 804 6 BULK
port 1 nsew
rlabel viali s 48 698 82 732 6 BULK
port 1 nsew
rlabel viali s 48 626 82 660 6 BULK
port 1 nsew
rlabel viali s 48 554 82 588 6 BULK
port 1 nsew
rlabel viali s 48 482 82 516 6 BULK
port 1 nsew
rlabel viali s 48 410 82 444 6 BULK
port 1 nsew
rlabel viali s 48 338 82 372 6 BULK
port 1 nsew
rlabel viali s 48 266 82 300 6 BULK
port 1 nsew
rlabel viali s 48 194 82 228 6 BULK
port 1 nsew
rlabel locali s 774 122 808 1092 6 BULK
port 1 nsew
rlabel locali s 48 122 82 1092 6 BULK
port 1 nsew
rlabel metal1 s 762 110 820 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 846 1104 6 DRAIN
port 2 nsew
rlabel viali s 627 1160 661 1194 6 GATE
port 3 nsew
rlabel viali s 627 20 661 54 6 GATE
port 3 nsew
rlabel viali s 555 1160 589 1194 6 GATE
port 3 nsew
rlabel viali s 555 20 589 54 6 GATE
port 3 nsew
rlabel viali s 483 1160 517 1194 6 GATE
port 3 nsew
rlabel viali s 483 20 517 54 6 GATE
port 3 nsew
rlabel viali s 411 1160 445 1194 6 GATE
port 3 nsew
rlabel viali s 411 20 445 54 6 GATE
port 3 nsew
rlabel viali s 339 1160 373 1194 6 GATE
port 3 nsew
rlabel viali s 339 20 373 54 6 GATE
port 3 nsew
rlabel viali s 267 1160 301 1194 6 GATE
port 3 nsew
rlabel viali s 267 20 301 54 6 GATE
port 3 nsew
rlabel viali s 195 1160 229 1194 6 GATE
port 3 nsew
rlabel viali s 195 20 229 54 6 GATE
port 3 nsew
rlabel locali s 191 1160 665 1194 6 GATE
port 3 nsew
rlabel locali s 191 20 665 54 6 GATE
port 3 nsew
rlabel metal1 s 183 1148 673 1214 6 GATE
port 3 nsew
rlabel metal1 s 183 0 673 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 846 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 856 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10422700
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10400732
<< end >>
