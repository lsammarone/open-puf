magic
tech sky130A
magscale 1 2
timestamp 1656544606
<< nwell >>
rect -406 636 388 882
rect -574 -766 -356 -198
rect -62 -278 382 -258
rect -62 -444 416 -278
rect 690 -416 1048 -200
rect -62 -452 434 -444
rect 202 -594 434 -452
<< locali >>
rect 92 452 142 456
rect 460 452 526 484
rect 92 446 526 452
rect 92 406 98 446
rect 136 436 526 446
rect 136 406 580 436
rect 92 402 580 406
rect 92 400 142 402
rect 276 -596 334 -590
rect 276 -636 282 -596
rect 320 -602 334 -596
rect 464 -602 530 -522
rect 320 -636 588 -602
rect 276 -642 334 -636
rect -384 -766 -288 -764
rect -384 -806 -374 -766
rect -336 -806 -288 -766
rect -384 -810 -288 -806
rect -176 -768 10 -764
rect -176 -808 -64 -768
rect -26 -808 10 -768
rect -176 -810 10 -808
<< viali >>
rect 98 406 136 446
rect -342 282 -304 322
rect -164 282 -124 318
rect -252 180 -208 224
rect -248 -102 -204 -58
rect -342 -198 -304 -158
rect -164 -198 -126 -158
rect 1044 -202 1082 -162
rect 1218 -394 1256 -354
rect 282 -636 320 -596
rect -374 -806 -336 -766
rect -64 -808 -26 -768
rect 1040 -818 1078 -778
rect 80 -886 118 -846
<< metal1 >>
rect -574 1120 1322 1192
rect -574 1004 961 1120
rect 1269 1004 1322 1120
rect -574 938 1322 1004
rect -366 634 -300 938
rect 92 456 146 458
rect -16 454 146 456
rect -16 402 -6 454
rect 46 446 146 454
rect 46 406 98 446
rect 136 406 146 446
rect 46 402 146 406
rect -16 400 146 402
rect 92 394 146 400
rect -178 338 -102 344
rect -428 330 -296 338
rect -428 274 -424 330
rect -368 322 -296 330
rect -368 282 -342 322
rect -304 282 -296 322
rect -368 274 -296 282
rect -178 282 -170 338
rect -114 332 -102 338
rect 258 342 406 350
rect -114 282 -60 332
rect -178 276 -60 282
rect 258 290 270 342
rect 322 290 406 342
rect 258 280 406 290
rect -428 266 -296 274
rect -266 230 94 234
rect -266 224 20 230
rect -266 180 -252 224
rect -208 180 20 224
rect -266 178 20 180
rect 72 178 94 230
rect -266 168 94 178
rect -118 34 432 110
rect -262 -52 98 -48
rect -262 -58 24 -52
rect -262 -102 -248 -58
rect -204 -102 24 -58
rect -262 -104 24 -102
rect 76 -104 98 -52
rect 850 -64 920 938
rect -262 -114 98 -104
rect 206 -140 920 -64
rect -428 -150 -296 -142
rect -428 -206 -424 -150
rect -368 -158 -296 -150
rect -368 -198 -342 -158
rect -304 -198 -296 -158
rect -368 -206 -296 -198
rect -428 -214 -296 -206
rect -178 -158 -96 -152
rect -178 -164 -164 -158
rect -126 -164 -96 -158
rect -178 -220 -168 -164
rect -112 -220 -96 -164
rect -178 -230 -96 -220
rect 206 -176 282 -140
rect 258 -228 282 -176
rect 800 -228 810 -176
rect 206 -434 282 -228
rect 792 -236 810 -228
rect 186 -448 282 -434
rect 186 -520 196 -448
rect 272 -520 282 -448
rect 186 -530 282 -520
rect 844 -454 920 -140
rect 986 -150 1096 -134
rect 986 -202 998 -150
rect 1050 -162 1096 -150
rect 1082 -202 1096 -162
rect 986 -210 1096 -202
rect 1202 -354 1298 -326
rect 1202 -394 1218 -354
rect 1256 -394 1298 -354
rect 1202 -404 1298 -394
rect 844 -530 1052 -454
rect 268 -596 334 -590
rect 268 -600 282 -596
rect -50 -632 282 -600
rect -50 -730 -18 -632
rect 268 -636 282 -632
rect 320 -636 334 -596
rect 268 -642 334 -636
rect -534 -766 -320 -754
rect -56 -760 -12 -730
rect -534 -818 -526 -766
rect -474 -806 -374 -766
rect -336 -806 -320 -766
rect -474 -818 -320 -806
rect -80 -762 -12 -760
rect -80 -814 -70 -762
rect -18 -814 -12 -762
rect 972 -772 1096 -756
rect -534 -826 -320 -818
rect 972 -824 982 -772
rect 1034 -778 1096 -772
rect 1034 -818 1040 -778
rect 1078 -818 1096 -778
rect 1034 -824 1096 -818
rect 972 -830 1096 -824
rect 68 -846 134 -834
rect 68 -886 80 -846
rect 118 -850 134 -846
rect 118 -886 500 -850
rect 68 -894 500 -886
rect -566 -970 1224 -930
rect -566 -1022 -264 -970
rect -212 -1022 -186 -970
rect -134 -1004 1224 -970
rect 1284 -1004 1322 -930
rect -134 -1022 961 -1004
rect -566 -1120 961 -1022
rect 1269 -1120 1322 -1004
rect -566 -1184 1322 -1120
<< via1 >>
rect 961 1004 1269 1120
rect -6 402 46 454
rect -424 274 -368 330
rect -170 318 -114 338
rect -170 282 -164 318
rect -164 282 -124 318
rect -124 282 -114 318
rect 270 290 322 342
rect 642 252 694 304
rect 20 178 72 230
rect 746 156 798 208
rect -266 38 -214 90
rect 24 -104 76 -52
rect 1112 28 1164 80
rect -424 -206 -368 -150
rect -168 -198 -164 -164
rect -164 -198 -126 -164
rect -126 -198 -112 -164
rect -168 -220 -112 -198
rect 206 -228 258 -176
rect 748 -228 800 -176
rect 392 -354 462 -286
rect 628 -340 686 -282
rect 196 -520 272 -448
rect 998 -162 1050 -150
rect 998 -202 1044 -162
rect 1044 -202 1050 -162
rect -526 -818 -474 -766
rect -70 -768 -18 -762
rect -70 -808 -64 -768
rect -64 -808 -26 -768
rect -26 -808 -18 -768
rect -70 -814 -18 -808
rect 982 -824 1034 -772
rect -264 -1022 -212 -970
rect -186 -1022 -134 -970
rect 961 -1120 1269 -1004
<< metal2 >>
rect 940 1120 1290 1134
rect 940 1004 961 1120
rect 1269 1004 1290 1120
rect 940 990 1290 1004
rect -566 816 1322 844
rect -436 332 -364 346
rect -124 344 -96 816
rect 528 512 600 520
rect -574 330 -364 332
rect -574 274 -424 330
rect -368 274 -364 330
rect -178 338 -96 344
rect -178 282 -170 338
rect -114 282 -96 338
rect -178 276 -96 282
rect -574 270 -364 274
rect -436 260 -364 270
rect -266 90 -214 110
rect -436 -144 -396 -134
rect -436 -148 -364 -144
rect -574 -150 -364 -148
rect -574 -206 -424 -150
rect -368 -206 -364 -150
rect -574 -210 -364 -206
rect -436 -220 -364 -210
rect -554 -754 -510 -398
rect -554 -766 -462 -754
rect -554 -818 -526 -766
rect -474 -818 -462 -766
rect -554 -826 -462 -818
rect -554 -1014 -510 -826
rect -266 -962 -214 38
rect -124 -152 -96 276
rect -178 -164 -96 -152
rect -178 -220 -168 -164
rect -112 -220 -96 -164
rect -178 -230 -96 -220
rect -36 454 46 464
rect -36 402 -6 454
rect 528 456 530 512
rect 590 456 600 512
rect 528 450 600 456
rect 1002 512 1082 528
rect 1002 456 1012 512
rect 1072 456 1082 512
rect 1002 450 1082 456
rect 1196 512 1272 522
rect 1196 456 1206 512
rect 1266 456 1272 512
rect -36 396 46 402
rect -36 -748 -8 396
rect 258 342 344 350
rect 258 290 270 342
rect 322 290 344 342
rect 20 230 30 236
rect 20 170 30 178
rect 96 170 122 236
rect 24 -52 34 -46
rect 24 -112 34 -104
rect 100 -112 126 -46
rect 316 -52 344 290
rect 622 304 710 306
rect 622 252 642 304
rect 694 252 710 304
rect 622 238 710 252
rect 384 232 470 236
rect 384 176 394 232
rect 454 176 470 232
rect 258 -108 270 -52
rect 330 -108 344 -52
rect 258 -112 344 -108
rect 206 -176 258 -166
rect 206 -448 258 -228
rect 442 -286 470 176
rect 622 182 638 238
rect 698 182 710 238
rect 622 172 710 182
rect 742 208 808 214
rect 742 156 746 208
rect 798 156 808 208
rect 742 144 808 156
rect 384 -354 392 -286
rect 462 -354 470 -286
rect 622 -48 696 -33
rect 622 -104 628 -48
rect 690 -104 696 -48
rect 622 -282 696 -104
rect 742 -170 796 144
rect 1022 -134 1050 450
rect 1196 448 1272 456
rect 1244 332 1272 448
rect 1244 270 1322 332
rect 1112 80 1164 116
rect 986 -150 1058 -134
rect 742 -176 808 -170
rect 742 -228 748 -176
rect 800 -228 808 -176
rect 986 -202 998 -150
rect 1050 -202 1058 -150
rect 986 -210 1058 -202
rect 742 -236 808 -228
rect 622 -340 628 -282
rect 686 -340 696 -282
rect 622 -344 696 -340
rect 384 -360 470 -354
rect 578 -440 614 -420
rect 188 -520 196 -448
rect 272 -520 282 -448
rect 596 -496 614 -440
rect 578 -506 614 -496
rect 996 -440 1076 -424
rect 996 -496 1006 -440
rect 1066 -496 1076 -440
rect 996 -502 1076 -496
rect 188 -530 282 -520
rect -80 -762 -8 -748
rect 1016 -754 1044 -502
rect -80 -814 -70 -762
rect -18 -814 -8 -762
rect 970 -772 1046 -754
rect 970 -824 982 -772
rect 1034 -824 1046 -772
rect 970 -832 1046 -824
rect -276 -970 -124 -962
rect -276 -1022 -264 -970
rect -212 -1022 -186 -970
rect -134 -1022 -124 -970
rect 1112 -990 1164 28
rect 1218 -210 1322 -148
rect 1218 -430 1246 -210
rect 1206 -440 1276 -430
rect 1266 -496 1276 -440
rect 1206 -506 1276 -496
rect -276 -1028 -124 -1022
rect 940 -1004 1290 -990
rect 940 -1120 961 -1004
rect 1269 -1120 1290 -1004
rect 940 -1134 1290 -1120
<< via2 >>
rect 967 1034 1023 1090
rect 1047 1034 1103 1090
rect 1127 1034 1183 1090
rect 1207 1034 1263 1090
rect 530 456 590 512
rect 1012 456 1072 512
rect 1206 456 1266 512
rect 30 230 96 236
rect 30 178 72 230
rect 72 178 96 230
rect 30 170 96 178
rect 34 -52 100 -46
rect 34 -104 76 -52
rect 76 -104 100 -52
rect 34 -112 100 -104
rect 394 176 454 232
rect 270 -108 330 -52
rect 638 182 698 238
rect 628 -104 690 -48
rect 536 -496 596 -440
rect 1006 -496 1066 -440
rect 1206 -496 1266 -440
rect 967 -1090 1023 -1034
rect 1047 -1090 1103 -1034
rect 1127 -1090 1183 -1034
rect 1207 -1090 1263 -1034
<< metal3 >>
rect -574 1090 1322 1192
rect -574 1034 967 1090
rect 1023 1034 1047 1090
rect 1103 1034 1127 1090
rect 1183 1034 1207 1090
rect 1263 1034 1322 1090
rect -574 938 1322 1034
rect 514 512 1278 520
rect 514 456 530 512
rect 590 456 1012 512
rect 1072 456 1206 512
rect 1266 456 1278 512
rect 514 450 1278 456
rect 10 237 162 250
rect 626 238 706 244
rect 626 237 638 238
rect 10 236 638 237
rect 10 170 30 236
rect 96 232 638 236
rect 96 176 394 232
rect 454 182 638 232
rect 698 237 706 238
rect 698 182 717 237
rect 454 176 717 182
rect 96 171 717 176
rect 96 170 162 171
rect 10 158 162 170
rect 14 -45 166 -32
rect 622 -45 696 -32
rect 14 -46 721 -45
rect 14 -112 34 -46
rect 100 -48 721 -46
rect 100 -52 628 -48
rect 100 -108 270 -52
rect 330 -104 628 -52
rect 690 -104 721 -48
rect 330 -108 721 -104
rect 100 -111 721 -108
rect 100 -112 166 -111
rect 14 -124 166 -112
rect 258 -118 344 -111
rect 526 -440 1276 -420
rect 526 -496 536 -440
rect 596 -496 1006 -440
rect 1066 -496 1206 -440
rect 1266 -496 1276 -440
rect 526 -506 1276 -496
rect -566 -1034 1322 -930
rect -566 -1090 967 -1034
rect 1023 -1090 1047 -1034
rect 1103 -1090 1127 -1034
rect 1183 -1090 1207 -1034
rect 1263 -1090 1322 -1034
rect -566 -1185 1322 -1090
use mux  mux_0
timestamp 1654402208
transform 1 0 432 0 1 146
box -54 -122 366 878
use mux  mux_1
timestamp 1654402208
transform 1 0 436 0 1 -892
box -54 -122 366 878
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0
timestamp 1654402208
transform 1 0 1008 0 1 -1027
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_1
timestamp 1654402208
transform 1 0 1008 0 -1 61
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1_0
timestamp 1654402208
transform 1 0 -90 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1#0  sky130_fd_sc_hd__inv_1_1
timestamp 1654402208
transform 1 0 -366 0 1 -1026
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0
timestamp 1654402208
transform 1 0 -366 0 1 62
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1654402208
transform 1 0 -366 0 -1 62
box -38 -48 314 592
<< labels >>
flabel metal2 -574 270 -424 332 1 FreeSans 800 0 0 0 IN1
port 1 n
flabel metal2 -554 -1014 -510 -818 1 FreeSans 800 0 0 0 C
port 2 n
flabel metal2 -566 816 1322 844 1 FreeSans 800 0 0 0 RESET
port 3 n
flabel metal3 -134 -1184 961 -930 1 FreeSans 800 0 0 0 VSS
port 4 n
flabel metal3 -574 938 967 1192 1 FreeSans 800 0 0 0 VDD
port 5 n
flabel metal2 1218 -210 1322 -148 1 FreeSans 800 0 0 0 OUT2
port 6 n
flabel metal1 1256 -404 1298 -326 1 FreeSans 800 0 0 0 buf_out
port 7 n
flabel metal2 1244 270 1322 332 1 FreeSans 800 0 0 0 OUT1
port 8 n
flabel metal2 -574 -210 -424 -148 1 FreeSans 800 0 0 0 IN2
port 9 n
<< end >>
