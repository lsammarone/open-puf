magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 157 275 203
rect 1 21 827 157
rect 27 -17 61 21
<< scnmos >>
rect 84 47 114 177
rect 168 47 198 177
rect 264 47 294 131
rect 357 47 387 131
rect 551 47 581 131
rect 635 47 665 131
rect 719 47 749 131
<< scpmoshvt >>
rect 84 297 114 497
rect 168 297 198 497
rect 265 369 295 497
rect 375 369 405 497
rect 547 369 577 497
rect 635 369 665 497
rect 719 369 749 497
<< ndiff >>
rect 27 159 84 177
rect 27 125 39 159
rect 73 125 84 159
rect 27 91 84 125
rect 27 57 39 91
rect 73 57 84 91
rect 27 47 84 57
rect 114 159 168 177
rect 114 125 124 159
rect 158 125 168 159
rect 114 91 168 125
rect 114 57 124 91
rect 158 57 168 91
rect 114 47 168 57
rect 198 131 249 177
rect 198 122 264 131
rect 198 88 213 122
rect 247 88 264 122
rect 198 47 264 88
rect 294 47 357 131
rect 387 113 439 131
rect 387 79 397 113
rect 431 79 439 113
rect 387 47 439 79
rect 499 114 551 131
rect 499 80 507 114
rect 541 80 551 114
rect 499 47 551 80
rect 581 114 635 131
rect 581 80 591 114
rect 625 80 635 114
rect 581 47 635 80
rect 665 95 719 131
rect 665 61 675 95
rect 709 61 719 95
rect 665 47 719 61
rect 749 104 801 131
rect 749 70 759 104
rect 793 70 801 104
rect 749 47 801 70
<< pdiff >>
rect 27 477 84 497
rect 27 443 39 477
rect 73 443 84 477
rect 27 409 84 443
rect 27 375 39 409
rect 73 375 84 409
rect 27 341 84 375
rect 27 307 39 341
rect 73 307 84 341
rect 27 297 84 307
rect 114 477 168 497
rect 114 443 124 477
rect 158 443 168 477
rect 114 409 168 443
rect 114 375 124 409
rect 158 375 168 409
rect 114 297 168 375
rect 198 481 265 497
rect 198 447 208 481
rect 242 447 265 481
rect 198 369 265 447
rect 295 369 375 497
rect 405 481 547 497
rect 405 447 456 481
rect 490 447 547 481
rect 405 369 547 447
rect 577 485 635 497
rect 577 451 587 485
rect 621 451 635 485
rect 577 417 635 451
rect 577 383 587 417
rect 621 383 635 417
rect 577 369 635 383
rect 665 369 719 497
rect 749 485 801 497
rect 749 451 759 485
rect 793 451 801 485
rect 749 417 801 451
rect 749 383 759 417
rect 793 383 801 417
rect 749 369 801 383
rect 198 297 250 369
rect 310 343 360 369
rect 310 309 318 343
rect 352 309 360 343
rect 310 297 360 309
<< ndiffc >>
rect 39 125 73 159
rect 39 57 73 91
rect 124 125 158 159
rect 124 57 158 91
rect 213 88 247 122
rect 397 79 431 113
rect 507 80 541 114
rect 591 80 625 114
rect 675 61 709 95
rect 759 70 793 104
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 124 443 158 477
rect 124 375 158 409
rect 208 447 242 481
rect 456 447 490 481
rect 587 451 621 485
rect 587 383 621 417
rect 759 451 793 485
rect 759 383 793 417
rect 318 309 352 343
<< poly >>
rect 84 497 114 523
rect 168 497 198 523
rect 265 497 295 523
rect 375 497 405 523
rect 547 497 577 523
rect 635 497 665 523
rect 719 497 749 523
rect 84 265 114 297
rect 168 265 198 297
rect 265 265 295 369
rect 84 249 219 265
rect 84 215 175 249
rect 209 215 219 249
rect 84 199 219 215
rect 261 249 315 265
rect 261 215 271 249
rect 305 215 315 249
rect 375 220 405 369
rect 547 337 577 369
rect 448 321 581 337
rect 448 287 458 321
rect 492 287 581 321
rect 448 271 581 287
rect 261 199 315 215
rect 357 204 415 220
rect 84 177 114 199
rect 168 177 198 199
rect 264 131 294 199
rect 357 170 371 204
rect 405 170 415 204
rect 357 154 415 170
rect 357 131 387 154
rect 551 131 581 271
rect 635 265 665 369
rect 719 265 749 369
rect 623 249 677 265
rect 623 215 633 249
rect 667 215 677 249
rect 623 199 677 215
rect 719 249 805 265
rect 719 215 756 249
rect 790 215 805 249
rect 719 199 805 215
rect 635 131 665 199
rect 719 131 749 199
rect 84 21 114 47
rect 168 21 198 47
rect 264 21 294 47
rect 357 21 387 47
rect 551 21 581 47
rect 635 21 665 47
rect 719 21 749 47
<< polycont >>
rect 175 215 209 249
rect 271 215 305 249
rect 458 287 492 321
rect 371 170 405 204
rect 633 215 667 249
rect 756 215 790 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 22 477 73 527
rect 22 443 39 477
rect 22 409 73 443
rect 22 375 39 409
rect 22 341 73 375
rect 22 307 39 341
rect 22 282 73 307
rect 107 477 158 493
rect 107 443 124 477
rect 192 481 258 527
rect 192 447 208 481
rect 242 447 258 481
rect 432 481 513 527
rect 746 485 809 527
rect 432 447 456 481
rect 490 447 513 481
rect 567 451 587 485
rect 621 451 637 485
rect 107 409 158 443
rect 567 417 637 451
rect 567 411 587 417
rect 107 375 124 409
rect 107 359 158 375
rect 220 383 587 411
rect 621 383 637 417
rect 220 377 637 383
rect 22 159 73 182
rect 22 125 39 159
rect 22 91 73 125
rect 22 57 39 91
rect 22 17 73 57
rect 107 165 141 359
rect 220 323 254 377
rect 175 289 254 323
rect 288 309 318 343
rect 352 321 492 343
rect 352 309 458 321
rect 288 299 458 309
rect 175 249 209 289
rect 439 287 458 299
rect 439 271 492 287
rect 526 299 637 377
rect 243 249 337 255
rect 243 215 271 249
rect 305 215 337 249
rect 175 199 209 215
rect 371 204 405 220
rect 303 170 371 181
rect 107 159 174 165
rect 107 125 124 159
rect 158 125 174 159
rect 303 154 405 170
rect 107 91 174 125
rect 107 57 124 91
rect 158 57 174 91
rect 107 51 174 57
rect 213 122 247 150
rect 213 17 247 88
rect 303 147 404 154
rect 303 76 347 147
rect 439 113 473 271
rect 526 249 560 299
rect 671 265 705 485
rect 746 451 759 485
rect 793 451 809 485
rect 746 417 809 451
rect 746 383 759 417
rect 793 383 809 417
rect 746 363 809 383
rect 522 215 560 249
rect 594 249 705 265
rect 594 215 633 249
rect 667 215 705 249
rect 740 249 809 329
rect 740 215 756 249
rect 790 215 809 249
rect 522 138 556 215
rect 381 79 397 113
rect 431 79 473 113
rect 507 114 556 138
rect 541 80 556 114
rect 507 64 556 80
rect 591 145 809 181
rect 591 114 637 145
rect 625 80 637 114
rect 591 64 637 80
rect 675 95 709 111
rect 743 104 809 145
rect 743 70 759 104
rect 793 70 809 104
rect 743 64 809 70
rect 675 17 709 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 303 221 337 255 0 FreeSans 400 0 0 0 A1_N
port 1 nsew signal input
flabel locali s 119 425 153 459 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 303 85 337 119 0 FreeSans 400 0 0 0 A2_N
port 2 nsew signal input
flabel locali s 671 289 705 323 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 763 221 797 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel pwell s 27 -17 61 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 27 527 61 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 27 -17 61 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 27 527 61 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o2bb2a_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1242556
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1235508
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.140 0.000 
<< end >>
