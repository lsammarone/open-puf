.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

