magic
tech sky130A
magscale 1 2
timestamp 1654151215
<< error_s >>
rect 4610 5343 4683 5354
rect 19739 5352 19799 5355
rect 19739 5349 19807 5352
rect 19739 5347 19799 5349
rect 19799 5291 19803 5347
<< locali >>
rect 4626 5009 4668 5012
rect 2742 5005 2784 5008
rect 2742 4971 2746 5005
rect 2780 4971 2784 5005
rect 2742 4968 2784 4971
rect 4626 4975 4630 5009
rect 4664 4975 4668 5009
rect 19724 5009 19766 5012
rect 4626 4972 4668 4975
rect 17840 5005 17882 5008
rect 17840 4971 17844 5005
rect 17878 4971 17882 5005
rect 17840 4968 17882 4971
rect 19724 4975 19728 5009
rect 19762 4975 19766 5009
rect 19724 4972 19766 4975
<< viali >>
rect 2268 5068 2302 5102
rect 2381 5068 2415 5102
rect 2494 5068 2528 5102
rect 2607 5068 2641 5102
rect 2720 5068 2754 5102
rect 2833 5068 2867 5102
rect 2946 5068 2980 5102
rect 3062 5068 3096 5102
rect 3166 5068 3200 5102
rect 4022 5068 4056 5102
rect 4141 5068 4175 5102
rect 4260 5068 4294 5102
rect 4379 5068 4413 5102
rect 4498 5068 4532 5102
rect 4617 5068 4651 5102
rect 4736 5068 4770 5102
rect 17434 5068 17468 5102
rect 17531 5068 17565 5102
rect 17628 5068 17662 5102
rect 17725 5068 17759 5102
rect 17822 5068 17856 5102
rect 17919 5068 17953 5102
rect 18016 5068 18050 5102
rect 18113 5068 18147 5102
rect 18264 5068 18298 5102
rect 19120 5068 19154 5102
rect 19228 5068 19262 5102
rect 19336 5068 19370 5102
rect 19444 5068 19478 5102
rect 19552 5068 19586 5102
rect 19660 5068 19694 5102
rect 19768 5068 19802 5102
rect 19876 5068 19910 5102
rect 2245 4973 2279 5007
rect 2411 4971 2445 5005
rect 2575 4969 2609 5003
rect 2746 4971 2780 5005
rect 2915 4967 2949 5001
rect 3084 4966 3118 5000
rect 3250 4972 3284 5006
rect 3420 4974 3454 5008
rect 4134 4971 4168 5005
rect 4294 4971 4328 5005
rect 4461 4965 4495 4999
rect 4630 4975 4664 5009
rect 4794 4962 4828 4996
rect 4964 4968 4998 5002
rect 5134 4970 5168 5004
rect 5293 4972 5327 5006
rect 17343 4967 17377 5001
rect 17506 4962 17540 4996
rect 17679 4966 17713 5000
rect 17844 4971 17878 5005
rect 18011 4958 18045 4992
rect 18179 4956 18213 4990
rect 18349 4965 18383 4999
rect 19222 4966 19256 5000
rect 19395 4967 19429 5001
rect 19557 4972 19591 5006
rect 19728 4975 19762 5009
rect 19897 4961 19931 4995
rect 20062 4961 20096 4995
rect 20232 4959 20266 4993
rect 20395 4963 20429 4997
<< metal1 >>
rect 3584 5274 3994 5367
rect 18682 5274 19103 5365
rect 3688 5108 3894 5220
rect 18800 5108 18998 5222
rect 2218 5102 5022 5108
rect 2218 5068 2268 5102
rect 2302 5068 2381 5102
rect 2415 5068 2494 5102
rect 2528 5068 2607 5102
rect 2641 5068 2720 5102
rect 2754 5068 2833 5102
rect 2867 5068 2946 5102
rect 2980 5068 3062 5102
rect 3096 5068 3166 5102
rect 3200 5068 4022 5102
rect 4056 5068 4141 5102
rect 4175 5068 4260 5102
rect 4294 5068 4379 5102
rect 4413 5068 4498 5102
rect 4532 5068 4617 5102
rect 4651 5068 4736 5102
rect 4770 5068 5022 5102
rect 2218 5062 5022 5068
rect 17369 5102 20060 5108
rect 17369 5068 17434 5102
rect 17468 5068 17531 5102
rect 17565 5068 17628 5102
rect 17662 5068 17725 5102
rect 17759 5068 17822 5102
rect 17856 5068 17919 5102
rect 17953 5068 18016 5102
rect 18050 5068 18113 5102
rect 18147 5068 18264 5102
rect 18298 5068 19120 5102
rect 19154 5068 19228 5102
rect 19262 5068 19336 5102
rect 19370 5068 19444 5102
rect 19478 5068 19552 5102
rect 19586 5068 19660 5102
rect 19694 5068 19768 5102
rect 19802 5068 19876 5102
rect 19910 5068 20060 5102
rect 17369 5062 20060 5068
rect 2230 5008 3467 5020
rect 2230 5007 3420 5008
rect 2230 4973 2245 5007
rect 2279 5006 3420 5007
rect 2279 5005 3250 5006
rect 2279 5002 2411 5005
rect 2445 5004 2746 5005
rect 2780 5004 3250 5005
rect 2445 5003 2740 5004
rect 2445 5002 2575 5003
rect 2279 4973 2282 5002
rect 2230 4950 2282 4973
rect 2334 4950 2389 5002
rect 2445 4971 2495 5002
rect 2441 4950 2495 4971
rect 2547 4969 2575 5002
rect 2609 5002 2740 5003
rect 2609 4969 2611 5002
rect 2547 4950 2611 4969
rect 2663 4952 2740 5002
rect 2792 5003 3250 5004
rect 3284 5003 3420 5006
rect 2792 4952 2874 5003
rect 2926 5001 2991 5003
rect 2949 4967 2991 5001
rect 2663 4951 2874 4952
rect 2926 4951 2991 4967
rect 3043 5000 3096 5003
rect 3043 4966 3084 5000
rect 3043 4951 3096 4966
rect 3148 4951 3202 5003
rect 3284 4972 3299 5003
rect 3254 4951 3299 4972
rect 3351 4951 3396 5003
rect 3454 4974 3467 5008
rect 3448 4951 3467 4974
rect 2663 4950 3467 4951
rect 2230 4936 3467 4950
rect 4120 5009 5346 5018
rect 4120 5005 4630 5009
rect 4120 4971 4134 5005
rect 4168 4999 4294 5005
rect 4328 5002 4630 5005
rect 4664 5006 5346 5009
rect 4664 5004 5293 5006
rect 4664 5002 5134 5004
rect 4328 4999 4622 5002
rect 4168 4971 4171 4999
rect 4120 4947 4171 4971
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4965 4461 4999
rect 4495 4965 4500 4999
rect 4436 4947 4500 4965
rect 4552 4950 4622 4999
rect 4674 5001 4964 5002
rect 4681 5000 4964 5001
rect 4998 5000 5134 5002
rect 5168 5000 5293 5004
rect 5327 5000 5346 5006
rect 4552 4949 4629 4950
rect 4681 4949 4763 5000
rect 4815 4996 4880 5000
rect 4828 4962 4880 4996
rect 4552 4948 4763 4949
rect 4815 4948 4880 4962
rect 4932 4968 4964 5000
rect 4932 4948 4985 4968
rect 5037 4948 5091 5000
rect 5168 4970 5188 5000
rect 5143 4948 5188 4970
rect 5240 4948 5285 5000
rect 5337 4948 5346 5000
rect 4552 4947 5346 4948
rect 4120 4934 5346 4947
rect 17321 5008 18588 5020
rect 17321 5001 17391 5008
rect 17321 4967 17343 5001
rect 17377 4967 17391 5001
rect 17321 4956 17391 4967
rect 17443 5006 18588 5008
rect 17443 4956 17503 5006
rect 17321 4954 17503 4956
rect 17555 4954 17610 5006
rect 17662 5000 17712 5006
rect 17764 5005 18588 5006
rect 17764 5004 17844 5005
rect 17878 5004 18588 5005
rect 17662 4966 17679 5000
rect 17662 4954 17712 4966
rect 17764 4954 17838 5004
rect 17321 4952 17838 4954
rect 17890 4952 17992 5004
rect 18044 4992 18129 5004
rect 18045 4958 18129 4992
rect 18181 4990 18226 5004
rect 18044 4952 18129 4958
rect 18213 4956 18226 4990
rect 18181 4952 18226 4956
rect 18278 4952 18326 5004
rect 18378 5003 18588 5004
rect 18378 4999 18415 5003
rect 18383 4965 18415 4999
rect 18378 4952 18415 4965
rect 17321 4951 18415 4952
rect 18467 4951 18511 5003
rect 18563 4951 18588 5003
rect 17321 4936 18588 4951
rect 19207 5009 20463 5018
rect 19207 5006 19728 5009
rect 19207 5002 19557 5006
rect 19591 5002 19728 5006
rect 19762 5002 20463 5009
rect 19207 5000 19225 5002
rect 19207 4966 19222 5000
rect 19207 4950 19225 4966
rect 19277 4950 19319 5002
rect 19371 5001 19418 5002
rect 19371 4967 19395 5001
rect 19371 4950 19418 4967
rect 19470 4950 19526 5002
rect 19591 4972 19622 5002
rect 19578 4950 19622 4972
rect 19674 4950 19720 5002
rect 19772 5001 20463 5002
rect 19772 4950 19839 5001
rect 19207 4949 19839 4950
rect 19891 4995 19953 5001
rect 19891 4961 19897 4995
rect 19931 4961 19953 4995
rect 19891 4949 19953 4961
rect 20005 4995 20070 5001
rect 20005 4961 20062 4995
rect 20005 4949 20070 4961
rect 20122 4949 20197 5001
rect 20249 4993 20312 5001
rect 20266 4959 20312 4993
rect 20249 4949 20312 4959
rect 20364 4997 20463 5001
rect 20364 4963 20395 4997
rect 20429 4963 20463 4997
rect 20364 4949 20463 4963
rect 19207 4934 20463 4949
rect 26631 3308 26744 3386
<< via1 >>
rect 4610 5290 4683 5343
rect 19704 5289 19780 5343
rect 2282 4950 2334 5002
rect 2389 4971 2411 5002
rect 2411 4971 2441 5002
rect 2389 4950 2441 4971
rect 2495 4950 2547 5002
rect 2611 4950 2663 5002
rect 2740 4971 2746 5004
rect 2746 4971 2780 5004
rect 2780 4971 2792 5004
rect 2740 4952 2792 4971
rect 2874 5001 2926 5003
rect 2874 4967 2915 5001
rect 2915 4967 2926 5001
rect 2874 4951 2926 4967
rect 2991 4951 3043 5003
rect 3096 5000 3148 5003
rect 3096 4966 3118 5000
rect 3118 4966 3148 5000
rect 3096 4951 3148 4966
rect 3202 4972 3250 5003
rect 3250 4972 3254 5003
rect 3202 4951 3254 4972
rect 3299 4951 3351 5003
rect 3396 4974 3420 5003
rect 3420 4974 3448 5003
rect 3396 4951 3448 4974
rect 4171 4947 4223 4999
rect 4278 4971 4294 4999
rect 4294 4971 4328 4999
rect 4328 4971 4330 4999
rect 4278 4947 4330 4971
rect 4384 4947 4436 4999
rect 4500 4947 4552 4999
rect 4622 4975 4630 5002
rect 4630 4975 4664 5002
rect 4664 5001 4674 5002
rect 4664 4975 4681 5001
rect 4622 4950 4681 4975
rect 4629 4949 4681 4950
rect 4763 4996 4815 5000
rect 4763 4962 4794 4996
rect 4794 4962 4815 4996
rect 4763 4948 4815 4962
rect 4880 4948 4932 5000
rect 4985 4968 4998 5000
rect 4998 4968 5037 5000
rect 4985 4948 5037 4968
rect 5091 4970 5134 5000
rect 5134 4970 5143 5000
rect 5091 4948 5143 4970
rect 5188 4948 5240 5000
rect 5285 4972 5293 5000
rect 5293 4972 5327 5000
rect 5327 4972 5337 5000
rect 5285 4948 5337 4972
rect 17391 4956 17443 5008
rect 17503 4996 17555 5006
rect 17503 4962 17506 4996
rect 17506 4962 17540 4996
rect 17540 4962 17555 4996
rect 17503 4954 17555 4962
rect 17610 4954 17662 5006
rect 17712 5000 17764 5006
rect 17712 4966 17713 5000
rect 17713 4966 17764 5000
rect 17712 4954 17764 4966
rect 17838 4971 17844 5004
rect 17844 4971 17878 5004
rect 17878 4971 17890 5004
rect 17838 4952 17890 4971
rect 17992 4992 18044 5004
rect 17992 4958 18011 4992
rect 18011 4958 18044 4992
rect 18129 4990 18181 5004
rect 17992 4952 18044 4958
rect 18129 4956 18179 4990
rect 18179 4956 18181 4990
rect 18129 4952 18181 4956
rect 18226 4952 18278 5004
rect 18326 4999 18378 5004
rect 18326 4965 18349 4999
rect 18349 4965 18378 4999
rect 18326 4952 18378 4965
rect 18415 4951 18467 5003
rect 18511 4951 18563 5003
rect 19225 5000 19277 5002
rect 19225 4966 19256 5000
rect 19256 4966 19277 5000
rect 19225 4950 19277 4966
rect 19319 4950 19371 5002
rect 19418 5001 19470 5002
rect 19418 4967 19429 5001
rect 19429 4967 19470 5001
rect 19418 4950 19470 4967
rect 19526 4972 19557 5002
rect 19557 4972 19578 5002
rect 19526 4950 19578 4972
rect 19622 4950 19674 5002
rect 19720 4975 19728 5002
rect 19728 4975 19762 5002
rect 19762 4975 19772 5002
rect 19720 4950 19772 4975
rect 19839 4949 19891 5001
rect 19953 4949 20005 5001
rect 20070 4995 20122 5001
rect 20070 4961 20096 4995
rect 20096 4961 20122 4995
rect 20070 4949 20122 4961
rect 20197 4993 20249 5001
rect 20197 4959 20232 4993
rect 20232 4959 20249 4993
rect 20197 4949 20249 4959
rect 20312 4949 20364 5001
<< metal2 >>
rect 4475 5343 4844 5373
rect 4475 5290 4610 5343
rect 4683 5290 4844 5343
rect 4475 5272 4844 5290
rect 19621 5349 19892 5371
rect 19621 5343 19740 5349
rect 19621 5289 19704 5343
rect 19807 5296 19892 5349
rect 19780 5289 19892 5296
rect 19621 5271 19892 5289
rect -1439 5082 -413 5083
rect 446 5082 1472 5084
rect 13643 5082 14669 5084
rect 15544 5082 16570 5083
rect 21211 5082 22237 5086
rect 23115 5082 24141 5083
rect -3546 5020 11208 5082
rect 11562 5020 26308 5082
rect -3544 5004 11208 5020
rect -3544 5002 2740 5004
rect -3544 4950 2282 5002
rect 2334 4950 2389 5002
rect 2441 4950 2495 5002
rect 2547 4950 2611 5002
rect 2663 4952 2740 5002
rect 2792 5003 11208 5004
rect 2792 4952 2874 5003
rect 2663 4951 2874 4952
rect 2926 4951 2991 5003
rect 3043 4951 3096 5003
rect 3148 4951 3202 5003
rect 3254 4951 3299 5003
rect 3351 4951 3396 5003
rect 3448 5002 11208 5003
rect 3448 4999 4622 5002
rect 4674 5001 11208 5002
rect 3448 4951 4171 4999
rect 2663 4950 4171 4951
rect -3544 4947 4171 4950
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4947 4500 4999
rect 4552 4950 4622 4999
rect 4681 5000 11208 5001
rect 4552 4949 4629 4950
rect 4681 4949 4763 5000
rect 4552 4948 4763 4949
rect 4815 4948 4880 5000
rect 4932 4948 4985 5000
rect 5037 4948 5091 5000
rect 5143 4948 5188 5000
rect 5240 4948 5285 5000
rect 5337 4948 11208 5000
rect 11563 5008 26308 5020
rect 11563 4956 17391 5008
rect 17443 5006 26308 5008
rect 17443 4956 17503 5006
rect 4552 4947 11208 4948
rect -3544 4894 11208 4947
rect 11562 4954 17503 4956
rect 17555 4954 17610 5006
rect 17662 4954 17712 5006
rect 17764 5004 26308 5006
rect 17764 4954 17838 5004
rect 11562 4952 17838 4954
rect 17890 4952 17992 5004
rect 18044 4952 18129 5004
rect 18181 4952 18226 5004
rect 18278 4952 18326 5004
rect 18378 5003 26308 5004
rect 18378 4952 18415 5003
rect 11562 4951 18415 4952
rect 18467 4951 18511 5003
rect 18563 5002 26308 5003
rect 18563 4951 19225 5002
rect 11562 4950 19225 4951
rect 19277 4950 19319 5002
rect 19371 4950 19418 5002
rect 19470 4950 19526 5002
rect 19578 4950 19622 5002
rect 19674 4950 19720 5002
rect 19772 5001 26308 5002
rect 19772 4950 19839 5001
rect 11562 4949 19839 4950
rect 19891 4949 19953 5001
rect 20005 4949 20070 5001
rect 20122 4949 20197 5001
rect 20249 4949 20312 5001
rect 20364 4949 26308 5001
rect 11562 4894 26308 4949
rect -3326 4637 -2300 4894
rect -1439 4637 -413 4894
rect 446 4637 1472 4894
rect 2150 4886 5358 4894
rect 2150 4637 3470 4886
rect -3544 4590 3470 4637
rect 4034 4633 5358 4886
rect 6115 4633 7141 4894
rect 8010 4633 9036 4894
rect 9879 4633 10905 4894
rect 11756 4637 12782 4894
rect 13643 4637 14669 4894
rect 15544 4637 16570 4894
rect 17248 4886 20456 4894
rect 17248 4637 18568 4886
rect 19132 4637 20456 4886
rect 21211 4637 22237 4894
rect 23115 4637 24141 4894
rect 24991 4637 26017 4894
rect 4034 4590 11208 4633
rect -3544 4528 11208 4590
rect 11562 4590 26307 4637
rect 11562 4528 26306 4590
rect 2150 4524 3470 4528
rect 4034 4524 11208 4528
rect 17248 4524 18568 4528
rect 19132 4524 20456 4528
rect -3544 4002 -3352 4038
<< via2 >>
rect 4610 5290 4683 5343
rect 19740 5343 19807 5349
rect 19740 5296 19780 5343
rect 19780 5296 19807 5343
<< metal3 >>
rect 4475 5343 4844 5373
rect 4475 5290 4610 5343
rect 4683 5290 4844 5343
rect 4475 5272 4844 5290
rect 19618 5349 19894 5374
rect 19618 5347 19740 5349
rect 19618 5291 19739 5347
rect 19807 5296 19894 5349
rect 19799 5291 19894 5296
rect 19618 5270 19894 5291
rect -3552 4650 -2011 4904
rect -3544 2527 -2011 2782
<< via3 >>
rect 4610 5290 4683 5343
rect 19739 5296 19740 5347
rect 19740 5296 19799 5347
rect 19739 5291 19799 5296
rect 4606 2570 4673 2653
rect 19699 2572 19780 2656
<< metal4 >>
rect 4486 5343 4812 5412
rect 4486 5290 4610 5343
rect 4683 5290 4812 5343
rect 4486 2653 4812 5290
rect 4486 2570 4606 2653
rect 4673 2570 4812 2653
rect 4486 2535 4812 2570
rect 19628 5347 19893 5374
rect 19628 5291 19739 5347
rect 19799 5291 19893 5347
rect 19628 2656 19893 5291
rect 19628 2572 19699 2656
rect 19780 2572 19893 2656
rect 19628 2507 19893 2572
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654066915
transform 1 0 19092 0 -1 5320
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654066915
transform 1 0 17210 0 -1 5322
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1654066915
transform 1 0 3994 0 -1 5320
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1654066915
transform 1 0 2112 0 -1 5322
box -38 -48 1510 592
use unitcell2buf  unitcell2buf_0
timestamp 1654115785
transform 1 0 23448 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_1
timestamp 1654115785
transform 1 0 21560 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_2
timestamp 1654115785
transform 1 0 19672 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_3
timestamp 1654115785
transform 1 0 17784 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_4
timestamp 1654115785
transform 1 0 15896 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_5
timestamp 1654115785
transform 1 0 14008 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_6
timestamp 1654115785
transform 1 0 12120 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_7
timestamp 1654115785
transform 1 0 8350 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_8
timestamp 1654115785
transform 1 0 6462 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_9
timestamp 1654115785
transform 1 0 4574 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_10
timestamp 1654115785
transform 1 0 2686 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_11
timestamp 1654115785
transform 1 0 798 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_12
timestamp 1654115785
transform 1 0 -1090 0 1 3712
box -574 -1185 1322 1192
use unitcell2buf  unitcell2buf_13
timestamp 1654115785
transform 1 0 -2978 0 1 3712
box -574 -1185 1322 1192
use unitcell2bufcut  unitcell2bufcut_0
timestamp 1654116291
transform 1 0 25336 0 1 3712
box -574 -1184 1322 1192
use unitcell2bufcut  unitcell2bufcut_1
timestamp 1654116291
transform 1 0 10238 0 1 3712
box -574 -1184 1322 1192
<< labels >>
flabel metal1 3688 5062 3894 5220 1 FreeSans 400 0 0 0 RESET1
flabel metal1 18800 5062 18998 5222 1 FreeSans 800 0 0 0 RESET2
flabel metal3 -3552 4650 -2011 4904 1 FreeSans 800 0 0 0 VDD
flabel metal2 -3544 4002 -3352 4038 1 FreeSans 800 0 0 0 IN
flabel metal1 26631 3308 26744 3386 1 FreeSans 400 0 0 0 OUT
flabel metal3 -3544 2527 -2011 2782 1 FreeSans 800 0 0 0 VSS
<< end >>
