magic
tech sky130A
magscale 1 2
timestamp 1649788711
<< nmoslvt >>
rect -200 -900 200 900
<< ndiff >>
rect -258 888 -200 900
rect -258 -888 -246 888
rect -212 -888 -200 888
rect -258 -900 -200 -888
rect 200 888 258 900
rect 200 -888 212 888
rect 246 -888 258 888
rect 200 -900 258 -888
<< ndiffc >>
rect -246 -888 -212 888
rect 212 -888 246 888
<< poly >>
rect -126 972 126 988
rect -126 955 -110 972
rect -200 938 -110 955
rect 110 955 126 972
rect 110 938 200 955
rect -200 900 200 938
rect -200 -938 200 -900
rect -200 -955 -110 -938
rect -126 -972 -110 -955
rect 110 -955 200 -938
rect 110 -972 126 -955
rect -126 -988 126 -972
<< polycont >>
rect -110 938 110 972
rect -110 -972 110 -938
<< locali >>
rect -126 938 -110 972
rect 110 938 126 972
rect -246 888 -212 904
rect -246 -904 -212 -888
rect 212 888 246 904
rect 212 -904 246 -888
rect -126 -972 -110 -938
rect 110 -972 126 -938
<< viali >>
rect -74 938 74 972
rect -246 -888 -212 888
rect 212 -888 246 888
rect -74 -972 74 -938
<< metal1 >>
rect -86 972 86 978
rect -86 938 -74 972
rect 74 938 86 972
rect -86 932 86 938
rect -252 888 -206 900
rect -252 -888 -246 888
rect -212 -888 -206 888
rect -252 -900 -206 -888
rect 206 888 252 900
rect 206 -888 212 888
rect 246 -888 252 888
rect 206 -900 252 -888
rect -86 -938 86 -932
rect -86 -972 -74 -938
rect 74 -972 86 -938
rect -86 -978 86 -972
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 9 l 2 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
