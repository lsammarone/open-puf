magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 183
rect 29 -17 63 21
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 459 719 493
rect 17 425 29 459
rect 63 425 121 459
rect 155 425 213 459
rect 247 425 305 459
rect 339 425 397 459
rect 431 425 489 459
rect 523 425 581 459
rect 615 425 673 459
rect 707 425 719 459
rect 17 309 719 425
rect 17 171 347 275
rect 381 205 719 309
rect 17 17 719 171
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 425 63 459
rect 121 425 155 459
rect 213 425 247 459
rect 305 425 339 459
rect 397 425 431 459
rect 489 425 523 459
rect 581 425 615 459
rect 673 425 707 459
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 14 459 722 468
rect 14 428 29 459
rect 17 425 29 428
rect 63 425 121 459
rect 155 425 213 459
rect 247 425 305 459
rect 339 425 397 459
rect 431 425 489 459
rect 523 425 581 459
rect 615 425 673 459
rect 707 428 722 459
rect 707 425 719 428
rect 17 416 719 425
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel metal1 s 17 416 719 428 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 14 428 722 468 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 735 183 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2348336
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2344084
<< end >>
