magic
tech sky130B
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_0
timestamp 1648127584
transform -1 0 -165 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_1
timestamp 1648127584
transform 1 0 471 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_2
timestamp 1648127584
transform 1 0 1307 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_3
timestamp 1648127584
transform 1 0 2143 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_4
timestamp 1648127584
transform 1 0 2979 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_5
timestamp 1648127584
transform 1 0 3815 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_6
timestamp 1648127584
transform 1 0 4651 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_7
timestamp 1648127584
transform 1 0 5487 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_8
timestamp 1648127584
transform 1 0 6323 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_9
timestamp 1648127584
transform 1 0 7159 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_10
timestamp 1648127584
transform 1 0 7995 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_11
timestamp 1648127584
transform 1 0 8831 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808702  sky130_fd_pr__dftpl1s2__example_55959141808702_12
timestamp 1648127584
transform 1 0 9667 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 9767 675 9767 675 0 FreeSans 300 0 0 0 S
flabel comment s 9349 700 9349 700 0 FreeSans 300 0 0 0 D
flabel comment s 8931 675 8931 675 0 FreeSans 300 0 0 0 S
flabel comment s 8513 700 8513 700 0 FreeSans 300 0 0 0 D
flabel comment s 8095 675 8095 675 0 FreeSans 300 0 0 0 S
flabel comment s 7677 700 7677 700 0 FreeSans 300 0 0 0 D
flabel comment s 7259 675 7259 675 0 FreeSans 300 0 0 0 S
flabel comment s 6841 700 6841 700 0 FreeSans 300 0 0 0 D
flabel comment s 6423 675 6423 675 0 FreeSans 300 0 0 0 S
flabel comment s 6005 700 6005 700 0 FreeSans 300 0 0 0 D
flabel comment s 5587 675 5587 675 0 FreeSans 300 0 0 0 S
flabel comment s 5169 700 5169 700 0 FreeSans 300 0 0 0 D
flabel comment s 4751 675 4751 675 0 FreeSans 300 0 0 0 S
flabel comment s 4333 700 4333 700 0 FreeSans 300 0 0 0 D
flabel comment s 3915 675 3915 675 0 FreeSans 300 0 0 0 S
flabel comment s 3497 700 3497 700 0 FreeSans 300 0 0 0 D
flabel comment s 3079 675 3079 675 0 FreeSans 300 0 0 0 S
flabel comment s 2661 700 2661 700 0 FreeSans 300 0 0 0 D
flabel comment s 2243 675 2243 675 0 FreeSans 300 0 0 0 S
flabel comment s 1825 700 1825 700 0 FreeSans 300 0 0 0 D
flabel comment s 1407 675 1407 675 0 FreeSans 300 0 0 0 S
flabel comment s 989 700 989 700 0 FreeSans 300 0 0 0 D
flabel comment s 571 675 571 675 0 FreeSans 300 0 0 0 S
flabel comment s 153 700 153 700 0 FreeSans 300 0 0 0 D
flabel comment s -265 675 -265 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 15403846
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15391188
<< end >>
