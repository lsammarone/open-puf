magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 779 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 503 297 533 497
rect 587 297 617 497
rect 671 297 701 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 95 167 129
rect 113 61 123 95
rect 157 61 167 95
rect 113 47 167 61
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 95 335 129
rect 281 61 291 95
rect 325 61 335 95
rect 281 47 335 61
rect 365 95 419 177
rect 365 61 375 95
rect 409 61 419 95
rect 365 47 419 61
rect 449 163 503 177
rect 449 129 459 163
rect 493 129 503 163
rect 449 95 503 129
rect 449 61 459 95
rect 493 61 503 95
rect 449 47 503 61
rect 533 95 587 177
rect 533 61 543 95
rect 577 61 587 95
rect 533 47 587 61
rect 617 163 671 177
rect 617 129 627 163
rect 661 129 671 163
rect 617 95 671 129
rect 617 61 627 95
rect 661 61 671 95
rect 617 47 671 61
rect 701 95 753 177
rect 701 61 711 95
rect 745 61 753 95
rect 701 47 753 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 485 167 497
rect 113 451 123 485
rect 157 451 167 485
rect 113 417 167 451
rect 113 383 123 417
rect 157 383 167 417
rect 113 297 167 383
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 485 335 497
rect 281 451 291 485
rect 325 451 335 485
rect 281 417 335 451
rect 281 383 291 417
rect 325 383 335 417
rect 281 297 335 383
rect 365 485 419 497
rect 365 451 375 485
rect 409 451 419 485
rect 365 417 419 451
rect 365 383 375 417
rect 409 383 419 417
rect 365 341 419 383
rect 365 307 375 341
rect 409 307 419 341
rect 365 297 419 307
rect 449 409 503 497
rect 449 375 459 409
rect 493 375 503 409
rect 449 341 503 375
rect 449 307 459 341
rect 493 307 503 341
rect 449 297 503 307
rect 533 489 587 497
rect 533 455 543 489
rect 577 455 587 489
rect 533 421 587 455
rect 533 387 543 421
rect 577 387 587 421
rect 533 297 587 387
rect 617 409 671 497
rect 617 375 627 409
rect 661 375 671 409
rect 617 341 671 375
rect 617 307 627 341
rect 661 307 671 341
rect 617 297 671 307
rect 701 485 755 497
rect 701 451 711 485
rect 745 451 755 485
rect 701 417 755 451
rect 701 383 711 417
rect 745 383 755 417
rect 701 297 755 383
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 123 61 157 95
rect 207 61 241 95
rect 291 129 325 163
rect 291 61 325 95
rect 375 61 409 95
rect 459 129 493 163
rect 459 61 493 95
rect 543 61 577 95
rect 627 129 661 163
rect 627 61 661 95
rect 711 61 745 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 451 157 485
rect 123 383 157 417
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 451 325 485
rect 291 383 325 417
rect 375 451 409 485
rect 375 383 409 417
rect 375 307 409 341
rect 459 375 493 409
rect 459 307 493 341
rect 543 455 577 489
rect 543 387 577 421
rect 627 375 661 409
rect 627 307 661 341
rect 711 451 745 485
rect 711 383 745 417
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 419 497 449 523
rect 503 497 533 523
rect 587 497 617 523
rect 671 497 701 523
rect 83 265 113 297
rect 167 265 197 297
rect 251 265 281 297
rect 335 265 365 297
rect 83 249 365 265
rect 83 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 365 249
rect 83 199 365 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 177 281 199
rect 335 177 365 199
rect 419 265 449 297
rect 503 265 533 297
rect 587 265 617 297
rect 671 265 701 297
rect 419 249 701 265
rect 419 215 442 249
rect 476 215 510 249
rect 544 215 578 249
rect 612 215 646 249
rect 680 215 701 249
rect 419 199 701 215
rect 419 177 449 199
rect 503 177 533 199
rect 587 177 617 199
rect 671 177 701 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
<< polycont >>
rect 103 215 137 249
rect 171 215 205 249
rect 239 215 273 249
rect 307 215 341 249
rect 442 215 476 249
rect 510 215 544 249
rect 578 215 612 249
rect 646 215 680 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 477 73 493
rect 18 443 39 477
rect 18 409 73 443
rect 18 375 39 409
rect 18 341 73 375
rect 107 485 173 527
rect 107 451 123 485
rect 157 451 173 485
rect 107 417 173 451
rect 107 383 123 417
rect 157 383 173 417
rect 107 367 173 383
rect 207 477 241 493
rect 207 409 241 443
rect 18 307 39 341
rect 207 341 241 375
rect 275 485 325 527
rect 275 451 291 485
rect 275 417 325 451
rect 275 383 291 417
rect 275 367 325 383
rect 359 489 778 493
rect 359 485 543 489
rect 359 451 375 485
rect 409 459 543 485
rect 409 451 425 459
rect 359 417 425 451
rect 527 455 543 459
rect 577 485 778 489
rect 577 459 711 485
rect 577 455 593 459
rect 359 383 375 417
rect 409 383 425 417
rect 73 307 207 333
rect 359 341 425 383
rect 359 333 375 341
rect 241 307 375 333
rect 409 307 425 341
rect 18 291 425 307
rect 459 409 493 425
rect 527 421 593 455
rect 695 451 711 459
rect 745 451 778 485
rect 527 387 543 421
rect 577 387 593 421
rect 627 409 661 425
rect 459 349 493 375
rect 695 417 778 451
rect 695 383 711 417
rect 745 383 778 417
rect 627 349 661 375
rect 459 341 811 349
rect 493 307 627 341
rect 661 307 811 341
rect 459 289 811 307
rect 28 249 360 255
rect 28 215 103 249
rect 137 215 171 249
rect 205 215 239 249
rect 273 215 307 249
rect 341 215 360 249
rect 424 249 697 255
rect 424 215 442 249
rect 476 215 510 249
rect 544 215 578 249
rect 612 215 646 249
rect 680 215 697 249
rect 731 181 811 289
rect 18 163 73 181
rect 18 129 39 163
rect 18 95 73 129
rect 18 61 39 95
rect 18 17 73 61
rect 107 163 811 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 107 95 173 129
rect 275 129 291 145
rect 325 145 459 163
rect 325 129 341 145
rect 107 61 123 95
rect 157 61 173 95
rect 107 51 173 61
rect 207 95 241 111
rect 207 17 241 61
rect 275 95 341 129
rect 443 129 459 145
rect 493 145 627 163
rect 493 129 509 145
rect 275 61 291 95
rect 325 61 341 95
rect 275 51 341 61
rect 375 95 409 111
rect 375 17 409 61
rect 443 95 509 129
rect 611 129 627 145
rect 661 145 811 163
rect 661 129 677 145
rect 443 61 459 95
rect 493 61 509 95
rect 443 51 509 61
rect 543 95 577 111
rect 543 17 577 61
rect 611 95 677 129
rect 611 61 627 95
rect 661 61 677 95
rect 611 51 677 61
rect 711 95 768 111
rect 745 61 768 95
rect 711 17 768 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 765 289 799 323 0 FreeSans 400 0 0 0 Y
port 7 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor2_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1963870
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1956824
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
