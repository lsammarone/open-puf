magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 37 67 504 203
rect 37 21 407 67
rect 37 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 131 47 161 177
rect 215 47 245 177
rect 299 47 329 177
rect 396 93 426 177
<< scpmoshvt >>
rect 131 297 161 497
rect 215 297 245 497
rect 299 297 329 497
rect 396 330 426 414
<< ndiff >>
rect 63 163 131 177
rect 63 129 71 163
rect 105 129 131 163
rect 63 95 131 129
rect 63 61 71 95
rect 105 61 131 95
rect 63 47 131 61
rect 161 95 215 177
rect 161 61 171 95
rect 205 61 215 95
rect 161 47 215 61
rect 245 116 299 177
rect 245 82 255 116
rect 289 82 299 116
rect 245 47 299 82
rect 329 163 396 177
rect 329 129 339 163
rect 373 129 396 163
rect 329 95 396 129
rect 329 61 339 95
rect 373 93 396 95
rect 426 149 478 177
rect 426 115 436 149
rect 470 115 478 149
rect 426 93 478 115
rect 373 61 381 93
rect 329 47 381 61
<< pdiff >>
rect 67 475 131 497
rect 67 441 75 475
rect 109 441 131 475
rect 67 347 131 441
rect 67 313 75 347
rect 109 313 131 347
rect 67 297 131 313
rect 161 297 215 497
rect 245 297 299 497
rect 329 459 381 497
rect 329 425 339 459
rect 373 425 381 459
rect 329 414 381 425
rect 329 330 396 414
rect 426 391 478 414
rect 426 357 436 391
rect 470 357 478 391
rect 426 330 478 357
rect 329 297 381 330
<< ndiffc >>
rect 71 129 105 163
rect 71 61 105 95
rect 171 61 205 95
rect 255 82 289 116
rect 339 129 373 163
rect 339 61 373 95
rect 436 115 470 149
<< pdiffc >>
rect 75 441 109 475
rect 75 313 109 347
rect 339 425 373 459
rect 436 357 470 391
<< poly >>
rect 131 497 161 523
rect 215 497 245 523
rect 299 497 329 523
rect 396 414 426 440
rect 131 265 161 297
rect 215 265 245 297
rect 299 265 329 297
rect 396 265 426 330
rect 91 249 161 265
rect 91 215 101 249
rect 135 215 161 249
rect 91 199 161 215
rect 203 249 257 265
rect 203 215 213 249
rect 247 215 257 249
rect 203 199 257 215
rect 299 249 353 265
rect 299 215 309 249
rect 343 215 353 249
rect 299 199 353 215
rect 395 249 449 265
rect 395 215 405 249
rect 439 215 449 249
rect 395 199 449 215
rect 131 177 161 199
rect 215 177 245 199
rect 299 177 329 199
rect 396 177 426 199
rect 396 67 426 93
rect 131 21 161 47
rect 215 21 245 47
rect 299 21 329 47
<< polycont >>
rect 101 215 135 249
rect 213 215 247 249
rect 309 215 343 249
rect 405 215 439 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 475 109 491
rect 17 441 75 475
rect 17 347 109 441
rect 323 459 389 527
rect 323 425 339 459
rect 373 425 389 459
rect 17 313 75 347
rect 17 289 109 313
rect 143 357 436 391
rect 470 357 535 391
rect 17 165 51 289
rect 143 249 177 357
rect 85 215 101 249
rect 135 215 177 249
rect 213 249 261 323
rect 247 215 261 249
rect 213 199 261 215
rect 295 249 363 323
rect 295 215 309 249
rect 343 215 363 249
rect 295 199 363 215
rect 397 249 467 323
rect 397 215 405 249
rect 439 215 467 249
rect 397 199 467 215
rect 501 165 535 357
rect 17 163 289 165
rect 17 129 71 163
rect 105 131 289 163
rect 105 129 121 131
rect 17 95 121 129
rect 255 116 289 131
rect 17 61 71 95
rect 105 61 121 95
rect 17 51 121 61
rect 155 95 221 97
rect 155 61 171 95
rect 205 61 221 95
rect 255 62 289 82
rect 323 163 389 165
rect 323 129 339 163
rect 373 129 389 163
rect 323 95 389 129
rect 155 17 221 61
rect 323 61 339 95
rect 373 61 389 95
rect 436 149 535 165
rect 470 131 535 149
rect 436 81 470 115
rect 323 17 389 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 29 357 63 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 305 221 339 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor3b_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 1128596
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1123852
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 2.760 0.000 
<< end >>
