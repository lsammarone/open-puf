magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 1 293 1415 625
<< pwell >>
rect 41 19 1375 155
<< mvnmos >>
rect 120 45 240 129
rect 296 45 416 129
rect 472 45 592 129
rect 648 45 768 129
rect 824 45 944 129
rect 1000 45 1120 129
rect 1176 45 1296 129
<< mvpmos >>
rect 120 359 240 559
rect 296 359 416 559
rect 472 359 592 559
rect 648 359 768 559
rect 824 359 944 559
rect 1000 359 1120 559
rect 1176 359 1296 559
<< mvndiff >>
rect 67 91 120 129
rect 67 57 75 91
rect 109 57 120 91
rect 67 45 120 57
rect 240 91 296 129
rect 240 57 251 91
rect 285 57 296 91
rect 240 45 296 57
rect 416 91 472 129
rect 416 57 427 91
rect 461 57 472 91
rect 416 45 472 57
rect 592 91 648 129
rect 592 57 603 91
rect 637 57 648 91
rect 592 45 648 57
rect 768 91 824 129
rect 768 57 779 91
rect 813 57 824 91
rect 768 45 824 57
rect 944 91 1000 129
rect 944 57 955 91
rect 989 57 1000 91
rect 944 45 1000 57
rect 1120 91 1176 129
rect 1120 57 1131 91
rect 1165 57 1176 91
rect 1120 45 1176 57
rect 1296 91 1349 129
rect 1296 57 1307 91
rect 1341 57 1349 91
rect 1296 45 1349 57
<< mvpdiff >>
rect 67 541 120 559
rect 67 507 75 541
rect 109 507 120 541
rect 67 473 120 507
rect 67 439 75 473
rect 109 439 120 473
rect 67 405 120 439
rect 67 371 75 405
rect 109 371 120 405
rect 67 359 120 371
rect 240 541 296 559
rect 240 507 251 541
rect 285 507 296 541
rect 240 473 296 507
rect 240 439 251 473
rect 285 439 296 473
rect 240 405 296 439
rect 240 371 251 405
rect 285 371 296 405
rect 240 359 296 371
rect 416 541 472 559
rect 416 507 427 541
rect 461 507 472 541
rect 416 473 472 507
rect 416 439 427 473
rect 461 439 472 473
rect 416 405 472 439
rect 416 371 427 405
rect 461 371 472 405
rect 416 359 472 371
rect 592 541 648 559
rect 592 507 603 541
rect 637 507 648 541
rect 592 473 648 507
rect 592 439 603 473
rect 637 439 648 473
rect 592 405 648 439
rect 592 371 603 405
rect 637 371 648 405
rect 592 359 648 371
rect 768 541 824 559
rect 768 507 779 541
rect 813 507 824 541
rect 768 473 824 507
rect 768 439 779 473
rect 813 439 824 473
rect 768 405 824 439
rect 768 371 779 405
rect 813 371 824 405
rect 768 359 824 371
rect 944 541 1000 559
rect 944 507 955 541
rect 989 507 1000 541
rect 944 473 1000 507
rect 944 439 955 473
rect 989 439 1000 473
rect 944 405 1000 439
rect 944 371 955 405
rect 989 371 1000 405
rect 944 359 1000 371
rect 1120 541 1176 559
rect 1120 507 1131 541
rect 1165 507 1176 541
rect 1120 473 1176 507
rect 1120 439 1131 473
rect 1165 439 1176 473
rect 1120 405 1176 439
rect 1120 371 1131 405
rect 1165 371 1176 405
rect 1120 359 1176 371
rect 1296 541 1349 559
rect 1296 507 1307 541
rect 1341 507 1349 541
rect 1296 473 1349 507
rect 1296 439 1307 473
rect 1341 439 1349 473
rect 1296 405 1349 439
rect 1296 371 1307 405
rect 1341 371 1349 405
rect 1296 359 1349 371
<< mvndiffc >>
rect 75 57 109 91
rect 251 57 285 91
rect 427 57 461 91
rect 603 57 637 91
rect 779 57 813 91
rect 955 57 989 91
rect 1131 57 1165 91
rect 1307 57 1341 91
<< mvpdiffc >>
rect 75 507 109 541
rect 75 439 109 473
rect 75 371 109 405
rect 251 507 285 541
rect 251 439 285 473
rect 251 371 285 405
rect 427 507 461 541
rect 427 439 461 473
rect 427 371 461 405
rect 603 507 637 541
rect 603 439 637 473
rect 603 371 637 405
rect 779 507 813 541
rect 779 439 813 473
rect 779 371 813 405
rect 955 507 989 541
rect 955 439 989 473
rect 955 371 989 405
rect 1131 507 1165 541
rect 1131 439 1165 473
rect 1131 371 1165 405
rect 1307 507 1341 541
rect 1307 439 1341 473
rect 1307 371 1341 405
<< poly >>
rect 120 559 240 585
rect 296 559 416 585
rect 472 559 592 585
rect 648 559 768 585
rect 824 559 944 585
rect 1000 559 1120 585
rect 1176 559 1296 585
rect 120 333 240 359
rect 296 333 416 359
rect 472 333 592 359
rect 648 333 768 359
rect 824 333 944 359
rect 1000 333 1120 359
rect 1176 333 1296 359
rect 120 295 1296 333
rect 120 261 156 295
rect 190 261 1296 295
rect 120 258 1296 261
rect 120 227 340 258
rect 120 193 156 227
rect 190 224 340 227
rect 374 224 409 258
rect 443 224 478 258
rect 512 224 722 258
rect 756 224 835 258
rect 869 224 1094 258
rect 1128 224 1223 258
rect 1257 224 1296 258
rect 190 193 1296 224
rect 120 155 1296 193
rect 120 129 240 155
rect 296 129 416 155
rect 472 129 592 155
rect 648 129 768 155
rect 824 129 944 155
rect 1000 129 1120 155
rect 1176 129 1296 155
rect 120 19 240 45
rect 296 19 416 45
rect 472 19 592 45
rect 648 19 768 45
rect 824 19 944 45
rect 1000 19 1120 45
rect 1176 19 1296 45
<< polycont >>
rect 156 261 190 295
rect 156 193 190 227
rect 340 224 374 258
rect 409 224 443 258
rect 478 224 512 258
rect 722 224 756 258
rect 835 224 869 258
rect 1094 224 1128 258
rect 1223 224 1257 258
<< locali >>
rect 75 495 109 507
rect 75 405 109 439
rect 241 541 285 559
rect 241 507 251 541
rect 241 473 285 507
rect 241 439 251 473
rect 241 405 285 439
rect 241 378 251 405
rect 427 495 461 507
rect 427 405 461 439
rect 75 355 109 371
rect 285 371 291 378
rect 253 344 291 371
rect 427 355 461 371
rect 566 541 672 557
rect 566 507 603 541
rect 637 507 672 541
rect 566 473 672 507
rect 566 439 603 473
rect 637 439 672 473
rect 566 405 672 439
rect 566 378 603 405
rect 600 371 603 378
rect 637 378 672 405
rect 637 371 638 378
rect 600 344 638 371
rect 779 495 813 507
rect 779 405 813 439
rect 779 355 813 371
rect 919 541 1025 557
rect 919 507 955 541
rect 989 507 1025 541
rect 919 473 1025 507
rect 919 439 955 473
rect 989 439 1025 473
rect 919 405 1025 439
rect 919 378 955 405
rect 156 295 190 311
rect 156 258 190 261
rect 122 227 160 258
rect 122 224 156 227
rect 156 177 190 193
rect 75 91 109 103
rect 241 91 285 344
rect 324 258 528 276
rect 324 224 340 258
rect 374 224 382 258
rect 443 224 454 258
rect 512 224 528 258
rect 324 206 528 224
rect 241 57 251 91
rect 241 41 285 57
rect 427 91 461 103
rect 566 91 672 344
rect 953 371 955 378
rect 989 378 1025 405
rect 989 371 991 378
rect 953 344 991 371
rect 1131 495 1165 507
rect 1131 405 1165 439
rect 1307 541 1349 557
rect 1341 507 1349 541
rect 1307 473 1349 507
rect 1341 439 1349 473
rect 1307 405 1349 439
rect 1341 378 1349 405
rect 1131 355 1165 371
rect 1278 371 1307 378
rect 1278 344 1316 371
rect 706 258 885 276
rect 706 224 722 258
rect 786 224 824 258
rect 869 224 885 258
rect 706 206 885 224
rect 566 57 603 91
rect 637 57 672 91
rect 566 41 672 57
rect 779 91 813 103
rect 919 91 1025 344
rect 1078 258 1273 276
rect 1078 224 1094 258
rect 1143 224 1181 258
rect 1215 224 1223 258
rect 1257 224 1273 258
rect 1078 206 1273 224
rect 919 57 955 91
rect 989 57 1025 91
rect 919 41 1025 57
rect 1131 91 1165 103
rect 1307 91 1349 344
rect 1341 57 1349 91
rect 1307 41 1349 57
<< viali >>
rect 75 541 109 567
rect 75 533 109 541
rect 75 473 109 495
rect 75 461 109 473
rect 427 541 461 567
rect 427 533 461 541
rect 427 473 461 495
rect 427 461 461 473
rect 219 371 251 378
rect 251 371 253 378
rect 219 344 253 371
rect 291 344 325 378
rect 566 344 600 378
rect 638 344 672 378
rect 779 541 813 567
rect 779 533 813 541
rect 779 473 813 495
rect 779 461 813 473
rect 88 224 122 258
rect 160 227 194 258
rect 160 224 190 227
rect 190 224 194 227
rect 75 103 109 137
rect 75 57 109 65
rect 75 31 109 57
rect 382 224 409 258
rect 409 224 416 258
rect 454 224 478 258
rect 478 224 488 258
rect 427 103 461 137
rect 427 57 461 65
rect 427 31 461 57
rect 919 344 953 378
rect 991 344 1025 378
rect 1131 541 1165 567
rect 1131 533 1165 541
rect 1131 473 1165 495
rect 1131 461 1165 473
rect 1244 344 1278 378
rect 1316 371 1341 378
rect 1341 371 1350 378
rect 1316 344 1350 371
rect 752 224 756 258
rect 756 224 786 258
rect 824 224 835 258
rect 835 224 858 258
rect 779 103 813 137
rect 779 57 813 65
rect 779 31 813 57
rect 1109 224 1128 258
rect 1128 224 1143 258
rect 1181 224 1215 258
rect 1131 103 1165 137
rect 1131 57 1165 65
rect 1131 31 1165 57
<< metal1 >>
rect 69 567 1171 579
rect 69 533 75 567
rect 109 533 427 567
rect 461 533 779 567
rect 813 533 1131 567
rect 1165 533 1171 567
rect 69 495 1171 533
rect 69 461 75 495
rect 109 461 427 495
rect 461 461 779 495
rect 813 461 1131 495
rect 1165 461 1171 495
rect 69 449 1171 461
rect 207 378 1362 384
rect 207 344 219 378
rect 253 344 291 378
rect 325 344 566 378
rect 600 344 638 378
rect 672 344 919 378
rect 953 344 991 378
rect 1025 344 1244 378
rect 1278 344 1316 378
rect 1350 344 1362 378
rect 207 338 1362 344
rect 76 258 1227 264
rect 76 224 88 258
rect 122 224 160 258
rect 194 224 382 258
rect 416 224 454 258
rect 488 224 752 258
rect 786 224 824 258
rect 858 224 1109 258
rect 1143 224 1181 258
rect 1215 224 1227 258
rect 76 218 1227 224
rect 69 137 1171 149
rect 69 103 75 137
rect 109 103 427 137
rect 461 103 779 137
rect 813 103 1131 137
rect 1165 103 1171 137
rect 69 65 1171 103
rect 69 31 75 65
rect 109 31 427 65
rect 461 31 779 65
rect 813 31 1131 65
rect 1165 31 1171 65
rect 69 19 1171 31
use sky130_fd_pr__nfet_01v8__example_55959141808565  sky130_fd_pr__nfet_01v8__example_55959141808565_0
timestamp 1648127584
transform 1 0 120 0 1 45
box -28 0 1204 29
use sky130_fd_pr__pfet_01v8__example_55959141808566  sky130_fd_pr__pfet_01v8__example_55959141808566_0
timestamp 1648127584
transform 1 0 120 0 1 359
box -28 0 1204 97
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1648127584
transform -1 0 206 0 -1 311
box 0 0 1 1
<< labels >>
flabel metal1 s 147 42 243 99 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal1 s 146 490 233 554 3 FreeSans 520 0 0 0 VDA
port 2 nsew
flabel metal1 s 265 348 323 375 3 FreeSans 520 90 0 0 Y
port 3 nsew
flabel metal1 s 195 71 195 71 3 FreeSans 520 0 0 0 VSSA
port 1 nsew
flabel metal1 s 189 522 189 522 3 FreeSans 520 0 0 0 VDA
port 2 nsew
flabel metal1 s 121 227 190 253 3 FreeSans 520 0 0 0 A
port 4 nsew
<< properties >>
string GDS_END 8192054
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8185346
<< end >>
