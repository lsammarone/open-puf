magic
tech sky130A
magscale 1 2
timestamp 1652999729
<< nwell >>
rect 4402 3714 4966 3840
rect 4430 2798 5178 2838
rect 4428 2688 5178 2798
rect 4866 2558 5178 2688
rect 11040 2557 11361 2733
rect 11040 2325 11576 2557
rect 16734 2446 17055 4129
rect 24873 3223 25194 3756
rect 11038 2004 11576 2325
<< pwell >>
rect 4454 4181 4636 4561
<< psubdiff >>
rect 4534 4500 4630 4522
rect 4534 4464 4560 4500
rect 4604 4464 4630 4500
rect 4534 4438 4630 4464
<< nsubdiff >>
rect 4608 3796 4652 3832
rect 4688 3796 4712 3832
rect 25058 3642 25124 3666
rect 25058 3608 25074 3642
rect 25108 3608 25124 3642
rect 25058 3584 25124 3608
rect 11346 3466 11386 3506
rect 11346 3432 11350 3466
rect 11384 3432 11386 3466
rect 11346 3382 11386 3432
rect 16840 2824 16946 2826
rect 16840 2790 16868 2824
rect 16902 2790 16946 2824
rect 4598 2748 4674 2788
rect 4720 2748 4812 2788
rect 16840 2784 16946 2790
rect 4598 2742 4812 2748
<< psubdiffcont >>
rect 4560 4464 4604 4500
<< nsubdiffcont >>
rect 4652 3796 4688 3832
rect 25074 3608 25108 3642
rect 11350 3432 11384 3466
rect 16868 2790 16902 2824
rect 4674 2748 4720 2788
<< locali >>
rect 12274 5236 12342 5242
rect 12274 5168 12564 5236
rect 18465 5193 18751 5255
rect 12274 4558 12342 5168
rect 4534 4500 4634 4522
rect 4534 4464 4560 4500
rect 4604 4464 4634 4500
rect 4534 4434 4634 4464
rect 4440 4433 4634 4434
rect 4089 4398 4634 4433
rect 4089 4355 4521 4398
rect 4534 4370 4634 4398
rect 12168 4490 12342 4558
rect 4089 3543 4167 4355
rect 12168 4290 12236 4490
rect 18465 4485 18527 5193
rect 18355 4423 18527 4485
rect 18171 4404 18268 4405
rect 18355 4404 18417 4423
rect 18171 4343 18417 4404
rect 11822 4222 12236 4290
rect 4298 4170 4367 4182
rect 16632 4174 16790 4176
rect 4298 4122 4540 4170
rect 16628 4128 16790 4174
rect 4298 3707 4367 4122
rect 16628 4056 16692 4128
rect 5984 3980 11168 4049
rect 11829 3992 16692 4056
rect 4608 3796 4652 3824
rect 4688 3796 4710 3824
rect 4608 3776 4710 3796
rect 5984 3707 6053 3980
rect 4298 3638 6053 3707
rect 4089 3465 4275 3543
rect 4197 2220 4275 3465
rect 11334 3466 11490 3516
rect 11334 3432 11350 3466
rect 11384 3432 11490 3466
rect 11334 3376 11490 3432
rect 11354 3374 11490 3376
rect 11168 3298 11204 3326
rect 4328 3129 4397 3134
rect 6108 3129 6177 3132
rect 4326 3060 6177 3129
rect 4328 2452 4397 3060
rect 6108 2809 6177 3060
rect 16838 2824 16954 2838
rect 4648 2748 4674 2788
rect 4720 2748 4750 2788
rect 4648 2726 4750 2748
rect 6108 2740 11164 2809
rect 11825 2734 16696 2798
rect 4648 2722 4744 2726
rect 4328 2406 4550 2452
rect 16632 2446 16696 2734
rect 16838 2790 16868 2824
rect 16902 2790 16954 2824
rect 16838 2712 16954 2790
rect 16632 2404 16824 2446
rect 16634 2400 16824 2404
rect 4197 2142 4548 2220
rect 18355 2202 18417 4343
rect 25056 3642 25124 3654
rect 25056 3608 25074 3642
rect 25108 3608 25124 3642
rect 25056 3604 25124 3608
rect 25056 3523 25090 3604
rect 25056 3496 25088 3523
rect 25110 3200 25130 3228
rect 4467 1511 4545 2142
rect 18192 2140 18422 2202
rect 18351 1521 18413 2140
rect 4309 1433 4545 1511
rect 18199 1459 18413 1521
<< viali >>
rect 5744 4122 5790 4168
rect 18076 4124 18120 4164
rect 5768 2388 5814 2446
rect 18098 2398 18150 2444
rect 24916 3176 24960 3214
<< metal1 >>
rect 5732 4172 5802 4186
rect 5732 4120 5740 4172
rect 5794 4120 5802 4172
rect 5732 4108 5802 4120
rect 4440 2686 4544 3888
rect 5974 3884 6056 4683
rect 11797 4185 12085 4283
rect 5845 3803 6056 3884
rect 5870 3792 5901 3803
rect 5974 3802 6056 3803
rect 10887 3600 11140 3694
rect 5892 2762 5923 2782
rect 5870 2687 6055 2762
rect 5756 2446 5830 2458
rect 5756 2444 5768 2446
rect 5814 2444 5830 2446
rect 5756 2384 5764 2444
rect 5818 2384 5830 2444
rect 5756 2378 5830 2384
rect 5758 2376 5828 2378
rect 4416 2229 4478 2236
rect 4402 2150 4495 2229
rect 4416 2142 4478 2150
rect 18 2042 70 2050
rect 18 1990 82 2042
rect 34 1986 82 1990
rect 4178 1978 4258 2068
rect 5980 1983 6054 2687
rect 10887 2503 10981 3600
rect 11987 3086 12085 4185
rect 16627 3878 16701 4677
rect 24512 4622 24952 4718
rect 24856 4494 24952 4622
rect 24852 4452 24952 4494
rect 18187 4370 18254 4433
rect 18062 4174 18132 4178
rect 18062 4122 18072 4174
rect 18126 4122 18132 4174
rect 18062 4112 18132 4122
rect 16627 3804 16827 3878
rect 16775 3798 16806 3804
rect 11830 2988 12085 3086
rect 16809 2766 16840 2776
rect 16669 2691 16862 2766
rect 10887 2409 11175 2503
rect 10887 2067 10981 2409
rect 10887 1973 11033 2067
rect 16669 2066 16744 2691
rect 18166 2680 18268 3894
rect 24852 3462 24948 4452
rect 24902 3224 24972 3230
rect 24902 3172 24910 3224
rect 24966 3172 24972 3224
rect 24902 3166 24972 3172
rect 24902 3162 24970 3166
rect 18086 2444 18162 2456
rect 18086 2392 18096 2444
rect 18154 2392 18162 2444
rect 18086 2382 18162 2392
rect 18258 2223 18304 2232
rect 18241 2160 18308 2223
rect 18258 2138 18304 2160
rect 16621 1991 16744 2066
rect 24865 106 24947 3003
rect 34 40 76 76
rect 132 34 190 84
rect 24575 24 24947 106
<< via1 >>
rect 5740 4168 5794 4172
rect 5740 4122 5744 4168
rect 5744 4122 5790 4168
rect 5790 4122 5794 4168
rect 5740 4120 5794 4122
rect 5764 2388 5768 2444
rect 5768 2388 5814 2444
rect 5814 2388 5818 2444
rect 5764 2384 5818 2388
rect 18072 4164 18126 4174
rect 18072 4124 18076 4164
rect 18076 4124 18120 4164
rect 18120 4124 18126 4164
rect 18072 4122 18126 4124
rect 24910 3214 24966 3224
rect 24910 3176 24916 3214
rect 24916 3176 24960 3214
rect 24960 3176 24966 3214
rect 24910 3172 24966 3176
rect 18096 2398 18098 2444
rect 18098 2398 18150 2444
rect 18150 2398 18154 2444
rect 18096 2392 18154 2398
<< metal2 >>
rect 1438 6608 1454 6634
rect 2982 6620 2998 6646
rect 4524 6612 4540 6638
rect 6062 6616 6078 6642
rect 7604 6614 7620 6640
rect 9144 6614 9160 6640
rect 10692 6620 10708 6646
rect 12206 6624 12222 6650
rect 13754 6624 13770 6650
rect 15314 6602 15330 6628
rect 16856 6612 16872 6638
rect 18396 6622 18412 6648
rect 19942 6608 19958 6634
rect 21484 6602 21500 6628
rect 23026 6614 23042 6640
rect 24562 6614 24578 6640
rect -148 5330 20 5366
rect -148 4494 -112 5330
rect 24568 5326 24798 5362
rect -150 4390 -112 4494
rect -150 1362 -114 4390
rect 5768 4178 5800 4834
rect 10658 4812 10920 4840
rect 13692 4812 13912 4840
rect 5732 4172 5800 4178
rect 5732 4120 5740 4172
rect 5794 4120 5800 4172
rect 18060 4182 18090 4812
rect 18060 4174 18132 4182
rect 18060 4168 18072 4174
rect 5732 4114 5800 4120
rect 18062 4122 18072 4168
rect 18126 4122 18132 4174
rect 18062 4112 18132 4122
rect 24762 3196 24798 5326
rect 24902 3224 24972 3230
rect 24902 3196 24910 3224
rect 24762 3172 24910 3196
rect 24966 3172 24972 3224
rect 24762 3166 24972 3172
rect 5758 2444 5828 2450
rect 5758 2396 5764 2444
rect 5756 2384 5764 2396
rect 5818 2384 5828 2444
rect 18086 2444 18162 2458
rect 18086 2408 18096 2444
rect 5756 2376 5828 2384
rect 18084 2392 18096 2408
rect 18154 2392 18162 2444
rect 18084 2382 18162 2392
rect 5756 1852 5798 2376
rect 10752 1852 10952 1880
rect 13736 1852 13926 1880
rect 18084 1852 18134 2382
rect 24762 1362 24798 3166
rect -150 1326 58 1362
rect 24588 1326 24798 1362
rect 26 50 42 76
rect 1570 48 1586 74
rect 3108 52 3124 78
rect 4652 58 4668 84
rect 6198 54 6214 80
rect 7740 58 7756 84
rect 9274 50 9290 76
rect 10846 54 10862 80
rect 12386 50 12402 76
rect 13908 54 13924 80
rect 15448 54 15464 80
rect 16982 64 16998 90
rect 18534 50 18550 76
rect 20080 48 20096 74
rect 21612 54 21628 80
rect 23152 64 23168 90
use 8inv  8inv_0
timestamp 1652772933
transform 1 0 8738 0 1 -2200
box 2302 4602 3210 6484
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 24880 0 1 2962
box -38 -48 314 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 4466 0 1 2190
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1650294714
transform 1 0 16798 0 1 2184
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1650294714
transform 1 0 4440 0 -1 4384
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1650294714
transform 1 0 16772 0 -1 4390
box -38 -48 1510 592
use unitcell2  unitcell2_0
timestamp 1652990473
transform 1 0 566 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_1
timestamp 1652990473
transform 1 0 2108 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_2
timestamp 1652990473
transform 1 0 3650 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_3
timestamp 1652990473
transform 1 0 5192 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_4
timestamp 1652990473
transform 1 0 6734 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_5
timestamp 1652990473
transform 1 0 8276 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_6
timestamp 1652990473
transform 1 0 9818 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_7
timestamp 1652990473
transform -1 0 24042 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_8
timestamp 1652990473
transform -1 0 22500 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_9
timestamp 1652990473
transform 1 0 14444 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_10
timestamp 1652990473
transform 1 0 15986 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_11
timestamp 1652990473
transform 1 0 17528 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_12
timestamp 1652990473
transform 1 0 19070 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_13
timestamp 1652990473
transform 1 0 20612 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_14
timestamp 1652990473
transform 1 0 22154 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_15
timestamp 1652990473
transform 1 0 23696 0 1 1036
box -566 -1036 976 1034
use unitcell2  unitcell2_16
timestamp 1652990473
transform -1 0 20958 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_17
timestamp 1652990473
transform -1 0 19416 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_18
timestamp 1652990473
transform -1 0 17874 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_19
timestamp 1652990473
transform -1 0 16332 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_20
timestamp 1652990473
transform -1 0 14790 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_21
timestamp 1652990473
transform -1 0 10164 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_22
timestamp 1652990473
transform -1 0 8622 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_23
timestamp 1652990473
transform -1 0 7080 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_24
timestamp 1652990473
transform -1 0 5538 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_25
timestamp 1652990473
transform -1 0 3996 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_26
timestamp 1652990473
transform -1 0 2454 0 -1 5656
box -566 -1036 976 1034
use unitcell2  unitcell2_27
timestamp 1652990473
transform -1 0 912 0 -1 5656
box -566 -1036 976 1034
use unitcell2_cut  unitcell2_cut_0
timestamp 1652832150
transform 1 0 11360 0 1 1036
box -566 -1036 976 1034
use unitcell2_cut  unitcell2_cut_1
timestamp 1652832150
transform 1 0 12902 0 1 1036
box -566 -1036 976 1034
use unitcell2_cut  unitcell2_cut_2
timestamp 1652832150
transform -1 0 13248 0 -1 5656
box -566 -1036 976 1034
use unitcell2_cut  unitcell2_cut_3
timestamp 1652832150
transform -1 0 11706 0 -1 5656
box -566 -1036 976 1034
<< labels >>
flabel locali 11168 3298 11204 3326 1 FreeSans 160 0 0 0 RESET
port 36 n
flabel locali 25110 3200 25130 3228 1 FreeSans 160 0 0 0 OUT
port 3 n
flabel metal1 132 34 190 84 1 FreeSans 160 0 0 0 VSS
port 2 n
flabel metal1 18 1990 70 2050 1 FreeSans 160 0 0 0 VDD
port 1 n
flabel metal2 24562 6614 24578 6640 1 FreeSans 160 0 0 0 C1
port 28 n
flabel metal2 23026 6614 23042 6640 1 FreeSans 160 0 0 0 C2
port 29 n
flabel metal2 21484 6602 21500 6628 1 FreeSans 160 0 0 0 C3
port 30 n
flabel metal2 19942 6608 19958 6634 1 FreeSans 160 0 0 0 C4
port 31 n
flabel metal2 18396 6622 18412 6648 1 FreeSans 160 0 0 0 C5
port 32 n
flabel metal2 16856 6612 16872 6638 1 FreeSans 160 0 0 0 C6
port 33 n
flabel metal2 15314 6602 15330 6628 1 FreeSans 160 0 0 0 C7
port 34 n
flabel metal2 13754 6624 13770 6650 1 FreeSans 160 0 0 0 C8
port 35 n
flabel metal2 12206 6624 12222 6650 1 FreeSans 160 0 0 0 C9
port 4 n
flabel metal2 10692 6620 10708 6646 1 FreeSans 160 0 0 0 C10
port 5 n
flabel metal2 9144 6614 9160 6640 1 FreeSans 160 0 0 0 C11
port 6 n
flabel metal2 7604 6614 7620 6640 1 FreeSans 160 0 0 0 C12
port 7 n
flabel metal2 6062 6616 6078 6642 1 FreeSans 160 0 0 0 C13
port 8 n
flabel metal2 4524 6612 4540 6638 1 FreeSans 160 0 0 0 C14
port 9 n
flabel metal2 2982 6620 2998 6646 1 FreeSans 160 0 0 0 C15
port 10 n
flabel metal2 1438 6608 1454 6634 1 FreeSans 160 0 0 0 C16
port 11 n
flabel metal2 26 50 42 76 1 FreeSans 160 0 0 0 C17
port 12 n
flabel metal2 1570 48 1586 74 1 FreeSans 160 0 0 0 C18
port 13 n
flabel metal2 3108 52 3124 78 1 FreeSans 160 0 0 0 C19
port 14 n
flabel metal2 4652 58 4668 84 1 FreeSans 160 0 0 0 C20
port 15 n
flabel metal2 6198 54 6214 80 1 FreeSans 160 0 0 0 C21
port 16 n
flabel metal2 7740 58 7756 84 1 FreeSans 160 0 0 0 C22
port 17 n
flabel metal2 9274 50 9290 76 1 FreeSans 160 0 0 0 C23
port 18 n
flabel metal2 10846 54 10862 80 1 FreeSans 160 0 0 0 C24
port 19 n
flabel metal2 12386 50 12402 76 1 FreeSans 160 0 0 0 C25
port 20 n
flabel metal2 13908 54 13924 80 1 FreeSans 160 0 0 0 C26
port 21 n
flabel metal2 15448 54 15464 80 1 FreeSans 160 0 0 0 C27
port 22 n
flabel metal2 16982 64 16998 90 1 FreeSans 160 0 0 0 C28
port 23 n
flabel metal2 18534 50 18550 76 1 FreeSans 160 0 0 0 C29
port 24 n
flabel metal2 20080 48 20096 74 1 FreeSans 160 0 0 0 C30
port 25 n
flabel metal2 21612 54 21628 80 1 FreeSans 160 0 0 0 C31
port 26 n
flabel metal2 23152 64 23168 90 1 FreeSans 160 0 0 0 C32
port 27 n
<< end >>
