magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1174 157 1356 201
rect 1659 157 2023 203
rect 1 145 824 157
rect 1028 145 2023 157
rect 1 21 2023 145
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 355 47 385 131
rect 456 47 486 131
rect 534 47 564 131
rect 630 47 660 131
rect 706 47 736 131
rect 910 47 940 119
rect 1006 47 1036 119
rect 1104 47 1134 131
rect 1250 47 1280 175
rect 1351 47 1381 119
rect 1454 47 1484 119
rect 1549 47 1579 131
rect 1737 47 1767 177
rect 1828 47 1858 177
rect 1912 47 1942 177
<< scpmoshvt >>
rect 80 363 110 491
rect 164 363 194 491
rect 352 369 382 497
rect 437 369 467 497
rect 529 369 559 497
rect 613 369 643 497
rect 706 369 736 497
rect 909 413 939 497
rect 1002 413 1032 497
rect 1098 413 1128 497
rect 1230 347 1260 497
rect 1325 413 1355 497
rect 1409 413 1439 497
rect 1526 413 1556 497
rect 1737 297 1767 497
rect 1828 297 1858 497
rect 1912 297 1942 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 89 355 131
rect 299 55 311 89
rect 345 55 355 89
rect 299 47 355 55
rect 385 89 456 131
rect 385 55 411 89
rect 445 55 456 89
rect 385 47 456 55
rect 486 47 534 131
rect 564 89 630 131
rect 564 55 585 89
rect 619 55 630 89
rect 564 47 630 55
rect 660 47 706 131
rect 736 89 798 131
rect 1200 131 1250 175
rect 1054 119 1104 131
rect 736 55 752 89
rect 786 55 798 89
rect 736 47 798 55
rect 854 107 910 119
rect 854 73 862 107
rect 896 73 910 107
rect 854 47 910 73
rect 940 107 1006 119
rect 940 73 962 107
rect 996 73 1006 107
rect 940 47 1006 73
rect 1036 47 1104 119
rect 1134 101 1250 131
rect 1134 67 1178 101
rect 1212 67 1250 101
rect 1134 47 1250 67
rect 1280 119 1330 175
rect 1685 162 1737 177
rect 1499 119 1549 131
rect 1280 107 1351 119
rect 1280 73 1296 107
rect 1330 73 1351 107
rect 1280 47 1351 73
rect 1381 107 1454 119
rect 1381 73 1408 107
rect 1442 73 1454 107
rect 1381 47 1454 73
rect 1484 47 1549 119
rect 1579 107 1631 131
rect 1579 73 1589 107
rect 1623 73 1631 107
rect 1579 47 1631 73
rect 1685 128 1693 162
rect 1727 128 1737 162
rect 1685 94 1737 128
rect 1685 60 1693 94
rect 1727 60 1737 94
rect 1685 47 1737 60
rect 1767 123 1828 177
rect 1767 89 1781 123
rect 1815 89 1828 123
rect 1767 47 1828 89
rect 1858 164 1912 177
rect 1858 130 1868 164
rect 1902 130 1912 164
rect 1858 96 1912 130
rect 1858 62 1868 96
rect 1902 62 1912 96
rect 1858 47 1912 62
rect 1942 164 1997 177
rect 1942 130 1955 164
rect 1989 130 1997 164
rect 1942 96 1997 130
rect 1942 62 1955 96
rect 1989 62 1997 96
rect 1942 47 1997 62
<< pdiff >>
rect 28 477 80 491
rect 28 443 36 477
rect 70 443 80 477
rect 28 409 80 443
rect 28 375 36 409
rect 70 375 80 409
rect 28 363 80 375
rect 110 461 164 491
rect 110 427 120 461
rect 154 427 164 461
rect 110 363 164 427
rect 194 477 246 491
rect 194 443 204 477
rect 238 443 246 477
rect 194 409 246 443
rect 194 375 204 409
rect 238 375 246 409
rect 194 363 246 375
rect 300 452 352 497
rect 300 418 308 452
rect 342 418 352 452
rect 300 369 352 418
rect 382 483 437 497
rect 382 449 392 483
rect 426 449 437 483
rect 382 369 437 449
rect 467 369 529 497
rect 559 483 613 497
rect 559 449 569 483
rect 603 449 613 483
rect 559 369 613 449
rect 643 369 706 497
rect 736 483 793 497
rect 736 449 751 483
rect 785 449 793 483
rect 736 369 793 449
rect 847 472 909 497
rect 847 438 855 472
rect 889 438 909 472
rect 847 413 909 438
rect 939 472 1002 497
rect 939 438 954 472
rect 988 438 1002 472
rect 939 413 1002 438
rect 1032 413 1098 497
rect 1128 485 1230 497
rect 1128 451 1186 485
rect 1220 451 1230 485
rect 1128 417 1230 451
rect 1128 413 1186 417
rect 1143 383 1186 413
rect 1220 383 1230 417
rect 1143 347 1230 383
rect 1260 477 1325 497
rect 1260 443 1270 477
rect 1304 443 1325 477
rect 1260 413 1325 443
rect 1355 467 1409 497
rect 1355 433 1365 467
rect 1399 433 1409 467
rect 1355 413 1409 433
rect 1439 413 1526 497
rect 1556 477 1631 497
rect 1556 443 1588 477
rect 1622 443 1631 477
rect 1556 413 1631 443
rect 1685 475 1737 497
rect 1685 441 1693 475
rect 1727 441 1737 475
rect 1260 347 1310 413
rect 1685 353 1737 441
rect 1685 319 1693 353
rect 1727 319 1737 353
rect 1685 297 1737 319
rect 1767 455 1828 497
rect 1767 421 1781 455
rect 1815 421 1828 455
rect 1767 375 1828 421
rect 1767 341 1781 375
rect 1815 341 1828 375
rect 1767 297 1828 341
rect 1858 479 1912 497
rect 1858 445 1868 479
rect 1902 445 1912 479
rect 1858 411 1912 445
rect 1858 377 1868 411
rect 1902 377 1912 411
rect 1858 343 1912 377
rect 1858 309 1868 343
rect 1902 309 1912 343
rect 1858 297 1912 309
rect 1942 479 1997 497
rect 1942 445 1955 479
rect 1989 445 1997 479
rect 1942 411 1997 445
rect 1942 377 1955 411
rect 1989 377 1997 411
rect 1942 343 1997 377
rect 1942 309 1955 343
rect 1989 309 1997 343
rect 1942 297 1997 309
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 311 55 345 89
rect 411 55 445 89
rect 585 55 619 89
rect 752 55 786 89
rect 862 73 896 107
rect 962 73 996 107
rect 1178 67 1212 101
rect 1296 73 1330 107
rect 1408 73 1442 107
rect 1589 73 1623 107
rect 1693 128 1727 162
rect 1693 60 1727 94
rect 1781 89 1815 123
rect 1868 130 1902 164
rect 1868 62 1902 96
rect 1955 130 1989 164
rect 1955 62 1989 96
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 120 427 154 461
rect 204 443 238 477
rect 204 375 238 409
rect 308 418 342 452
rect 392 449 426 483
rect 569 449 603 483
rect 751 449 785 483
rect 855 438 889 472
rect 954 438 988 472
rect 1186 451 1220 485
rect 1186 383 1220 417
rect 1270 443 1304 477
rect 1365 433 1399 467
rect 1588 443 1622 477
rect 1693 441 1727 475
rect 1693 319 1727 353
rect 1781 421 1815 455
rect 1781 341 1815 375
rect 1868 445 1902 479
rect 1868 377 1902 411
rect 1868 309 1902 343
rect 1955 445 1989 479
rect 1955 377 1989 411
rect 1955 309 1989 343
<< poly >>
rect 80 491 110 517
rect 164 491 194 517
rect 352 497 382 523
rect 437 497 467 523
rect 529 497 559 523
rect 613 497 643 523
rect 706 497 736 523
rect 909 497 939 523
rect 1002 497 1032 523
rect 1098 497 1128 523
rect 1230 497 1260 523
rect 1325 497 1355 523
rect 1409 497 1439 523
rect 1526 497 1556 523
rect 1737 497 1767 523
rect 1828 497 1858 523
rect 1912 497 1942 523
rect 909 375 939 413
rect 1002 381 1032 413
rect 80 348 110 363
rect 47 318 110 348
rect 47 265 77 318
rect 164 274 194 363
rect 352 331 382 369
rect 437 331 467 369
rect 529 337 559 369
rect 613 337 643 369
rect 340 321 467 331
rect 340 287 356 321
rect 390 301 467 321
rect 514 321 568 337
rect 390 287 406 301
rect 340 277 406 287
rect 514 287 524 321
rect 558 287 568 321
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 119 264 194 274
rect 119 230 135 264
rect 169 230 194 264
rect 119 220 194 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 354 166 384 277
rect 514 271 568 287
rect 610 321 664 337
rect 610 287 620 321
rect 654 287 664 321
rect 610 271 664 287
rect 706 304 736 369
rect 894 365 960 375
rect 894 331 910 365
rect 944 331 960 365
rect 894 321 960 331
rect 1002 365 1056 381
rect 1002 331 1012 365
rect 1046 331 1056 365
rect 1002 315 1056 331
rect 706 288 760 304
rect 426 225 492 235
rect 426 191 442 225
rect 476 191 492 225
rect 426 181 492 191
rect 354 157 385 166
rect 355 131 385 157
rect 456 131 486 181
rect 534 131 564 271
rect 706 254 716 288
rect 750 254 760 288
rect 1002 279 1032 315
rect 706 238 760 254
rect 910 249 1032 279
rect 606 207 660 223
rect 606 173 616 207
rect 650 173 660 207
rect 606 157 660 173
rect 630 131 660 157
rect 706 131 736 238
rect 910 119 940 249
rect 1098 213 1128 413
rect 1230 309 1260 347
rect 1325 315 1355 413
rect 1409 375 1439 413
rect 1526 381 1556 413
rect 1408 365 1474 375
rect 1408 331 1424 365
rect 1458 331 1474 365
rect 1408 321 1474 331
rect 1526 365 1604 381
rect 1526 331 1560 365
rect 1594 331 1604 365
rect 1526 315 1604 331
rect 1170 299 1260 309
rect 1170 265 1186 299
rect 1220 265 1260 299
rect 1170 255 1260 265
rect 1230 220 1260 255
rect 1312 299 1366 315
rect 1312 265 1322 299
rect 1356 279 1366 299
rect 1356 265 1484 279
rect 1312 249 1484 265
rect 982 191 1036 207
rect 982 157 992 191
rect 1026 157 1036 191
rect 1098 203 1178 213
rect 1098 183 1128 203
rect 982 141 1036 157
rect 1006 119 1036 141
rect 1104 169 1128 183
rect 1162 169 1178 203
rect 1230 190 1280 220
rect 1250 175 1280 190
rect 1351 191 1412 207
rect 1104 159 1178 169
rect 1104 131 1134 159
rect 1351 157 1368 191
rect 1402 157 1412 191
rect 1351 141 1412 157
rect 1351 119 1381 141
rect 1454 119 1484 249
rect 1549 131 1579 315
rect 1737 265 1767 297
rect 1828 265 1858 297
rect 1912 265 1942 297
rect 1635 249 1767 265
rect 1635 215 1645 249
rect 1679 215 1767 249
rect 1635 199 1767 215
rect 1809 249 1942 265
rect 1809 215 1819 249
rect 1853 215 1942 249
rect 1809 199 1942 215
rect 1737 177 1767 199
rect 1828 177 1858 199
rect 1912 177 1942 199
rect 79 21 109 47
rect 163 21 193 47
rect 355 21 385 47
rect 456 21 486 47
rect 534 21 564 47
rect 630 21 660 47
rect 706 21 736 47
rect 910 21 940 47
rect 1006 21 1036 47
rect 1104 21 1134 47
rect 1250 21 1280 47
rect 1351 21 1381 47
rect 1454 21 1484 47
rect 1549 21 1579 47
rect 1737 21 1767 47
rect 1828 21 1858 47
rect 1912 21 1942 47
<< polycont >>
rect 356 287 390 321
rect 524 287 558 321
rect 33 215 67 249
rect 135 230 169 264
rect 620 287 654 321
rect 910 331 944 365
rect 1012 331 1046 365
rect 442 191 476 225
rect 716 254 750 288
rect 616 173 650 207
rect 1424 331 1458 365
rect 1560 331 1594 365
rect 1186 265 1220 299
rect 1322 265 1356 299
rect 992 157 1026 191
rect 1128 169 1162 203
rect 1368 157 1402 191
rect 1645 215 1679 249
rect 1819 215 1853 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 36 477 70 493
rect 36 409 70 443
rect 104 461 170 527
rect 104 427 120 461
rect 154 427 170 461
rect 204 477 249 493
rect 238 443 249 477
rect 204 409 249 443
rect 70 391 169 393
rect 70 375 128 391
rect 36 359 128 375
rect 123 357 128 359
rect 162 357 169 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 123 264 169 357
rect 123 230 135 264
rect 123 194 169 230
rect 238 375 249 409
rect 123 161 162 194
rect 35 127 162 161
rect 204 187 249 375
rect 204 153 210 187
rect 244 153 249 187
rect 204 143 249 153
rect 35 119 69 127
rect 203 119 249 143
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 249 119
rect 203 69 249 85
rect 287 452 342 489
rect 287 418 308 452
rect 376 483 442 527
rect 751 483 785 527
rect 376 449 392 483
rect 426 449 442 483
rect 538 449 569 483
rect 603 449 717 483
rect 287 415 342 418
rect 287 372 649 415
rect 287 89 321 372
rect 356 321 390 337
rect 356 157 390 287
rect 424 225 458 372
rect 615 337 649 372
rect 683 399 717 449
rect 751 433 785 449
rect 842 472 889 488
rect 1186 485 1220 527
rect 842 438 855 472
rect 938 438 954 472
rect 988 438 1152 472
rect 842 413 889 438
rect 842 399 876 413
rect 683 365 876 399
rect 996 391 1084 402
rect 492 321 558 337
rect 492 287 524 321
rect 492 271 558 287
rect 615 321 654 337
rect 615 287 620 321
rect 615 271 654 287
rect 706 288 804 331
rect 706 254 716 288
rect 750 254 804 288
rect 424 191 442 225
rect 476 191 492 225
rect 616 207 650 223
rect 706 207 804 254
rect 842 173 876 365
rect 616 157 650 173
rect 356 123 650 157
rect 684 139 876 173
rect 910 365 958 381
rect 944 331 958 365
rect 996 365 1041 391
rect 996 331 1012 365
rect 1075 357 1084 391
rect 1046 331 1084 357
rect 910 207 958 331
rect 1118 315 1152 438
rect 1186 417 1220 451
rect 1186 367 1220 383
rect 1254 477 1304 493
rect 1254 443 1270 477
rect 1562 477 1623 527
rect 1254 427 1304 443
rect 1349 433 1365 467
rect 1399 433 1526 467
rect 1118 299 1220 315
rect 1118 297 1186 299
rect 1060 265 1186 297
rect 1060 263 1220 265
rect 910 191 1026 207
rect 910 187 992 191
rect 910 153 949 187
rect 983 157 992 187
rect 983 153 1026 157
rect 910 141 1026 153
rect 103 17 169 59
rect 287 55 311 89
rect 345 55 361 89
rect 395 55 411 89
rect 445 55 461 89
rect 495 61 530 123
rect 684 89 718 139
rect 842 107 876 139
rect 1060 107 1094 263
rect 1186 249 1220 263
rect 1128 213 1162 219
rect 1254 213 1288 427
rect 1322 391 1360 393
rect 1322 357 1324 391
rect 1358 357 1360 391
rect 1322 299 1360 357
rect 1356 265 1360 299
rect 1322 249 1360 265
rect 1394 365 1458 381
rect 1394 331 1424 365
rect 1394 315 1458 331
rect 1128 203 1288 213
rect 1394 207 1432 315
rect 1492 281 1526 433
rect 1562 443 1588 477
rect 1622 443 1623 477
rect 1562 427 1623 443
rect 1693 475 1747 491
rect 1727 441 1747 475
rect 1693 381 1747 441
rect 1560 365 1747 381
rect 1594 353 1747 365
rect 1594 331 1693 353
rect 1560 319 1693 331
rect 1727 319 1747 353
rect 1781 455 1816 527
rect 1955 479 1989 527
rect 1815 421 1816 455
rect 1781 375 1816 421
rect 1815 341 1816 375
rect 1781 325 1816 341
rect 1852 445 1868 479
rect 1902 445 1921 479
rect 1852 411 1921 445
rect 1852 377 1868 411
rect 1902 377 1921 411
rect 1852 343 1921 377
rect 1560 315 1747 319
rect 1162 169 1288 203
rect 1128 153 1288 169
rect 564 55 585 89
rect 619 55 718 89
rect 752 89 792 105
rect 786 55 792 89
rect 842 73 862 107
rect 896 73 912 107
rect 946 73 962 107
rect 996 73 1094 107
rect 1144 101 1218 117
rect 395 17 461 55
rect 752 17 792 55
rect 1144 67 1178 101
rect 1212 67 1218 101
rect 1254 107 1288 153
rect 1322 191 1432 207
rect 1322 187 1368 191
rect 1322 153 1326 187
rect 1360 157 1368 187
rect 1402 157 1432 191
rect 1360 153 1432 157
rect 1322 141 1432 153
rect 1466 265 1526 281
rect 1713 265 1747 315
rect 1852 309 1868 343
rect 1902 309 1921 343
rect 1852 301 1921 309
rect 1466 249 1679 265
rect 1466 215 1645 249
rect 1466 199 1679 215
rect 1713 249 1853 265
rect 1713 215 1819 249
rect 1713 199 1853 215
rect 1466 107 1500 199
rect 1713 165 1747 199
rect 1677 162 1747 165
rect 1887 164 1921 301
rect 1955 411 1989 445
rect 1955 343 1989 377
rect 1955 281 1989 309
rect 1677 128 1693 162
rect 1727 128 1747 162
rect 1254 73 1296 107
rect 1330 73 1346 107
rect 1392 73 1408 107
rect 1442 73 1500 107
rect 1549 107 1623 123
rect 1549 73 1589 107
rect 1144 17 1218 67
rect 1549 17 1623 73
rect 1677 94 1747 128
rect 1677 60 1693 94
rect 1727 60 1747 94
rect 1781 123 1815 139
rect 1781 17 1815 89
rect 1852 130 1868 164
rect 1902 130 1921 164
rect 1852 96 1921 130
rect 1852 62 1868 96
rect 1902 62 1921 96
rect 1852 61 1921 62
rect 1955 164 1989 186
rect 1955 96 1989 130
rect 1955 17 1989 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 128 357 162 391
rect 210 153 244 187
rect 1041 365 1075 391
rect 1041 357 1046 365
rect 1046 357 1075 365
rect 949 153 983 187
rect 1324 357 1358 391
rect 1326 153 1360 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 116 391 174 397
rect 116 357 128 391
rect 162 388 174 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 162 360 1041 388
rect 162 357 174 360
rect 116 351 174 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1312 391 1370 397
rect 1312 388 1324 391
rect 1075 360 1324 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1312 357 1324 360
rect 1358 357 1370 391
rect 1312 351 1370 357
rect 198 187 256 193
rect 198 153 210 187
rect 244 184 256 187
rect 937 187 995 193
rect 937 184 949 187
rect 244 156 949 184
rect 244 153 256 156
rect 198 147 256 153
rect 937 153 949 156
rect 983 184 995 187
rect 1314 187 1372 193
rect 1314 184 1326 187
rect 983 156 1326 184
rect 983 153 995 156
rect 937 147 995 153
rect 1314 153 1326 156
rect 1360 153 1372 187
rect 1314 147 1372 153
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 765 221 799 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew signal input
flabel locali s 501 289 535 323 0 FreeSans 300 0 0 0 D
port 2 nsew signal input
flabel locali s 495 85 529 119 0 FreeSans 300 0 0 0 SCE
port 4 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1869 85 1903 119 0 FreeSans 200 0 0 0 Q
port 9 nsew signal output
flabel locali s 1869 357 1903 391 0 FreeSans 200 0 0 0 Q
port 9 nsew signal output
flabel locali s 1869 425 1903 459 0 FreeSans 200 0 0 0 Q
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
port 7 nsew
rlabel comment s 0 0 0 0 4 sdfxtp_2
rlabel metal1 s 0 -48 2024 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 392160
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 376362
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 10.120 0.000 
<< end >>
