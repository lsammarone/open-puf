magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 67 1074 203
rect 1 21 886 67
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 526 47 556 177
rect 610 47 640 177
rect 694 47 724 177
rect 778 47 808 177
rect 966 93 996 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 526 297 556 497
rect 610 297 640 497
rect 694 297 724 497
rect 778 297 808 497
rect 966 413 996 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 163 177
rect 109 129 119 163
rect 153 129 163 163
rect 109 95 163 129
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 95 247 177
rect 193 61 203 95
rect 237 61 247 95
rect 193 47 247 61
rect 277 163 331 177
rect 277 129 287 163
rect 321 129 331 163
rect 277 95 331 129
rect 277 61 287 95
rect 321 61 331 95
rect 277 47 331 61
rect 361 95 413 177
rect 361 61 371 95
rect 405 61 413 95
rect 361 47 413 61
rect 474 95 526 177
rect 474 61 482 95
rect 516 61 526 95
rect 474 47 526 61
rect 556 163 610 177
rect 556 129 566 163
rect 600 129 610 163
rect 556 95 610 129
rect 556 61 566 95
rect 600 61 610 95
rect 556 47 610 61
rect 640 95 694 177
rect 640 61 650 95
rect 684 61 694 95
rect 640 47 694 61
rect 724 163 778 177
rect 724 129 734 163
rect 768 129 778 163
rect 724 95 778 129
rect 724 61 734 95
rect 768 61 778 95
rect 724 47 778 61
rect 808 163 860 177
rect 808 129 818 163
rect 852 129 860 163
rect 808 95 860 129
rect 808 61 818 95
rect 852 61 860 95
rect 914 149 966 177
rect 914 115 922 149
rect 956 115 966 149
rect 914 93 966 115
rect 996 149 1048 177
rect 996 115 1006 149
rect 1040 115 1048 149
rect 996 93 1048 115
rect 808 47 860 61
<< pdiff >>
rect 27 479 79 497
rect 27 445 35 479
rect 69 445 79 479
rect 27 411 79 445
rect 27 377 35 411
rect 69 377 79 411
rect 27 343 79 377
rect 27 309 35 343
rect 69 309 79 343
rect 27 297 79 309
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 341 247 375
rect 193 307 203 341
rect 237 307 247 341
rect 193 297 247 307
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 411 413 497
rect 361 377 371 411
rect 405 377 413 411
rect 361 343 413 377
rect 361 309 371 343
rect 405 309 413 343
rect 361 297 413 309
rect 474 411 526 497
rect 474 377 482 411
rect 516 377 526 411
rect 474 343 526 377
rect 474 309 482 343
rect 516 309 526 343
rect 474 297 526 309
rect 556 477 610 497
rect 556 443 566 477
rect 600 443 610 477
rect 556 409 610 443
rect 556 375 566 409
rect 600 375 610 409
rect 556 297 610 375
rect 640 477 694 497
rect 640 443 650 477
rect 684 443 694 477
rect 640 409 694 443
rect 640 375 650 409
rect 684 375 694 409
rect 640 341 694 375
rect 640 307 650 341
rect 684 307 694 341
rect 640 297 694 307
rect 724 409 778 497
rect 724 375 734 409
rect 768 375 778 409
rect 724 341 778 375
rect 724 307 734 341
rect 768 307 778 341
rect 724 297 778 307
rect 808 477 860 497
rect 808 443 818 477
rect 852 443 860 477
rect 808 409 860 443
rect 914 474 966 497
rect 914 440 922 474
rect 956 440 966 474
rect 914 413 966 440
rect 996 477 1048 497
rect 996 443 1006 477
rect 1040 443 1048 477
rect 996 413 1048 443
rect 808 375 818 409
rect 852 375 860 409
rect 808 297 860 375
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 119 129 153 163
rect 119 61 153 95
rect 203 61 237 95
rect 287 129 321 163
rect 287 61 321 95
rect 371 61 405 95
rect 482 61 516 95
rect 566 129 600 163
rect 566 61 600 95
rect 650 61 684 95
rect 734 129 768 163
rect 734 61 768 95
rect 818 129 852 163
rect 818 61 852 95
rect 922 115 956 149
rect 1006 115 1040 149
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 119 443 153 477
rect 119 375 153 409
rect 203 443 237 477
rect 203 375 237 409
rect 203 307 237 341
rect 287 443 321 477
rect 287 375 321 409
rect 371 377 405 411
rect 371 309 405 343
rect 482 377 516 411
rect 482 309 516 343
rect 566 443 600 477
rect 566 375 600 409
rect 650 443 684 477
rect 650 375 684 409
rect 650 307 684 341
rect 734 375 768 409
rect 734 307 768 341
rect 818 443 852 477
rect 922 440 956 474
rect 1006 443 1040 477
rect 818 375 852 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 526 497 556 523
rect 610 497 640 523
rect 694 497 724 523
rect 778 497 808 523
rect 966 497 996 523
rect 79 265 109 297
rect 163 265 193 297
rect 79 249 193 265
rect 79 215 108 249
rect 142 215 193 249
rect 79 199 193 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 265 277 297
rect 331 265 361 297
rect 247 249 361 265
rect 247 215 300 249
rect 334 215 361 249
rect 247 199 361 215
rect 247 177 277 199
rect 331 177 361 199
rect 526 265 556 297
rect 610 265 640 297
rect 526 249 640 265
rect 526 215 579 249
rect 613 215 640 249
rect 526 199 640 215
rect 526 177 556 199
rect 610 177 640 199
rect 694 265 724 297
rect 778 265 808 297
rect 966 265 996 413
rect 694 249 924 265
rect 694 215 880 249
rect 914 215 924 249
rect 694 199 924 215
rect 966 249 1021 265
rect 966 215 977 249
rect 1011 215 1021 249
rect 966 199 1021 215
rect 694 177 724 199
rect 778 177 808 199
rect 966 177 996 199
rect 966 67 996 93
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 526 21 556 47
rect 610 21 640 47
rect 694 21 724 47
rect 778 21 808 47
<< polycont >>
rect 108 215 142 249
rect 300 215 334 249
rect 579 215 613 249
rect 880 215 914 249
rect 977 215 1011 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 17 479 85 493
rect 17 445 35 479
rect 69 445 85 479
rect 17 411 85 445
rect 17 377 35 411
rect 69 377 85 411
rect 17 343 85 377
rect 119 477 161 527
rect 153 443 161 477
rect 119 409 161 443
rect 153 375 161 409
rect 119 359 161 375
rect 195 477 245 493
rect 195 443 203 477
rect 237 443 245 477
rect 195 409 245 443
rect 195 375 203 409
rect 237 375 245 409
rect 17 309 35 343
rect 69 325 85 343
rect 195 341 245 375
rect 279 477 608 493
rect 279 443 287 477
rect 321 459 566 477
rect 279 409 321 443
rect 600 443 608 477
rect 279 375 287 409
rect 279 359 321 375
rect 355 411 421 425
rect 355 377 371 411
rect 405 377 421 411
rect 195 325 203 341
rect 69 309 203 325
rect 17 307 203 309
rect 237 325 245 341
rect 355 343 421 377
rect 355 325 371 343
rect 237 309 371 325
rect 405 309 421 343
rect 237 307 421 309
rect 17 291 421 307
rect 455 411 532 425
rect 455 377 482 411
rect 516 377 532 411
rect 455 343 532 377
rect 566 409 608 443
rect 600 375 608 409
rect 566 359 608 375
rect 642 477 859 493
rect 642 443 650 477
rect 684 459 818 477
rect 684 443 692 459
rect 642 409 692 443
rect 810 443 818 459
rect 852 443 859 477
rect 642 375 650 409
rect 684 375 692 409
rect 455 309 482 343
rect 516 325 532 343
rect 642 341 692 375
rect 642 325 650 341
rect 516 309 650 325
rect 455 307 650 309
rect 684 307 692 341
rect 455 291 692 307
rect 726 409 776 425
rect 726 375 734 409
rect 768 375 776 409
rect 726 341 776 375
rect 810 409 859 443
rect 810 375 818 409
rect 852 375 859 409
rect 810 359 859 375
rect 893 474 964 490
rect 893 440 922 474
rect 956 440 964 474
rect 893 407 964 440
rect 998 477 1048 527
rect 998 443 1006 477
rect 1040 443 1048 477
rect 998 427 1048 443
rect 726 307 734 341
rect 768 325 776 341
rect 768 307 807 325
rect 726 291 807 307
rect 20 249 248 257
rect 20 215 108 249
rect 142 215 248 249
rect 284 249 527 257
rect 284 215 300 249
rect 334 215 527 249
rect 563 249 707 257
rect 563 215 579 249
rect 613 215 707 249
rect 743 215 807 291
rect 893 249 927 407
rect 1037 257 1087 391
rect 864 215 880 249
rect 914 215 927 249
rect 961 249 1087 257
rect 961 215 977 249
rect 1011 215 1087 249
rect 743 181 784 215
rect 17 163 69 181
rect 17 129 35 163
rect 17 95 69 129
rect 17 61 35 95
rect 17 17 69 61
rect 103 163 784 181
rect 893 181 927 215
rect 103 129 119 163
rect 153 145 287 163
rect 153 129 169 145
rect 103 95 169 129
rect 271 129 287 145
rect 321 145 566 163
rect 321 129 337 145
rect 103 61 119 95
rect 153 61 169 95
rect 103 51 169 61
rect 203 95 237 111
rect 203 17 237 61
rect 271 95 337 129
rect 550 129 566 145
rect 600 145 734 163
rect 600 129 616 145
rect 271 61 287 95
rect 321 61 337 95
rect 271 51 337 61
rect 371 95 516 111
rect 405 61 482 95
rect 371 17 516 61
rect 550 95 616 129
rect 718 129 734 145
rect 768 129 784 163
rect 550 61 566 95
rect 600 61 616 95
rect 550 51 616 61
rect 650 95 684 111
rect 650 17 684 61
rect 718 95 784 129
rect 718 61 734 95
rect 768 61 784 95
rect 718 51 784 61
rect 818 163 859 179
rect 852 129 859 163
rect 818 95 859 129
rect 852 61 859 95
rect 893 149 964 181
rect 893 115 922 149
rect 956 115 964 149
rect 893 76 964 115
rect 998 149 1048 165
rect 998 115 1006 149
rect 1040 115 1048 149
rect 818 17 859 61
rect 998 17 1048 115
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
flabel locali s 1041 221 1075 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 765 289 799 323 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 581 221 615 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 118 221 152 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 302 221 336 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor4b_2
rlabel metal1 s 0 -48 1104 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1104 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string GDS_END 1186068
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1176798
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.520 0.000 
<< end >>
