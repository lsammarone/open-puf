/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/cdl/sky130_fd_sc_hvl.cdl