magic
tech sky130A
magscale 1 2
timestamp 1649788711
<< nwell >>
rect -294 -1390 294 1390
<< pmoslvt >>
rect -200 -1290 200 1290
<< pdiff >>
rect -258 1278 -200 1290
rect -258 -1278 -246 1278
rect -212 -1278 -200 1278
rect -258 -1290 -200 -1278
rect 200 1278 258 1290
rect 200 -1278 212 1278
rect 246 -1278 258 1278
rect 200 -1290 258 -1278
<< pdiffc >>
rect -246 -1278 -212 1278
rect 212 -1278 246 1278
<< poly >>
rect -126 1371 126 1387
rect -126 1354 -110 1371
rect -200 1337 -110 1354
rect 110 1354 126 1371
rect 110 1337 200 1354
rect -200 1290 200 1337
rect -200 -1337 200 -1290
rect -200 -1354 -110 -1337
rect -126 -1371 -110 -1354
rect 110 -1354 200 -1337
rect 110 -1371 126 -1354
rect -126 -1387 126 -1371
<< polycont >>
rect -110 1337 110 1371
rect -110 -1371 110 -1337
<< locali >>
rect -126 1337 -110 1371
rect 110 1337 126 1371
rect -246 1278 -212 1294
rect -246 -1294 -212 -1278
rect 212 1278 246 1294
rect 212 -1294 246 -1278
rect -126 -1371 -110 -1337
rect 110 -1371 126 -1337
<< viali >>
rect -74 1337 74 1371
rect -246 -1278 -212 1278
rect 212 -1278 246 1278
rect -74 -1371 74 -1337
<< metal1 >>
rect -86 1371 86 1377
rect -86 1337 -74 1371
rect 74 1337 86 1371
rect -86 1331 86 1337
rect -252 1278 -206 1290
rect -252 -1278 -246 1278
rect -212 -1278 -206 1278
rect -252 -1290 -206 -1278
rect 206 1278 252 1290
rect 206 -1278 212 1278
rect 246 -1278 252 1278
rect 206 -1290 252 -1278
rect -86 -1337 86 -1331
rect -86 -1371 -74 -1337
rect 74 -1371 86 -1337
rect -86 -1377 86 -1371
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 12.9 l 2 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
