magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1063 203
rect 29 -17 63 21
<< locali >>
rect 125 351 159 437
rect 297 351 347 437
rect 29 317 347 351
rect 29 157 126 317
rect 479 199 541 305
rect 729 302 987 336
rect 729 255 764 302
rect 937 258 987 302
rect 685 202 764 255
rect 798 202 903 255
rect 937 211 1020 258
rect 29 123 347 157
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 23 387 89 527
rect 195 387 261 527
rect 383 303 433 527
rect 491 459 693 493
rect 491 339 525 459
rect 160 199 441 265
rect 407 157 441 199
rect 575 168 609 425
rect 657 404 693 459
rect 727 455 793 527
rect 827 404 861 493
rect 895 455 961 527
rect 1006 404 1072 479
rect 657 370 1072 404
rect 657 289 693 370
rect 1021 292 1072 370
rect 575 157 873 168
rect 407 134 873 157
rect 407 123 609 134
rect 21 17 89 89
rect 195 17 261 89
rect 382 17 537 89
rect 575 51 609 123
rect 651 17 717 89
rect 817 81 873 134
rect 989 17 1045 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 798 202 903 255 6 A1
port 1 nsew signal input
rlabel locali s 937 211 1020 258 6 A2
port 2 nsew signal input
rlabel locali s 937 258 987 302 6 A2
port 2 nsew signal input
rlabel locali s 685 202 764 255 6 A2
port 2 nsew signal input
rlabel locali s 729 255 764 302 6 A2
port 2 nsew signal input
rlabel locali s 729 302 987 336 6 A2
port 2 nsew signal input
rlabel locali s 479 199 541 305 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1063 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 29 123 347 157 6 X
port 8 nsew signal output
rlabel locali s 29 157 126 317 6 X
port 8 nsew signal output
rlabel locali s 29 317 347 351 6 X
port 8 nsew signal output
rlabel locali s 297 351 347 437 6 X
port 8 nsew signal output
rlabel locali s 125 351 159 437 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4096876
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4088712
<< end >>
