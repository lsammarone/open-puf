magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -83 34709 16087 35795
rect -83 34095 1503 34709
rect 13394 34095 16087 34709
rect -83 34046 16087 34095
rect -83 33703 16088 34046
rect -83 29338 1277 33703
rect 15726 29338 16088 33703
rect -83 28976 16088 29338
rect 9208 28076 16088 28077
rect -83 26133 16088 28076
rect 9388 18849 16134 19033
rect 12530 18747 16134 18849
rect -83 18364 559 18480
rect -83 17697 1195 18364
rect -24 17656 1195 17697
rect -24 17548 1684 17656
rect -24 17332 1699 17548
rect -24 17116 906 17332
rect 15848 16869 16134 18747
rect 9388 16633 16134 16869
rect -143 15961 4963 16247
rect -143 12468 143 15961
rect 15848 14755 16134 16633
rect 12530 14653 16134 14755
rect 9388 14519 16134 14653
rect 15825 13209 16134 14519
rect 14067 13039 16134 13209
rect -143 12204 762 12468
rect -143 12154 2707 12204
rect -143 12036 2092 12154
rect -143 11604 143 12036
rect -143 11318 4703 11604
rect 15825 10410 16134 13039
rect 14067 10124 16134 10410
rect 9783 6853 16090 7211
rect 11655 6482 16090 6853
rect 12966 5957 16090 6482
rect 12966 4616 16090 5069
rect 916 3831 16090 4616
rect -83 1133 622 1865
<< pwell >>
rect -58 28137 16058 28913
rect -43 25863 8049 26071
rect 13382 25863 16058 26071
rect -43 25027 16058 25863
rect -43 20710 1147 25027
rect 15573 20710 16058 25027
rect -43 20393 16058 20710
rect -43 19251 1043 20393
rect 7877 20164 16058 20393
rect 10576 19904 16058 20164
rect 15354 19597 16058 19904
rect 7877 19251 16058 19597
rect -43 19195 16058 19251
rect -43 19052 9168 19195
rect -43 18991 9318 19052
rect -43 18587 1860 18991
<< obsli1 >>
rect 0 35729 16000 39941
rect -17 34018 16021 35729
rect -23 29043 16021 34018
rect -23 29031 16000 29043
rect 0 28887 16000 29031
rect -32 28163 16032 28887
rect 0 28030 16000 28163
rect -23 28011 16000 28030
rect -23 26255 16017 28011
rect -17 26199 16017 26255
rect 0 26045 16000 26199
rect -17 26044 16032 26045
rect -23 19221 16032 26044
rect -23 19179 16000 19221
rect -17 18916 16000 19179
rect -17 18613 16017 18916
rect 0 18414 16017 18613
rect -17 17763 16017 18414
rect 0 16121 16017 17763
rect -17 11444 16017 16121
rect 0 10250 16017 11444
rect 0 7145 16000 10250
rect 0 6023 16024 7145
rect 0 5003 16000 6023
rect 0 3897 16024 5003
rect 0 1799 16000 3897
rect -17 1199 16000 1799
rect 0 46 16000 1199
<< metal1 >>
rect 12486 0 12538 261
<< obsm1 >>
rect 0 36195 16000 40000
rect 0 35780 16004 36195
rect 0 34018 16000 35780
rect -23 26255 16029 34018
rect 0 26044 16000 26255
rect -23 19179 16029 26044
rect 0 18916 16000 19179
rect 0 18296 16012 18916
rect -29 17950 16012 18296
rect 0 16127 16012 17950
rect -23 14586 16012 16127
tri 16012 14586 16023 14597 sw
rect -23 11438 16023 14586
rect 0 10244 16023 11438
rect 0 7145 16000 10244
rect 0 6024 16023 7145
rect 0 5003 16000 6024
rect 0 3897 16023 5003
rect 0 317 16000 3897
rect 0 52 12430 317
rect 12594 52 16000 317
<< metal2 >>
rect 675 0 721 895
rect 1084 0 1130 895
rect 1226 0 1278 310
rect 2551 0 2603 1070
rect 3262 0 3314 464
rect 4471 0 4523 1285
rect 5320 0 5372 541
rect 5698 0 5750 814
rect 6150 0 6202 453
rect 6363 0 6415 668
rect 7092 0 7144 310
rect 7678 0 7730 618
rect 9049 0 9101 1018
rect 9971 0 10023 109
rect 13367 0 13419 239
rect 13655 0 13785 454
rect 15256 0 15384 411
rect 15522 0 15574 237
rect 15741 0 15781 243
rect 15943 0 15983 35574
<< obsm2 >>
rect 42 35630 15983 40000
rect 42 1341 15887 35630
rect 42 1126 4415 1341
rect 42 951 2495 1126
rect 42 50 619 951
rect 777 50 1028 951
rect 1186 366 2495 951
rect 1334 50 2495 366
rect 2659 520 4415 1126
rect 2659 50 3206 520
rect 3370 50 4415 520
rect 4579 1074 15887 1341
rect 4579 870 8993 1074
rect 4579 597 5642 870
rect 4579 50 5264 597
rect 5428 50 5642 597
rect 5806 724 8993 870
rect 5806 509 6307 724
rect 6471 674 8993 724
rect 5806 50 6094 509
rect 6258 50 6307 509
rect 6471 366 7622 674
rect 6471 50 7036 366
rect 7200 50 7622 366
rect 7786 50 8993 674
rect 9157 510 15887 1074
rect 9157 295 13599 510
rect 13841 467 15887 510
rect 9157 165 13311 295
rect 9157 50 9915 165
rect 10079 50 13311 165
rect 13475 50 13599 295
rect 13841 50 15200 467
rect 15440 299 15887 467
rect 15440 293 15685 299
rect 15440 50 15466 293
rect 15630 50 15685 293
rect 15837 50 15887 299
<< metal3 >>
rect 80 0 204 35697
rect 9173 0 9239 7361
rect 12564 0 12778 1941
rect 15716 0 15782 36955
rect 15848 0 15914 37912
<< obsm3 >>
rect 80 37992 15914 40000
rect 80 37035 15768 37992
rect 80 35777 15636 37035
rect 284 7441 15636 35777
rect 284 49 9093 7441
rect 9319 2021 15636 7441
rect 9319 49 12484 2021
rect 12858 49 15636 2021
<< metal4 >>
rect 0 35157 5110 40000
rect 13246 35157 16000 40000
rect 1714 24002 1960 24248
rect 1962 24241 2500 24250
rect 400 21317 1094 23791
rect 1503 23791 1714 24002
rect 1566 21006 1960 21317
rect 1566 20923 2500 21006
rect 0 14007 292 19000
rect 13606 14007 16000 19000
rect 0 12817 1372 13707
rect 12189 12817 16000 13707
rect 0 11647 13969 12537
rect 14315 11647 16000 12537
rect 0 11281 522 11347
rect 0 10625 7288 11221
rect 0 10329 522 10565
rect 9418 11281 16000 11347
rect 7752 10625 16000 11221
rect 9418 10329 16000 10565
rect 0 9673 10429 10269
rect 10893 9673 16000 10269
rect 0 9547 522 9613
rect 9418 9547 16000 9613
rect 0 8317 2782 9247
rect 11141 8317 16000 9247
rect 0 7347 1087 8037
rect 13462 7347 16000 8037
rect 0 6377 4454 7067
rect 4770 6377 16000 7067
rect 0 5167 3866 6097
rect 4306 5167 16000 6097
rect 0 3957 1486 4887
rect 14347 3957 16000 4887
rect 0 2987 4918 3677
rect 10314 2987 16000 3677
rect 0 1777 6847 2707
rect 14053 1777 16000 2707
rect 0 407 2230 1497
rect 15362 407 16000 1497
<< obsm4 >>
rect 5190 35077 13166 40000
rect 269 24330 15633 35077
rect 269 24328 1882 24330
rect 269 24082 1634 24328
rect 269 23871 1423 24082
rect 2580 24161 15633 24330
rect 269 21237 320 23871
rect 1174 23711 1423 23871
rect 2040 23922 15633 24161
rect 1794 23711 15633 23922
rect 1174 21397 15633 23711
rect 1174 21237 1486 21397
rect 269 20843 1486 21237
rect 2040 21086 15633 21397
rect 2580 20843 15633 21086
rect 269 19080 15633 20843
rect 372 13927 13526 19080
rect 269 13787 15633 13927
rect 1452 12737 12109 13787
rect 269 12617 15633 12737
rect 14049 11567 14235 12617
rect 269 11427 15633 11567
rect 602 11301 9338 11427
rect 7368 10545 7672 11301
rect 602 10349 9338 10545
rect 10509 9693 10813 10249
rect 602 9467 9338 9593
rect 269 9327 15633 9467
rect 2862 8237 11061 9327
rect 269 8117 15633 8237
rect 1167 7267 13382 8117
rect 269 7147 15633 7267
rect 4534 6297 4690 7147
rect 269 6177 15633 6297
rect 3946 5087 4226 6177
rect 269 4967 15633 5087
rect 1566 3877 14267 4967
rect 269 3757 15633 3877
rect 4998 2907 10234 3757
rect 269 2787 15633 2907
rect 6927 1697 13973 2787
rect 269 1577 15633 1697
rect 2310 327 15282 1577
rect 269 107 15633 327
<< metal5 >>
rect 2240 20912 14760 33402
<< obsm5 >>
rect 1960 33722 15040 34697
rect 1960 19617 15040 20592
<< labels >>
rlabel metal5 s 2240 20912 14760 33402 6 PAD
port 1 nsew signal bidirectional
rlabel metal4 s 0 8317 2782 9247 6 VSSD
port 2 nsew ground bidirectional
rlabel metal4 s 11141 8317 16000 9247 6 VSSD
port 2 nsew ground bidirectional
rlabel metal4 s 0 9673 10429 10269 6 AMUXBUS_B
port 3 nsew signal bidirectional
rlabel metal4 s 10893 9673 16000 10269 6 AMUXBUS_B
port 3 nsew signal bidirectional
rlabel metal4 s 0 10625 7288 11221 6 AMUXBUS_A
port 4 nsew signal bidirectional
rlabel metal4 s 7752 10625 16000 11221 6 AMUXBUS_A
port 4 nsew signal bidirectional
rlabel metal4 s 0 12817 1372 13707 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal4 s 12189 12817 16000 13707 6 VDDIO_Q
port 5 nsew power bidirectional
rlabel metal4 s 0 14007 292 19000 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 0 3957 1486 4887 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 13606 14007 16000 19000 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 14347 3957 16000 4887 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 0 6377 4454 7067 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal4 s 4770 6377 16000 7067 6 VSWITCH
port 7 nsew power bidirectional
rlabel metal4 s 0 5167 3866 6097 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal4 s 4306 5167 16000 6097 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal4 s 13246 35157 16000 40000 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal4 s 0 35157 5110 40000 6 VSSIO
port 8 nsew ground bidirectional
rlabel metal4 s 0 2987 4918 3677 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 10314 2987 16000 3677 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 0 1777 6847 2707 6 VCCD
port 10 nsew power bidirectional
rlabel metal4 s 14053 1777 16000 2707 6 VCCD
port 10 nsew power bidirectional
rlabel metal4 s 0 407 2230 1497 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 15362 407 16000 1497 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 0 11281 522 11347 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 0 9547 522 9613 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 0 10329 522 10565 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 0 7347 1087 8037 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 13462 7347 16000 8037 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 9418 11281 16000 11347 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 9418 9547 16000 9613 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 9418 10329 16000 10565 6 VSSA
port 12 nsew ground bidirectional
rlabel metal4 s 0 11647 13969 12537 6 VSSIO_Q
port 13 nsew ground bidirectional
rlabel metal4 s 14315 11647 16000 12537 6 VSSIO_Q
port 13 nsew ground bidirectional
rlabel metal4 s 400 21317 1094 23791 6 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal3 s 12564 0 12778 1941 6 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1962 24241 2500 24250 6 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1960 20923 2500 21006 6 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1714 24002 1960 24248 6 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1566 20923 1960 21317 6 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal4 s 1503 23791 1714 24002 6 PAD_A_NOESD_H
port 14 nsew signal bidirectional
rlabel metal3 s 9173 0 9239 7361 6 ANALOG_POL
port 15 nsew signal input
rlabel metal3 s 15716 0 15782 36955 6 ENABLE_VDDIO
port 16 nsew signal input
rlabel metal3 s 80 0 204 35697 6 IN_H
port 17 nsew signal output
rlabel metal3 s 15848 0 15914 37912 6 IN
port 18 nsew signal output
rlabel metal1 s 12486 0 12538 261 6 ANALOG_EN
port 19 nsew signal input
rlabel metal2 s 4471 0 4523 1285 6 OUT
port 20 nsew signal input
rlabel metal2 s 15741 0 15781 243 6 TIE_HI_ESD
port 21 nsew signal output
rlabel metal2 s 13655 0 13785 454 6 PAD_A_ESD_1_H
port 22 nsew signal bidirectional
rlabel metal2 s 9971 0 10023 109 6 DM[0]
port 23 nsew signal input
rlabel metal2 s 13367 0 13419 239 6 DM[1]
port 24 nsew signal input
rlabel metal2 s 5698 0 5750 814 6 DM[2]
port 25 nsew signal input
rlabel metal2 s 6363 0 6415 668 6 HLD_H_N
port 26 nsew signal input
rlabel metal2 s 5320 0 5372 541 6 HLD_OVR
port 27 nsew signal input
rlabel metal2 s 9049 0 9101 1018 6 INP_DIS
port 28 nsew signal input
rlabel metal2 s 2551 0 2603 1070 6 ENABLE_VDDA_H
port 29 nsew signal input
rlabel metal2 s 1226 0 1278 310 6 VTRIP_SEL
port 30 nsew signal input
rlabel metal2 s 675 0 721 895 6 OE_N
port 31 nsew signal input
rlabel metal2 s 15522 0 15574 237 6 SLOW
port 32 nsew signal input
rlabel metal2 s 15943 0 15983 35574 6 TIE_LO_ESD
port 33 nsew signal output
rlabel metal2 s 15256 0 15384 411 6 PAD_A_ESD_0_H
port 34 nsew signal bidirectional
rlabel metal2 s 6150 0 6202 453 6 ANALOG_SEL
port 35 nsew signal input
rlabel metal2 s 7678 0 7730 618 6 ENABLE_INP_H
port 36 nsew signal input
rlabel metal2 s 7092 0 7144 310 6 ENABLE_H
port 37 nsew signal input
rlabel metal2 s 1084 0 1130 895 6 IB_MODE_SEL
port 38 nsew signal input
rlabel metal2 s 3262 0 3314 464 6 ENABLE_VSWITCH_H
port 39 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 11194436
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 9423270
<< end >>
