/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/sonos_see/end_of_life.spice