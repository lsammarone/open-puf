magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 710 157 892 201
rect 1200 157 1741 203
rect 1 21 1741 157
rect 29 -17 63 21
<< locali >>
rect 18 195 88 325
rect 288 213 344 333
rect 1397 327 1464 479
rect 1568 327 1634 479
rect 1397 293 1731 327
rect 1682 180 1731 293
rect 1397 146 1731 180
rect 1397 61 1464 146
rect 1568 61 1635 146
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 248 493
rect 288 435 341 527
rect 378 413 425 488
rect 474 438 688 472
rect 291 17 341 109
rect 378 107 412 413
rect 446 207 494 381
rect 532 331 620 402
rect 654 315 688 438
rect 722 367 756 527
rect 790 427 840 493
rect 885 433 1062 467
rect 654 297 756 315
rect 596 263 756 297
rect 446 141 562 207
rect 596 107 630 263
rect 722 249 756 263
rect 664 213 698 219
rect 790 213 824 427
rect 858 249 896 393
rect 930 315 994 381
rect 664 153 824 213
rect 930 207 968 315
rect 378 73 444 107
rect 480 73 630 107
rect 680 17 754 117
rect 790 107 824 153
rect 858 141 968 207
rect 1028 249 1062 433
rect 1098 427 1141 527
rect 1234 366 1268 491
rect 1325 371 1361 527
rect 1096 334 1268 366
rect 1096 300 1318 334
rect 1284 249 1318 300
rect 1500 361 1534 527
rect 1668 361 1702 527
rect 1028 215 1246 249
rect 1284 215 1648 249
rect 1028 107 1062 215
rect 1284 181 1318 215
rect 1218 147 1318 181
rect 790 73 882 107
rect 928 73 1062 107
rect 1125 17 1159 123
rect 1218 59 1290 147
rect 1325 17 1359 113
rect 1499 17 1533 112
rect 1669 17 1703 112
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< obsm1 >>
rect 110 388 168 397
rect 574 388 632 397
rect 850 388 908 397
rect 110 360 908 388
rect 110 351 168 360
rect 574 351 632 360
rect 850 351 908 360
rect 202 184 260 193
rect 482 184 540 193
rect 850 184 908 193
rect 202 156 908 184
rect 202 147 260 156
rect 482 147 540 156
rect 850 147 908 156
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 288 213 344 333 6 D
port 2 nsew signal input
rlabel metal1 s 0 -48 1748 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1741 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1200 157 1741 203 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 710 157 892 201 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1786 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1748 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1568 61 1635 146 6 Q
port 7 nsew signal output
rlabel locali s 1397 61 1464 146 6 Q
port 7 nsew signal output
rlabel locali s 1397 146 1731 180 6 Q
port 7 nsew signal output
rlabel locali s 1682 180 1731 293 6 Q
port 7 nsew signal output
rlabel locali s 1397 293 1731 327 6 Q
port 7 nsew signal output
rlabel locali s 1568 327 1634 479 6 Q
port 7 nsew signal output
rlabel locali s 1397 327 1464 479 6 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1748 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2696512
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2682412
<< end >>
