magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< metal3 >>
rect 10151 2588 14931 3276
<< obsm3 >>
rect 120 2588 4900 3276
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 208 3208 272 3272
rect 290 3208 354 3272
rect 372 3208 436 3272
rect 454 3208 518 3272
rect 536 3208 600 3272
rect 618 3208 682 3272
rect 699 3208 763 3272
rect 780 3208 844 3272
rect 861 3208 925 3272
rect 942 3208 1006 3272
rect 1023 3208 1087 3272
rect 1104 3208 1168 3272
rect 1185 3208 1249 3272
rect 1266 3208 1330 3272
rect 1347 3208 1411 3272
rect 1428 3208 1492 3272
rect 1509 3208 1573 3272
rect 1590 3208 1654 3272
rect 1671 3208 1735 3272
rect 1752 3208 1816 3272
rect 1833 3208 1897 3272
rect 1914 3208 1978 3272
rect 1995 3208 2059 3272
rect 2076 3208 2140 3272
rect 2157 3208 2221 3272
rect 2238 3208 2302 3272
rect 2319 3208 2383 3272
rect 2400 3208 2464 3272
rect 2481 3208 2545 3272
rect 2562 3208 2626 3272
rect 2643 3208 2707 3272
rect 2724 3208 2788 3272
rect 2805 3208 2869 3272
rect 2886 3208 2950 3272
rect 2967 3208 3031 3272
rect 3048 3208 3112 3272
rect 3129 3208 3193 3272
rect 3210 3208 3274 3272
rect 3291 3208 3355 3272
rect 3372 3208 3436 3272
rect 3453 3208 3517 3272
rect 3534 3208 3598 3272
rect 3615 3208 3679 3272
rect 3696 3208 3760 3272
rect 3777 3208 3841 3272
rect 3858 3208 3922 3272
rect 3939 3208 4003 3272
rect 4020 3208 4084 3272
rect 4101 3208 4165 3272
rect 4182 3208 4246 3272
rect 4263 3208 4327 3272
rect 4344 3208 4408 3272
rect 4425 3208 4489 3272
rect 4506 3208 4570 3272
rect 4587 3208 4651 3272
rect 4668 3208 4732 3272
rect 4749 3208 4813 3272
rect 4830 3208 4894 3272
rect 208 3120 272 3184
rect 290 3120 354 3184
rect 372 3120 436 3184
rect 454 3120 518 3184
rect 536 3120 600 3184
rect 618 3120 682 3184
rect 699 3120 763 3184
rect 780 3120 844 3184
rect 861 3120 925 3184
rect 942 3120 1006 3184
rect 1023 3120 1087 3184
rect 1104 3120 1168 3184
rect 1185 3120 1249 3184
rect 1266 3120 1330 3184
rect 1347 3120 1411 3184
rect 1428 3120 1492 3184
rect 1509 3120 1573 3184
rect 1590 3120 1654 3184
rect 1671 3120 1735 3184
rect 1752 3120 1816 3184
rect 1833 3120 1897 3184
rect 1914 3120 1978 3184
rect 1995 3120 2059 3184
rect 2076 3120 2140 3184
rect 2157 3120 2221 3184
rect 2238 3120 2302 3184
rect 2319 3120 2383 3184
rect 2400 3120 2464 3184
rect 2481 3120 2545 3184
rect 2562 3120 2626 3184
rect 2643 3120 2707 3184
rect 2724 3120 2788 3184
rect 2805 3120 2869 3184
rect 2886 3120 2950 3184
rect 2967 3120 3031 3184
rect 3048 3120 3112 3184
rect 3129 3120 3193 3184
rect 3210 3120 3274 3184
rect 3291 3120 3355 3184
rect 3372 3120 3436 3184
rect 3453 3120 3517 3184
rect 3534 3120 3598 3184
rect 3615 3120 3679 3184
rect 3696 3120 3760 3184
rect 3777 3120 3841 3184
rect 3858 3120 3922 3184
rect 3939 3120 4003 3184
rect 4020 3120 4084 3184
rect 4101 3120 4165 3184
rect 4182 3120 4246 3184
rect 4263 3120 4327 3184
rect 4344 3120 4408 3184
rect 4425 3120 4489 3184
rect 4506 3120 4570 3184
rect 4587 3120 4651 3184
rect 4668 3120 4732 3184
rect 4749 3120 4813 3184
rect 4830 3120 4894 3184
rect 208 3032 272 3096
rect 290 3032 354 3096
rect 372 3032 436 3096
rect 454 3032 518 3096
rect 536 3032 600 3096
rect 618 3032 682 3096
rect 699 3032 763 3096
rect 780 3032 844 3096
rect 861 3032 925 3096
rect 942 3032 1006 3096
rect 1023 3032 1087 3096
rect 1104 3032 1168 3096
rect 1185 3032 1249 3096
rect 1266 3032 1330 3096
rect 1347 3032 1411 3096
rect 1428 3032 1492 3096
rect 1509 3032 1573 3096
rect 1590 3032 1654 3096
rect 1671 3032 1735 3096
rect 1752 3032 1816 3096
rect 1833 3032 1897 3096
rect 1914 3032 1978 3096
rect 1995 3032 2059 3096
rect 2076 3032 2140 3096
rect 2157 3032 2221 3096
rect 2238 3032 2302 3096
rect 2319 3032 2383 3096
rect 2400 3032 2464 3096
rect 2481 3032 2545 3096
rect 2562 3032 2626 3096
rect 2643 3032 2707 3096
rect 2724 3032 2788 3096
rect 2805 3032 2869 3096
rect 2886 3032 2950 3096
rect 2967 3032 3031 3096
rect 3048 3032 3112 3096
rect 3129 3032 3193 3096
rect 3210 3032 3274 3096
rect 3291 3032 3355 3096
rect 3372 3032 3436 3096
rect 3453 3032 3517 3096
rect 3534 3032 3598 3096
rect 3615 3032 3679 3096
rect 3696 3032 3760 3096
rect 3777 3032 3841 3096
rect 3858 3032 3922 3096
rect 3939 3032 4003 3096
rect 4020 3032 4084 3096
rect 4101 3032 4165 3096
rect 4182 3032 4246 3096
rect 4263 3032 4327 3096
rect 4344 3032 4408 3096
rect 4425 3032 4489 3096
rect 4506 3032 4570 3096
rect 4587 3032 4651 3096
rect 4668 3032 4732 3096
rect 4749 3032 4813 3096
rect 4830 3032 4894 3096
rect 208 2944 272 3008
rect 290 2944 354 3008
rect 372 2944 436 3008
rect 454 2944 518 3008
rect 536 2944 600 3008
rect 618 2944 682 3008
rect 699 2944 763 3008
rect 780 2944 844 3008
rect 861 2944 925 3008
rect 942 2944 1006 3008
rect 1023 2944 1087 3008
rect 1104 2944 1168 3008
rect 1185 2944 1249 3008
rect 1266 2944 1330 3008
rect 1347 2944 1411 3008
rect 1428 2944 1492 3008
rect 1509 2944 1573 3008
rect 1590 2944 1654 3008
rect 1671 2944 1735 3008
rect 1752 2944 1816 3008
rect 1833 2944 1897 3008
rect 1914 2944 1978 3008
rect 1995 2944 2059 3008
rect 2076 2944 2140 3008
rect 2157 2944 2221 3008
rect 2238 2944 2302 3008
rect 2319 2944 2383 3008
rect 2400 2944 2464 3008
rect 2481 2944 2545 3008
rect 2562 2944 2626 3008
rect 2643 2944 2707 3008
rect 2724 2944 2788 3008
rect 2805 2944 2869 3008
rect 2886 2944 2950 3008
rect 2967 2944 3031 3008
rect 3048 2944 3112 3008
rect 3129 2944 3193 3008
rect 3210 2944 3274 3008
rect 3291 2944 3355 3008
rect 3372 2944 3436 3008
rect 3453 2944 3517 3008
rect 3534 2944 3598 3008
rect 3615 2944 3679 3008
rect 3696 2944 3760 3008
rect 3777 2944 3841 3008
rect 3858 2944 3922 3008
rect 3939 2944 4003 3008
rect 4020 2944 4084 3008
rect 4101 2944 4165 3008
rect 4182 2944 4246 3008
rect 4263 2944 4327 3008
rect 4344 2944 4408 3008
rect 4425 2944 4489 3008
rect 4506 2944 4570 3008
rect 4587 2944 4651 3008
rect 4668 2944 4732 3008
rect 4749 2944 4813 3008
rect 4830 2944 4894 3008
rect 208 2856 272 2920
rect 290 2856 354 2920
rect 372 2856 436 2920
rect 454 2856 518 2920
rect 536 2856 600 2920
rect 618 2856 682 2920
rect 699 2856 763 2920
rect 780 2856 844 2920
rect 861 2856 925 2920
rect 942 2856 1006 2920
rect 1023 2856 1087 2920
rect 1104 2856 1168 2920
rect 1185 2856 1249 2920
rect 1266 2856 1330 2920
rect 1347 2856 1411 2920
rect 1428 2856 1492 2920
rect 1509 2856 1573 2920
rect 1590 2856 1654 2920
rect 1671 2856 1735 2920
rect 1752 2856 1816 2920
rect 1833 2856 1897 2920
rect 1914 2856 1978 2920
rect 1995 2856 2059 2920
rect 2076 2856 2140 2920
rect 2157 2856 2221 2920
rect 2238 2856 2302 2920
rect 2319 2856 2383 2920
rect 2400 2856 2464 2920
rect 2481 2856 2545 2920
rect 2562 2856 2626 2920
rect 2643 2856 2707 2920
rect 2724 2856 2788 2920
rect 2805 2856 2869 2920
rect 2886 2856 2950 2920
rect 2967 2856 3031 2920
rect 3048 2856 3112 2920
rect 3129 2856 3193 2920
rect 3210 2856 3274 2920
rect 3291 2856 3355 2920
rect 3372 2856 3436 2920
rect 3453 2856 3517 2920
rect 3534 2856 3598 2920
rect 3615 2856 3679 2920
rect 3696 2856 3760 2920
rect 3777 2856 3841 2920
rect 3858 2856 3922 2920
rect 3939 2856 4003 2920
rect 4020 2856 4084 2920
rect 4101 2856 4165 2920
rect 4182 2856 4246 2920
rect 4263 2856 4327 2920
rect 4344 2856 4408 2920
rect 4425 2856 4489 2920
rect 4506 2856 4570 2920
rect 4587 2856 4651 2920
rect 4668 2856 4732 2920
rect 4749 2856 4813 2920
rect 4830 2856 4894 2920
rect 208 2768 272 2832
rect 290 2768 354 2832
rect 372 2768 436 2832
rect 454 2768 518 2832
rect 536 2768 600 2832
rect 618 2768 682 2832
rect 699 2768 763 2832
rect 780 2768 844 2832
rect 861 2768 925 2832
rect 942 2768 1006 2832
rect 1023 2768 1087 2832
rect 1104 2768 1168 2832
rect 1185 2768 1249 2832
rect 1266 2768 1330 2832
rect 1347 2768 1411 2832
rect 1428 2768 1492 2832
rect 1509 2768 1573 2832
rect 1590 2768 1654 2832
rect 1671 2768 1735 2832
rect 1752 2768 1816 2832
rect 1833 2768 1897 2832
rect 1914 2768 1978 2832
rect 1995 2768 2059 2832
rect 2076 2768 2140 2832
rect 2157 2768 2221 2832
rect 2238 2768 2302 2832
rect 2319 2768 2383 2832
rect 2400 2768 2464 2832
rect 2481 2768 2545 2832
rect 2562 2768 2626 2832
rect 2643 2768 2707 2832
rect 2724 2768 2788 2832
rect 2805 2768 2869 2832
rect 2886 2768 2950 2832
rect 2967 2768 3031 2832
rect 3048 2768 3112 2832
rect 3129 2768 3193 2832
rect 3210 2768 3274 2832
rect 3291 2768 3355 2832
rect 3372 2768 3436 2832
rect 3453 2768 3517 2832
rect 3534 2768 3598 2832
rect 3615 2768 3679 2832
rect 3696 2768 3760 2832
rect 3777 2768 3841 2832
rect 3858 2768 3922 2832
rect 3939 2768 4003 2832
rect 4020 2768 4084 2832
rect 4101 2768 4165 2832
rect 4182 2768 4246 2832
rect 4263 2768 4327 2832
rect 4344 2768 4408 2832
rect 4425 2768 4489 2832
rect 4506 2768 4570 2832
rect 4587 2768 4651 2832
rect 4668 2768 4732 2832
rect 4749 2768 4813 2832
rect 4830 2768 4894 2832
rect 208 2680 272 2744
rect 290 2680 354 2744
rect 372 2680 436 2744
rect 454 2680 518 2744
rect 536 2680 600 2744
rect 618 2680 682 2744
rect 699 2680 763 2744
rect 780 2680 844 2744
rect 861 2680 925 2744
rect 942 2680 1006 2744
rect 1023 2680 1087 2744
rect 1104 2680 1168 2744
rect 1185 2680 1249 2744
rect 1266 2680 1330 2744
rect 1347 2680 1411 2744
rect 1428 2680 1492 2744
rect 1509 2680 1573 2744
rect 1590 2680 1654 2744
rect 1671 2680 1735 2744
rect 1752 2680 1816 2744
rect 1833 2680 1897 2744
rect 1914 2680 1978 2744
rect 1995 2680 2059 2744
rect 2076 2680 2140 2744
rect 2157 2680 2221 2744
rect 2238 2680 2302 2744
rect 2319 2680 2383 2744
rect 2400 2680 2464 2744
rect 2481 2680 2545 2744
rect 2562 2680 2626 2744
rect 2643 2680 2707 2744
rect 2724 2680 2788 2744
rect 2805 2680 2869 2744
rect 2886 2680 2950 2744
rect 2967 2680 3031 2744
rect 3048 2680 3112 2744
rect 3129 2680 3193 2744
rect 3210 2680 3274 2744
rect 3291 2680 3355 2744
rect 3372 2680 3436 2744
rect 3453 2680 3517 2744
rect 3534 2680 3598 2744
rect 3615 2680 3679 2744
rect 3696 2680 3760 2744
rect 3777 2680 3841 2744
rect 3858 2680 3922 2744
rect 3939 2680 4003 2744
rect 4020 2680 4084 2744
rect 4101 2680 4165 2744
rect 4182 2680 4246 2744
rect 4263 2680 4327 2744
rect 4344 2680 4408 2744
rect 4425 2680 4489 2744
rect 4506 2680 4570 2744
rect 4587 2680 4651 2744
rect 4668 2680 4732 2744
rect 4749 2680 4813 2744
rect 4830 2680 4894 2744
rect 208 2592 272 2656
rect 290 2592 354 2656
rect 372 2592 436 2656
rect 454 2592 518 2656
rect 536 2592 600 2656
rect 618 2592 682 2656
rect 699 2592 763 2656
rect 780 2592 844 2656
rect 861 2592 925 2656
rect 942 2592 1006 2656
rect 1023 2592 1087 2656
rect 1104 2592 1168 2656
rect 1185 2592 1249 2656
rect 1266 2592 1330 2656
rect 1347 2592 1411 2656
rect 1428 2592 1492 2656
rect 1509 2592 1573 2656
rect 1590 2592 1654 2656
rect 1671 2592 1735 2656
rect 1752 2592 1816 2656
rect 1833 2592 1897 2656
rect 1914 2592 1978 2656
rect 1995 2592 2059 2656
rect 2076 2592 2140 2656
rect 2157 2592 2221 2656
rect 2238 2592 2302 2656
rect 2319 2592 2383 2656
rect 2400 2592 2464 2656
rect 2481 2592 2545 2656
rect 2562 2592 2626 2656
rect 2643 2592 2707 2656
rect 2724 2592 2788 2656
rect 2805 2592 2869 2656
rect 2886 2592 2950 2656
rect 2967 2592 3031 2656
rect 3048 2592 3112 2656
rect 3129 2592 3193 2656
rect 3210 2592 3274 2656
rect 3291 2592 3355 2656
rect 3372 2592 3436 2656
rect 3453 2592 3517 2656
rect 3534 2592 3598 2656
rect 3615 2592 3679 2656
rect 3696 2592 3760 2656
rect 3777 2592 3841 2656
rect 3858 2592 3922 2656
rect 3939 2592 4003 2656
rect 4020 2592 4084 2656
rect 4101 2592 4165 2656
rect 4182 2592 4246 2656
rect 4263 2592 4327 2656
rect 4344 2592 4408 2656
rect 4425 2592 4489 2656
rect 4506 2592 4570 2656
rect 4587 2592 4651 2656
rect 4668 2592 4732 2656
rect 4749 2592 4813 2656
rect 4830 2592 4894 2656
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 3272 14727 3357
rect 273 3208 290 3272
rect 354 3208 372 3272
rect 436 3208 454 3272
rect 518 3208 536 3272
rect 600 3208 618 3272
rect 682 3208 699 3272
rect 763 3208 780 3272
rect 844 3208 861 3272
rect 925 3208 942 3272
rect 1006 3208 1023 3272
rect 1087 3208 1104 3272
rect 1168 3208 1185 3272
rect 1249 3208 1266 3272
rect 1330 3208 1347 3272
rect 1411 3208 1428 3272
rect 1492 3208 1509 3272
rect 1573 3208 1590 3272
rect 1654 3208 1671 3272
rect 1735 3208 1752 3272
rect 1816 3208 1833 3272
rect 1897 3208 1914 3272
rect 1978 3208 1995 3272
rect 2059 3208 2076 3272
rect 2140 3208 2157 3272
rect 2221 3208 2238 3272
rect 2302 3208 2319 3272
rect 2383 3208 2400 3272
rect 2464 3208 2481 3272
rect 2545 3208 2562 3272
rect 2626 3208 2643 3272
rect 2707 3208 2724 3272
rect 2788 3208 2805 3272
rect 2869 3208 2886 3272
rect 2950 3208 2967 3272
rect 3031 3208 3048 3272
rect 3112 3208 3129 3272
rect 3193 3208 3210 3272
rect 3274 3208 3291 3272
rect 3355 3208 3372 3272
rect 3436 3208 3453 3272
rect 3517 3208 3534 3272
rect 3598 3208 3615 3272
rect 3679 3208 3696 3272
rect 3760 3208 3777 3272
rect 3841 3208 3858 3272
rect 3922 3208 3939 3272
rect 4003 3208 4020 3272
rect 4084 3208 4101 3272
rect 4165 3208 4182 3272
rect 4246 3208 4263 3272
rect 4327 3208 4344 3272
rect 4408 3208 4425 3272
rect 4489 3208 4506 3272
rect 4570 3208 4587 3272
rect 4651 3208 4668 3272
rect 4732 3208 4749 3272
rect 4813 3208 4830 3272
rect 4894 3208 14727 3272
rect 273 3184 14727 3208
rect 273 3120 290 3184
rect 354 3120 372 3184
rect 436 3120 454 3184
rect 518 3120 536 3184
rect 600 3120 618 3184
rect 682 3120 699 3184
rect 763 3120 780 3184
rect 844 3120 861 3184
rect 925 3120 942 3184
rect 1006 3120 1023 3184
rect 1087 3120 1104 3184
rect 1168 3120 1185 3184
rect 1249 3120 1266 3184
rect 1330 3120 1347 3184
rect 1411 3120 1428 3184
rect 1492 3120 1509 3184
rect 1573 3120 1590 3184
rect 1654 3120 1671 3184
rect 1735 3120 1752 3184
rect 1816 3120 1833 3184
rect 1897 3120 1914 3184
rect 1978 3120 1995 3184
rect 2059 3120 2076 3184
rect 2140 3120 2157 3184
rect 2221 3120 2238 3184
rect 2302 3120 2319 3184
rect 2383 3120 2400 3184
rect 2464 3120 2481 3184
rect 2545 3120 2562 3184
rect 2626 3120 2643 3184
rect 2707 3120 2724 3184
rect 2788 3120 2805 3184
rect 2869 3120 2886 3184
rect 2950 3120 2967 3184
rect 3031 3120 3048 3184
rect 3112 3120 3129 3184
rect 3193 3120 3210 3184
rect 3274 3120 3291 3184
rect 3355 3120 3372 3184
rect 3436 3120 3453 3184
rect 3517 3120 3534 3184
rect 3598 3120 3615 3184
rect 3679 3120 3696 3184
rect 3760 3120 3777 3184
rect 3841 3120 3858 3184
rect 3922 3120 3939 3184
rect 4003 3120 4020 3184
rect 4084 3120 4101 3184
rect 4165 3120 4182 3184
rect 4246 3120 4263 3184
rect 4327 3120 4344 3184
rect 4408 3120 4425 3184
rect 4489 3120 4506 3184
rect 4570 3120 4587 3184
rect 4651 3120 4668 3184
rect 4732 3120 4749 3184
rect 4813 3120 4830 3184
rect 4894 3120 14727 3184
rect 273 3096 14727 3120
rect 273 3032 290 3096
rect 354 3032 372 3096
rect 436 3032 454 3096
rect 518 3032 536 3096
rect 600 3032 618 3096
rect 682 3032 699 3096
rect 763 3032 780 3096
rect 844 3032 861 3096
rect 925 3032 942 3096
rect 1006 3032 1023 3096
rect 1087 3032 1104 3096
rect 1168 3032 1185 3096
rect 1249 3032 1266 3096
rect 1330 3032 1347 3096
rect 1411 3032 1428 3096
rect 1492 3032 1509 3096
rect 1573 3032 1590 3096
rect 1654 3032 1671 3096
rect 1735 3032 1752 3096
rect 1816 3032 1833 3096
rect 1897 3032 1914 3096
rect 1978 3032 1995 3096
rect 2059 3032 2076 3096
rect 2140 3032 2157 3096
rect 2221 3032 2238 3096
rect 2302 3032 2319 3096
rect 2383 3032 2400 3096
rect 2464 3032 2481 3096
rect 2545 3032 2562 3096
rect 2626 3032 2643 3096
rect 2707 3032 2724 3096
rect 2788 3032 2805 3096
rect 2869 3032 2886 3096
rect 2950 3032 2967 3096
rect 3031 3032 3048 3096
rect 3112 3032 3129 3096
rect 3193 3032 3210 3096
rect 3274 3032 3291 3096
rect 3355 3032 3372 3096
rect 3436 3032 3453 3096
rect 3517 3032 3534 3096
rect 3598 3032 3615 3096
rect 3679 3032 3696 3096
rect 3760 3032 3777 3096
rect 3841 3032 3858 3096
rect 3922 3032 3939 3096
rect 4003 3032 4020 3096
rect 4084 3032 4101 3096
rect 4165 3032 4182 3096
rect 4246 3032 4263 3096
rect 4327 3032 4344 3096
rect 4408 3032 4425 3096
rect 4489 3032 4506 3096
rect 4570 3032 4587 3096
rect 4651 3032 4668 3096
rect 4732 3032 4749 3096
rect 4813 3032 4830 3096
rect 4894 3032 14727 3096
rect 273 3008 14727 3032
rect 273 2944 290 3008
rect 354 2944 372 3008
rect 436 2944 454 3008
rect 518 2944 536 3008
rect 600 2944 618 3008
rect 682 2944 699 3008
rect 763 2944 780 3008
rect 844 2944 861 3008
rect 925 2944 942 3008
rect 1006 2944 1023 3008
rect 1087 2944 1104 3008
rect 1168 2944 1185 3008
rect 1249 2944 1266 3008
rect 1330 2944 1347 3008
rect 1411 2944 1428 3008
rect 1492 2944 1509 3008
rect 1573 2944 1590 3008
rect 1654 2944 1671 3008
rect 1735 2944 1752 3008
rect 1816 2944 1833 3008
rect 1897 2944 1914 3008
rect 1978 2944 1995 3008
rect 2059 2944 2076 3008
rect 2140 2944 2157 3008
rect 2221 2944 2238 3008
rect 2302 2944 2319 3008
rect 2383 2944 2400 3008
rect 2464 2944 2481 3008
rect 2545 2944 2562 3008
rect 2626 2944 2643 3008
rect 2707 2944 2724 3008
rect 2788 2944 2805 3008
rect 2869 2944 2886 3008
rect 2950 2944 2967 3008
rect 3031 2944 3048 3008
rect 3112 2944 3129 3008
rect 3193 2944 3210 3008
rect 3274 2944 3291 3008
rect 3355 2944 3372 3008
rect 3436 2944 3453 3008
rect 3517 2944 3534 3008
rect 3598 2944 3615 3008
rect 3679 2944 3696 3008
rect 3760 2944 3777 3008
rect 3841 2944 3858 3008
rect 3922 2944 3939 3008
rect 4003 2944 4020 3008
rect 4084 2944 4101 3008
rect 4165 2944 4182 3008
rect 4246 2944 4263 3008
rect 4327 2944 4344 3008
rect 4408 2944 4425 3008
rect 4489 2944 4506 3008
rect 4570 2944 4587 3008
rect 4651 2944 4668 3008
rect 4732 2944 4749 3008
rect 4813 2944 4830 3008
rect 4894 2944 14727 3008
rect 273 2920 14727 2944
rect 273 2856 290 2920
rect 354 2856 372 2920
rect 436 2856 454 2920
rect 518 2856 536 2920
rect 600 2856 618 2920
rect 682 2856 699 2920
rect 763 2856 780 2920
rect 844 2856 861 2920
rect 925 2856 942 2920
rect 1006 2856 1023 2920
rect 1087 2856 1104 2920
rect 1168 2856 1185 2920
rect 1249 2856 1266 2920
rect 1330 2856 1347 2920
rect 1411 2856 1428 2920
rect 1492 2856 1509 2920
rect 1573 2856 1590 2920
rect 1654 2856 1671 2920
rect 1735 2856 1752 2920
rect 1816 2856 1833 2920
rect 1897 2856 1914 2920
rect 1978 2856 1995 2920
rect 2059 2856 2076 2920
rect 2140 2856 2157 2920
rect 2221 2856 2238 2920
rect 2302 2856 2319 2920
rect 2383 2856 2400 2920
rect 2464 2856 2481 2920
rect 2545 2856 2562 2920
rect 2626 2856 2643 2920
rect 2707 2856 2724 2920
rect 2788 2856 2805 2920
rect 2869 2856 2886 2920
rect 2950 2856 2967 2920
rect 3031 2856 3048 2920
rect 3112 2856 3129 2920
rect 3193 2856 3210 2920
rect 3274 2856 3291 2920
rect 3355 2856 3372 2920
rect 3436 2856 3453 2920
rect 3517 2856 3534 2920
rect 3598 2856 3615 2920
rect 3679 2856 3696 2920
rect 3760 2856 3777 2920
rect 3841 2856 3858 2920
rect 3922 2856 3939 2920
rect 4003 2856 4020 2920
rect 4084 2856 4101 2920
rect 4165 2856 4182 2920
rect 4246 2856 4263 2920
rect 4327 2856 4344 2920
rect 4408 2856 4425 2920
rect 4489 2856 4506 2920
rect 4570 2856 4587 2920
rect 4651 2856 4668 2920
rect 4732 2856 4749 2920
rect 4813 2856 4830 2920
rect 4894 2856 14727 2920
rect 273 2832 14727 2856
rect 273 2768 290 2832
rect 354 2768 372 2832
rect 436 2768 454 2832
rect 518 2768 536 2832
rect 600 2768 618 2832
rect 682 2768 699 2832
rect 763 2768 780 2832
rect 844 2768 861 2832
rect 925 2768 942 2832
rect 1006 2768 1023 2832
rect 1087 2768 1104 2832
rect 1168 2768 1185 2832
rect 1249 2768 1266 2832
rect 1330 2768 1347 2832
rect 1411 2768 1428 2832
rect 1492 2768 1509 2832
rect 1573 2768 1590 2832
rect 1654 2768 1671 2832
rect 1735 2768 1752 2832
rect 1816 2768 1833 2832
rect 1897 2768 1914 2832
rect 1978 2768 1995 2832
rect 2059 2768 2076 2832
rect 2140 2768 2157 2832
rect 2221 2768 2238 2832
rect 2302 2768 2319 2832
rect 2383 2768 2400 2832
rect 2464 2768 2481 2832
rect 2545 2768 2562 2832
rect 2626 2768 2643 2832
rect 2707 2768 2724 2832
rect 2788 2768 2805 2832
rect 2869 2768 2886 2832
rect 2950 2768 2967 2832
rect 3031 2768 3048 2832
rect 3112 2768 3129 2832
rect 3193 2768 3210 2832
rect 3274 2768 3291 2832
rect 3355 2768 3372 2832
rect 3436 2768 3453 2832
rect 3517 2768 3534 2832
rect 3598 2768 3615 2832
rect 3679 2768 3696 2832
rect 3760 2768 3777 2832
rect 3841 2768 3858 2832
rect 3922 2768 3939 2832
rect 4003 2768 4020 2832
rect 4084 2768 4101 2832
rect 4165 2768 4182 2832
rect 4246 2768 4263 2832
rect 4327 2768 4344 2832
rect 4408 2768 4425 2832
rect 4489 2768 4506 2832
rect 4570 2768 4587 2832
rect 4651 2768 4668 2832
rect 4732 2768 4749 2832
rect 4813 2768 4830 2832
rect 4894 2768 14727 2832
rect 273 2744 14727 2768
rect 273 2680 290 2744
rect 354 2680 372 2744
rect 436 2680 454 2744
rect 518 2680 536 2744
rect 600 2680 618 2744
rect 682 2680 699 2744
rect 763 2680 780 2744
rect 844 2680 861 2744
rect 925 2680 942 2744
rect 1006 2680 1023 2744
rect 1087 2680 1104 2744
rect 1168 2680 1185 2744
rect 1249 2680 1266 2744
rect 1330 2680 1347 2744
rect 1411 2680 1428 2744
rect 1492 2680 1509 2744
rect 1573 2680 1590 2744
rect 1654 2680 1671 2744
rect 1735 2680 1752 2744
rect 1816 2680 1833 2744
rect 1897 2680 1914 2744
rect 1978 2680 1995 2744
rect 2059 2680 2076 2744
rect 2140 2680 2157 2744
rect 2221 2680 2238 2744
rect 2302 2680 2319 2744
rect 2383 2680 2400 2744
rect 2464 2680 2481 2744
rect 2545 2680 2562 2744
rect 2626 2680 2643 2744
rect 2707 2680 2724 2744
rect 2788 2680 2805 2744
rect 2869 2680 2886 2744
rect 2950 2680 2967 2744
rect 3031 2680 3048 2744
rect 3112 2680 3129 2744
rect 3193 2680 3210 2744
rect 3274 2680 3291 2744
rect 3355 2680 3372 2744
rect 3436 2680 3453 2744
rect 3517 2680 3534 2744
rect 3598 2680 3615 2744
rect 3679 2680 3696 2744
rect 3760 2680 3777 2744
rect 3841 2680 3858 2744
rect 3922 2680 3939 2744
rect 4003 2680 4020 2744
rect 4084 2680 4101 2744
rect 4165 2680 4182 2744
rect 4246 2680 4263 2744
rect 4327 2680 4344 2744
rect 4408 2680 4425 2744
rect 4489 2680 4506 2744
rect 4570 2680 4587 2744
rect 4651 2680 4668 2744
rect 4732 2680 4749 2744
rect 4813 2680 4830 2744
rect 4894 2680 14727 2744
rect 273 2656 14727 2680
rect 273 2592 290 2656
rect 354 2592 372 2656
rect 436 2592 454 2656
rect 518 2592 536 2656
rect 600 2592 618 2656
rect 682 2592 699 2656
rect 763 2592 780 2656
rect 844 2592 861 2656
rect 925 2592 942 2656
rect 1006 2592 1023 2656
rect 1087 2592 1104 2656
rect 1168 2592 1185 2656
rect 1249 2592 1266 2656
rect 1330 2592 1347 2656
rect 1411 2592 1428 2656
rect 1492 2592 1509 2656
rect 1573 2592 1590 2656
rect 1654 2592 1671 2656
rect 1735 2592 1752 2656
rect 1816 2592 1833 2656
rect 1897 2592 1914 2656
rect 1978 2592 1995 2656
rect 2059 2592 2076 2656
rect 2140 2592 2157 2656
rect 2221 2592 2238 2656
rect 2302 2592 2319 2656
rect 2383 2592 2400 2656
rect 2464 2592 2481 2656
rect 2545 2592 2562 2656
rect 2626 2592 2643 2656
rect 2707 2592 2724 2656
rect 2788 2592 2805 2656
rect 2869 2592 2886 2656
rect 2950 2592 2967 2656
rect 3031 2592 3048 2656
rect 3112 2592 3129 2656
rect 3193 2592 3210 2656
rect 3274 2592 3291 2656
rect 3355 2592 3372 2656
rect 3436 2592 3453 2656
rect 3517 2592 3534 2656
rect 3598 2592 3615 2656
rect 3679 2592 3696 2656
rect 3760 2592 3777 2656
rect 3841 2592 3858 2656
rect 3922 2592 3939 2656
rect 4003 2592 4020 2656
rect 4084 2592 4101 2656
rect 4165 2592 4182 2656
rect 4246 2592 4263 2656
rect 4327 2592 4344 2656
rect 4408 2592 4425 2656
rect 4489 2592 4506 2656
rect 4570 2592 4587 2656
rect 4651 2592 4668 2656
rect 4732 2592 4749 2656
rect 4813 2592 4830 2656
rect 4894 2592 14727 2656
rect 273 2507 14727 2592
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 2 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 2 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 3 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10151 2588 14931 3276 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 3220 14913 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 3132 14913 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 3044 14913 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 2956 14913 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 2868 14913 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 2780 14913 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 2692 14913 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14873 2604 14913 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 3220 14832 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 3132 14832 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 3044 14832 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 2956 14832 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 2868 14832 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 2780 14832 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 2692 14832 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14792 2604 14832 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 3220 14751 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 3132 14751 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 3044 14751 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 2956 14751 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 2868 14751 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 2780 14751 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 2692 14751 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14711 2604 14751 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 3220 14670 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 3132 14670 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 3044 14670 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 2956 14670 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 2868 14670 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 2780 14670 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 2692 14670 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14630 2604 14670 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 3220 14589 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 3132 14589 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 3044 14589 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 2956 14589 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 2868 14589 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 2780 14589 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 2692 14589 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14549 2604 14589 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 3220 14508 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 3132 14508 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 3044 14508 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 2956 14508 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 2868 14508 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 2780 14508 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 2692 14508 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14468 2604 14508 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 3220 14427 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 3132 14427 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 3044 14427 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 2956 14427 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 2868 14427 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 2780 14427 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 2692 14427 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14387 2604 14427 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 3220 14346 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 3132 14346 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 3044 14346 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 2956 14346 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 2868 14346 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 2780 14346 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 2692 14346 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14306 2604 14346 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 3220 14265 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 3132 14265 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 3044 14265 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 2956 14265 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 2868 14265 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 2780 14265 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 2692 14265 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14225 2604 14265 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 3220 14184 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 3132 14184 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 3044 14184 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 2956 14184 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 2868 14184 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 2780 14184 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 2692 14184 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14144 2604 14184 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 3220 14103 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 3132 14103 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 3044 14103 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 2956 14103 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 2868 14103 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 2780 14103 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 2692 14103 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 14063 2604 14103 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 3220 14022 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 3132 14022 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 3044 14022 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 2956 14022 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 2868 14022 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 2780 14022 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 2692 14022 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13982 2604 14022 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 3220 13941 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 3132 13941 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 3044 13941 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 2956 13941 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 2868 13941 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 2780 13941 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 2692 13941 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13901 2604 13941 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 3220 13860 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 3132 13860 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 3044 13860 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 2956 13860 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 2868 13860 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 2780 13860 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 2692 13860 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13820 2604 13860 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 3220 13779 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 3132 13779 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 3044 13779 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 2956 13779 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 2868 13779 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 2780 13779 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 2692 13779 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13739 2604 13779 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 3220 13698 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 3132 13698 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 3044 13698 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 2956 13698 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 2868 13698 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 2780 13698 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 2692 13698 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13658 2604 13698 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 3220 13617 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 3132 13617 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 3044 13617 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 2956 13617 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 2868 13617 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 2780 13617 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 2692 13617 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13577 2604 13617 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 3220 13536 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 3132 13536 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 3044 13536 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 2956 13536 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 2868 13536 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 2780 13536 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 2692 13536 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13496 2604 13536 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 3220 13455 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 3132 13455 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 3044 13455 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 2956 13455 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 2868 13455 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 2780 13455 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 2692 13455 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13415 2604 13455 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 3220 13374 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 3132 13374 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 3044 13374 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 2956 13374 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 2868 13374 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 2780 13374 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 2692 13374 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13334 2604 13374 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 3220 13293 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 3132 13293 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 3044 13293 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 2956 13293 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 2868 13293 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 2780 13293 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 2692 13293 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13253 2604 13293 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 3220 13212 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 3132 13212 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 3044 13212 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 2956 13212 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 2868 13212 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 2780 13212 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 2692 13212 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13172 2604 13212 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 3220 13131 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 3132 13131 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 3044 13131 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 2956 13131 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 2868 13131 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 2780 13131 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 2692 13131 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13091 2604 13131 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 3220 13050 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 3132 13050 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 3044 13050 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 2956 13050 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 2868 13050 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 2780 13050 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 2692 13050 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 13010 2604 13050 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 3220 12969 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 3132 12969 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 3044 12969 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 2956 12969 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 2868 12969 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 2780 12969 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 2692 12969 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12929 2604 12969 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 3220 12888 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 3132 12888 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 3044 12888 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 2956 12888 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 2868 12888 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 2780 12888 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 2692 12888 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12848 2604 12888 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 3220 12807 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 3132 12807 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 3044 12807 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 2956 12807 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 2868 12807 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 2780 12807 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 2692 12807 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12767 2604 12807 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 3220 12726 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 3132 12726 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 3044 12726 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 2956 12726 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 2868 12726 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 2780 12726 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 2692 12726 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12686 2604 12726 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 3220 12645 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 3132 12645 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 3044 12645 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 2956 12645 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 2868 12645 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 2780 12645 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 2692 12645 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12605 2604 12645 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 3220 12564 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 3132 12564 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 3044 12564 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 2956 12564 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 2868 12564 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 2780 12564 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 2692 12564 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12524 2604 12564 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 3220 12483 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 3132 12483 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 3044 12483 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 2956 12483 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 2868 12483 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 2780 12483 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 2692 12483 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12443 2604 12483 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 3220 12402 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 3132 12402 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 3044 12402 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 2956 12402 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 2868 12402 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 2780 12402 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 2692 12402 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12362 2604 12402 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 3220 12321 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 3132 12321 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 3044 12321 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 2956 12321 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 2868 12321 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 2780 12321 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 2692 12321 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12281 2604 12321 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 3220 12240 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 3132 12240 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 3044 12240 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 2956 12240 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 2868 12240 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 2780 12240 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 2692 12240 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12200 2604 12240 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 3220 12159 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 3132 12159 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 3044 12159 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 2956 12159 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 2868 12159 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 2780 12159 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 2692 12159 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12119 2604 12159 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 3220 12078 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 3132 12078 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 3044 12078 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 2956 12078 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 2868 12078 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 2780 12078 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 2692 12078 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 12038 2604 12078 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 3220 11997 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 3132 11997 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 3044 11997 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 2956 11997 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 2868 11997 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 2780 11997 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 2692 11997 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11957 2604 11997 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 3220 11916 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 3132 11916 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 3044 11916 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 2956 11916 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 2868 11916 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 2780 11916 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 2692 11916 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11876 2604 11916 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 3220 11835 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 3132 11835 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 3044 11835 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 2956 11835 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 2868 11835 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 2780 11835 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 2692 11835 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11795 2604 11835 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 3220 11754 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 3132 11754 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 3044 11754 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 2956 11754 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 2868 11754 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 2780 11754 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 2692 11754 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11714 2604 11754 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 3220 11673 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 3132 11673 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 3044 11673 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 2956 11673 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 2868 11673 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 2780 11673 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 2692 11673 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11633 2604 11673 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 3220 11592 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 3132 11592 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 3044 11592 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 2956 11592 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 2868 11592 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 2780 11592 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 2692 11592 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11552 2604 11592 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 3220 11511 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 3132 11511 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 3044 11511 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 2956 11511 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 2868 11511 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 2780 11511 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 2692 11511 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11471 2604 11511 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 3220 11430 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 3132 11430 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 3044 11430 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 2956 11430 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 2868 11430 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 2780 11430 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 2692 11430 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11390 2604 11430 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 3220 11349 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 3132 11349 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 3044 11349 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 2956 11349 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 2868 11349 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 2780 11349 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 2692 11349 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11309 2604 11349 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 3220 11268 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 3132 11268 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 3044 11268 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 2956 11268 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 2868 11268 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 2780 11268 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 2692 11268 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11228 2604 11268 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 3220 11187 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 3132 11187 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 3044 11187 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 2956 11187 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 2868 11187 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 2780 11187 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 2692 11187 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11147 2604 11187 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 3220 11106 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 3132 11106 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 3044 11106 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 2956 11106 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 2868 11106 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 2780 11106 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 2692 11106 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 11066 2604 11106 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 3220 11025 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 3132 11025 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 3044 11025 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 2956 11025 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 2868 11025 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 2780 11025 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 2692 11025 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10985 2604 11025 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 3220 10944 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 3132 10944 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 3044 10944 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 2956 10944 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 2868 10944 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 2780 10944 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 2692 10944 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10904 2604 10944 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 3220 10863 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 3132 10863 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 3044 10863 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 2956 10863 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 2868 10863 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 2780 10863 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 2692 10863 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10823 2604 10863 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 3220 10782 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 3132 10782 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 3044 10782 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 2956 10782 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 2868 10782 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 2780 10782 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 2692 10782 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10742 2604 10782 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 3220 10701 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 3132 10701 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 3044 10701 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 2956 10701 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 2868 10701 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 2780 10701 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 2692 10701 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10661 2604 10701 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 3220 10619 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 3132 10619 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 3044 10619 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 2956 10619 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 2868 10619 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 2780 10619 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 2692 10619 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10579 2604 10619 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 3220 10537 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 3132 10537 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 3044 10537 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 2956 10537 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 2868 10537 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 2780 10537 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 2692 10537 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10497 2604 10537 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 3220 10455 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 3132 10455 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 3044 10455 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 2956 10455 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 2868 10455 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 2780 10455 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 2692 10455 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10415 2604 10455 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 3220 10373 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 3132 10373 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 3044 10373 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 2956 10373 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 2868 10373 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 2780 10373 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 2692 10373 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10333 2604 10373 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 3220 10291 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 3132 10291 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 3044 10291 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 2956 10291 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 2868 10291 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 2780 10291 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 2692 10291 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10251 2604 10291 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 3220 10209 3260 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 3132 10209 3172 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 3044 10209 3084 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 2956 10209 2996 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 2868 10209 2908 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 2780 10209 2820 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 2692 10209 2732 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 10169 2604 10209 2644 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 3208 4894 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 3208 4894 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 3120 4894 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 3120 4894 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 3032 4894 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 3032 4894 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 2944 4894 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 2944 4894 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 2856 4894 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 2856 4894 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 2768 4894 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 2768 4894 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 2680 4894 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 2680 4894 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4830 2592 4894 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4830 2592 4894 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 3208 4813 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 3208 4813 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 3120 4813 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 3120 4813 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 3032 4813 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 3032 4813 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 2944 4813 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 2944 4813 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 2856 4813 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 2856 4813 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 2768 4813 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 2768 4813 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 2680 4813 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 2680 4813 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4749 2592 4813 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4749 2592 4813 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 3208 4732 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 3208 4732 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 3120 4732 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 3120 4732 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 3032 4732 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 3032 4732 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 2944 4732 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 2944 4732 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 2856 4732 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 2856 4732 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 2768 4732 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 2768 4732 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 2680 4732 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 2680 4732 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4668 2592 4732 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4668 2592 4732 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 3208 4651 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 3208 4651 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 3120 4651 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 3120 4651 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 3032 4651 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 3032 4651 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 2944 4651 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 2944 4651 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 2856 4651 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 2856 4651 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 2768 4651 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 2768 4651 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 2680 4651 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 2680 4651 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4587 2592 4651 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4587 2592 4651 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 3208 4570 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 3208 4570 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 3120 4570 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 3120 4570 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 3032 4570 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 3032 4570 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 2944 4570 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 2944 4570 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 2856 4570 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 2856 4570 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 2768 4570 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 2768 4570 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 2680 4570 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 2680 4570 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4506 2592 4570 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4506 2592 4570 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 3208 4489 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 3208 4489 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 3120 4489 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 3120 4489 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 3032 4489 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 3032 4489 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 2944 4489 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 2944 4489 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 2856 4489 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 2856 4489 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 2768 4489 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 2768 4489 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 2680 4489 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 2680 4489 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4425 2592 4489 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4425 2592 4489 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 3208 4408 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 3208 4408 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 3120 4408 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 3120 4408 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 3032 4408 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 3032 4408 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 2944 4408 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 2944 4408 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 2856 4408 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 2856 4408 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 2768 4408 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 2768 4408 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 2680 4408 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 2680 4408 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4344 2592 4408 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4344 2592 4408 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 3208 4327 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 3208 4327 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 3120 4327 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 3120 4327 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 3032 4327 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 3032 4327 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 2944 4327 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 2944 4327 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 2856 4327 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 2856 4327 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 2768 4327 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 2768 4327 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 2680 4327 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 2680 4327 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4263 2592 4327 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4263 2592 4327 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 3208 4246 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 3208 4246 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 3120 4246 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 3120 4246 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 3032 4246 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 3032 4246 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 2944 4246 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 2944 4246 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 2856 4246 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 2856 4246 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 2768 4246 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 2768 4246 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 2680 4246 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 2680 4246 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4182 2592 4246 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4182 2592 4246 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 3208 4165 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 3208 4165 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 3120 4165 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 3120 4165 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 3032 4165 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 3032 4165 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 2944 4165 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 2944 4165 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 2856 4165 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 2856 4165 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 2768 4165 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 2768 4165 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 2680 4165 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 2680 4165 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4101 2592 4165 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4101 2592 4165 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 3208 4084 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 3208 4084 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 3120 4084 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 3120 4084 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 3032 4084 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 3032 4084 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 2944 4084 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 2944 4084 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 2856 4084 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 2856 4084 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 2768 4084 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 2768 4084 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 2680 4084 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 2680 4084 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 4020 2592 4084 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 4020 2592 4084 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 3208 4003 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 3208 4003 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 3120 4003 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 3120 4003 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 3032 4003 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 3032 4003 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 2944 4003 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 2944 4003 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 2856 4003 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 2856 4003 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 2768 4003 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 2768 4003 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 2680 4003 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 2680 4003 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3939 2592 4003 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3939 2592 4003 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 3208 3922 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 3208 3922 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 3120 3922 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 3120 3922 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 3032 3922 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 3032 3922 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 2944 3922 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 2944 3922 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 2856 3922 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 2856 3922 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 2768 3922 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 2768 3922 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 2680 3922 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 2680 3922 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3858 2592 3922 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3858 2592 3922 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 3208 3841 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 3208 3841 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 3120 3841 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 3120 3841 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 3032 3841 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 3032 3841 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 2944 3841 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 2944 3841 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 2856 3841 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 2856 3841 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 2768 3841 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 2768 3841 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 2680 3841 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 2680 3841 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3777 2592 3841 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3777 2592 3841 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 3208 3760 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 3208 3760 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 3120 3760 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 3120 3760 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 3032 3760 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 3032 3760 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 2944 3760 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 2944 3760 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 2856 3760 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 2856 3760 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 2768 3760 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 2768 3760 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 2680 3760 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 2680 3760 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3696 2592 3760 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3696 2592 3760 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 3208 3679 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 3208 3679 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 3120 3679 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 3120 3679 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 3032 3679 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 3032 3679 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 2944 3679 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 2944 3679 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 2856 3679 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 2856 3679 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 2768 3679 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 2768 3679 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 2680 3679 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 2680 3679 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3615 2592 3679 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3615 2592 3679 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 3208 3598 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 3208 3598 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 3120 3598 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 3120 3598 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 3032 3598 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 3032 3598 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 2944 3598 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 2944 3598 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 2856 3598 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 2856 3598 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 2768 3598 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 2768 3598 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 2680 3598 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 2680 3598 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3534 2592 3598 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3534 2592 3598 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 3208 3517 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 3208 3517 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 3120 3517 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 3120 3517 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 3032 3517 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 3032 3517 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 2944 3517 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 2944 3517 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 2856 3517 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 2856 3517 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 2768 3517 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 2768 3517 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 2680 3517 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 2680 3517 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3453 2592 3517 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3453 2592 3517 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 3208 3436 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 3208 3436 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 3120 3436 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 3120 3436 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 3032 3436 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 3032 3436 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 2944 3436 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 2944 3436 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 2856 3436 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 2856 3436 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 2768 3436 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 2768 3436 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 2680 3436 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 2680 3436 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3372 2592 3436 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3372 2592 3436 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 3208 3355 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 3208 3355 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 3120 3355 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 3120 3355 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 3032 3355 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 3032 3355 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 2944 3355 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 2944 3355 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 2856 3355 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 2856 3355 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 2768 3355 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 2768 3355 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 2680 3355 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 2680 3355 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3291 2592 3355 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3291 2592 3355 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 3208 3274 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 3208 3274 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 3120 3274 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 3120 3274 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 3032 3274 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 3032 3274 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 2944 3274 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 2944 3274 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 2856 3274 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 2856 3274 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 2768 3274 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 2768 3274 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 2680 3274 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 2680 3274 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3210 2592 3274 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3210 2592 3274 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 3208 3193 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 3208 3193 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 3120 3193 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 3120 3193 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 3032 3193 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 3032 3193 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 2944 3193 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 2944 3193 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 2856 3193 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 2856 3193 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 2768 3193 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 2768 3193 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 2680 3193 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 2680 3193 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3129 2592 3193 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3129 2592 3193 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 3208 3112 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 3208 3112 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 3120 3112 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 3120 3112 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 3032 3112 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 3032 3112 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 2944 3112 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 2944 3112 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 2856 3112 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 2856 3112 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 2768 3112 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 2768 3112 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 2680 3112 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 2680 3112 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 3048 2592 3112 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 3048 2592 3112 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 3208 3031 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 3208 3031 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 3120 3031 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 3120 3031 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 3032 3031 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 3032 3031 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 2944 3031 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 2944 3031 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 2856 3031 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 2856 3031 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 2768 3031 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 2768 3031 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 2680 3031 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 2680 3031 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2967 2592 3031 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2967 2592 3031 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 3208 2950 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 3208 2950 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 3120 2950 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 3120 2950 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 3032 2950 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 3032 2950 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 2944 2950 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 2944 2950 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 2856 2950 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 2856 2950 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 2768 2950 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 2768 2950 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 2680 2950 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 2680 2950 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2886 2592 2950 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2886 2592 2950 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 3208 2869 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 3208 2869 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 3120 2869 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 3120 2869 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 3032 2869 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 3032 2869 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 2944 2869 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 2944 2869 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 2856 2869 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 2856 2869 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 2768 2869 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 2768 2869 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 2680 2869 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 2680 2869 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2805 2592 2869 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2805 2592 2869 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 3208 2788 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 3208 2788 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 3120 2788 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 3120 2788 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 3032 2788 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 3032 2788 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 2944 2788 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 2944 2788 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 2856 2788 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 2856 2788 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 2768 2788 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 2768 2788 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 2680 2788 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 2680 2788 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2724 2592 2788 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2724 2592 2788 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 3208 2707 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 3208 2707 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 3120 2707 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 3120 2707 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 3032 2707 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 3032 2707 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 2944 2707 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 2944 2707 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 2856 2707 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 2856 2707 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 2768 2707 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 2768 2707 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 2680 2707 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 2680 2707 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2643 2592 2707 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2643 2592 2707 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 3208 2626 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 3208 2626 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 3120 2626 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 3120 2626 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 3032 2626 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 3032 2626 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 2944 2626 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 2944 2626 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 2856 2626 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 2856 2626 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 2768 2626 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 2768 2626 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 2680 2626 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 2680 2626 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2562 2592 2626 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2562 2592 2626 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 3208 2545 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 3208 2545 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 3120 2545 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 3120 2545 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 3032 2545 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 3032 2545 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 2944 2545 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 2944 2545 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 2856 2545 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 2856 2545 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 2768 2545 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 2768 2545 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 2680 2545 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 2680 2545 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2481 2592 2545 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2481 2592 2545 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 3208 2464 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 3208 2464 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 3120 2464 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 3120 2464 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 3032 2464 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 3032 2464 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 2944 2464 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 2944 2464 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 2856 2464 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 2856 2464 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 2768 2464 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 2768 2464 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 2680 2464 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 2680 2464 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2400 2592 2464 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2400 2592 2464 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 3208 2383 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 3208 2383 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 3120 2383 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 3120 2383 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 3032 2383 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 3032 2383 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 2944 2383 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 2944 2383 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 2856 2383 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 2856 2383 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 2768 2383 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 2768 2383 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 2680 2383 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 2680 2383 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2319 2592 2383 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2319 2592 2383 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 3208 2302 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 3208 2302 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 3120 2302 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 3120 2302 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 3032 2302 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 3032 2302 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 2944 2302 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 2944 2302 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 2856 2302 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 2856 2302 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 2768 2302 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 2768 2302 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 2680 2302 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 2680 2302 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2238 2592 2302 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2238 2592 2302 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 3208 2221 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 3208 2221 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 3120 2221 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 3120 2221 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 3032 2221 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 3032 2221 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 2944 2221 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 2944 2221 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 2856 2221 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 2856 2221 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 2768 2221 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 2768 2221 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 2680 2221 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 2680 2221 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2157 2592 2221 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2157 2592 2221 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 3208 2140 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 3208 2140 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 3120 2140 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 3120 2140 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 3032 2140 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 3032 2140 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 2944 2140 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 2944 2140 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 2856 2140 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 2856 2140 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 2768 2140 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 2768 2140 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 2680 2140 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 2680 2140 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 2076 2592 2140 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 2076 2592 2140 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 3208 2059 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 3208 2059 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 3120 2059 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 3120 2059 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 3032 2059 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 3032 2059 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 2944 2059 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 2944 2059 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 2856 2059 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 2856 2059 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 2768 2059 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 2768 2059 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 2680 2059 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 2680 2059 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1995 2592 2059 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1995 2592 2059 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 3208 1978 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 3208 1978 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 3120 1978 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 3120 1978 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 3032 1978 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 3032 1978 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 2944 1978 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 2944 1978 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 2856 1978 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 2856 1978 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 2768 1978 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 2768 1978 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 2680 1978 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 2680 1978 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1914 2592 1978 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1914 2592 1978 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 3208 1897 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 3208 1897 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 3120 1897 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 3120 1897 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 3032 1897 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 3032 1897 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 2944 1897 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 2944 1897 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 2856 1897 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 2856 1897 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 2768 1897 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 2768 1897 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 2680 1897 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 2680 1897 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1833 2592 1897 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1833 2592 1897 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 3208 1816 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 3208 1816 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 3120 1816 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 3120 1816 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 3032 1816 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 3032 1816 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 2944 1816 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 2944 1816 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 2856 1816 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 2856 1816 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 2768 1816 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 2768 1816 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 2680 1816 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 2680 1816 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1752 2592 1816 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1752 2592 1816 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 3208 1735 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 3208 1735 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 3120 1735 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 3120 1735 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 3032 1735 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 3032 1735 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 2944 1735 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 2944 1735 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 2856 1735 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 2856 1735 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 2768 1735 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 2768 1735 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 2680 1735 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 2680 1735 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1671 2592 1735 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1671 2592 1735 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 3208 1654 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 3208 1654 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 3120 1654 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 3120 1654 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 3032 1654 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 3032 1654 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 2944 1654 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 2944 1654 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 2856 1654 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 2856 1654 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 2768 1654 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 2768 1654 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 2680 1654 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 2680 1654 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1590 2592 1654 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1590 2592 1654 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 3208 1573 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 3208 1573 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 3120 1573 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 3120 1573 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 3032 1573 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 3032 1573 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 2944 1573 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 2944 1573 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 2856 1573 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 2856 1573 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 2768 1573 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 2768 1573 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 2680 1573 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 2680 1573 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1509 2592 1573 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1509 2592 1573 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 3208 1492 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 3208 1492 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 3120 1492 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 3120 1492 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 3032 1492 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 3032 1492 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 2944 1492 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 2944 1492 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 2856 1492 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 2856 1492 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 2768 1492 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 2768 1492 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 2680 1492 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 2680 1492 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1428 2592 1492 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1428 2592 1492 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 3208 1411 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 3208 1411 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 3120 1411 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 3120 1411 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 3032 1411 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 3032 1411 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 2944 1411 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 2944 1411 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 2856 1411 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 2856 1411 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 2768 1411 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 2768 1411 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 2680 1411 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 2680 1411 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1347 2592 1411 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1347 2592 1411 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 3208 1330 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 3208 1330 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 3120 1330 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 3120 1330 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 3032 1330 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 3032 1330 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 2944 1330 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 2944 1330 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 2856 1330 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 2856 1330 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 2768 1330 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 2768 1330 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 2680 1330 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 2680 1330 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1266 2592 1330 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1266 2592 1330 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 3208 1249 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 3208 1249 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 3120 1249 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 3120 1249 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 3032 1249 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 3032 1249 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 2944 1249 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 2944 1249 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 2856 1249 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 2856 1249 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 2768 1249 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 2768 1249 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 2680 1249 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 2680 1249 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1185 2592 1249 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1185 2592 1249 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 3208 1168 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 3208 1168 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 3120 1168 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 3120 1168 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 3032 1168 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 3032 1168 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 2944 1168 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 2944 1168 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 2856 1168 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 2856 1168 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 2768 1168 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 2768 1168 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 2680 1168 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 2680 1168 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1104 2592 1168 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1104 2592 1168 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 3208 1087 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 3208 1087 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 3120 1087 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 3120 1087 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 3032 1087 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 3032 1087 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 2944 1087 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 2944 1087 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 2856 1087 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 2856 1087 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 2768 1087 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 2768 1087 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 2680 1087 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 2680 1087 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 1023 2592 1087 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 1023 2592 1087 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 3208 1006 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 3208 1006 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 3120 1006 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 3120 1006 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 3032 1006 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 3032 1006 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 2944 1006 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 2944 1006 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 2856 1006 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 2856 1006 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 2768 1006 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 2768 1006 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 2680 1006 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 2680 1006 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 942 2592 1006 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 942 2592 1006 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 3208 925 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 3208 925 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 3120 925 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 3120 925 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 3032 925 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 3032 925 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 2944 925 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 2944 925 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 2856 925 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 2856 925 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 2768 925 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 2768 925 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 2680 925 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 2680 925 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 861 2592 925 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 861 2592 925 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 3208 844 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 3208 844 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 3120 844 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 3120 844 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 3032 844 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 3032 844 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 2944 844 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 2944 844 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 2856 844 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 2856 844 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 2768 844 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 2768 844 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 2680 844 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 2680 844 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 780 2592 844 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 780 2592 844 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 3208 763 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 3208 763 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 3120 763 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 3120 763 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 3032 763 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 3032 763 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 2944 763 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 2944 763 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 2856 763 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 2856 763 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 2768 763 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 2768 763 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 2680 763 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 2680 763 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 699 2592 763 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 699 2592 763 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 3208 682 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 3208 682 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 3120 682 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 3120 682 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 3032 682 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 3032 682 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 2944 682 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 2944 682 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 2856 682 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 2856 682 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 2768 682 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 2768 682 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 2680 682 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 2680 682 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 618 2592 682 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 618 2592 682 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 3208 600 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 3208 600 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 3120 600 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 3120 600 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 3032 600 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 3032 600 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 2944 600 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 2944 600 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 2856 600 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 2856 600 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 2768 600 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 2768 600 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 2680 600 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 2680 600 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 536 2592 600 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 536 2592 600 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 3208 518 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 3208 518 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 3120 518 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 3120 518 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 3032 518 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 3032 518 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 2944 518 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 2944 518 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 2856 518 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 2856 518 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 2768 518 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 2768 518 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 2680 518 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 2680 518 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 454 2592 518 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 454 2592 518 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 3208 436 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 3208 436 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 3120 436 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 3120 436 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 3032 436 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 3032 436 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 2944 436 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 2944 436 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 2856 436 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 2856 436 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 2768 436 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 2768 436 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 2680 436 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 2680 436 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 372 2592 436 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 372 2592 436 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 3208 354 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 3208 354 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 3120 354 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 3120 354 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 3032 354 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 3032 354 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 2944 354 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 2944 354 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 2856 354 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 2856 354 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 2768 354 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 2768 354 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 2680 354 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 2680 354 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 290 2592 354 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 290 2592 354 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 3208 272 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 3208 272 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 3120 272 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 3120 272 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 3032 272 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 3032 272 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 2944 272 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 2944 272 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 2856 272 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 2856 272 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 2768 272 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 2768 272 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 2680 272 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 2680 272 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal4 s 208 2592 272 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 208 2592 272 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 3208 190 3272 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 3120 190 3184 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 3032 190 3096 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 2944 190 3008 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 2856 190 2920 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 2768 190 2832 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 2680 190 2744 6 VDDA
port 4 nsew power bidirectional
rlabel metal3 s 126 2592 190 2656 6 VDDA
port 4 nsew power bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 5 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 5 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 5 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 5 nsew ground bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 6 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 6 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 7 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 8 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 8 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 10 nsew ground bidirectional
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 675976
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 607096
<< end >>
