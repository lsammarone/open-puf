magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 833 157 1287 203
rect 1 21 1287 157
rect 30 -17 64 21
<< locali >>
rect 17 197 66 325
rect 292 191 358 265
rect 1131 375 1185 493
rect 1151 300 1185 375
rect 1151 285 1271 300
rect 1152 283 1271 285
rect 1153 282 1271 283
rect 1155 277 1271 282
rect 896 199 1034 265
rect 1157 178 1271 277
rect 1154 173 1271 178
rect 1151 153 1271 173
rect 1151 97 1185 153
rect 1119 51 1185 97
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 156 393
rect 122 280 156 359
rect 203 337 248 493
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 237 337
rect 291 333 357 483
rect 391 367 454 527
rect 555 451 721 485
rect 291 299 428 333
rect 392 219 428 299
rect 494 271 551 401
rect 585 283 653 399
rect 585 229 619 283
rect 687 265 721 451
rect 760 427 822 527
rect 856 427 912 527
rect 946 373 984 493
rect 1018 375 1092 527
rect 764 341 984 373
rect 764 307 1117 341
rect 1083 265 1117 307
rect 1219 334 1271 527
rect 687 249 862 265
rect 392 157 468 219
rect 307 153 468 157
rect 307 123 428 153
rect 535 141 619 229
rect 666 205 862 249
rect 307 69 341 123
rect 666 107 700 205
rect 1070 199 1123 265
rect 1083 165 1117 199
rect 375 17 441 89
rect 562 73 700 107
rect 848 131 1117 165
rect 747 17 814 106
rect 848 51 918 131
rect 1019 17 1085 97
rect 1219 17 1271 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< obsm1 >>
rect 202 388 260 397
rect 482 388 540 397
rect 202 360 540 388
rect 202 351 260 360
rect 482 351 540 360
rect 110 320 168 329
rect 574 320 632 329
rect 110 292 632 320
rect 110 283 168 292
rect 574 283 632 292
<< labels >>
rlabel locali s 292 191 358 265 6 D
port 1 nsew signal input
rlabel locali s 17 197 66 325 6 GATE_N
port 2 nsew clock input
rlabel locali s 896 199 1034 265 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 1288 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1287 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 833 157 1287 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1326 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1288 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1119 51 1185 97 6 Q
port 8 nsew signal output
rlabel locali s 1151 97 1185 153 6 Q
port 8 nsew signal output
rlabel locali s 1151 153 1271 173 6 Q
port 8 nsew signal output
rlabel locali s 1154 173 1271 178 6 Q
port 8 nsew signal output
rlabel locali s 1157 178 1271 277 6 Q
port 8 nsew signal output
rlabel locali s 1155 277 1271 282 6 Q
port 8 nsew signal output
rlabel locali s 1153 282 1271 283 6 Q
port 8 nsew signal output
rlabel locali s 1152 283 1271 285 6 Q
port 8 nsew signal output
rlabel locali s 1151 285 1271 300 6 Q
port 8 nsew signal output
rlabel locali s 1151 300 1185 375 6 Q
port 8 nsew signal output
rlabel locali s 1131 375 1185 493 6 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1288 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2747906
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2736500
<< end >>
