magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 9 67 1195 203
rect 29 -17 63 67
rect 294 21 1195 67
<< locali >>
rect 85 199 156 339
rect 190 199 247 265
rect 580 289 799 341
rect 715 181 799 289
rect 833 215 992 255
rect 1026 215 1179 255
rect 412 145 1090 181
rect 412 51 478 145
rect 580 51 646 145
rect 856 51 922 145
rect 1024 51 1090 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 411 69 491
rect 103 448 169 527
rect 328 459 730 493
rect 328 445 394 459
rect 496 443 730 459
rect 772 443 998 493
rect 17 377 383 411
rect 17 165 51 377
rect 199 305 315 343
rect 281 249 315 305
rect 349 317 383 377
rect 428 409 462 425
rect 428 375 922 409
rect 428 359 462 375
rect 349 283 546 317
rect 864 291 922 375
rect 956 325 998 443
rect 1032 359 1074 527
rect 1108 325 1174 493
rect 956 291 1174 325
rect 512 255 546 283
rect 281 215 478 249
rect 512 215 681 255
rect 281 165 315 215
rect 17 90 93 165
rect 127 17 161 165
rect 211 131 315 165
rect 211 90 250 131
rect 312 17 378 96
rect 512 17 546 111
rect 680 17 822 111
rect 956 17 990 111
rect 1124 17 1179 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 1026 215 1179 255 6 A
port 1 nsew signal input
rlabel locali s 833 215 992 255 6 B
port 2 nsew signal input
rlabel locali s 190 199 247 265 6 C_N
port 3 nsew signal input
rlabel locali s 85 199 156 339 6 D_N
port 4 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 294 21 1195 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 29 -17 63 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 9 67 1195 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1024 51 1090 145 6 Y
port 9 nsew signal output
rlabel locali s 856 51 922 145 6 Y
port 9 nsew signal output
rlabel locali s 580 51 646 145 6 Y
port 9 nsew signal output
rlabel locali s 412 51 478 145 6 Y
port 9 nsew signal output
rlabel locali s 412 145 1090 181 6 Y
port 9 nsew signal output
rlabel locali s 715 181 799 289 6 Y
port 9 nsew signal output
rlabel locali s 580 289 799 341 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1215418
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1206094
<< end >>
