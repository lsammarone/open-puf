* NGSPICE file created from BR128_lvs_tap_flat.ext - technology: sky130A

.subckt BR128_lvs_tap_flat VDD VSS OUT C[127] C[126] C[125] C[124] C[123] C[122] C[121] C[120]
+ C[119] C[118] C[117] C[116] C[115] C[114] C[113] C[112] C[111] C[110] C[109] C[108]
+ C[107] C[106] C[105] C[104] C[103] C[102] C[101] C[100] C[99] C[98] C[97] C[96]
+ C[95] C[94] C[93] C[92] C[91] C[90] C[89] C[88] C[87] C[86] C[85] C[84] C[83] C[82]
+ C[81] C[80] C[79] C[78] C[77] C[76] C[75] C[74] C[73] C[72] C[71] C[70] C[69] C[68]
+ C[67] C[66] C[65] C[64] C[63] C[62] C[61] C[60] C[59] C[58] C[57] C[56] C[55] C[54]
+ C[53] C[52] C[51] C[50] C[49] C[48] C[47] C[46] C[45] C[44] C[43] C[42] C[41] C[40]
+ C[39] C[38] C[37] C[36] C[35] C[34] C[33] C[32] C[31] C[30] C[29] C[28] C[27] C[26]
+ C[25] C[24] C[23] C[22] C[21] C[20] C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12]
+ C[11] C[10] C[9] C[8] C[7] C[6] C[5] C[4] C[3] C[2] C[1] C[0] RESET
X0 a_58650_6655# a_57775_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=3.37905e+14p ps=3.18564e+09u w=790000u l=150000u
X1 a_29545_1829# a_28953_690# a_27559_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2 a_10802_n5622# a_10308_n5789# a_10363_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3 a_55834_n5879# a_55608_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=2.14887e+14p ps=2.29896e+09u w=650000u l=150000u
X4 a_12573_7009# a_12571_5953# a_12874_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X5 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X6 VSS a_25900_n5622# a_26825_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X7 a_14676_n6678# a_14310_n5879# a_12690_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X8 VDD C[6] a_47717_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X9 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X10 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X11 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X12 a_48321_773# a_49715_690# a_49765_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X13 VSS a_53985_773# a_54910_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X14 a_20236_n5622# a_21856_n5879# a_21680_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X15 a_37685_n6843# a_37326_n6678# a_37324_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X16 VDD a_34341_n11370# a_34291_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X17 VDD a_4909_773# a_5834_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X18 VDD a_44283_836# a_44107_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X19 a_37338_n10732# a_36572_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X20 a_25685_5953# a_25067_6408# a_25285_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X21 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_6532_n5789# C[35] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X23 a_22222_n6678# a_21630_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X24 VSS a_37228_n5622# a_38153_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X25 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X26 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X27 VDD a_818_1932# a_776_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X28 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X29 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X30 a_2228_696# a_2058_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X31 a_37641_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X32 a_47908_5708# a_47935_6449# a_47920_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X33 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_20649_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X35 VSS a_44780_n5622# a_45705_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X36 a_52193_773# a_51603_690# a_52097_773# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X37 a_48149_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X38 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_33237_5953# a_34507_6408# a_34698_5708# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X40 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X41 VSS a_54874_6655# a_54824_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X42 a_40873_1829# a_40507_836# a_38887_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X43 VDD a_20896_6655# a_20846_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X44 a_29461_5953# a_28791_6434# a_29061_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X45 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X46 VDD a_36229_n11370# a_36179_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X47 VDD a_39776_6655# a_39726_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X48 a_39226_n10732# a_38460_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X49 VDD a_2022_6655# a_1972_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X50 a_5005_773# a_4415_690# a_4909_773# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X51 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X52 a_20103_773# a_19739_836# a_20007_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X53 a_41102_n6678# a_40510_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X54 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X55 a_52193_773# a_52195_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X56 VSS a_49605_6408# a_49553_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X57 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X58 a_32729_690# C[113] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X59 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X60 VDD a_51722_n11559# a_51940_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X61 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 a_22537_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X63 a_55663_n6843# a_55658_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X64 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X65 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X66 VDD a_20007_773# a_20932_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X67 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X68 a_51829_836# a_51603_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X69 a_24108_n5622# a_24110_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X70 VDD a_31249_n6869# a_32021_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X71 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X72 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X73 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X74 VDD a_31249_n6869# a_33909_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X75 a_35524_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X76 VDD a_21125_n11370# a_21075_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X77 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X78 VSS a_818_1932# a_14445_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X79 VDD a_15627_6408# a_15845_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X80 a_18229_5953# a_17515_6408# a_18133_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X81 VSS a_46347_n6869# a_50534_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X82 a_3133_7009# a_2417_6408# a_1147_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X83 a_16558_n6678# a_15966_n5789# a_14578_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X84 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X85 a_47964_1994# a_47877_1896# a_47882_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X86 a_14459_5953# a_13693_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X87 VDD a_53610_n11559# a_53828_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X88 a_42677_5953# a_42059_6408# a_42277_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X89 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X90 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X91 a_53985_773# a_55379_690# a_55429_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X92 a_14139_n6843# a_14134_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X93 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X94 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X95 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X96 a_31748_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X97 VSS a_40885_5953# a_40887_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X98 a_42988_n5622# a_42990_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X99 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X100 a_7122_n5622# a_6758_n5879# a_7026_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X101 VSS a_51493_6408# a_51441_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X102 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X103 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X104 a_9010_n5622# a_8646_n5879# a_8914_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X105 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X106 a_35221_5953# a_34455_6434# a_35125_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X107 a_4909_773# a_4641_836# a_4470_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X108 VDD a_23013_n11370# a_22963_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X109 VSS a_29557_5953# a_29559_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X110 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X111 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 a_34547_n5795# a_34377_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X113 a_26010_n10732# a_25244_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X114 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 a_31564_n5622# a_31296_n5879# a_31125_n6843# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X116 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X117 VSS a_818_1932# a_13910_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X118 VDD a_39116_n5622# a_40041_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X119 VDD a_41004_n5622# a_41929_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X120 a_35438_n6678# a_34846_n5789# a_33452_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X121 VDD a_55498_n11559# a_55716_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X122 a_39130_n10732# a_40400_n11559# a_40591_n10487# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X123 a_37888_6655# a_37013_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X124 a_14578_n5622# a_14084_n5789# a_14139_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X125 a_1147_5953# a_2417_6408# a_2608_5708# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X126 VSS a_13350_6655# a_13300_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X127 VDD a_18080_n5879# a_17904_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X128 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X129 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X130 VDD a_19968_n5879# a_19792_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X131 a_41102_n6678# a_40510_n5789# a_39116_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X132 a_42990_n6678# a_42398_n5789# a_41004_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X133 a_11215_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X134 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X135 a_9780_696# a_9610_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X136 VDD a_36395_6408# a_36613_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X137 a_31445_5953# a_30679_6434# a_31349_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X138 a_12573_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X139 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X141 a_43758_696# a_43588_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X142 a_7026_n5622# a_6532_n5789# a_6587_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X143 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X144 a_7210_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X145 a_10669_773# a_10671_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X146 a_52783_n6843# a_52424_n6678# a_52422_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X147 a_3035_5953# a_4253_6434# a_4496_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X148 a_8191_690# C[100] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X149 a_27898_n10732# a_27132_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X150 a_13579_n11370# a_12704_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X151 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X152 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X153 VDD a_9969_6408# a_9917_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X154 a_37111_7009# a_37109_5953# a_37412_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X155 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X156 VSS a_52326_n5622# a_53251_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X157 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X158 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X160 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X161 a_18348_n5622# a_19742_n5789# a_19792_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X162 VDD a_57386_n11559# a_57604_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X163 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X164 VSS C[18] a_25067_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X165 VSS a_29447_773# a_30372_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X166 a_33550_n6678# a_32958_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X167 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X168 a_35221_5953# a_34507_6408# a_35125_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X169 VDD a_38848_n5879# a_38672_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X170 VDD a_46347_n6869# a_48193_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X171 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X172 VSS a_31445_5953# a_31447_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X173 VSS a_59878_n5622# a_60803_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X174 a_13103_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X175 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X176 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X177 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X178 a_29559_7009# a_28791_6434# a_27573_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X179 a_3434_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X180 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X181 a_17625_690# C[105] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X182 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X183 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X184 a_12048_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X185 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X186 VDD a_16145_n6869# a_18805_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X187 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X188 a_42775_7009# a_42059_6408# a_40789_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X189 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X190 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X191 VDD a_46347_n6869# a_55745_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X192 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X193 a_18444_n5622# a_17854_n5789# a_18348_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X194 a_37013_5953# a_36343_6434# a_36613_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X195 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X196 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X197 a_12461_773# a_13855_690# a_13905_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X198 VSS a_15916_1932# a_18215_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X199 VDD a_59274_n11559# a_59492_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X200 a_18229_5953# a_17463_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X201 a_9574_6655# a_8699_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X202 a_46447_5953# a_45829_6408# a_46047_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X203 a_24108_n5622# a_23518_n5789# a_24012_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X204 a_25996_n5622# a_25406_n5789# a_25900_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X205 a_1474_n11788# a_706_n11533# a_453_n11561# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X206 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X207 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X208 VSS a_52097_773# a_53022_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X209 OUT a_60574_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X210 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X211 a_13785_n5795# a_13615_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X212 VSS a_16145_n6869# a_17909_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X213 VSS a_16145_n6869# a_19797_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X214 a_22005_5953# a_21239_6434# a_21909_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X215 a_3131_5953# a_2365_6434# a_3035_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X216 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X217 VDD a_18348_n5622# a_19273_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X218 VDD a_32848_n11559# a_32796_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X219 VDD a_31249_n6869# a_37685_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X220 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X221 VSS a_16145_n6869# a_25461_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X222 VSS a_19621_6449# a_19594_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X223 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X224 a_37324_n5622# a_36734_n5789# a_37228_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X225 a_7439_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X226 a_37456_1994# a_37097_1829# a_37095_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X227 VDD a_46118_1932# a_51740_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X228 a_16460_n5622# a_16192_n5879# a_16021_n6843# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X229 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X230 a_52986_6655# a_52111_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X231 VDD a_25900_n5622# a_26825_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X232 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 a_8797_7009# a_8795_5953# a_9098_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X234 a_25270_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X235 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X236 a_4923_5953# a_4305_6408# a_4523_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X237 a_25781_5953# a_25067_6408# a_25685_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X238 a_52195_1829# a_51603_690# a_50209_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X239 a_44876_n5622# a_44286_n5789# a_44780_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X240 a_3362_n11788# a_2594_n11533# a_1376_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X241 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 VSS a_17120_6655# a_17070_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X243 a_24012_n5622# a_23744_n5879# a_23573_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X244 a_31660_n5622# a_31296_n5879# a_31564_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X245 VSS a_31249_n6869# a_38677_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X246 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X247 VDD C[24] a_13745_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X248 a_55887_5953# a_57105_6434# a_57348_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X249 VDD a_6027_n11370# a_5977_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X250 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X251 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X252 VSS C[9] a_42059_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X253 a_16343_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X254 VDD a_37228_n5622# a_38153_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X255 VDD a_34736_n11559# a_34684_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X256 VSS C[64] a_59274_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X257 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X258 VSS a_2864_n11298# a_2837_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X259 VSS a_31249_n6869# a_44341_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X260 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X261 a_35340_n5622# a_35072_n5879# a_34901_n6843# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X262 a_52438_n11788# a_51670_n11533# a_50452_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X263 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X264 a_8699_5953# a_8029_6434# a_8299_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X265 a_47827_690# C[121] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X266 VDD a_44780_n5622# a_45705_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X267 a_52438_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X268 a_27294_n5789# C[46] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X269 a_50536_n6678# a_49944_n5789# a_48550_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X270 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X271 a_13936_5708# a_13963_6449# a_13948_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X272 a_56286_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X273 VDD a_46058_n11559# a_46276_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X274 a_29690_n10732# a_30960_n11559# a_31151_n10487# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X275 a_5250_n11788# a_4482_n11533# a_3264_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X276 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X277 VSS a_31020_1932# a_35207_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X278 a_42892_n5622# a_42624_n5879# a_42453_n6843# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X279 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X280 VDD a_15916_1932# a_24240_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X281 VSS a_51940_n11298# a_51913_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X282 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X283 a_35221_5953# a_34455_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X284 a_2753_836# a_2527_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X285 VDD a_36624_n11559# a_36572_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X286 a_52111_5953# a_51441_6434# a_51711_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X287 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X288 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X289 a_4923_5953# a_4253_6434# a_4523_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X290 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X291 a_56559_n6843# a_56200_n6678# a_56198_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X292 a_46545_7009# a_45829_6408# a_44565_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X293 a_28016_1994# a_27657_1829# a_27655_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X294 a_9142_1994# a_8783_1829# a_8781_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X295 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 VDD a_46394_n5879# a_46218_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X297 a_54326_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X298 VDD a_15916_1932# a_20464_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X299 a_12559_1829# a_11967_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X300 a_27520_n5879# a_27294_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X301 a_55103_n11370# a_54228_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X302 a_1472_n10732# a_706_n11533# a_1376_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X303 a_37111_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X304 VDD a_47946_n11559# a_48164_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X305 a_27146_5708# a_27173_6449# a_27158_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X306 VSS a_53828_n11298# a_53801_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X307 a_42262_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X308 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X309 VDD a_52058_n5879# a_51882_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X310 VDD a_53946_n5879# a_53770_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X311 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X312 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X313 VDD a_38512_n11559# a_38460_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X314 a_29788_n11788# a_29020_n11533# a_27802_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X315 a_42773_5953# a_42059_6408# a_42677_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X316 a_2837_n10487# a_2864_n11298# a_2849_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X317 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X318 VSS a_34112_6655# a_34062_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X319 a_50548_n10732# a_49782_n11533# a_50452_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X320 a_57859_1829# a_57267_690# a_55873_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X321 VDD a_44551_773# a_45476_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X322 VDD a_57157_6408# a_57375_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X323 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X324 a_13992_1994# a_13905_1896# a_13910_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X325 VDD a_34843_836# a_34667_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X326 a_41116_n11788# a_40348_n11533# a_39130_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X327 a_56214_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X328 a_21331_n5795# a_21161_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X329 a_56991_n11370# a_56116_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X330 a_3360_n10732# a_2594_n11533# a_3264_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X331 a_29772_n5622# a_29182_n5789# a_29676_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X332 a_16556_n5622# a_16192_n5879# a_16460_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X333 a_51913_n10487# a_51940_n11298# a_51925_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X334 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X335 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X336 VSS a_55716_n11298# a_55689_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X337 VDD C[22] a_17515_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X338 a_25781_5953# a_25015_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X339 a_57873_7009# a_57871_5953# a_58174_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X340 a_53999_5953# a_53381_6408# a_53599_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X341 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X342 a_45939_690# C[120] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X343 a_58856_696# a_58686_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X344 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X345 a_10389_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X346 a_6907_5953# a_6141_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X347 VSS a_8914_n5622# a_9839_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X348 VSS C[7] a_45829_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X349 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X350 a_36731_836# a_36505_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X351 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X352 a_52436_n10732# a_51670_n11533# a_52340_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X353 VDD a_31020_1932# a_41232_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X354 VDD a_23408_n11559# a_23356_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X355 VSS a_52207_5953# a_52209_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X356 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X357 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X358 a_10009_n5795# a_9839_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X359 VDD a_46347_n6869# a_52783_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X360 a_44647_773# a_44057_690# a_44551_773# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X361 a_58102_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X362 VDD a_15916_1932# a_29904_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X363 a_45008_1994# a_44649_1829# a_44647_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X364 a_27349_n6843# a_27344_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X365 a_17706_5708# a_17733_6449# a_17718_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X366 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X367 a_865_836# a_639_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X368 VSS a_8299_6449# a_8272_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X369 a_32822_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X370 VSS a_15916_1932# a_25232_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X371 a_35436_n5622# a_35072_n5879# a_35340_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X372 a_53801_n10487# a_53828_n11298# a_53813_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X373 a_134_6655# a_224_6410# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X374 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X375 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X376 a_18362_n10732# a_19632_n11559# a_19823_n10487# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X377 VSS a_57604_n11298# a_57577_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X378 a_33013_n6843# a_33008_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X379 a_27898_n10732# a_27132_n11533# a_27802_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X380 VSS a_46347_n6869# a_51887_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X381 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X382 a_34901_n6843# a_34896_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X383 a_12277_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X384 a_57990_n5622# a_59384_n5789# a_59434_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X385 VSS a_46347_n6869# a_53775_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X386 VSS a_24672_6655# a_24622_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X387 a_10671_1829# a_10305_836# a_8685_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X388 a_42988_n5622# a_42624_n5879# a_42892_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X389 VDD a_52326_n5622# a_53251_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X390 VSS C[69] a_49834_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X391 a_8797_7009# a_8029_6434# a_6811_5953# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X392 a_4415_690# C[98] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X393 VSS a_16145_n6869# a_22220_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X394 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X395 VDD a_47717_6408# a_47935_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X396 VDD a_10198_n11559# a_10146_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X397 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X398 a_50438_n5622# a_50170_n5879# a_49999_n6843# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X399 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X400 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X401 a_21991_773# a_21993_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X402 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X403 VSS a_19403_6408# a_19351_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X404 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X405 VDD a_59878_n5622# a_60803_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X406 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X407 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X408 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X409 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X410 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X411 VSS C[31] a_529_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X412 a_48433_7009# a_48431_5953# a_48734_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X413 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X414 a_24878_696# a_24708_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X415 a_20250_n10732# a_21520_n11559# a_21711_n10487# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X416 a_55689_n10487# a_55716_n11298# a_55701_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X417 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X418 a_14674_n5622# a_14676_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X419 VSS C[82] a_25296_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X420 a_29786_n10732# a_29020_n11533# a_29690_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X421 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X422 a_46032_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X423 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X424 a_14165_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X425 a_52209_7009# a_51441_6434# a_50223_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X426 a_23289_690# C[108] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X427 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X428 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X429 a_46543_5953# a_45829_6408# a_46447_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X430 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X431 VSS a_4909_773# a_5834_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X432 VSS a_31249_n6869# a_41100_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X433 VDD a_56991_n11370# a_56941_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X434 VDD C[13] a_34507_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X435 a_7122_n5622# a_7124_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X436 VDD a_12086_n11559# a_12034_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X437 a_41114_n10732# a_40348_n11533# a_41018_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X438 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X439 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X440 a_44551_773# a_44283_836# a_44112_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X441 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X442 a_17762_1994# a_17675_1896# a_17680_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X443 a_13785_n5795# a_13615_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X444 VSS a_17962_n11298# a_17935_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X445 a_12475_5953# a_11857_6408# a_12075_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X446 a_14676_n6678# a_14084_n5789# a_12690_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X447 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X448 a_23783_773# a_25177_690# a_25227_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X449 a_47528_696# a_47358_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X450 a_57577_n10487# a_57604_n11298# a_57589_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X451 a_12461_773# a_11967_690# a_12022_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X452 VSS C[81] a_27184_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X453 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X454 a_38848_n5879# a_38622_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X455 VDD C[28] a_6193_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X456 a_34698_5708# a_34725_6449# a_34710_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X457 VSS a_21291_6408# a_21239_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X458 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X459 a_42759_773# a_42761_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X460 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X461 VDD a_58879_n11370# a_58829_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X462 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X463 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X464 a_60106_1994# a_59747_1829# a_59745_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X465 a_32021_n6843# a_31662_n6678# a_31660_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X466 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X467 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X468 VSS a_41664_6655# a_41614_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X469 a_453_n11561# a_758_n11559# a_949_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X470 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X471 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X472 a_20250_n10732# a_19632_n11559# a_19850_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X473 a_46774_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X474 VSS a_19850_n11298# a_19823_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X475 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X476 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X477 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X478 a_48778_1994# a_48419_1829# a_48417_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X479 a_59384_n5789# C[63] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X480 VSS a_31564_n5622# a_32489_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X481 a_10802_n5622# a_12422_n5879# a_12246_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X482 a_52111_5953# a_53381_6408# a_53572_5708# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X483 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X484 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X485 a_35111_773# a_34617_690# a_34672_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X486 a_32659_n5795# a_32489_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X487 VSS a_46276_n11298# a_46249_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X488 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X489 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X490 VSS a_20007_773# a_20932_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X491 a_10900_n6678# a_10308_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X492 a_19797_n6843# a_19792_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X493 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X494 VDD a_16145_n6869# a_27431_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X495 a_57873_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X496 VDD a_10305_836# a_10129_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X497 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X498 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X499 a_36999_773# a_36505_690# a_36560_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X500 VSS C[3] a_53381_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X501 a_27657_1829# a_27065_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X502 a_868_n5789# C[32] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X503 a_1376_n10732# a_2646_n11559# a_2837_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X504 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X505 VDD a_31020_1932# a_30978_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X506 a_17935_n10487# a_17962_n11298# a_17947_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X507 a_9012_n6678# a_8420_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X508 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X509 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X510 a_12193_836# a_11967_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X511 a_1005_n6843# a_918_n6611# a_923_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X512 a_1362_n5622# a_2756_n5789# a_2806_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X513 a_34754_1994# a_34667_1896# a_34672_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X514 a_50534_n5622# a_50170_n5879# a_50438_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X515 a_38677_n6843# a_38672_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X516 a_18458_n10732# a_17692_n11533# a_18362_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X517 a_35125_5953# a_36343_6434# a_36586_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X518 VSS a_33066_n11298# a_33039_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X519 a_49210_6655# a_48335_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X520 VSS a_46118_1932# a_46529_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X521 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X522 VDD a_23179_6408# a_23127_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X523 a_40775_773# a_42169_690# a_42219_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X524 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X525 VDD a_1047_n6869# a_15035_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X526 VDD a_45663_n11370# a_45613_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X527 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X528 a_48660_n10732# a_47894_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X529 a_3264_n10732# a_4534_n11559# a_4725_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X530 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X531 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X532 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X533 a_19823_n10487# a_19850_n11298# a_19835_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X534 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X535 a_639_690# C[96] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X536 a_46168_n5789# C[56] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X537 a_16245_5953# a_15627_6408# a_15845_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X538 a_48963_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X539 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X540 VSS a_26955_6408# a_26903_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X541 a_59988_n10732# a_59222_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X542 a_46249_n10487# a_46276_n11298# a_46261_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X543 a_29772_n5622# a_29774_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X544 VSS C[87] a_15856_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X545 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X546 a_48433_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X547 a_9780_696# a_9610_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X548 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X549 a_46305_n6843# a_46218_n6611# a_46223_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X550 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X551 a_53584_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X552 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X553 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X554 a_21331_n5795# a_21161_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X555 a_60291_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X556 VSS a_31020_1932# a_32784_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X557 a_59745_773# a_59155_690# a_59649_773# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X558 a_1376_n10732# a_758_n11559# a_976_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X559 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X560 VDD a_15916_1932# a_21538_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X561 a_16917_n6843# a_16558_n6678# a_16556_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X562 VDD a_47551_n11370# a_47501_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X563 a_5152_n10732# a_6422_n11559# a_6613_n10487# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X564 VSS a_45434_6655# a_45384_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X565 a_31433_1829# a_31067_836# a_29447_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X566 a_14578_n5622# a_14310_n5879# a_14139_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X567 a_46394_n5879# a_46168_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X568 VDD a_8914_n5622# a_9839_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X569 VSS a_16460_n5622# a_17385_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X570 a_25685_5953# a_26903_6434# a_27146_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X571 a_6440_1994# a_6353_1896# a_6358_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X572 a_15737_690# C[104] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X573 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_12557_773# a_12193_836# a_12461_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X575 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X576 a_10009_n5795# a_9839_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X577 a_28245_n6843# a_27886_n6678# a_27884_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X578 VSS C[25] a_11857_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X579 VDD a_10573_773# a_11498_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X580 a_53946_n5879# a_53720_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X581 a_33039_n10487# a_33066_n11298# a_33051_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X582 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X583 VSS a_24012_n5622# a_24937_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X584 a_12788_n6678# a_12422_n5879# a_10802_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X585 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X586 a_3119_1829# a_2753_836# a_1133_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X587 a_42395_836# a_42169_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X588 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X589 a_3264_n10732# a_2646_n11559# a_2864_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X590 VDD a_49439_n11370# a_49389_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X591 VSS a_1472_n10732# a_1474_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X592 a_18348_n5622# a_19968_n5879# a_19792_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X593 a_35797_n6843# a_35438_n6678# a_35436_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X594 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X595 VDD a_46118_1932# a_52554_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X596 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X597 a_4644_n5789# C[34] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X598 a_26084_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X599 a_20334_n6678# a_19742_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X600 a_59236_5708# a_59263_6449# a_59248_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X601 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X602 VDD a_25632_n5879# a_25456_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X603 VSS a_35340_n5622# a_36265_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X604 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X605 a_1229_773# a_1231_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X606 OUT a_60574_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X607 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X608 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X609 a_36999_773# a_38619_836# a_38443_1896# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X610 a_35207_773# a_34843_836# a_35111_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X611 a_33237_5953# a_32619_6408# a_32837_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X612 a_453_n11561# a_865_836# a_689_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X613 VSS a_42892_n5622# a_43817_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X614 a_44551_773# a_45939_690# a_45989_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X615 VSS a_43947_6408# a_43895_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X616 a_59649_773# a_59381_836# a_59210_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X617 a_5152_n10732# a_4534_n11559# a_4752_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X618 a_21993_1829# a_21627_836# a_20007_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X619 VSS a_30960_n11559# a_30908_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X620 VSS a_3360_n10732# a_3362_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X621 a_55460_5708# a_55487_6449# a_55472_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X622 a_4870_n5879# a_4644_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X623 VDD a_44512_n5879# a_44336_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X624 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X625 a_2608_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X626 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X627 a_12060_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X628 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X629 a_12571_5953# a_11857_6408# a_12475_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X630 a_3021_773# a_4415_690# a_4465_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X631 VDD a_16145_n6869# a_24469_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X632 a_53775_n6843# a_53770_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X633 a_28448_6655# a_27573_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X634 a_2251_n11370# a_1376_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X635 a_7040_n10732# a_6422_n11559# a_6640_n11298# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X636 a_42677_5953# a_43895_6434# a_44138_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X637 a_1474_n11788# a_1472_n10732# a_1775_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X638 a_56762_6655# a_55887_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X639 a_27657_1829# a_27065_690# a_25671_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X640 VDD a_26955_6408# a_27173_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X641 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X642 VDD a_16145_n6869# a_30133_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X643 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X644 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X645 a_59292_1994# a_59205_1896# a_59210_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X646 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X647 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X648 a_51327_n11370# a_50452_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X649 a_27671_7009# a_27669_5953# a_27972_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X650 a_23797_5953# a_23179_6408# a_23397_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X651 VDD a_25403_836# a_25227_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X652 a_14674_n5622# a_14310_n5879# a_14578_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X653 a_43076_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X654 a_25769_1829# a_25177_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X655 a_24425_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X656 a_38448_1994# a_38443_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X657 VSS a_31249_n6869# a_31125_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X658 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X659 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X660 VDD a_818_1932# a_11030_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X661 VSS a_22005_5953# a_22007_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X662 a_22124_n5622# a_21856_n5879# a_21685_n6843# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X663 a_3362_n11788# a_3360_n10732# a_3663_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X664 a_44057_690# C[119] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X665 VDD a_31564_n5622# a_32489_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X666 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X667 a_26789_n11370# a_25914_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X668 a_14806_1994# a_14447_1829# a_14445_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X669 a_32659_n5795# a_32489_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X670 a_33335_7009# a_32619_6408# a_31349_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X671 a_27291_836# a_27065_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X672 VDD a_30731_6408# a_30679_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X673 VSS a_52986_6655# a_52936_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X674 a_27573_5953# a_26903_6434# a_27173_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X675 a_33550_n6678# a_32958_n5789# a_31564_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X676 a_20334_n6678# a_19968_n5879# a_18348_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X677 a_53215_n11370# a_52340_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X678 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X679 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X680 VDD a_48053_836# a_47877_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X681 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X682 VSS a_1047_n6869# a_12786_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X683 a_26313_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X684 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X685 a_50305_773# a_50307_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X686 a_43004_n11788# a_42288_n11559# a_41018_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X687 VSS a_41114_n10732# a_41116_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X688 VSS a_47717_6408# a_47665_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X689 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X690 VDD a_17515_6408# a_17733_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X691 VSS a_44551_773# a_45476_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X692 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X693 VDD a_49941_836# a_49765_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X694 a_28677_n11370# a_27802_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X695 a_50895_n6843# a_50536_n6678# a_50534_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X696 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X697 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X698 a_24110_n6678# a_23518_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X699 VDD a_29408_n5879# a_29232_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X700 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 a_18231_7009# a_18229_5953# a_18532_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X702 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X703 a_44649_1829# a_44057_690# a_42663_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X704 VSS a_50438_n5622# a_51363_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X705 VDD a_43947_6408# a_44165_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X706 a_40510_n5789# C[53] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X707 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X708 VSS a_818_1932# a_12557_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X709 a_40005_n11370# a_39130_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X710 a_28201_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X711 VDD a_36960_n5879# a_36784_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X712 a_16341_5953# a_15627_6408# a_16245_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X713 VDD a_46347_n6869# a_46305_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X714 VSS a_43002_n10732# a_43004_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X715 a_12571_5953# a_11805_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X716 a_44663_7009# a_44661_5953# a_44964_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X717 a_39982_696# a_39812_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X718 a_46447_5953# a_47665_6434# a_47908_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X719 a_40789_5953# a_40171_6408# a_40389_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X720 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X721 a_52097_773# a_53491_690# a_53541_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X722 VSS a_21520_n11559# a_21468_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X723 a_23895_7009# a_23179_6408# a_21909_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X724 VDD a_16145_n6869# a_16917_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 VDD a_46347_n6869# a_53857_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X726 a_38393_690# C[116] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X727 a_16556_n5622# a_15966_n5789# a_16460_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X728 a_55460_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X729 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X730 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X731 a_27655_773# a_27291_836# a_27559_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X732 VDD a_9574_6655# a_9524_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X733 a_38622_n5789# C[52] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X734 a_57493_836# a_57267_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X735 a_34927_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X736 a_694_1994# a_689_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X737 VSS a_818_1932# a_12022_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X738 a_11897_n5795# a_11727_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X739 VSS a_16145_n6869# a_16021_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X740 VSS a_44890_n10732# a_44892_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X741 a_41116_n11788# a_41114_n10732# a_41417_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X742 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X743 a_363_n11370# a_453_n11561# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X744 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X745 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X746 VDD a_47946_n11559# a_47894_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X747 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X748 a_52195_1829# a_51603_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X749 a_224_6410# a_529_6408# a_720_5708# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X750 VSS a_11462_6655# a_11412_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X751 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X752 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X753 a_57761_773# a_59381_836# a_59205_1896# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X754 VDD a_16460_n5622# a_17385_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X755 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X756 VDD a_31249_n6869# a_35797_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X757 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X758 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X759 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X760 a_18576_1994# a_18217_1829# a_18215_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X761 a_35436_n5622# a_34846_n5789# a_35340_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X762 VDD a_34507_6408# a_34725_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X763 a_10685_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X764 a_37109_5953# a_36395_6408# a_37013_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X765 a_19008_6655# a_18133_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X766 a_24878_696# a_24708_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X767 VDD a_24012_n5622# a_24937_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X768 a_5322_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X769 a_41100_n5622# a_40510_n5789# a_41004_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X770 a_42988_n5622# a_42398_n5789# a_42892_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X771 a_36815_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X772 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X773 VSS a_31249_n6869# a_34901_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X774 a_43004_n11788# a_43002_n10732# a_43305_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X775 a_35223_7009# a_35221_5953# a_35524_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X776 VSS a_31249_n6869# a_36789_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X777 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X778 a_10669_773# a_10079_690# a_10573_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X779 VDD a_49834_n11559# a_49782_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X780 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X781 a_31676_n11788# a_30960_n11559# a_29690_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X782 VSS C[19] a_23179_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X783 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X784 VDD a_35340_n5622# a_36265_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X785 a_19742_n5789# C[42] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X786 VSS a_31249_n6869# a_42453_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X787 a_33333_5953# a_32619_6408# a_33237_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X788 a_46020_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X789 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X790 a_33452_n5622# a_33184_n5879# a_33013_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X791 a_17349_n11370# a_16474_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X792 a_1546_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X793 a_20236_n5622# a_19742_n5789# a_19797_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X794 a_9327_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X795 a_48419_1829# a_47827_690# a_46433_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X796 VDD a_42892_n5622# a_43817_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X797 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X798 a_27559_773# a_27065_690# a_27120_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X799 a_47528_696# a_47358_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X800 a_25406_n5789# C[45] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X801 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X802 a_40887_7009# a_40171_6408# a_38901_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X803 a_18217_1829# a_17625_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X804 a_11691_n11370# a_10816_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X805 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X806 a_38703_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X807 VSS a_15916_1932# a_16327_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X808 VSS a_2646_n11559# a_2594_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X809 a_44892_n11788# a_44890_n10732# a_45193_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X810 a_10573_773# a_11967_690# a_12017_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X811 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X812 VSS a_31674_n10732# a_31676_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X813 a_33564_n11788# a_32848_n11559# a_31578_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X814 a_7686_6655# a_6811_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X815 a_16341_5953# a_15575_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X817 a_18080_n5879# a_17854_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X818 VSS a_1047_n6869# a_9010_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X819 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X820 a_38997_5953# a_38231_6434# a_38901_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X821 a_19968_n5879# a_19742_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X822 a_19237_n11370# a_18362_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X823 a_6895_1829# a_6303_690# a_4909_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X824 VSS a_41893_n11370# a_41843_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X825 a_54326_n11788# a_53558_n11533# a_52340_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X826 a_1243_5953# a_477_6434# a_1147_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X827 a_25632_n5879# a_25406_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X828 a_44286_n5789# C[55] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X829 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X830 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X831 a_18231_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X832 a_35568_1994# a_35209_1829# a_35207_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X833 VSS a_4534_n11559# a_4482_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X834 a_51098_6655# a_50223_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X835 VDD a_50170_n5879# a_49994_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X836 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X837 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X838 a_38901_5953# a_40171_6408# a_40362_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X839 a_6909_7009# a_6907_5953# a_7210_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X840 a_23382_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X841 a_59155_690# C[127] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X842 a_10573_773# a_10305_836# a_10134_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X843 a_44423_n6843# a_44336_n6611# a_44341_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X844 a_23599_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X845 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X846 a_50307_1829# a_49715_690# a_48321_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X847 a_32955_836# a_32729_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X848 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X849 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X850 VSS a_15232_6655# a_15182_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X851 a_23893_5953# a_23179_6408# a_23797_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X852 a_5019_5953# a_4305_6408# a_4923_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X853 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X854 a_53999_5953# a_55217_6434# a_55460_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X855 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X856 VSS a_43781_n11370# a_43731_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X857 a_56214_n11788# a_55446_n11533# a_54228_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X858 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X859 VSS C[10] a_40171_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X860 a_44512_n5879# a_44286_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X861 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X862 a_15444_696# a_15274_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X863 VSS a_14578_n5622# a_15503_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X864 a_53720_n5789# C[60] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X865 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X866 VSS a_6422_n11559# a_6370_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X867 a_6811_5953# a_6141_6434# a_6411_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X868 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X869 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X870 a_31676_n11788# a_31674_n10732# a_31977_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X871 a_31674_n10732# a_30960_n11559# a_31578_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X872 a_25487_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X873 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X874 a_54398_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X875 a_49770_1994# a_49765_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X876 a_20348_n11788# a_19632_n11559# a_18362_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X877 VDD a_15916_1932# a_22352_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X878 VSS a_31020_1932# a_33319_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X879 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X880 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X881 VDD a_46347_n6869# a_50895_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X882 a_58102_n11788# a_57334_n11533# a_56116_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X883 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X884 a_50534_n5622# a_49944_n5789# a_50438_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X885 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X886 VDD a_865_836# a_689_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X887 a_25461_n6843# a_25456_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X888 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X889 a_38094_696# a_37924_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X890 VSS a_8310_n11559# a_8258_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X891 a_7254_1994# a_6895_1829# a_6893_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X892 a_53985_773# a_53491_690# a_53546_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X893 a_33548_n5622# a_33184_n5879# a_33452_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X894 VSS a_59759_5953# a_59761_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X895 a_14349_773# a_15737_690# a_15787_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X896 a_27375_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X897 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X898 a_54214_n5622# a_55608_n5789# a_55658_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X899 VSS a_46347_n6869# a_49999_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X900 VSS a_13745_6408# a_13693_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X901 a_31125_n6843# a_31120_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X902 a_56102_n5622# a_57496_n5789# a_57546_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X903 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X904 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X905 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X906 a_54095_5953# a_53329_6434# a_53999_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X907 a_35223_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X908 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X909 a_22236_n11788# a_21520_n11559# a_20250_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X910 a_25258_5708# a_25285_6449# a_25270_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X911 VDD a_50438_n5622# a_51363_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X912 a_11967_690# C[102] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X913 VSS a_16145_n6869# a_20332_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X914 VDD a_25296_n11559# a_25244_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X915 a_54324_n10732# a_53558_n11533# a_54228_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X916 a_40374_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X917 VSS a_30565_n11370# a_30515_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X918 VSS a_32224_6655# a_32174_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X919 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X920 VSS a_42288_n11559# a_42236_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X921 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X922 a_41018_n10732# a_42236_n11533# a_42479_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X923 a_55971_1829# a_55379_690# a_53985_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X924 VDD a_25671_773# a_26596_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X925 VDD a_55269_6408# a_55487_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X926 a_31447_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X927 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X928 VSS a_10573_773# a_11498_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X929 VDD a_15963_836# a_15787_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 a_12786_n5622# a_12788_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X931 a_29263_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X932 a_12475_5953# a_13693_6434# a_13936_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X933 a_29319_n6843# a_29232_n6611# a_29237_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X934 a_26560_6655# a_25685_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X935 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X936 VDD a_51829_836# a_51653_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X937 a_24124_n11788# a_23408_n11559# a_22138_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X938 VDD C[77] a_34736_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X939 VSS a_818_1932# a_5005_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X940 a_29090_1994# a_29003_1896# a_29008_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X941 VDD a_27184_n11559# a_27132_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X942 a_56212_n10732# a_55446_n11533# a_56116_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X943 VDD C[23] a_15627_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X944 a_34617_690# C[114] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X945 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X946 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X947 a_55985_7009# a_55983_5953# a_56286_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X948 a_5234_n5622# a_5236_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X949 a_5019_5953# a_4253_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X950 VSS a_32453_n11370# a_32403_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X951 a_17851_836# a_17625_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X952 a_11897_n5795# a_11727_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X953 VSS a_44176_n11559# a_44124_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X954 a_42906_n10732# a_44124_n11533# a_44367_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X955 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X956 VSS a_50319_5953# a_50321_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X957 a_53717_836# a_53491_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X958 a_12788_n6678# a_12196_n5789# a_10802_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X959 VDD a_48321_773# a_49246_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X960 a_25767_773# a_25177_690# a_25671_773# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X961 a_41870_696# a_41700_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X962 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X963 a_22581_n6843# a_22222_n6678# a_22220_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X964 a_20346_n10732# a_19632_n11559# a_20250_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X965 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X966 a_15818_5708# a_15845_6449# a_15830_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X967 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X968 VDD C[76] a_36624_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X969 VSS a_6411_6449# a_6384_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X970 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X971 a_40281_690# C[117] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X972 VDD C[85] a_19632_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X973 VDD a_29072_n11559# a_29020_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X974 a_58100_n10732# a_57334_n11533# a_58004_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X975 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X976 VSS a_22124_n5622# a_23049_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X977 VSS a_22784_6655# a_22734_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X978 VSS a_34341_n11370# a_34291_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X979 a_40603_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X980 a_42250_5708# a_42277_6449# a_42262_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X981 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X982 a_59381_836# a_59155_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X983 a_57496_n5789# C[62] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X984 a_59610_n5879# a_59384_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X985 VDD a_16145_n6869# a_17991_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X986 a_6909_7009# a_6141_6434# a_4923_5953# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X987 VSS a_29676_n5622# a_30601_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X988 VDD a_16145_n6869# a_19879_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X989 a_59759_5953# a_58993_6434# a_59649_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X990 a_5007_1829# a_4415_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X991 a_3362_n11788# a_2646_n11559# a_1376_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X992 a_20103_773# a_20105_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X993 VSS a_17515_6408# a_17463_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X994 VDD C[12] a_36395_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X995 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X996 a_38983_773# a_38985_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X997 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X998 a_41461_n6843# a_41102_n6678# a_41100_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X999 a_22234_n10732# a_21520_n11559# a_22138_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1000 a_16047_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1001 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1002 VDD a_16145_n6869# a_25543_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1003 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1004 VDD C[84] a_21520_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1005 a_46545_7009# a_46543_5953# a_46846_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1006 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1007 a_5138_n5622# a_6758_n5879# a_6582_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1008 a_7026_n5622# a_8646_n5879# a_8470_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1009 VSS a_36229_n11370# a_36179_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1010 a_43552_6655# a_42677_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1011 a_14447_1829# a_13855_690# a_12461_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1012 a_52193_773# a_51829_836# a_52097_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1013 a_42491_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1014 VDD a_13745_6408# a_13963_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1015 a_42906_n10732# a_42236_n11533# a_42506_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1016 VSS a_747_6449# a_720_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1017 a_7124_n6678# a_6532_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1018 VDD C[14] a_32619_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1019 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1020 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1021 a_57722_n5879# a_57496_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1022 VDD a_31249_n6869# a_38759_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1023 a_25671_773# a_25403_836# a_25232_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1024 a_29690_n10732# a_30908_n11533# a_31151_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1025 a_5250_n11788# a_4534_n11559# a_3264_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1026 VSS a_20346_n10732# a_20348_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1027 VSS a_46118_1932# a_57857_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1028 a_224_6410# a_868_n5789# a_918_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1029 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1030 a_15874_1994# a_15787_1896# a_15792_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1031 a_48053_836# a_47827_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1032 VSS a_48164_n11298# a_48137_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1033 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1034 a_16245_5953# a_17463_6434# a_17706_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1035 a_57871_5953# a_57105_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1036 a_10587_5953# a_9969_6408# a_10187_6449# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1037 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1038 VDD a_31249_n6869# a_44423_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1039 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1040 a_21895_773# a_23289_690# a_23339_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1041 VDD C[83] a_23408_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1042 a_2620_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1043 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 VDD a_1047_n6869# a_13147_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1045 a_32810_5708# a_32837_6449# a_32822_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1046 a_20105_1829# a_19513_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1047 a_14674_n5622# a_14084_n5789# a_14578_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1048 a_44794_n10732# a_44124_n11533# a_44394_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1049 VSS a_38283_6408# a_38231_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1050 VSS a_21125_n11370# a_21075_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1051 a_1472_n10732# a_758_n11559# a_1376_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1052 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1053 a_31578_n10732# a_32796_n11533# a_33039_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 a_7138_n11788# a_6422_n11559# a_5152_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1055 a_29543_773# a_29545_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1056 a_14363_5953# a_13693_6434# a_13963_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1057 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1058 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1059 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1060 VSS a_1047_n6869# a_14139_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1061 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1062 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1063 a_27559_773# a_29179_836# a_29003_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1064 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1065 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1066 a_17947_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1067 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1068 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1069 VDD a_14578_n5622# a_15503_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1070 VDD C[90] a_10198_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1071 VSS a_34507_6408# a_34455_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1072 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1073 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1074 a_52097_773# a_51603_690# a_51658_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1075 a_20334_n6678# a_19742_n5789# a_18348_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1076 a_55985_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1077 a_12690_n5622# a_12422_n5879# a_12251_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1078 VSS a_23013_n11370# a_22963_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1079 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1080 a_3360_n10732# a_2646_n11559# a_3264_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1081 a_57633_n6843# a_57546_n6611# a_57551_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1082 VDD C[29] a_4305_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1083 a_33466_n10732# a_34684_n11533# a_34927_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1084 a_9026_n11788# a_8310_n11559# a_7040_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1085 a_20348_n11788# a_20346_n10732# a_20649_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1086 VSS C[4] a_51493_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1087 a_48137_n10487# a_48164_n11298# a_48149_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1088 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1089 a_10079_690# C[101] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1090 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1091 a_52058_n5879# a_51832_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1092 a_26357_n6843# a_25998_n6678# a_25996_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1093 a_36229_n11370# a_35354_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1094 a_39982_696# a_39812_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1095 a_54228_n10732# a_55498_n11559# a_55689_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1096 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1097 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1098 VDD a_15916_1932# a_17762_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 a_9012_n6678# a_8420_n5789# a_7026_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1100 a_19835_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1101 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1102 a_32866_1994# a_32779_1896# a_32784_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1103 a_29179_836# a_28953_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1104 VDD a_16192_n5879# a_16016_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1105 VDD C[89] a_12086_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1106 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1107 a_33909_n6843# a_33550_n6678# a_33548_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1108 a_33237_5953# a_34455_6434# a_34698_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1109 a_4496_5708# a_4523_6449# a_4508_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1110 a_18217_1829# a_17625_690# a_16231_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1111 a_47322_6655# a_46447_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1112 a_38887_773# a_40281_690# a_40331_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1113 a_59761_7009# a_58993_6434# a_57775_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1114 a_10685_7009# a_9969_6408# a_8699_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1115 a_2756_n5789# C[33] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1116 a_3250_n5622# a_2756_n5789# a_2811_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1117 a_31578_n10732# a_30908_n11533# a_31178_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1118 a_31163_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1119 a_5248_n10732# a_4534_n11559# a_5152_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1120 VDD a_23744_n5879# a_23568_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1121 VSS a_33452_n5622# a_34377_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1122 a_35354_n10732# a_36572_n11533# a_36815_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1123 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1124 a_42250_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1125 a_8420_n5789# C[36] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1126 a_18362_n10732# a_19580_n11533# a_19823_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1127 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1128 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1129 a_8417_836# a_8191_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1130 VDD a_46118_1932# a_60106_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1131 a_45237_n6843# a_44878_n6678# a_44876_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1132 a_38117_n11370# a_37242_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1133 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1134 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1135 VSS a_14459_5953# a_14461_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1136 a_33321_1829# a_32955_836# a_31335_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1137 a_18119_773# a_19739_836# a_19563_1896# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1138 VDD a_2753_836# a_2577_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1139 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 a_49715_690# C[122] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1141 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1142 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1143 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1144 VDD C[88] a_13974_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1145 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1146 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1147 a_1094_n5879# a_868_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1148 a_51696_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1149 a_2982_n5879# a_2756_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1150 a_33466_n10732# a_32796_n11533# a_33066_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1151 a_33051_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1152 a_7136_n10732# a_6422_n11559# a_7040_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1153 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1154 VDD a_42624_n5879# a_42448_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1155 a_4641_836# a_4415_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1156 VDD C[92] a_6422_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1157 VDD a_46347_n6869# a_51969_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1158 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1159 VDD a_31020_1932# a_38530_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1160 a_18133_5953# a_17463_6434# a_17733_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1161 VSS a_49823_6449# a_49796_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1162 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1163 a_20250_n10732# a_21468_n11533# a_21711_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1164 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1165 a_54228_n10732# a_53610_n11559# a_53828_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1166 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1167 a_20105_1829# a_19513_690# a_18119_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1168 VDD a_16145_n6869# a_22581_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1169 a_51887_n6843# a_51882_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1170 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1171 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1172 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1173 a_4552_1994# a_4465_1896# a_4470_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1174 a_23797_5953# a_25015_6434# a_25258_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1175 VDD C[1] a_57157_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1176 VSS a_5248_n10732# a_5250_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1177 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1178 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X1179 VSS C[26] a_9969_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1180 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 a_23515_836# a_23289_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1182 a_35354_n10732# a_34684_n11533# a_34954_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1183 a_9024_n10732# a_8310_n11559# a_8928_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1184 a_32810_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1185 a_35125_5953# a_34507_6408# a_34725_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1186 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1187 VDD C[91] a_8310_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1188 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1189 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1190 a_46433_773# a_47827_690# a_47877_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1191 a_22138_n10732# a_23356_n11533# a_23599_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1192 a_12786_n5622# a_12422_n5879# a_12690_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1193 VDD a_22124_n5622# a_23049_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1194 a_56116_n10732# a_55498_n11559# a_55716_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1195 a_24196_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1196 VSS a_54324_n10732# a_54326_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1197 a_19568_1994# a_19563_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1198 VDD a_31249_n6869# a_41461_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1199 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1200 VSS a_6027_n11370# a_5977_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1201 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1202 a_20236_n5622# a_19968_n5879# a_19797_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1203 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1204 VSS a_7136_n10732# a_7138_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1205 a_35111_773# a_36731_836# a_36555_1896# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1206 a_16327_773# a_15963_836# a_16231_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1207 VDD a_29676_n5622# a_30601_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1208 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1209 a_31349_5953# a_30731_6408# a_30949_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1210 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1211 VDD a_50209_773# a_51134_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1212 a_20250_n10732# a_19580_n11533# a_19850_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1213 a_38985_1829# a_38619_836# a_36999_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1214 a_31662_n6678# a_31070_n5789# a_29676_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1215 a_53572_5708# a_53599_6449# a_53584_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1216 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1217 a_1231_1829# a_865_836# a_453_n11561# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1218 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1219 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1220 VSS a_59045_6408# a_58993_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1221 a_5005_773# a_4641_836# a_4909_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1222 a_10912_n10732# a_10146_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1223 VSS a_56212_n10732# a_56214_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1224 VSS a_1047_n6869# a_10898_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1225 a_10172_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1226 a_5250_n11788# a_5248_n10732# a_5551_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1227 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1228 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X1229 a_10683_5953# a_9969_6408# a_10587_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1230 a_1133_773# a_2527_690# a_2577_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1231 a_31070_n5789# C[48] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1232 VSS a_1047_n6869# a_3346_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1233 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1234 a_15444_696# a_15274_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1235 a_44649_1829# a_44057_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1236 a_22138_n10732# a_21468_n11533# a_21738_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1237 a_40789_5953# a_42007_6434# a_42250_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1238 a_25769_1829# a_25177_690# a_23783_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1239 a_50305_773# a_49715_690# a_50209_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1240 VDD a_27520_n5879# a_27344_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1241 VDD a_25067_6408# a_25285_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1242 a_54874_6655# a_53999_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1243 a_55103_n11370# a_54228_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1244 a_57404_1994# a_57317_1896# a_57322_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1245 VSS a_58100_n10732# a_58102_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1246 a_54326_n11788# a_54324_n10732# a_54627_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1247 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1248 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1249 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1250 a_60335_n6843# a_59976_n6678# a_59974_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1251 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1252 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 VDD a_16231_773# a_17156_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1254 a_7138_n11788# a_7136_n10732# a_7439_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1255 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1256 a_21909_5953# a_21291_6408# a_21509_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1257 a_25783_7009# a_25781_5953# a_26084_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1258 a_41188_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1259 a_6797_773# a_8417_836# a_8241_1896# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1260 a_3035_5953# a_2417_6408# a_2635_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1261 a_36560_1994# a_36555_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1262 a_29182_n5789# C[47] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1263 a_24026_n10732# a_23356_n11533# a_23626_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1264 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1265 VSS a_20117_5953# a_20119_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1266 VSS a_38997_5953# a_38999_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1267 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1268 a_38094_696# a_37924_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1269 a_25177_690# C[109] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1270 a_49941_836# a_49715_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1271 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1272 a_56991_n11370# a_56116_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1273 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1274 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 a_4909_773# a_4415_690# a_4470_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1276 a_56214_n11788# a_56212_n10732# a_56515_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1277 a_50025_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1278 a_31447_7009# a_30731_6408# a_29461_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1279 a_12918_1994# a_12559_1829# a_12557_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1280 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1281 a_50209_773# a_51829_836# a_51653_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1282 a_8246_1994# a_8241_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1283 VSS a_46118_1932# a_55434_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1284 a_16327_773# a_15737_690# a_16231_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1285 a_32430_696# a_32260_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1286 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1287 a_54083_1829# a_53717_836# a_52097_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1288 a_5152_n10732# a_6370_n11533# a_6613_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1289 VSS a_14192_n11298# a_14165_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1290 a_12048_5708# a_12075_6449# a_12060_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1291 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1292 a_33548_n5622# a_32958_n5789# a_33452_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1293 a_20332_n5622# a_19968_n5879# a_20236_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1294 VSS a_45829_6408# a_45777_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1295 a_50209_773# a_49941_836# a_49770_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1296 a_29557_5953# a_28791_6434# a_29461_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1297 VSS a_25671_773# a_26596_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1298 a_6233_n5795# a_6063_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1299 a_54214_n5622# a_55834_n5879# a_55658_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1300 a_24901_n11370# a_24026_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1301 a_58102_n11788# a_58100_n10732# a_58403_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1302 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1303 VSS a_31249_n6869# a_33013_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1304 a_37228_n5622# a_38622_n5789# a_38672_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1305 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1306 a_42761_1829# a_42169_690# a_40775_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1307 a_46774_n11788# a_46058_n11559# a_44794_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1308 VDD a_42059_6408# a_42277_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1309 a_16343_7009# a_16341_5953# a_16644_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1310 VDD a_46118_1932# a_59292_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1311 a_29461_5953# a_30731_6408# a_30922_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1312 a_20119_7009# a_19351_6434# a_18133_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1313 a_15963_836# a_15737_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1314 a_55080_696# a_54910_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1315 VDD a_33452_n5622# a_34377_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1316 a_13350_6655# a_12475_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1317 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1318 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1319 a_17854_n5789# C[41] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1320 a_42775_7009# a_42773_5953# a_43076_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1321 a_44565_5953# a_45777_6434# a_46020_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1322 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1323 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1324 a_10914_n11788# a_10146_n11533# a_8928_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1325 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1326 VSS a_15916_1932# a_27655_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1327 VSS a_48321_773# a_49246_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1328 a_23518_n5789# C[44] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1329 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1330 a_22007_7009# a_21291_6408# a_20021_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1331 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1332 a_56968_696# a_56798_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1333 a_16103_n6843# a_16016_n6611# a_16021_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1334 a_17991_n6843# a_17904_n6611# a_17909_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1335 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1336 a_19513_690# C[106] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1337 a_41870_696# a_41700_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1338 a_53572_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1339 a_55379_690# C[125] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1340 VSS a_46772_n10732# a_46774_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1341 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1342 VDD a_7686_6655# a_7636_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1343 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1344 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1345 VDD a_818_1932# a_14806_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1346 a_16231_773# a_15963_836# a_15792_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1347 VDD a_40005_n11370# a_39955_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1348 a_5152_n10732# a_4482_n11533# a_4752_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1349 a_16192_n5879# a_15966_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1350 a_14165_n10487# a_14192_n11298# a_14177_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1351 a_36734_n5789# C[51] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1352 VSS a_1047_n6869# a_7122_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1353 VSS a_56991_n11370# a_56941_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1354 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1355 VSS a_29061_6449# a_29034_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1356 a_12802_n11788# a_12034_n11533# a_10816_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1357 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1358 a_42398_n5789# C[54] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1359 a_55873_773# a_57493_836# a_57317_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1360 a_23744_n5879# a_23518_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1361 a_36871_n6843# a_36784_n6611# a_36789_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1362 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1363 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1364 a_44551_773# a_44057_690# a_44112_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1365 a_16688_1994# a_16329_1829# a_16327_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1366 a_51603_690# C[123] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1367 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1368 VDD a_32619_6408# a_32837_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1369 VDD a_46118_1932# a_49852_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1370 VSS a_48660_n10732# a_48662_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1371 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 a_20021_5953# a_21291_6408# a_21482_5708# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1373 a_59747_1829# a_59381_836# a_57761_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1374 a_7040_n10732# a_6370_n11533# a_6640_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1375 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1376 a_35072_n5879# a_34846_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1377 a_25783_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1378 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1379 a_36960_n5879# a_36734_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1380 VSS a_58879_n11370# a_58829_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1381 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1382 a_19739_836# a_19513_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1383 a_33335_7009# a_33333_5953# a_33636_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1384 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1385 a_3117_773# a_2753_836# a_3021_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1386 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1387 a_14690_n11788# a_13922_n11533# a_12704_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1388 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1389 VSS C[20] a_21291_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1390 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1391 a_42624_n5879# a_42398_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1392 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1393 VSS a_12690_n5622# a_13615_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1394 a_46774_n11788# a_46772_n10732# a_47075_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1395 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1396 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1397 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1398 VSS a_31020_1932# a_44647_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1399 a_46531_1829# a_45939_690# a_44551_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1400 VDD a_3021_773# a_3946_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1401 a_56200_n6678# a_55834_n5879# a_54214_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1402 VDD a_45829_6408# a_46047_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1403 VDD a_51098_6655# a_51048_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1404 VDD a_42395_836# a_42219_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1405 a_9371_n6843# a_9012_n6678# a_9010_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1406 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1407 a_42761_1829# a_42169_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1408 a_17120_6655# a_16245_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1409 a_8685_773# a_10079_690# a_10129_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1410 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1411 a_10912_n10732# a_10146_n11533# a_10816_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1412 a_224_6410# a_1094_n5879# a_918_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1413 VDD a_53381_6408# a_53329_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1414 VSS a_55498_n11559# a_55446_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1415 a_5798_6655# a_4923_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1416 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1417 a_23573_n6843# a_23568_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1418 a_46662_n5622# a_48056_n5789# a_48106_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1419 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1420 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1421 a_44283_836# a_44057_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1422 a_15461_n11370# a_14592_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1423 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1424 a_5007_1829# a_4415_690# a_3021_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1425 a_48662_n11788# a_48660_n10732# a_48963_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1426 VDD a_4305_6408# a_4523_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1427 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1428 a_52326_n5622# a_53720_n5789# a_53770_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1429 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1430 VDD a_15916_1932# a_18576_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1431 VDD a_14081_836# a_13905_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1432 a_9803_n11370# a_8928_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1433 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1434 a_5021_7009# a_5019_5953# a_5322_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1435 a_21494_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1436 a_12800_n10732# a_12034_n11533# a_12704_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1437 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1438 VSS a_45663_n11370# a_45613_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1439 VDD C[64] a_59274_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1440 VSS a_57386_n11559# a_57334_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1441 a_51925_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1442 a_56116_n10732# a_57334_n11533# a_57577_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1443 a_16572_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1444 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1445 a_42775_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1446 a_42453_n6843# a_42448_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1447 a_3131_5953# a_2417_6408# a_3035_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1448 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1449 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1450 a_52111_5953# a_53329_6434# a_53572_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1451 a_58879_n11370# a_58004_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1452 VSS C[95] a_758_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1453 a_10898_n5622# a_10900_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1454 VDD C[17] a_26955_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1455 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1456 a_3117_773# a_2527_690# a_3021_773# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1457 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1458 a_51832_n5789# C[59] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1459 a_3346_n5622# a_3348_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1460 VSS a_47551_n11370# a_47501_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1461 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1463 VSS a_59274_n11559# a_59222_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1464 a_53813_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1465 a_16231_773# a_17625_690# a_17675_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1466 a_47882_1994# a_47877_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1467 a_58004_n10732# a_59222_n11533# a_59465_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1468 a_34112_6655# a_33237_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1469 VSS a_31020_1932# a_31431_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1470 VDD a_31020_1932# a_39344_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1471 a_50081_n6843# a_49994_n6611# a_49999_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1472 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1473 a_10900_n6678# a_10308_n5789# a_8914_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1474 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1475 a_8795_5953# a_8029_6434# a_8699_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1476 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1477 VSS C[94] a_2646_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1478 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1479 VDD a_42663_773# a_43588_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1480 a_44647_773# a_44283_836# a_44551_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1481 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1482 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1483 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1484 a_20693_n6843# a_20334_n6678# a_20332_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1485 a_19214_696# a_19044_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1486 VDD a_38512_n11559# a_38730_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1487 a_5366_1994# a_5007_1829# a_5005_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1488 a_6233_n5795# a_6063_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1489 a_48056_n5789# C[57] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1490 a_50170_n5879# a_49944_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1491 VSS a_11857_6408# a_11805_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1492 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1493 VSS a_20236_n5622# a_21161_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1494 a_49944_n5789# C[58] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1495 VSS a_49439_n11370# a_49389_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1496 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1497 a_7124_n6678# a_6532_n5789# a_5138_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1498 VSS C[68] a_51722_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1499 a_55701_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1500 a_52207_5953# a_51441_6434# a_52111_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1501 a_33335_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1502 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1503 a_23370_5708# a_23397_6449# a_23382_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1504 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1505 a_7892_696# a_7722_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1506 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1507 a_55608_n5789# C[61] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1508 VDD a_16145_n6869# a_16103_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1509 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1510 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1511 a_56102_n5622# a_55608_n5789# a_55663_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1512 a_57990_n5622# a_57496_n5789# a_57551_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1513 a_1460_n6678# a_1094_n5879# a_224_6410# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1514 VSS C[93] a_4534_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1515 VDD a_758_n11559# a_976_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1516 VSS a_30336_6655# a_30286_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1517 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 a_6303_690# C[99] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1519 VSS a_36613_6449# a_36586_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1520 VDD a_16145_n6869# a_23655_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1521 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1522 VDD a_53381_6408# a_53599_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1523 a_3021_773# a_2753_836# a_2582_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1524 a_48282_n5879# a_48056_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1525 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1526 a_3250_n5622# a_4870_n5879# a_4694_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1527 a_58004_n10732# a_57334_n11533# a_57604_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1528 a_10587_5953# a_11805_6434# a_12048_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1529 VDD C[8] a_43947_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1530 a_58650_6655# a_57775_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1531 a_52422_n5622# a_51832_n5789# a_52326_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1532 VSS C[67] a_53610_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1533 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1534 a_24672_6655# a_23797_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1535 VSS a_818_1932# a_3117_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1536 a_27202_1994# a_27115_1896# a_27120_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1537 VSS a_46058_n11559# a_46006_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1538 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1539 a_5236_n6678# a_4644_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1540 a_55834_n5879# a_55608_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1541 VDD a_31249_n6869# a_34983_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1542 VDD a_31249_n6869# a_36871_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1543 a_44794_n10732# a_46006_n11533# a_46249_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1544 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1545 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1546 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1547 a_31674_n10732# a_30908_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1548 a_3131_5953# a_2365_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1549 a_33223_773# a_34617_690# a_34667_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1550 a_35209_1829# a_34617_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1551 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1552 VDD a_31249_n6869# a_42535_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1553 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1554 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1555 a_44138_5708# a_44165_6449# a_44150_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1556 a_8928_n10732# a_10198_n11559# a_10389_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1557 a_22990_696# a_22820_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1558 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1559 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1560 VSS a_50209_773# a_51134_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1561 VDD C[69] a_49834_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1562 a_5021_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1563 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1564 a_21401_690# C[107] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1565 a_12786_n5622# a_12196_n5789# a_12690_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1566 VSS C[74] a_40400_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1567 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1568 a_29447_773# a_30841_690# a_30891_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1569 a_46676_n10732# a_47894_n11533# a_48137_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1570 VSS a_20896_6655# a_20846_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1571 a_58218_1994# a_57859_1829# a_57857_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1572 VDD a_57493_836# a_57317_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1573 a_33562_n10732# a_32796_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1574 VSS a_39776_6655# a_39726_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1575 a_57859_1829# a_57267_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1576 a_49439_n11370# a_48564_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1577 VSS a_2022_6655# a_1972_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1578 a_40362_5708# a_40389_6449# a_40374_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1579 VDD a_1047_n6869# a_9371_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1580 VSS a_1047_n6869# a_12251_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1581 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1582 a_57775_5953# a_57105_6434# a_57375_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1583 VDD C[82] a_25296_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1584 a_10816_n10732# a_12086_n11559# a_12277_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1585 a_1245_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1586 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1587 a_37095_773# a_37097_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1588 VDD a_12690_n5622# a_13615_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1589 a_59990_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1590 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1591 VSS a_15627_6408# a_15575_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1592 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1593 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1594 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1595 a_10802_n5622# a_10534_n5879# a_10363_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1596 VSS C[73] a_42288_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1597 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1598 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1599 a_55745_n6843# a_55658_n6611# a_55663_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1600 a_41664_6655# a_40789_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1601 a_12559_1829# a_11967_690# a_10573_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1602 VDD a_11857_6408# a_12075_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1603 VDD a_15916_1932# a_29090_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 VDD a_29179_836# a_29003_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1605 a_44194_1994# a_44107_1896# a_44112_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1606 VSS a_16231_773# a_17156_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1607 a_24469_n6843# a_24110_n6678# a_24108_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1608 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 VDD C[15] a_30731_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1610 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1611 VDD C[81] a_27184_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1612 VDD a_29072_n11559# a_29290_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1613 a_12704_n10732# a_13974_n11559# a_14165_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1614 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1615 VSS a_46118_1932# a_55969_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1616 a_7026_n5622# a_6758_n5879# a_6587_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1617 VSS a_46347_n6869# a_48646_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1618 a_8914_n5622# a_8646_n5879# a_8475_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1619 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1620 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1621 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1622 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1623 a_14084_n5789# C[39] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1624 a_14363_5953# a_15575_6434# a_15818_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1625 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1626 a_14081_836# a_13855_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1627 a_58102_n11788# a_57386_n11559# a_56116_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1628 a_46261_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1629 a_20007_773# a_21401_690# a_21451_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1630 VSS C[72] a_44176_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1631 a_46676_n10732# a_46006_n11533# a_46276_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1632 a_42773_5953# a_42007_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1633 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1634 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1635 a_1362_n5622# a_868_n5789# a_923_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1636 a_23370_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1637 VDD a_21856_n5879# a_21680_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1638 a_14221_n6843# a_14134_n6611# a_14139_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1639 a_30922_5708# a_30949_6449# a_30934_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1640 a_5236_n6678# a_4870_n5879# a_3250_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1641 a_20346_n10732# a_19580_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1642 VSS a_36395_6408# a_36343_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1643 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1644 VSS a_46118_1932# a_52193_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1645 a_43349_n6843# a_42990_n6678# a_42988_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1646 a_37340_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1647 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1648 a_10816_n10732# a_10198_n11559# a_10416_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1649 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1650 a_32430_696# a_32260_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1651 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1652 a_27655_773# a_27657_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1653 a_10671_1829# a_10079_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1654 VDD a_33184_n5879# a_33008_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1655 VSS a_36842_n11298# a_36815_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1656 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1657 a_8781_773# a_8783_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1658 a_14310_n5879# a_14084_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1659 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1660 VSS a_31020_1932# a_42224_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1661 a_48564_n10732# a_47894_n11533# a_48164_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1662 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1663 a_25671_773# a_27291_836# a_27115_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1664 VSS C[80] a_29072_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1665 VSS a_32619_6408# a_32567_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1666 a_59745_773# a_59381_836# a_59649_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1667 VDD a_40736_n5879# a_40560_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1668 VDD a_46347_n6869# a_50081_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1669 VDD a_15916_1932# a_19650_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1670 a_54097_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1671 a_22234_n10732# a_21468_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1672 a_29545_1829# a_29179_836# a_27559_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1673 a_38619_836# a_38393_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1674 a_39228_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1675 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1676 a_12704_n10732# a_12086_n11559# a_12304_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1677 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1678 VDD C[30] a_2417_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1679 VDD a_32955_836# a_32779_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1680 VDD a_16145_n6869# a_20693_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1681 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1682 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1683 a_55080_696# a_54910_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1684 a_363_n11370# a_453_n11561# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1685 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1686 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1687 a_56212_n10732# a_55498_n11559# a_56116_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1688 VSS a_38730_n11298# a_38703_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1689 VSS a_57375_6449# a_57348_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1690 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1691 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1692 a_13910_1994# a_13905_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1693 VDD a_15916_1932# a_15874_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1694 a_56968_696# a_56798_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1695 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1696 a_30978_1994# a_30891_1896# a_30896_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1697 VSS C[79] a_30960_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1698 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1699 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1700 a_34843_836# a_34617_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1701 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1702 VSS a_16145_n6869# a_21685_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1703 a_25900_n5622# a_27294_n5789# a_27344_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1704 a_31349_5953# a_32567_6434# a_32810_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1705 a_2608_5708# a_2635_6449# a_2620_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1706 a_16329_1829# a_15737_690# a_14349_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1707 a_59085_n5795# a_58915_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1708 a_24122_n10732# a_23356_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1709 a_45434_6655# a_44565_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1710 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1711 a_57873_7009# a_57105_6434# a_55887_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1712 VSS a_8081_6408# a_8029_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1713 a_9010_n5622# a_8420_n5789# a_8914_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1714 a_10898_n5622# a_10534_n5879# a_10802_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1715 VDD a_20236_n5622# a_21161_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1716 a_14592_n10732# a_13974_n11559# a_14192_n11298# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1717 VSS a_976_n11298# a_949_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1718 a_42759_773# a_42169_690# a_42663_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1719 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1720 a_40362_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1721 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1722 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1723 VDD C[87] a_15856_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1724 a_36815_n10487# a_36842_n11298# a_36827_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1725 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1726 a_58100_n10732# a_57386_n11559# a_58004_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1727 a_22222_n6678# a_21630_n5789# a_20236_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1728 VSS C[5] a_49605_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1729 VSS a_12571_5953# a_12573_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1730 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1731 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1732 a_44647_773# a_44649_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1733 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1734 a_46543_5953# a_45777_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1735 a_59649_773# a_59155_690# a_59210_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1736 VSS C[78] a_32848_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1737 a_37338_n10732# a_36572_n11533# a_37242_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1738 VSS a_4305_6408# a_4253_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1739 VSS a_31249_n6869# a_40565_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1740 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1741 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1742 a_2527_690# C[97] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1743 a_11691_n11370# a_10816_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1744 a_1775_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1745 a_42663_773# a_44283_836# a_44107_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1746 a_21102_696# a_20932_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1747 VDD a_31020_1932# a_36642_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1748 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1749 a_38703_n10487# a_38730_n11298# a_38715_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1750 VSS a_47935_6449# a_47908_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1751 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1752 VSS a_46118_1932# a_45994_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1753 a_37097_1829# a_36505_690# a_35111_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1754 VSS a_1047_n6869# a_1458_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1755 a_3360_n10732# a_2594_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1756 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1757 a_5138_n5622# a_4644_n5789# a_4699_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1758 a_21909_5953# a_23127_6434# a_23370_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1759 VDD C[2] a_55269_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1760 a_2664_1994# a_2577_1896# a_2582_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1761 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1762 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1763 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1764 VDD a_31020_1932# a_32866_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1765 VSS a_3021_773# a_3946_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1766 a_8783_1829# a_8191_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1767 a_3663_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1768 a_949_n10487# a_976_n11298# a_961_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1769 a_30922_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1770 a_42663_773# a_42395_836# a_42224_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1771 a_27900_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1772 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1773 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1774 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1775 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1776 a_33321_1829# a_32729_690# a_31335_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1777 a_22308_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1778 VSS a_27402_n11298# a_27375_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1779 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1780 a_17680_1994# a_17675_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1781 a_10573_773# a_10079_690# a_10134_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1782 a_27294_n5789# C[46] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1783 a_5248_n10732# a_4482_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1784 VDD a_2251_n11370# a_2201_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1785 a_52739_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1786 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1787 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1788 VDD a_30960_n11559# a_30908_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1789 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1790 VDD a_40171_6408# a_40119_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1791 a_5551_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1792 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1793 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1794 a_39214_n6678# a_38848_n5879# a_37228_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1795 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1796 VDD a_51327_n11370# a_51277_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1797 VDD a_28843_6408# a_28791_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1798 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1799 VDD a_818_1932# a_8328_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1800 a_51684_5708# a_51711_6449# a_51696_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1801 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1802 a_59745_773# a_59747_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1803 VSS a_57157_6408# a_57105_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1804 VDD a_33223_773# a_34148_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1805 VSS a_29290_n11298# a_29263_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1806 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1807 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1808 VDD a_4139_n11370# a_4089_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1809 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1810 a_33223_773# a_32729_690# a_32784_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1811 a_27520_n5879# a_27294_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1812 a_7136_n10732# a_6370_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1813 a_31660_n5622# a_31070_n5789# a_31564_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1814 a_48417_773# a_48419_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1815 a_59747_1829# a_59155_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1816 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1817 a_4345_n5795# a_4175_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1818 VDD a_1047_n6869# a_14221_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1819 a_50550_n11788# a_49782_n11533# a_48564_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1820 a_46433_773# a_48053_836# a_47877_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1821 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1822 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1823 a_38901_5953# a_40119_6434# a_40362_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1824 a_23881_1829# a_23289_690# a_21895_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1825 VDD a_53215_n11370# a_53165_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1826 VDD a_23179_6408# a_23397_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1827 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1828 VDD a_529_6408# a_477_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1829 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1830 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1831 a_55516_1994# a_55429_1896# a_55434_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1832 a_27375_n10487# a_27402_n11298# a_27387_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1833 a_10305_836# a_10079_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1834 a_15966_n5789# C[40] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1835 a_9024_n10732# a_8258_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1836 a_26012_n11788# a_25244_n11533# a_24026_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1837 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1838 a_23895_7009# a_23893_5953# a_24196_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1839 a_41417_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1840 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1841 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1842 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1843 a_4909_773# a_6529_836# a_6353_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1844 VDD a_31067_836# a_30891_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1845 VDD a_28677_n11370# a_28627_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1846 a_1147_5953# a_529_6408# a_747_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1847 a_34672_1994# a_34667_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1848 VDD a_57761_773# a_58686_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1849 VSS a_42663_773# a_43588_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1850 VSS a_37109_5953# a_37111_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1851 a_19214_696# a_19044_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1852 VDD a_55103_n11370# a_55053_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1853 a_58100_n10732# a_57334_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1854 a_8783_1829# a_8417_836# a_6797_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1855 VSS a_758_n11559# a_706_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1856 a_29263_n10487# a_29290_n11298# a_29275_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1857 a_134_6655# a_224_6410# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1858 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1859 a_34846_n5789# C[50] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1860 a_27431_n6843# a_27344_n6611# a_27349_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1861 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1862 a_48321_773# a_49941_836# a_49765_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1863 VSS a_1047_n6869# a_5234_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1864 a_27900_n11788# a_27132_n11533# a_25914_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1865 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1866 a_7892_696# a_7722_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1867 a_43305_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1868 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1869 VSS a_46118_1932# a_53546_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1870 a_21856_n5879# a_21630_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1871 a_33095_n6843# a_33008_n6611# a_33013_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1872 a_10160_5708# a_10187_6449# a_10172_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1873 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1874 a_52195_1829# a_51829_836# a_50209_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1875 a_57857_773# a_57267_690# a_57761_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1876 a_34983_n6843# a_34896_n6611# a_34901_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1877 VDD a_37888_6655# a_37838_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1878 a_27669_5953# a_26903_6434# a_27573_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1879 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1880 a_44890_n10732# a_44124_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1881 a_13948_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1882 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1883 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1884 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1885 a_33184_n5879# a_32958_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1886 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1887 a_40873_1829# a_40281_690# a_38887_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1888 a_59085_n5795# a_58915_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1889 VDD a_40171_6408# a_40389_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1890 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1891 VDD a_46118_1932# a_57404_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1892 a_10669_773# a_10305_836# a_10573_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1893 a_45193_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1894 a_15035_n6843# a_14676_n6678# a_14674_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1895 VDD a_21520_n11559# a_21468_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1896 a_11462_6655# a_10587_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1897 a_40507_836# a_40281_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1898 a_40736_n5879# a_40510_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1899 a_6358_1994# a_6353_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1900 VSS a_10802_n5622# a_11727_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1901 a_39116_n5622# a_38622_n5789# a_38677_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1902 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1904 VSS a_8795_5953# a_8797_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1905 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1906 VSS a_15916_1932# a_25767_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1907 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1908 a_54312_n6678# a_53946_n5879# a_52326_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1909 VSS C[16] a_28843_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1910 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1911 a_7483_n6843# a_7124_n6678# a_7122_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1912 a_38999_7009# a_38283_6408# a_37013_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1913 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1914 a_22990_696# a_22820_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1915 a_1245_7009# a_529_6408# a_224_6410# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1916 a_51684_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1917 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1918 a_26010_n10732# a_25244_n11533# a_25914_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1919 VDD a_12422_n5879# a_12246_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1920 VSS a_7026_n5622# a_7951_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1921 a_33319_773# a_32955_836# a_33223_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1922 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1923 a_57990_n5622# a_59610_n5879# a_59434_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1924 a_44780_n5622# a_46168_n5789# a_46218_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X1925 VSS a_13974_n11559# a_13922_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1926 a_30089_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1927 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1928 a_57761_773# a_57493_836# a_57322_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1929 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1930 a_38848_n5879# a_38622_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1931 a_21685_n6843# a_21680_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1932 VSS a_15916_1932# a_21991_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1933 VDD a_8417_836# a_8241_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1934 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1935 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1936 a_58088_n6678# a_57496_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1937 a_2837_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1938 VSS a_40400_n11559# a_40348_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1939 a_961_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1940 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1941 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1942 a_50438_n5622# a_51832_n5789# a_51882_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1943 VSS a_13963_6449# a_13936_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1944 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1945 a_9026_n11788# a_8258_n11533# a_7040_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1946 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1947 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1948 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1949 a_25671_773# a_25177_690# a_25232_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1950 a_44565_5953# a_43895_6434# a_44165_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1951 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1952 a_37013_5953# a_38283_6408# a_38474_5708# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1953 VDD a_49605_6408# a_49553_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1954 a_57859_1829# a_57493_836# a_55873_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1955 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1956 a_16572_n11788# a_15804_n11533# a_14592_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1957 a_23895_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1958 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1959 VDD a_1047_n6869# a_11259_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1960 a_40565_n6843# a_40560_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1961 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1962 VDD a_5798_6655# a_5748_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1963 a_19879_n6843# a_19792_n6611# a_19797_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1964 VDD a_19237_n11370# a_19187_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1965 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1966 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1967 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1968 a_38323_n5795# a_38153_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1969 VSS C[21] a_19403_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1970 VSS C[11] a_38283_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1971 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1972 a_868_n5789# C[32] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1973 VSS a_27173_6449# a_27146_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1974 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1975 a_48321_773# a_47827_690# a_47882_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1976 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1977 VDD a_2646_n11559# a_2594_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1978 a_59210_1994# a_59205_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1979 VSS a_31020_1932# a_42759_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1980 VDD a_23515_836# a_23339_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1981 a_1458_n5622# a_1460_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1982 a_18460_n11788# a_17692_n11533# a_16474_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1983 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1984 a_23881_1829# a_23289_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1985 a_49210_6655# a_48335_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1986 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1987 a_15232_6655# a_14363_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1988 a_38759_n6843# a_38672_n6611# a_38677_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1989 a_27671_7009# a_26903_6434# a_25685_5953# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1990 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1991 a_54097_7009# a_53381_6408# a_52111_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1992 a_42169_690# C[118] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1993 a_10160_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1994 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1995 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1996 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1997 VDD a_51493_6408# a_51441_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1998 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1999 a_25403_836# a_25177_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2000 a_36229_n11370# a_35354_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2001 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2002 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2003 VDD a_4534_n11559# a_4482_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2004 a_4345_n5795# a_4175_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2005 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2006 VDD a_2417_6408# a_2635_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2007 VSS a_57871_5953# a_57873_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2008 a_14445_773# a_14447_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2009 a_33319_773# a_32729_690# a_33223_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2010 a_46168_n5789# C[56] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2011 VDD a_46165_836# a_45989_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2012 a_48550_n5622# a_48056_n5789# a_48111_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2013 a_5236_n6678# a_4644_n5789# a_3250_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2014 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2015 a_50321_7009# a_49605_6408# a_48335_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2016 VDD a_8685_773# a_9610_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2017 a_30133_n6843# a_29774_n6678# a_29772_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2018 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2019 a_12461_773# a_14081_836# a_13905_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2020 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2021 a_3133_7009# a_3131_5953# a_3434_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2022 a_38486_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2023 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2024 a_54214_n5622# a_53720_n5789# a_53775_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2025 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2026 a_9024_n10732# a_8258_n11533# a_8928_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2027 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2028 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2029 a_59976_n6678# a_59610_n5879# a_57990_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2030 a_58088_n6678# a_57722_n5879# a_56102_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2031 a_40887_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2032 a_13855_690# C[103] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2033 a_38117_n11370# a_37242_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2034 a_1243_5953# a_529_6408# a_1147_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2035 VSS a_17733_6449# a_17706_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2036 a_22138_n10732# a_23408_n11559# a_23599_n10487# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=0p ps=0u w=650000u l=150000u
X2037 VDD a_6422_n11559# a_6370_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2038 a_36000_6655# a_35125_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2039 a_48335_5953# a_47665_6434# a_47935_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2040 VDD a_58650_6655# a_58600_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2041 a_29559_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2042 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2043 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2044 a_46394_n5879# a_46168_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2045 a_16570_n10732# a_15804_n11533# a_16474_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2046 a_48564_n10732# a_49834_n11559# a_50025_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2047 VDD C[18] a_25067_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2048 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2049 a_1362_n5622# a_2982_n5879# a_2806_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2050 a_42479_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2051 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2052 a_3348_n6678# a_2756_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2053 VDD a_31249_n6869# a_33095_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2054 a_46772_n10732# a_46006_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2055 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2056 VDD a_8646_n5879# a_8470_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2057 a_53946_n5879# a_53720_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2058 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2059 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2060 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2061 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2062 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2063 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2064 a_36505_690# C[115] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2065 a_32224_6655# a_31349_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2066 VDD a_31020_1932# a_37456_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2067 VDD a_31249_n6869# a_40647_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2068 VDD a_8310_n11559# a_8258_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2069 a_44663_7009# a_43895_6434# a_42677_5953# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2070 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2071 a_24026_n10732# a_25296_n11559# a_25487_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2072 a_6907_5953# a_6141_6434# a_6811_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2073 VSS a_48431_5953# a_48433_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2074 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2075 a_25767_773# a_25403_836# a_25671_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2076 a_33223_773# a_32955_836# a_32784_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2077 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2078 VDD a_23783_773# a_24708_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2079 a_50452_n10732# a_51722_n11559# a_51913_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2080 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2081 a_55605_836# a_55379_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2082 VDD a_59649_773# a_60574_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2083 VSS C[66] a_55498_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2084 a_59988_n10732# a_59222_n11533# a_59878_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2085 a_59761_7009# a_59045_6408# a_57775_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2086 a_3478_1994# a_3119_1829# a_3117_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2087 a_10898_n5622# a_10308_n5789# a_10802_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2088 a_12802_n11788# a_12086_n11559# a_10816_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2089 a_44367_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2090 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2091 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2092 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2093 a_33333_5953# a_32567_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2094 a_21102_696# a_20932_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2095 a_50319_5953# a_49553_6434# a_50223_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2096 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2097 a_53421_n5795# a_53251_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2098 VDD a_42288_n11559# a_42236_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2099 a_21482_5708# a_21509_6449# a_21494_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2100 VSS a_1047_n6869# a_10363_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2101 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2102 VDD a_1047_n6869# a_7483_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2103 a_25914_n10732# a_27184_n11559# a_27375_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2104 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2105 a_48417_773# a_48053_836# a_48321_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2106 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2107 VDD a_10802_n5622# a_11727_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2108 a_52340_n10732# a_53610_n11559# a_53801_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2109 VSS a_34725_6449# a_34698_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2110 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2111 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2112 a_18215_773# a_18217_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2113 VSS C[65] a_57386_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2114 a_14690_n11788# a_13974_n11559# a_12704_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2115 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2116 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2117 VDD a_51493_6408# a_51711_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2118 a_16231_773# a_17851_836# a_17675_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2119 a_8685_773# a_8417_836# a_8246_1994# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=0p ps=0u w=650000u l=150000u
X2120 a_53857_n6843# a_53770_n6611# a_53775_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2121 a_57775_5953# a_59045_6408# a_59236_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2122 a_40885_5953# a_40171_6408# a_40789_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2123 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2124 VSS a_1047_n6869# a_8475_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2125 a_41116_n11788# a_40400_n11559# a_39130_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2126 a_8699_5953# a_9917_6434# a_10160_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2127 VDD C[9] a_42059_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2128 a_56762_6655# a_55887_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2129 a_22784_6655# a_21909_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2130 VDD a_44176_n11559# a_44124_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2131 a_24026_n10732# a_23408_n11559# a_23626_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2132 a_59439_n6843# a_59434_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2133 VSS a_818_1932# a_1229_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2134 VDD a_7026_n5622# a_7951_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2135 a_3910_6655# a_3035_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2136 VDD a_818_1932# a_9142_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2137 a_25314_1994# a_25227_1896# a_25232_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2138 a_27802_n10732# a_29072_n11559# a_29263_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2139 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2140 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2141 a_5138_n5622# a_4870_n5879# a_4699_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2142 VSS a_46347_n6869# a_46758_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2143 a_50452_n10732# a_49834_n11559# a_50052_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2144 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2145 a_31335_773# a_32729_690# a_32779_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2146 a_16329_1829# a_15737_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2147 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2148 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2149 a_12196_n5789# C[38] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2150 a_10912_n10732# a_10198_n11559# a_10816_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2151 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2152 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2153 VDD a_818_1932# a_5366_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2154 a_21538_1994# a_21451_1896# a_21456_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2155 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2156 a_59878_n5622# a_59384_n5789# a_59439_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2157 a_3348_n6678# a_2982_n5879# a_1362_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2158 a_3133_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2159 a_25914_n10732# a_25296_n11559# a_25514_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2160 a_732_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2161 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2162 a_48433_7009# a_47665_6434# a_46447_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2163 VSS a_33223_773# a_34148_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2164 a_52340_n10732# a_51722_n11559# a_51940_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2165 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2166 VDD a_31296_n5879# a_31120_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2167 a_12422_n5879# a_12196_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2168 a_12800_n10732# a_12086_n11559# a_12704_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2169 a_55887_5953# a_55217_6434# a_55487_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2170 VSS a_15916_1932# a_23344_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2171 a_38323_n5795# a_38153_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2172 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2173 a_57267_690# C[126] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2174 a_33039_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2175 a_35207_773# a_35209_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2176 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2177 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2178 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2179 a_39228_n11788# a_38460_n11533# a_37242_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2180 a_27802_n10732# a_27184_n11559# a_27402_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2181 a_59248_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2182 a_48417_773# a_47827_690# a_48321_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2183 a_14592_n10732# a_15856_n11559# a_16047_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2184 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2185 a_10671_1829# a_10079_690# a_8685_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2186 VDD a_9969_6408# a_10187_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2187 VDD a_15916_1932# a_27202_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2188 a_13556_696# a_13386_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2189 a_16460_n5622# a_17854_n5789# a_17904_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2190 a_14688_n10732# a_13974_n11559# a_14592_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2191 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2192 a_42306_1994# a_42219_1896# a_42224_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2193 a_56330_1994# a_55971_1829# a_55969_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2194 a_40510_n5789# C[53] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2195 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2196 VSS C[71] a_46058_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2197 VSS a_46118_1932# a_54081_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2198 VSS a_57761_773# a_58686_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2199 a_41114_n10732# a_40400_n11559# a_41018_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2200 a_50321_7009# a_49553_6434# a_48335_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2201 a_24012_n5622# a_25406_n5789# a_25456_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X2202 a_10685_7009# a_10683_5953# a_10986_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2203 a_28953_690# C[111] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2204 a_24901_n11370# a_24026_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2205 VDD C[7] a_45829_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2206 a_57197_n5795# a_57027_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2207 a_29690_n10732# a_29072_n11559# a_29290_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2208 a_36999_773# a_38393_690# a_38443_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2209 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2210 a_453_n11561# a_639_690# a_689_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2211 a_31067_836# a_30841_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2212 a_21482_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2213 a_16474_n10732# a_17744_n11559# a_17935_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2214 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2215 VSS a_9574_6655# a_9524_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2216 a_36206_696# a_36036_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2217 a_12251_n6843# a_12246_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2218 a_35340_n5622# a_36734_n5789# a_36784_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2219 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2220 VSS C[70] a_47946_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2221 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2222 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2223 a_46020_5708# a_46047_6449# a_46032_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2224 a_5234_n5622# a_4870_n5879# a_5138_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2225 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2226 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2227 a_6893_773# a_6895_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2228 a_42892_n5622# a_44286_n5789# a_44336_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2229 VSS a_50052_n11298# a_50025_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2230 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2231 VSS a_31020_1932# a_40336_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2232 a_8781_773# a_8191_690# a_8685_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2233 a_4699_n6843# a_4694_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2234 a_34939_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2235 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2236 a_23783_773# a_25403_836# a_25227_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2237 a_49808_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2238 VSS a_59263_6449# a_59236_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2239 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2240 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2241 a_48321_773# a_48053_836# a_47882_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2242 a_21630_n5789# C[43] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2243 a_54095_5953# a_53329_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2244 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2245 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2246 a_19008_6655# a_18133_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2247 a_14459_5953# a_13693_6434# a_14363_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2248 a_52209_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2249 VSS a_40005_n11370# a_39955_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2250 VDD a_19403_6408# a_19351_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2251 a_27657_1829# a_27291_836# a_25671_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2252 a_46890_1994# a_46531_1829# a_46529_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2253 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2254 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2255 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2256 VDD C[31] a_529_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2257 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2258 a_16231_773# a_15737_690# a_15792_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2259 a_8928_n10732# a_8310_n11559# a_8528_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2260 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2261 VDD a_31020_1932# a_44194_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2262 a_39226_n10732# a_38460_n11533# a_39130_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2263 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2264 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2265 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2266 VSS a_55487_6449# a_55460_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2267 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2268 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2269 a_32729_690# C[113] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2270 a_16474_n10732# a_15856_n11559# a_16074_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2271 a_19742_n5789# C[42] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2272 a_29461_5953# a_30679_6434# a_30922_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2273 a_29008_1994# a_29003_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2274 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2275 a_55985_7009# a_55217_6434# a_53999_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2276 VSS a_6193_6408# a_6141_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2277 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2278 a_51829_836# a_51603_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2279 a_46076_1994# a_45989_1896# a_45994_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2280 a_23879_773# a_23289_690# a_23783_773# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2281 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2282 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2283 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2284 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2285 a_25406_n5789# C[45] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2286 a_53421_n5795# a_53251_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2287 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2288 a_50025_n10487# a_50052_n11298# a_50037_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2289 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2290 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2291 a_8646_n5879# a_8420_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2292 VDD a_21291_6408# a_21239_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2293 a_38985_1829# a_38393_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2294 a_18362_n10732# a_17744_n11559# a_17962_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2295 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2296 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2297 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2298 VSS a_16570_n10732# a_16572_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2299 VSS a_2417_6408# a_2365_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2300 a_18080_n5879# a_17854_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2301 a_37326_n6678# a_36960_n5879# a_35340_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2302 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2303 a_22220_n5622# a_21630_n5789# a_22124_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2304 VSS a_27669_5953# a_27671_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2305 a_44780_n5622# a_46394_n5879# a_46218_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2306 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2307 a_3119_1829# a_2527_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2308 a_25632_n5879# a_25406_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2309 a_44286_n5789# C[55] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2310 a_20119_7009# a_19403_6408# a_18133_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2311 VDD a_31020_1932# a_34754_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2312 VDD a_46118_1932# a_48778_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2313 a_54627_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2314 a_44649_1829# a_44283_836# a_42663_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2315 VSS a_16145_n6869# a_23573_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2316 a_27788_n5622# a_29182_n5789# a_29232_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X2317 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2318 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2319 a_2457_n5795# a_2287_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2320 a_35209_1829# a_34617_690# a_33223_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2321 VDD a_1047_n6869# a_12333_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2322 a_15461_n11370# a_14592_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2323 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2324 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2325 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2326 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2327 VSS a_18458_n10732# a_18460_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2328 a_20021_5953# a_21239_6434# a_21482_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2329 a_50305_773# a_49941_836# a_50209_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2330 VDD C[3] a_53381_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2331 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2332 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2333 a_1147_5953# a_2365_6434# a_2608_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2334 VDD a_28448_6655# a_28398_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2335 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2336 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2337 a_9803_n11370# a_8928_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2338 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2339 a_23783_773# a_23515_836# a_23344_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2340 a_44512_n5879# a_44286_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2341 VSS a_29786_n10732# a_29788_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2342 a_39130_n10732# a_40348_n11533# a_40591_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2343 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2344 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2345 a_31433_1829# a_30841_690# a_29447_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2346 a_8191_690# C[100] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2347 a_56515_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2348 VDD a_46118_1932# a_47964_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2349 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2350 VDD a_30731_6408# a_30949_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2351 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2352 a_15792_1994# a_15787_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2353 a_8475_n6843# a_8470_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2354 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2355 a_16572_n11788# a_16570_n10732# a_16873_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2356 a_14461_7009# a_13693_6434# a_12475_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2357 a_58879_n11370# a_58004_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2358 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2359 VSS a_18229_5953# a_18231_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2360 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2361 a_28654_696# a_28484_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2362 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2363 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2364 a_46758_n5622# a_46760_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2365 VDD a_134_6655# a_84_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2366 a_48646_n5622# a_48648_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2367 a_27065_690# C[110] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2368 a_21711_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2369 a_29559_7009# a_28843_6408# a_27573_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2370 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2371 a_32958_n5789# C[49] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2372 a_25543_n6843# a_25456_n6611# a_25461_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2373 VDD a_26955_6408# a_26903_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2374 VDD a_818_1932# a_6440_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2375 a_58403_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2376 VSS a_44661_5953# a_44663_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2377 VSS a_8685_773# a_9610_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2378 VSS a_55269_6408# a_55217_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2379 a_20117_5953# a_19351_6434# a_20021_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2380 a_31207_n6843# a_31120_n6611# a_31125_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2381 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2382 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2383 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2384 a_46165_836# a_45939_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2385 a_39212_n5622# a_38848_n5879# a_39116_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2386 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2387 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2388 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2389 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2390 VSS a_51722_n11559# a_51670_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2391 a_18460_n11788# a_18458_n10732# a_18761_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2392 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2393 a_50209_773# a_49715_690# a_49770_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2394 a_12289_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2395 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2396 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2397 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2398 VDD a_818_1932# a_2664_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2399 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2400 a_31296_n5879# a_31070_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2401 a_29788_n11788# a_29786_n10732# a_30089_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2402 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2403 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2404 a_3021_773# a_2527_690# a_2582_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2405 a_35125_5953# a_34455_6434# a_34725_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2406 VSS a_46118_1932# a_49770_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2407 a_21993_1829# a_21401_690# a_20007_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2408 a_57197_n5795# a_57027_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2409 VDD a_21291_6408# a_21509_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2410 a_3119_1829# a_2527_690# a_1133_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2411 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2412 a_27573_5953# a_28843_6408# a_29034_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2413 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2414 a_53628_1994# a_53541_1896# a_53546_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2415 a_58088_n6678# a_57496_n5789# a_56102_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2416 VDD C[25] a_11857_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2417 a_26560_6655# a_25685_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2418 a_59976_n6678# a_59384_n5789# a_57990_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2419 a_13147_n6843# a_12788_n6678# a_12786_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2420 a_46760_n6678# a_46394_n5879# a_44780_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2421 VDD a_13714_3465# a_36341_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2422 a_37228_n5622# a_36734_n5789# a_36789_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2423 VSS a_53610_n11559# a_53558_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2424 a_14592_n10732# a_13922_n11533# a_14192_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2425 a_14177_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2426 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2427 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2428 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2429 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2430 a_52424_n6678# a_52058_n5879# a_50438_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2431 a_32784_1994# a_32779_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2432 a_3021_773# a_4641_836# a_4465_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2433 a_5595_n6843# a_5236_n6678# a_5234_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2434 VSS a_23783_773# a_24708_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2435 VSS a_31249_n6869# a_44876_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2436 a_41018_n10732# a_40348_n11533# a_40618_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2437 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2438 VSS a_59649_773# a_60574_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2439 VDD a_10534_n5879# a_10358_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2440 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2441 VSS a_35221_5953# a_35223_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2442 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2443 a_6529_836# a_6303_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2444 VSS a_5138_n5622# a_6063_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2445 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2446 a_6895_1829# a_6529_836# a_4909_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2447 a_30841_690# C[112] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2448 a_47827_690# C[121] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2449 a_56102_n5622# a_57722_n5879# a_57546_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2450 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2451 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2452 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2453 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2454 VDD a_43947_6408# a_43895_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2455 a_29860_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2456 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2457 a_56200_n6678# a_55608_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2458 a_18231_7009# a_17463_6434# a_16245_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2459 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2460 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2461 a_26128_1994# a_25769_1829# a_25767_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2462 VSS a_46118_1932# a_51658_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2463 a_50307_1829# a_49941_836# a_48321_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2464 VDD a_1047_n6869# a_8557_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2465 a_2753_836# a_2527_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2466 a_25685_5953# a_25015_6434# a_25285_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2467 a_41893_n11370# a_41018_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2468 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2469 a_59610_n5879# a_59384_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2470 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2471 a_18133_5953# a_19403_6408# a_19594_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2472 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2473 a_53491_690# C[124] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2474 a_47075_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2475 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2476 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2477 VDD a_46118_1932# a_55516_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2478 VDD a_38619_836# a_38443_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2479 a_4725_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2480 a_29046_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2481 a_49439_n11370# a_48564_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2482 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2483 a_43552_6655# a_42677_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2484 a_8699_5953# a_8081_6408# a_8299_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2485 a_21627_836# a_21401_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2486 a_4470_1994# a_4465_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2487 VDD a_1047_n6869# a_1819_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2488 a_12104_1994# a_12017_1896# a_12022_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2489 a_43781_n11370# a_42906_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2490 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2491 VSS a_6907_5953# a_6909_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2492 VSS a_15916_1932# a_23879_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2493 VDD a_36624_n11559# a_36842_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2494 VDD a_49210_6655# a_49160_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2495 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2496 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2497 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2498 VSS a_15856_n11559# a_15804_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2499 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2500 a_10683_5953# a_9917_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2501 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2502 a_54310_n5622# a_53946_n5879# a_54214_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2503 a_6613_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2504 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2505 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2506 VSS a_15916_1932# a_20103_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2507 a_1474_n11788# a_758_n11559# a_453_n11561# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2508 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2509 VDD a_15916_1932# a_28016_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2510 a_2457_n5795# a_2287_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2511 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2512 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2513 a_59878_n5622# a_59610_n5879# a_59439_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2514 a_3348_n6678# a_2756_n5789# a_1362_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2515 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2516 a_46662_n5622# a_46168_n5789# a_46223_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2517 a_55689_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2518 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2519 VSS a_818_1932# a_10134_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2520 VSS a_17744_n11559# a_17692_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2521 a_42677_5953# a_42007_6434# a_42277_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2522 a_40873_1829# a_40281_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2523 a_35125_5953# a_36395_6408# a_36586_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2524 VDD a_47717_6408# a_47665_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2525 a_19606_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2526 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2527 a_52326_n5622# a_51832_n5789# a_51887_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2528 a_50550_n11788# a_49834_n11559# a_48564_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2529 a_8501_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2530 a_23893_5953# a_23127_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2531 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2532 a_22007_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2533 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2534 VDD a_3910_6655# a_3860_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2535 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2536 a_13556_696# a_13386_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2537 VDD a_14310_n5879# a_14134_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2538 a_30565_n11370# a_29690_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2539 VDD a_818_1932# a_13992_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2540 a_26012_n11788# a_25296_n11559# a_24026_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2541 a_57577_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2542 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2543 a_8797_7009# a_8081_6408# a_6811_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2544 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2545 VSS a_19632_n11559# a_19580_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2546 VSS a_25285_6449# a_25258_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2547 a_57322_1994# a_57317_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2548 a_1460_n6678# a_868_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2549 VDD a_31249_n6869# a_31207_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2550 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2551 VSS a_31020_1932# a_40871_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2552 VDD a_1133_773# a_2058_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2553 VDD a_38887_773# a_39812_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2554 VDD a_6758_n5879# a_6582_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2555 a_52058_n5879# a_51832_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2556 a_52438_n11788# a_51722_n11559# a_50452_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2557 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2558 VDD a_55498_n11559# a_55446_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2559 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2560 a_47322_6655# a_46447_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2561 a_31445_5953# a_30731_6408# a_31349_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2562 VSS a_15916_1932# a_29543_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2563 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2564 a_25783_7009# a_25015_6434# a_23797_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2565 a_36206_696# a_36036_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2566 a_23289_690# C[108] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2567 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2568 a_52209_7009# a_51493_6408# a_50223_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2569 a_31676_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2570 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2571 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2572 a_32453_n11370# a_31578_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2573 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2574 a_27900_n11788# a_27184_n11559# a_25914_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2575 a_59465_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2576 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2577 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2578 a_8420_n5789# C[36] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2579 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2580 VDD a_10198_n11559# a_10416_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2581 VSS a_55983_5953# a_55985_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2582 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2583 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2584 a_12557_773# a_12559_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2585 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2586 a_54326_n11788# a_53610_n11559# a_52340_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2587 a_6811_5953# a_8081_6408# a_8272_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2588 a_30542_696# a_30372_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2589 VDD a_57386_n11559# a_57334_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2590 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2591 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2592 a_10573_773# a_12193_836# a_12017_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2593 VDD a_1047_n6869# a_5595_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2594 VDD C[95] a_758_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2595 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2596 a_1245_7009# a_1243_5953# a_1546_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2597 a_36598_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2598 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2599 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2600 a_5234_n5622# a_4644_n5789# a_5138_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2601 a_33564_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2602 a_34341_n11370# a_33466_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2603 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2604 VSS C[27] a_8081_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2605 a_29788_n11788# a_29072_n11559# a_27802_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2606 a_50223_5953# a_51493_6408# a_51684_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2607 VSS a_15845_6449# a_15818_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2608 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2609 a_14447_1829# a_14081_836# a_12461_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2610 a_33680_1994# a_33321_1829# a_33319_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2611 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2612 a_46447_5953# a_45777_6434# a_46047_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2613 VDD a_12086_n11559# a_12304_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2614 a_50548_n10732# a_49834_n11559# a_50452_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2615 VDD a_56762_6655# a_56712_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2616 a_56214_n11788# a_55498_n11559# a_54228_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2617 a_58086_n5622# a_57722_n5879# a_57990_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2618 VSS a_1047_n6869# a_6587_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2619 VDD a_59274_n11559# a_59222_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2620 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2621 a_51969_n6843# a_51882_n6611# a_51887_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2622 a_22005_5953# a_21291_6408# a_21909_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2623 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2624 a_53192_696# a_53022_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2625 a_59974_n5622# a_59610_n5879# a_59878_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2626 VDD C[19] a_23179_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2627 VSS a_42277_6449# a_42250_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2628 VDD a_5138_n5622# a_6063_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2629 VDD C[94] a_2646_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2630 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2631 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2632 a_35452_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2633 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2634 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2635 a_3250_n5622# a_2982_n5879# a_2811_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2636 a_26010_n10732# a_25296_n11559# a_25914_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2637 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2638 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2639 a_30336_6655# a_29461_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2640 a_17625_690# C[105] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2641 a_10308_n5789# C[37] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2642 a_42775_7009# a_42007_6434# a_40789_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2643 a_5019_5953# a_4253_6434# a_4923_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2644 VSS a_46543_5953# a_46545_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2645 VDD a_13974_n11559# a_14192_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2646 a_52436_n10732# a_51722_n11559# a_52340_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2647 a_46249_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2648 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2649 a_52510_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2650 a_38887_773# a_38619_836# a_38448_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2651 VDD C[68] a_51722_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2652 a_39212_n5622# a_39214_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2653 VSS a_46347_n6869# a_58086_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2654 a_57873_7009# a_57157_6408# a_55887_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2655 a_13936_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2656 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2657 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2658 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2659 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2660 a_27559_773# a_28953_690# a_29003_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2661 VDD C[93] a_4534_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2662 a_31445_5953# a_30679_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2663 a_8284_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2664 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2665 a_27898_n10732# a_27184_n11559# a_27802_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2666 a_42663_773# a_42169_690# a_42224_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2667 VSS a_50548_n10732# a_50550_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2668 a_20348_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2669 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2670 a_10534_n5879# a_10308_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2671 a_21125_n11370# a_20250_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2672 VSS a_25067_6408# a_25015_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2673 a_38474_5708# a_38501_6449# a_38486_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2674 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2675 VSS a_2251_n11370# a_2201_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2676 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2677 a_16572_n11788# a_15856_n11559# a_14592_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2678 a_54324_n10732# a_53610_n11559# a_54228_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2679 a_48137_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2680 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2681 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2682 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2683 VDD a_31020_1932# a_35568_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2684 a_639_690# C[96] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2685 a_24110_n6678# a_23744_n5879# a_22124_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2686 VDD C[67] a_53610_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2687 a_16327_773# a_16329_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2688 VSS a_32837_6449# a_32810_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2689 VDD a_46058_n11559# a_46006_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2690 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2691 VSS a_31020_1932# a_30896_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2692 a_1229_773# a_865_836# a_1133_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2693 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2694 a_14349_773# a_15963_836# a_15787_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2695 a_31070_n5789# C[48] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2696 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2697 VSS a_51327_n11370# a_51277_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2698 a_55887_5953# a_57157_6408# a_57348_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2699 VDD C[10] a_40171_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2700 a_54874_6655# a_53999_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2701 a_29786_n10732# a_29072_n11559# a_29690_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2702 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2703 a_20896_6655# a_20021_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2704 VSS a_15916_1932# a_19568_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2705 VDD a_14349_773# a_15274_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2706 VSS a_52436_n10732# a_52438_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2707 a_39776_6655# a_38901_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2708 a_27788_n5622# a_29408_n5879# a_29232_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2709 a_14578_n5622# a_15966_n5789# a_16016_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2710 a_23013_n11370# a_22138_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2711 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2712 a_2022_6655# a_1147_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2713 VDD a_818_1932# a_7254_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2714 a_23426_1994# a_23339_1896# a_23344_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2715 VSS a_4139_n11370# a_4089_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2716 a_49645_n5795# a_49475_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2717 a_18460_n11788# a_17744_n11559# a_16474_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X2718 VDD a_40507_836# a_40331_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2719 a_27886_n6678# a_27294_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2720 VSS a_54214_n5622# a_55139_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2721 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2722 a_20236_n5622# a_21630_n5789# a_21680_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2723 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2724 a_22124_n5622# a_23518_n5789# a_23568_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2725 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2726 a_55309_n5795# a_55139_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2727 VDD C[74] a_40400_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2728 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2729 a_18119_773# a_19513_690# a_19563_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2730 a_15737_690# C[104] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2731 a_28654_696# a_28484_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2732 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2733 a_54097_7009# a_54095_5953# a_54398_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2734 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2735 VSS a_53215_n11370# a_53165_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2736 a_42395_836# a_42169_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2737 a_50550_n11788# a_50548_n10732# a_50851_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2738 a_33452_n5622# a_34846_n5789# a_34896_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2739 a_14445_773# a_13855_690# a_14349_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2740 a_10363_n6843# a_10358_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2741 a_46545_7009# a_45777_6434# a_44565_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X2742 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2743 a_3346_n5622# a_2982_n5879# a_3250_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2744 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2745 VDD a_13745_6408# a_13693_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2746 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2747 VSS a_4523_6449# a_4496_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2748 a_41004_n5622# a_42398_n5789# a_42448_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X2749 a_453_n11561# a_706_n11533# a_949_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2750 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2751 VSS a_42059_6408# a_42007_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2752 a_53999_5953# a_53329_6434# a_53599_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2753 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2754 VSS a_15916_1932# a_21456_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X2755 a_2811_n6843# a_2806_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2756 VSS a_28677_n11370# a_28627_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2757 VDD C[73] a_42288_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2758 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2759 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2760 a_20105_1829# a_19739_836# a_18119_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2761 VSS a_55103_n11370# a_55053_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2762 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2763 a_52438_n11788# a_52436_n10732# a_52739_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2764 a_16570_n10732# a_15856_n11559# a_16474_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2765 a_5021_7009# a_4253_6434# a_3035_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2766 a_36341_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2767 a_37095_773# a_36505_690# a_36999_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2768 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2769 a_57871_5953# a_57105_6434# a_57775_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2770 a_10914_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2771 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2772 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2773 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2774 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2775 VDD a_15916_1932# a_25314_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2776 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2777 a_1376_n10732# a_2594_n11533# a_2837_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2778 a_40418_1994# a_40331_1896# a_40336_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2779 a_54442_1994# a_54083_1829# a_54081_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2780 VDD C[72] a_44176_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2781 VSS a_10416_n11298# a_10389_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2782 a_13350_6655# a_12475_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2783 a_1229_773# a_639_690# a_1133_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2784 a_38983_773# a_38393_690# a_38887_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2785 a_36827_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2786 a_54310_n5622# a_54312_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2787 a_4139_n11370# a_3264_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2788 a_17854_n5789# C[41] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2789 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2790 VDD a_19008_6655# a_18958_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2791 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2792 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2793 a_45939_690# C[120] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2794 a_14349_773# a_14081_836# a_13910_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2795 a_18458_n10732# a_17744_n11559# a_18362_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2796 a_50452_n10732# a_51670_n11533# a_51913_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2797 a_12802_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2798 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2799 a_36731_836# a_36505_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2800 a_42759_773# a_42395_836# a_42663_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2801 a_23518_n5789# C[44] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2802 VSS C[0] a_59045_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2803 a_38474_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2804 VDD a_40775_773# a_41700_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2805 a_25900_n5622# a_25406_n5789# a_25461_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2806 VDD a_363_n11370# a_313_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2807 VSS a_7686_6655# a_7636_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2808 a_17326_696# a_17156_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2809 a_29774_n6678# a_29408_n5879# a_27788_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2810 a_3264_n10732# a_4482_n11533# a_4725_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2811 a_55983_5953# a_55217_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2812 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2813 VSS a_12304_n11298# a_12277_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2814 VSS C[6] a_47717_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2815 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2816 a_6758_n5879# a_6532_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2817 a_38715_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2818 a_865_836# a_639_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2819 VDD C[80] a_29072_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2820 a_5250_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2821 a_6027_n11370# a_5152_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2822 a_16192_n5879# a_15966_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2823 a_36734_n5789# C[51] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2824 VDD a_24901_n11370# a_24851_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2825 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2826 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2827 a_5005_773# a_5007_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2828 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2829 a_6004_696# a_5834_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2830 a_20332_n5622# a_19742_n5789# a_20236_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2831 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2832 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2833 a_52340_n10732# a_53558_n11533# a_53801_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2834 a_23744_n5879# a_23518_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2835 a_42398_n5789# C[54] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2836 a_52207_5953# a_51441_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2837 a_12475_5953# a_11805_6434# a_12075_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2838 a_4415_690# C[98] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2839 a_44780_n5622# a_44286_n5789# a_44341_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2840 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2841 a_1376_n10732# a_706_n11533# a_976_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2842 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2843 VDD a_17515_6408# a_17463_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2844 a_25769_1829# a_25403_836# a_23783_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2845 a_10389_n10487# a_10416_n11298# a_10401_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2846 a_1133_773# a_865_836# a_694_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2847 VDD a_1047_n6869# a_10445_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2848 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2849 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2850 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2851 VDD C[79] a_30960_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2852 a_7915_n11370# a_7040_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2853 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2854 VDD a_31020_1932# a_42306_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2855 a_35072_n5879# a_34846_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2856 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2857 a_57761_773# a_57267_690# a_57322_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2858 a_36960_n5879# a_36734_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2859 a_27802_n10732# a_29020_n11533# a_29263_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2860 VSS a_53599_6449# a_53572_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2861 VDD a_11691_n11370# a_11641_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2862 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2863 a_14688_n10732# a_13922_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2864 a_50452_n10732# a_49782_n11533# a_50052_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2865 a_50037_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2866 a_6797_773# a_8191_690# a_8241_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2867 a_54228_n10732# a_55446_n11533# a_55689_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2868 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2869 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2870 a_42624_n5879# a_42398_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2871 a_48550_n5622# a_49944_n5789# a_49994_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2872 a_33321_1829# a_32729_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2873 a_41114_n10732# a_40348_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2874 a_27120_1994# a_27115_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X2875 a_3264_n10732# a_2594_n11533# a_2864_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2876 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2877 VSS a_51098_6655# a_51048_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2878 VSS a_818_1932# a_10669_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2879 a_14991_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2880 VDD a_36000_6655# a_35950_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2881 a_12277_n10487# a_12304_n11298# a_12289_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2882 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2883 a_6587_n6843# a_6582_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2884 a_17120_6655# a_16245_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2885 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2886 VSS a_19237_n11370# a_19187_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2887 VDD C[78] a_32848_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2888 VSS C[75] a_38512_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2889 a_25499_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2890 a_50209_773# a_51603_690# a_51653_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2891 VDD a_46347_n6869# a_47119_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X2892 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2893 VDD a_13579_n11370# a_13529_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2894 VDD a_38283_6408# a_38231_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2895 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2896 a_52340_n10732# a_51670_n11533# a_51940_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2897 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2898 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2899 VDD a_55605_836# a_55429_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2900 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2901 a_23655_n6843# a_23568_n6611# a_23573_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2902 a_43002_n10732# a_42236_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2903 a_55971_1829# a_55379_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2904 a_40775_773# a_40507_836# a_40336_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2905 VSS a_25781_5953# a_25783_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2906 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2907 a_38393_690# C[116] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2908 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2909 a_57857_773# a_57859_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2910 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2911 a_37324_n5622# a_36960_n5879# a_37228_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2912 a_27802_n10732# a_27132_n11533# a_27402_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2913 a_27387_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2914 a_58086_n5622# a_58088_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2915 VDD a_46118_1932# a_46890_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2916 VDD a_34507_6408# a_34455_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2917 a_57493_836# a_57267_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2918 a_49645_n5795# a_49475_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2919 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2920 a_54228_n10732# a_53558_n11533# a_53828_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2921 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2922 VDD a_54214_n5622# a_55139_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2923 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2924 a_29408_n5879# a_29182_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2925 a_42535_n6843# a_42448_n6611# a_42453_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2926 a_37013_5953# a_38231_6434# a_38474_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2927 VDD C[4] a_51493_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2928 a_16245_5953# a_15575_6434# a_15845_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2929 a_55309_n5795# a_55139_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2930 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2931 a_224_6410# a_477_6434# a_720_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2932 VDD a_26560_6655# a_26510_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2933 a_29676_n5622# a_29182_n5789# a_29237_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X2934 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2935 VSS a_1133_773# a_2058_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2936 VSS a_38887_773# a_39812_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2937 VDD a_7915_n11370# a_7865_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2938 a_56200_n6678# a_55608_n5789# a_54214_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2939 a_11259_n6843# a_10900_n6678# a_10898_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2940 VSS a_12075_6449# a_12048_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2941 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2942 a_29275_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2943 a_44112_1994# a_44107_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2944 a_29690_n10732# a_29020_n11533# a_29290_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2945 a_12193_836# a_11967_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2946 VDD a_46118_1932# a_46076_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2947 a_51832_n5789# C[59] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2948 a_3707_n6843# a_3348_n6678# a_3346_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2949 a_56116_n10732# a_55446_n11533# a_55716_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2950 a_34112_6655# a_33237_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2951 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2952 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2953 a_46662_n5622# a_48282_n5879# a_48106_n6611# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2954 a_12573_7009# a_11805_6434# a_10587_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2955 VSS a_9969_6408# a_9917_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2956 VSS a_16341_5953# a_16343_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2957 VSS a_3250_n5622# a_4175_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2958 a_46760_n6678# a_46168_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2959 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2960 a_48648_n6678# a_48056_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2961 VDD a_9803_n11370# a_9753_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2962 a_30542_696# a_30372_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2963 a_27671_7009# a_26955_6408# a_25685_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2964 a_59236_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2965 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2966 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2967 VDD a_818_1932# a_4552_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2968 VSS a_42773_5953# a_42775_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2969 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2970 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2971 a_50170_n5879# a_49944_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2972 a_949_n10487# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2973 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2974 a_29447_773# a_29179_836# a_29008_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2975 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2976 a_37109_5953# a_36343_6434# a_37013_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2977 a_57857_773# a_57493_836# a_57761_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2978 VDD a_55873_773# a_56798_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2979 a_28883_n5795# a_28713_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2980 a_53192_696# a_53022_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2981 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2982 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2983 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2984 a_33237_5953# a_32567_6434# a_32837_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2985 a_4116_696# a_3946_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2986 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2987 VDD a_38283_6408# a_38501_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2988 VDD a_43552_6655# a_43502_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2989 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2990 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2991 a_1231_1829# a_639_690# a_453_n11561# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2992 a_16059_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2993 a_25685_5953# a_26955_6408# a_27146_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2994 VDD C[26] a_9969_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2995 a_24672_6655# a_23797_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2996 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2997 a_9098_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2998 a_43004_n11788# a_42236_n11533# a_41018_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2999 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3000 VDD a_46347_n6869# a_58447_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3001 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3002 a_32955_836# a_32729_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3003 VDD a_758_n11559# a_706_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3004 a_58086_n5622# a_57496_n5789# a_57990_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3005 a_12690_n5622# a_14084_n5789# a_14134_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3006 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3007 a_59974_n5622# a_59384_n5789# a_59878_n5622# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X3008 a_30896_1994# a_30891_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3009 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3010 a_40871_773# a_40281_690# a_40775_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3011 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3012 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3013 VSS C[24] a_13745_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3014 a_49796_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3015 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3016 VSS a_33333_5953# a_33335_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3017 a_5007_1829# a_4641_836# a_3021_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3018 a_52422_n5622# a_52058_n5879# a_52326_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3019 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3020 a_38901_5953# a_38283_6408# a_38501_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3021 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3022 a_18362_n10732# a_17692_n11533# a_17962_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3023 VSS a_46347_n6869# a_59439_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3024 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3025 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3026 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3027 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3028 a_44892_n11788# a_44124_n11533# a_42906_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X3029 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3030 a_44663_7009# a_43947_6408# a_42677_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3031 a_27972_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3032 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3033 a_51740_1994# a_51653_1896# a_51658_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3034 a_48419_1829# a_47827_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3035 VSS a_16145_n6869# a_27884_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X3036 a_16343_7009# a_15575_6434# a_14363_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3037 a_56102_n5622# a_55834_n5879# a_55663_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3038 a_57990_n5622# a_57722_n5879# a_57551_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X3039 a_1460_n6678# a_868_n5789# a_224_6410# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3040 VDD a_59045_6408# a_58993_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3041 VDD a_21520_n11559# a_21738_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3042 a_23797_5953# a_23127_6434# a_23397_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3043 a_48648_n6678# a_48282_n5879# a_46662_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3044 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3045 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3046 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3047 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3048 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3049 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3050 VSS a_14349_773# a_15274_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3051 VDD a_19739_836# a_19563_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3052 a_45663_n11370# a_44794_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3053 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3054 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3055 a_42677_5953# a_43947_6408# a_44138_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X3056 a_27158_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3057 a_41664_6655# a_40789_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3058 a_6895_1829# a_6303_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3059 a_2582_1994# a_2577_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3060 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3061 a_54083_1829# a_53491_690# a_52097_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3062 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3063 VDD a_23408_n11559# a_23626_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3064 a_10216_1994# a_10129_1896# a_10134_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3065 a_24240_1994# a_23881_1829# a_23879_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3066 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3067 VSS a_5019_5953# a_5021_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3068 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3069 VDD a_4870_n5879# a_4694_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3070 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3071 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3072 a_10914_n11788# a_10198_n11559# a_8928_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3073 VDD a_49834_n11559# a_50052_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3074 a_37111_7009# a_36343_6434# a_35125_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3075 VDD a_47322_6655# a_47272_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3076 VDD a_13974_n11559# a_13922_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3077 a_43002_n10732# a_42236_n11533# a_42906_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3078 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3079 a_14084_n5789# C[39] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3080 a_29543_773# a_28953_690# a_29447_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3081 a_40887_7009# a_40885_5953# a_41188_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3082 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3083 a_45646_696# a_45476_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3084 VDD a_40400_n11559# a_40348_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3085 a_47551_n11370# a_46676_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3086 a_31676_n11788# a_30908_n11533# a_29690_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3087 a_29559_7009# a_29557_5953# a_29860_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3088 a_44057_690# C[119] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3089 a_44964_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3090 VDD a_25296_n11559# a_25514_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3091 a_33335_7009# a_32567_6434# a_31349_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3092 VSS C[22] a_17515_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3093 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3094 VDD a_818_1932# a_12918_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3095 a_27291_836# a_27065_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3096 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3097 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3098 VDD a_31335_773# a_32260_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3099 a_44890_n10732# a_44124_n11533# a_44794_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X3100 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3101 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3102 a_40789_5953# a_40119_6434# a_40389_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3103 a_21993_1829# a_21401_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3104 VDD a_529_6408# a_747_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3105 a_48433_7009# a_47717_6408# a_46447_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3106 a_14310_n5879# a_14084_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3107 VDD a_45829_6408# a_45777_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3108 a_17718_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3109 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3110 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3111 VDD a_1047_n6869# a_3707_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3112 a_33564_n11788# a_32796_n11533# a_31578_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X3113 a_48662_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3114 a_3346_n5622# a_2756_n5789# a_3250_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3115 a_22005_5953# a_21239_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3116 a_53985_773# a_55605_836# a_55429_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3117 a_40281_690# C[117] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3118 a_41004_n5622# a_42624_n5879# a_42448_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3119 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3120 a_20119_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3121 a_38999_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3122 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3123 VDD a_27184_n11559# a_27402_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3124 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3125 a_44661_5953# a_43895_6434# a_44565_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3126 a_48111_n6843# a_48106_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X3127 a_59381_836# a_59155_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3128 a_56198_n5622# a_55834_n5879# a_56102_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3129 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3130 VDD a_818_1932# a_12104_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3131 VSS a_1047_n6869# a_4699_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3132 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3133 a_6909_7009# a_6193_6408# a_4923_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3134 VSS a_23397_6449# a_23370_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3135 a_41232_1994# a_40873_1829# a_40871_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3136 a_18444_n5622# a_18446_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3137 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3138 a_31447_7009# a_31445_5953# a_31748_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3139 a_55434_1994# a_55429_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3140 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3141 VDD a_3250_n5622# a_4175_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3142 a_8781_773# a_8417_836# a_8685_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3143 a_35452_n11788# a_34684_n11533# a_33466_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X3144 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3145 a_1362_n5622# a_1094_n5879# a_923_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X3146 a_46447_5953# a_47717_6408# a_47908_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3147 a_45434_6655# a_44565_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3148 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3149 VSS a_40775_773# a_41700_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3150 VDD a_38117_n11370# a_38067_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3151 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3152 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3153 a_23895_7009# a_23127_6434# a_21909_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3154 a_17326_696# a_17156_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3155 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3156 VSS a_34954_n11298# a_34927_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3157 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3158 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3159 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3160 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3161 VSS a_46347_n6869# a_56198_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X3162 a_37324_n5622# a_37326_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3163 VSS C[13] a_34507_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3164 a_31674_n10732# a_30908_n11533# a_31578_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3165 a_6004_696# a_5834_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3166 a_48053_836# a_47827_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3167 a_6532_n5789# C[35] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3168 a_37340_n11788# a_36572_n11533# a_35354_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X3169 a_4923_5953# a_6193_6408# a_6384_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3170 a_28883_n5795# a_28713_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3171 VDD a_6422_n11559# a_6640_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3172 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3173 a_59649_773# a_59045_6408# a_59263_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3174 a_60062_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3175 a_20348_n11788# a_19580_n11533# a_18362_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3176 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3177 a_55969_773# a_55379_690# a_55873_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3178 a_29774_n6678# a_29182_n5789# a_27788_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3179 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3180 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3181 a_19594_5708# a_19621_6449# a_19606_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3182 a_6139_2600# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3183 VSS a_44165_6449# a_44138_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3184 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3185 VSS C[86] a_17744_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3186 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3187 a_48734_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3188 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3189 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3190 VSS C[28] a_6193_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3191 VDD a_15916_1932# a_16688_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3192 a_22222_n6678# a_21856_n5879# a_20236_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3193 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3194 a_12559_1829# a_12193_836# a_10573_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3195 a_31792_1994# a_31433_1829# a_31431_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3196 a_31335_773# a_31067_836# a_30896_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3197 a_48335_5953# a_49605_6408# a_49796_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3198 a_7040_n10732# a_8310_n11559# a_8501_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3199 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3200 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3201 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3202 a_33562_n10732# a_32796_n11533# a_33466_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3203 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3204 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3205 VDD a_54874_6655# a_54824_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3206 a_8685_773# a_8191_690# a_8246_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3207 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3208 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3209 VDD a_8310_n11559# a_8528_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3210 a_22236_n11788# a_21468_n11533# a_20250_n10732# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X3211 VDD C[20] a_21291_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3212 a_38997_5953# a_38283_6408# a_38901_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3213 VSS a_40389_6449# a_40362_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3214 a_25900_n5622# a_27520_n5879# a_27344_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3215 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3216 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3217 a_22236_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3218 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3219 a_48431_5953# a_47665_6434# a_48335_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3220 a_25998_n6678# a_25406_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3221 a_47757_n5795# a_47587_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3222 VDD a_15856_n11559# a_16074_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3223 a_34927_n10487# a_34954_n11298# a_34939_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3224 a_41102_n6678# a_40736_n5879# a_39116_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3225 a_42990_n6678# a_42624_n5879# a_41004_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3226 VDD C[66] a_55498_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3227 VSS a_21738_n11298# a_21711_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3228 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3229 a_41018_n10732# a_42288_n11559# a_42479_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3230 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3231 a_40887_7009# a_40119_6434# a_38901_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3232 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3233 a_37228_n5622# a_38848_n5879# a_38672_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3234 a_35450_n10732# a_34684_n11533# a_35354_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3235 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3236 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3237 a_20007_773# a_19739_836# a_19568_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3238 a_50622_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3239 a_39214_n6678# a_38622_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3240 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3241 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3242 a_7122_n5622# a_6532_n5789# a_7026_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3243 VDD a_6529_836# a_6353_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3244 a_55873_773# a_55605_836# a_55434_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3245 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3246 a_31564_n5622# a_32958_n5789# a_33008_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3247 a_24124_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X3248 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3249 a_6396_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3250 a_44878_n6678# a_44286_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3251 VDD a_17744_n11559# a_17962_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3252 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3253 a_29034_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3254 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3255 a_1458_n5622# a_1094_n5879# a_1362_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3256 VSS a_23626_n11298# a_23599_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3257 a_23783_773# a_23289_690# a_23344_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3258 a_39116_n5622# a_40510_n5789# a_40560_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3259 a_42906_n10732# a_44176_n11559# a_44367_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3260 VDD C[65] a_57386_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3261 a_1472_n10732# a_706_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3262 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3263 VSS a_23179_6408# a_23127_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3264 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3265 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3266 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3267 a_8417_836# a_8191_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3268 a_50307_1829# a_49715_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3269 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3270 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3271 a_20346_n10732# a_19580_n11533# a_20250_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3272 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3273 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3274 VDD a_31020_1932# a_33680_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3275 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3276 VSS a_30949_6449# a_30922_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3277 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3278 a_59155_690# C[127] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3279 a_26012_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3280 a_50548_n10732# a_49782_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3281 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3282 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3283 a_53999_5953# a_55269_6408# a_55460_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3284 VDD a_46433_773# a_47358_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3285 a_41018_n10732# a_40400_n11559# a_40618_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3286 VSS a_15916_1932# a_17680_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3287 VSS a_25514_n11298# a_25487_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3288 a_21711_n10487# a_21738_n11298# a_21723_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3289 VDD a_13350_6655# a_13300_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3290 a_37888_6655# a_37013_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3291 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3292 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3293 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3294 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3295 a_50851_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3296 a_54095_5953# a_53381_6408# a_53999_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3297 VDD a_21627_836# a_21451_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3298 a_52422_n5622# a_52424_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3299 a_22234_n10732# a_21468_n11533# a_22138_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3300 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3301 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3302 a_29676_n5622# a_29408_n5879# a_29237_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X3303 a_15966_n5789# C[40] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3304 a_16460_n5622# a_15966_n5789# a_16021_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3305 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3306 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3307 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3308 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3309 a_52209_7009# a_52207_5953# a_52510_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3310 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3311 a_8928_n10732# a_10146_n11533# a_10389_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3312 a_52436_n10732# a_51670_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3313 a_1243_5953# a_477_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3314 a_19594_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3315 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3316 a_22124_n5622# a_21630_n5789# a_21685_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3317 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3318 a_23515_836# a_23289_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3319 a_24012_n5622# a_23518_n5789# a_23573_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3320 a_42906_n10732# a_42288_n11559# a_42506_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3321 a_23599_n10487# a_23626_n11298# a_23611_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3322 a_50319_5953# a_49605_6408# a_50223_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3323 VDD a_18119_773# a_19044_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3324 a_18133_5953# a_19351_6434# a_19594_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3325 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3326 a_27886_n6678# a_27520_n5879# a_25900_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3327 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3328 a_8272_5708# a_8299_6449# a_8284_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3329 a_31431_773# a_30841_690# a_31335_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3330 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3331 a_14461_7009# a_13745_6408# a_12475_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3332 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3333 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3334 VDD a_11857_6408# a_11805_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3335 a_33223_773# a_34843_836# a_34667_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3336 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3337 VSS a_55873_773# a_56798_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3338 a_34846_n5789# C[50] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3339 a_35340_n5622# a_34846_n5789# a_34901_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3340 VSS a_2635_6449# a_2608_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3341 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3342 VSS a_31020_1932# a_38448_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3343 VDD a_6797_773# a_7722_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3344 VSS a_4752_n11298# a_4725_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3345 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3346 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3347 a_37097_1829# a_36731_836# a_35111_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3348 a_54324_n10732# a_53558_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3349 VSS a_37888_6655# a_37838_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3350 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3351 a_21856_n5879# a_21630_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3352 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3353 a_11967_690# C[102] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3354 a_42892_n5622# a_42398_n5789# a_42453_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3355 a_44794_n10732# a_44176_n11559# a_44394_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3356 a_25487_n10487# a_25514_n11298# a_25499_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3357 a_4116_696# a_3946_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3358 VSS a_56102_n5622# a_57027_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3359 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3360 a_9574_6655# a_8699_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3361 VSS a_57990_n5622# a_58915_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3362 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3363 a_55983_5953# a_55217_6434# a_55887_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3364 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3365 VDD C[71] a_46058_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3366 a_31578_n10732# a_32848_n11559# a_33039_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3367 a_7138_n11788# a_6370_n11533# a_5152_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3368 a_54081_773# a_53491_690# a_53985_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3369 a_52326_n5622# a_53946_n5879# a_53770_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3370 a_7138_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3371 VSS a_31020_1932# a_34672_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3372 a_33184_n5879# a_32958_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3373 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3374 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3375 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3376 VDD a_15916_1932# a_23426_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3377 VDD a_26789_n11370# a_26739_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3378 a_29786_n10732# a_29020_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3379 a_12475_5953# a_13745_6408# a_13936_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3380 a_52554_1994# a_52195_1829# a_52193_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3381 a_11462_6655# a_10587_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3382 a_54312_n6678# a_53720_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3383 VSS a_6640_n11298# a_6613_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3384 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3385 a_52986_6655# a_52111_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3386 a_56212_n10732# a_55446_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3387 a_40736_n5879# a_40510_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3388 a_41893_n11370# a_41018_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3389 a_59976_n6678# a_59384_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3390 VDD a_1047_n6869# a_6669_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3391 a_27573_5953# a_28791_6434# a_29034_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3392 a_59759_5953# a_59045_6408# a_59649_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3393 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3394 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3395 a_34617_690# C[114] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3396 VDD a_17120_6655# a_17070_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3397 VDD C[70] a_47946_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3398 a_33466_n10732# a_34736_n11559# a_34927_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3399 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3400 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3401 a_17851_836# a_17625_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3402 a_23879_773# a_23515_836# a_23783_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3403 a_36586_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3404 VDD a_21895_773# a_22820_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3405 a_9026_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3406 a_53717_836# a_53491_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3407 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3408 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3409 VSS a_8528_n11298# a_8501_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3410 a_4725_n10487# a_4752_n11298# a_4737_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3411 a_10816_n10732# a_10146_n11533# a_10416_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3412 a_14762_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3413 a_21767_n6843# a_21680_n6611# a_21685_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3414 a_43781_n11370# a_42906_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3415 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3416 a_3117_773# a_3119_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3417 a_29772_n5622# a_29408_n5879# a_29676_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3418 VSS a_46118_1932# a_50305_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3419 a_5248_n10732# a_4482_n11533# a_5152_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3420 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3421 VDD a_46118_1932# a_58218_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3422 a_40211_n5795# a_40041_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3423 a_31578_n10732# a_30960_n11559# a_31178_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3424 VSS a_16074_n11298# a_16047_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3425 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3426 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3427 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3428 a_35354_n10732# a_36624_n11559# a_36815_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3429 a_1133_773# a_2753_836# a_2577_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3430 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3431 a_50319_5953# a_49553_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3432 a_10587_5953# a_9917_6434# a_10187_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3433 a_46529_773# a_46165_836# a_46433_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3434 a_49941_836# a_49715_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3435 a_56198_n5622# a_56200_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3436 a_18231_7009# a_17515_6408# a_16245_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3437 VDD a_15627_6408# a_15575_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3438 VSS a_16145_n6869# a_16556_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3439 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3440 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3441 a_47757_n5795# a_47587_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3442 a_16570_n10732# a_15804_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3443 a_6613_n10487# a_6640_n11298# a_6625_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3444 a_6797_773# a_6529_836# a_6358_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3445 VSS a_5798_6655# a_5748_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3446 a_48648_n6678# a_48056_n5789# a_46662_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3447 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3448 VSS a_30731_6408# a_30679_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3449 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3450 a_40647_n6843# a_40560_n6611# a_40565_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3451 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3452 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3453 VSS a_51711_6449# a_51684_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3454 a_27788_n5622# a_27294_n5789# a_27349_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3455 a_7136_n10732# a_6370_n11533# a_7040_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3456 a_16873_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3457 a_33466_n10732# a_32848_n11559# a_33066_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3458 a_4909_773# a_6303_690# a_6353_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3459 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3460 a_54312_n6678# a_53720_n5789# a_52326_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3461 a_37242_n10732# a_38512_n11559# a_38703_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3462 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3463 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3464 a_11030_1994# a_10671_1829# a_10669_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3465 VSS a_59492_n11298# a_59465_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3466 a_8272_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3467 a_25232_1994# a_25227_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3468 VSS a_31249_n6869# a_35436_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3469 VDD a_34112_6655# a_34062_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3470 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3471 VDD a_28843_6408# a_29061_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3472 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3473 a_45646_696# a_45476_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3474 VDD a_15461_n11370# a_15411_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3475 a_18458_n10732# a_17692_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3476 a_8501_n10487# a_8528_n11298# a_8513_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3477 a_16245_5953# a_17515_6408# a_17706_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3478 a_15232_6655# a_14363_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3479 a_1819_n6843# a_1460_n6678# a_1458_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3480 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3481 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3482 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3483 a_15963_836# a_15737_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3484 VSS a_818_1932# a_694_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3485 VSS a_1362_n5622# a_2287_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3486 a_30565_n11370# a_29690_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3487 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3488 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3489 a_35354_n10732# a_34736_n11559# a_34954_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3490 a_18761_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3491 a_16047_n10487# a_16074_n11298# a_16059_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3492 VDD a_36395_6408# a_36343_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3493 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3494 VSS a_33562_n10732# a_33564_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3495 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3496 a_21456_1994# a_21451_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3497 VSS a_31335_773# a_32260_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3498 a_59759_5953# a_58993_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3499 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3500 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3501 a_21895_773# a_21627_836# a_21456_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3502 VSS a_23893_5953# a_23895_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3503 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3504 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3505 a_19513_690# C[106] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3506 a_29461_5953# a_28843_6408# a_29061_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3507 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3508 VDD a_2982_n5879# a_2806_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3509 VDD a_17349_n11370# a_17299_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3510 a_18229_5953# a_17463_6434# a_18133_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3511 a_55379_690# C[125] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3512 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3513 a_19443_n5795# a_19273_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3514 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3515 a_35223_7009# a_34507_6408# a_33237_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3516 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3517 VDD a_32619_6408# a_32567_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3518 a_18532_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3519 a_32453_n11370# a_31578_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3520 a_40775_773# a_42395_836# a_42219_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3521 a_37242_n10732# a_36624_n11559# a_36842_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3522 VSS a_46118_1932# a_59210_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3523 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3524 a_25107_n5795# a_24937_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3525 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3526 a_46529_773# a_45939_690# a_46433_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3527 a_26995_n5795# a_26825_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3528 a_59465_n10487# a_59492_n11298# a_59477_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3529 a_36000_6655# a_35125_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3530 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3531 a_11668_696# a_11498_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3532 VDD a_24672_6655# a_24622_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3533 VSS a_58650_6655# a_58600_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3534 VDD a_46347_n6869# a_49007_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3535 VDD a_19403_6408# a_19621_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3536 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3537 a_10079_690# C[101] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3538 VSS a_10187_6449# a_10160_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3539 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3540 a_42224_1994# a_42219_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3541 a_55969_773# a_55971_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3542 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3543 a_10802_n5622# a_12196_n5789# a_12246_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3544 a_34341_n11370# a_33466_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3545 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3546 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3547 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3548 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3549 a_56198_n5622# a_55608_n5789# a_56102_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3550 a_39130_n10732# a_38512_n11559# a_38730_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3551 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3552 a_32224_6655# a_31349_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3553 a_29179_836# a_28953_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3554 a_33564_n11788# a_33562_n10732# a_33865_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X3555 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3556 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3557 VDD a_8081_6408# a_8029_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3558 a_45875_n5795# a_45705_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3559 a_22138_n10732# a_21520_n11559# a_21738_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3560 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3561 a_10685_7009# a_9917_6434# a_8699_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3562 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3563 a_34318_696# a_34148_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3564 a_20021_5953# a_19403_6408# a_19621_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3565 a_20420_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3566 a_39300_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3567 a_59990_n11788# a_59222_n11533# a_58004_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3568 VSS a_46347_n6869# a_57551_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3569 VDD C[5] a_49605_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3570 a_25783_7009# a_25067_6408# a_23797_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3571 a_48550_n5622# a_48282_n5879# a_48111_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3572 VDD a_51722_n11559# a_51670_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3573 a_57348_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3574 VDD a_56102_n5622# a_57027_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3575 VDD a_57990_n5622# a_58915_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3576 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3577 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3578 VDD a_4305_6408# a_4253_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3579 a_49715_690# C[122] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3580 a_6893_773# a_6303_690# a_6797_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3581 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3582 a_57761_773# a_59155_690# a_59205_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3583 a_48419_1829# a_48053_836# a_46433_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3584 a_46433_773# a_46165_836# a_45994_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3585 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3586 a_6811_5953# a_8029_6434# a_8272_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3587 VSS a_31249_n6869# a_39212_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3588 a_4641_836# a_4415_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3589 a_40591_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3590 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3591 a_31660_n5622# a_31662_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3592 VDD a_53610_n11559# a_53558_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3593 a_31349_5953# a_30679_6434# a_30949_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3594 a_46529_773# a_46531_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3595 VDD a_41664_6655# a_41614_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3596 a_59384_n5789# C[63] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3597 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3598 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3599 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3600 a_23797_5953# a_25067_6408# a_25258_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3601 a_22784_6655# a_21909_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3602 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3603 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3604 a_50223_5953# a_51441_6434# a_51684_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3605 a_44551_773# a_46165_836# a_45989_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3606 a_14447_1829# a_13855_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3607 VDD a_16145_n6869# a_21767_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3608 a_21125_n11370# a_20250_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3609 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3610 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3611 a_3910_6655# a_3035_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3612 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3613 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3614 a_59521_n6843# a_59434_n6611# a_59439_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3615 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3616 a_21991_773# a_21401_690# a_21895_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3617 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3618 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3619 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3620 a_46774_n11788# a_46006_n11533# a_44794_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3621 a_47908_5708# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3622 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3623 a_12196_n5789# C[38] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3624 a_40211_n5795# a_40041_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3625 a_22007_7009# a_22005_5953# a_22308_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3626 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3627 a_37013_5953# a_36395_6408# a_36613_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3628 a_45994_1994# a_45989_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3629 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3630 a_923_n6843# a_918_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3631 a_37097_1829# a_36505_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3632 a_23013_n11370# a_22138_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3633 a_20117_5953# a_19403_6408# a_20021_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3634 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3635 VSS a_10912_n10732# a_10914_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3636 VDD a_57157_6408# a_57105_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3637 a_1231_1829# a_639_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3638 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3639 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3640 a_31564_n5622# a_33184_n5879# a_33008_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3641 a_48662_n11788# a_47894_n11533# a_46676_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X3642 a_21909_5953# a_21239_6434# a_21509_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3643 a_12422_n5879# a_12196_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3644 a_3035_5953# a_2365_6434# a_2635_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3645 a_8783_1829# a_8191_690# a_6797_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3646 VDD a_8081_6408# a_8299_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3647 a_1458_n5622# a_868_n5789# a_1362_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3648 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3649 a_39116_n5622# a_40736_n5879# a_40560_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3650 VSS a_46433_773# a_47358_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3651 a_48646_n5622# a_48282_n5879# a_48550_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3652 a_17935_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3653 a_25781_5953# a_25015_6434# a_25685_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3654 a_60973_n5795# a_60803_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3655 a_46223_n6843# a_46218_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X3656 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3657 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3658 a_40789_5953# a_42059_6408# a_42250_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3659 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3660 VSS a_1047_n6869# a_923_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3661 VSS a_12800_n10732# a_12802_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3662 VSS a_1047_n6869# a_2811_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3663 a_7026_n5622# a_8420_n5789# a_8470_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3664 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3665 VDD a_15856_n11559# a_15804_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3666 a_39529_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3667 a_22352_1994# a_21993_1829# a_21991_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3668 a_16556_n5622# a_16558_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3669 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3670 a_6303_690# C[99] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3671 VDD a_1362_n5622# a_2287_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3672 VSS a_3131_5953# a_3133_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3673 VSS a_31020_1932# a_38983_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3674 a_35223_7009# a_34455_6434# a_33237_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3675 VDD a_45434_6655# a_45384_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3676 VSS a_32848_n11559# a_32796_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3677 a_29557_5953# a_28843_6408# a_29461_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3678 VSS a_18119_773# a_19044_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3679 a_26766_696# a_26596_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3680 a_27884_n5622# a_27886_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3681 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3682 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3683 VSS a_14688_n10732# a_14690_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3684 a_10914_n11788# a_10912_n10732# a_11215_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3685 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3686 a_19443_n5795# a_19273_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3687 a_25177_690# C[109] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3688 VDD a_17744_n11559# a_17692_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3689 a_46772_n10732# a_46006_n11533# a_46676_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3690 a_35436_n5622# a_35438_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3691 a_31151_n10487# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3692 VSS a_46347_n6869# a_54310_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3693 a_31447_7009# a_30679_6434# a_29461_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3694 a_52111_5953# a_51493_6408# a_51711_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3695 VDD a_31249_n6869# a_43349_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3696 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3697 VSS C[23] a_15627_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3698 VSS a_6797_773# a_7722_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3699 a_12333_n6843# a_12246_n6611# a_12251_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3700 a_4139_n11370# a_3264_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3701 a_4644_n5789# C[34] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3702 a_25107_n5795# a_24937_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3703 a_26995_n5795# a_26825_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3704 a_38983_773# a_38619_836# a_38887_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3705 VSS a_34736_n11559# a_34684_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3706 VSS a_46347_n6869# a_59974_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3707 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3708 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3709 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3710 a_27886_n6678# a_27294_n5789# a_25900_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3711 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3712 a_4781_n6843# a_4694_n6611# a_4699_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3713 a_43120_1994# a_42761_1829# a_42759_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3714 a_49416_696# a_49246_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3715 VSS a_363_n11370# a_313_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3716 a_20117_5953# a_19351_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3717 a_52097_773# a_53717_836# a_53541_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3718 a_12802_n11788# a_12800_n10732# a_13103_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3719 a_38997_5953# a_38231_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3720 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3721 a_21401_690# C[107] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3722 a_21630_n5789# C[43] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3723 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3724 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3725 VDD a_19632_n11559# a_19580_n11533# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3726 a_48660_n10732# a_47894_n11533# a_48564_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3727 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3728 a_42773_5953# a_42007_6434# a_42677_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3729 a_16460_n5622# a_18080_n5879# a_17904_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3730 a_39214_n6678# a_38622_n5789# a_37228_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3731 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3732 a_55971_1829# a_55605_836# a_53985_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3733 a_6027_n11370# a_5152_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3734 a_4870_n5879# a_4644_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3735 a_45875_n5795# a_45705_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3736 VSS a_24901_n11370# a_24851_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3737 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3738 VDD a_818_1932# a_10216_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3739 VSS a_36624_n11559# a_36572_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3740 a_18446_n6678# a_17854_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3741 VSS a_21509_6449# a_21482_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3742 a_33550_n6678# a_33184_n5879# a_31564_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3743 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3744 a_24012_n5622# a_25632_n5879# a_25456_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3745 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3746 a_53546_1994# a_53541_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3747 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3748 VSS C[12] a_36395_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3749 a_56116_n10732# a_57386_n11559# a_57577_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3750 a_14690_n11788# a_14688_n10732# a_14991_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3751 a_44565_5953# a_45829_6408# a_46020_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3752 VSS a_21895_773# a_22820_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3753 VDD C[16] a_28843_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3754 a_28448_6655# a_27573_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3755 a_15830_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3756 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3757 VDD a_12193_836# a_12017_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3758 a_22007_7009# a_21239_6434# a_20021_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3759 VSS a_818_1932# a_6893_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3760 a_35340_n5622# a_36960_n5879# a_36784_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3761 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3762 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3763 a_3133_7009# a_2365_6434# a_1147_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3764 a_7915_n11370# a_7040_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3765 a_44892_n11788# a_44176_n11559# a_42906_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3766 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3767 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3768 a_1133_773# a_639_690# a_694_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3769 a_38887_773# a_38393_690# a_38448_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3770 VSS a_38512_n11559# a_38460_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3771 a_29545_1829# a_28953_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3772 a_37326_n6678# a_36734_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3773 VSS a_11691_n11370# a_11641_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3774 a_24124_n11788# a_23356_n11533# a_22138_n10732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3775 a_40885_5953# a_40119_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3776 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3777 a_42892_n5622# a_44512_n5879# a_44336_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3778 a_29676_n5622# a_31070_n5789# a_31120_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3779 VSS C[14] a_32619_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3780 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3781 a_14081_836# a_13855_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3782 a_20103_773# a_19513_690# a_20007_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3783 a_8646_n5879# a_8420_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3784 a_42990_n6678# a_42398_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3785 a_3035_5953# a_4305_6408# a_4496_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3786 a_29557_5953# a_28791_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3787 a_58004_n10732# a_59274_n11559# a_59465_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3788 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3789 a_57775_5953# a_57157_6408# a_57375_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3790 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3791 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3792 VDD a_46347_n6869# a_59521_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3793 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3794 a_8797_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3795 VDD a_31020_1932# a_45008_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3796 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3797 a_25767_773# a_25769_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3798 a_46846_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3799 VDD a_16145_n6869# a_28245_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3800 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3801 a_51603_690# C[123] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3802 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3803 VSS a_13579_n11370# a_13529_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3804 VDD a_36731_836# a_36555_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X3805 VSS a_23408_n11559# a_23356_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3806 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3807 VSS a_15916_1932# a_29008_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3808 VDD a_52986_6655# a_52936_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3809 a_19739_836# a_19513_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3810 a_22220_n5622# a_21856_n5879# a_22124_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3811 VDD C[21] a_19403_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3812 VSS a_16145_n6869# a_29237_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3813 VSS a_28448_6655# a_28398_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3814 VDD C[11] a_38283_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X3815 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3816 a_8121_n5795# a_7951_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3817 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3818 a_46543_5953# a_45777_6434# a_46447_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3819 a_43002_n10732# a_42288_n11559# a_42906_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3820 a_50534_n5622# a_50536_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3821 a_27671_7009# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3822 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3823 a_38619_836# a_38393_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3824 a_12022_1994# a_12017_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3825 a_27788_n5622# a_27520_n5879# a_27349_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3826 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3827 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3828 VSS C[29] a_4305_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3829 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3830 VDD a_59381_836# a_59205_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3831 a_18446_n6678# a_18080_n5879# a_16460_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3832 a_24026_n10732# a_25244_n11533# a_25487_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3833 a_8557_n6843# a_8470_n6611# a_8475_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3834 VSS a_10198_n11559# a_10146_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3835 a_58004_n10732# a_57386_n11559# a_57604_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3836 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3837 a_41100_n5622# a_40736_n5879# a_41004_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3838 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3839 a_44794_n10732# a_46058_n11559# a_46249_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3840 VSS a_7915_n11370# a_7865_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3841 VSS a_134_6655# a_84_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3842 a_14445_773# a_14081_836# a_14349_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3843 a_39116_n5622# a_38848_n5879# a_38677_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3844 a_25998_n6678# a_25632_n5879# a_24012_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3845 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3846 a_4508_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3847 a_59761_7009# a_59759_5953# a_60062_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3848 a_44283_836# a_44057_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3849 a_44890_n10732# a_44176_n11559# a_44794_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3850 a_47119_n6843# a_46760_n6678# a_46758_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X3851 a_49007_n6843# a_48648_n6678# a_48646_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3852 a_27146_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3853 a_24122_n10732# a_23356_n11533# a_24026_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3854 VSS a_10683_5953# a_10685_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3855 a_32958_n5789# C[49] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3856 a_1590_1994# a_1231_1829# a_1229_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3857 a_33452_n5622# a_32958_n5789# a_33013_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3858 a_60973_n5795# a_60803_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3859 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3860 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3861 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3862 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3863 a_38622_n5789# C[52] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3864 VSS a_48550_n5622# a_49475_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3865 a_18217_1829# a_17851_836# a_16231_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3866 VSS a_12086_n11559# a_12034_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3867 a_59878_n5622# a_59274_n11559# a_59492_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3868 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3869 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3870 VDD a_31020_1932# a_31792_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3871 a_10816_n10732# a_12034_n11533# a_12277_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3872 a_41004_n5622# a_40510_n5789# a_40565_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3873 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3874 a_8795_5953# a_8081_6408# a_8699_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3875 VSS a_9803_n11370# a_9753_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3876 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3877 a_11668_696# a_11498_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3878 a_44878_n6678# a_44512_n5879# a_42892_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3879 a_46676_n10732# a_47946_n11559# a_48137_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3880 a_37095_773# a_36731_836# a_36999_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3881 a_13579_n11370# a_12704_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3882 VSS a_46047_6449# a_46020_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3883 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3884 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3885 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3886 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3887 VSS a_15916_1932# a_15792_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3888 a_50438_n5622# a_52058_n5879# a_51882_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3889 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3890 VDD a_11462_6655# a_11412_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3891 a_31296_n5879# a_31070_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X3892 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3893 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3894 a_35452_n11788# a_34736_n11559# a_33466_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3895 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3896 a_52424_n6678# a_51832_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3897 a_44663_7009# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3898 a_52207_5953# a_51493_6408# a_52111_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3899 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3900 VDD a_36999_773# a_37924_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3901 VDD a_57722_n5879# a_57546_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3902 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3903 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3904 a_12704_n10732# a_13922_n11533# a_14165_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3905 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3906 VDD a_1047_n6869# a_4781_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3907 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3908 a_14349_773# a_13855_690# a_13910_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3909 a_14690_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3910 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3911 a_50321_7009# a_50319_5953# a_50622_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3912 a_34318_696# a_34148_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3913 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3914 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3915 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3916 VSS C[1] a_57157_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X3917 a_17706_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3918 a_37340_n11788# a_36624_n11559# a_35354_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3919 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3920 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3921 a_6384_5708# a_6411_6449# a_6396_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X3922 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3923 a_25914_n10732# a_25244_n11533# a_25514_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3924 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3925 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3926 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3927 a_12573_7009# a_11857_6408# a_10587_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3928 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3929 a_10401_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3930 a_44138_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3931 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3932 VDD a_818_1932# a_3478_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3933 a_38530_1994# a_38443_1896# a_38448_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3934 a_39212_n5622# a_38622_n5789# a_39116_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3935 a_46676_n10732# a_46058_n11559# a_46276_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3936 a_27884_n5622# a_27520_n5879# a_27788_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3937 VSS a_31020_1932# a_36560_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3938 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3939 VDD a_46347_n6869# a_56559_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3940 a_35209_1829# a_34843_836# a_33223_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3941 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3942 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3943 a_2849_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3944 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3945 a_7040_n10732# a_8258_n11533# a_8501_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3946 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3947 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3948 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3949 a_40871_773# a_40507_836# a_40775_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3950 a_33562_n10732# a_32848_n11559# a_33466_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3951 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3952 a_7686_6655# a_6811_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3953 a_19968_n5879# a_19742_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3954 a_39228_n11788# a_38512_n11559# a_37242_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X3955 a_18348_n5622# a_17854_n5789# a_17909_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3956 a_12704_n10732# a_12034_n11533# a_12304_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3957 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3958 a_33319_773# a_33321_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3959 a_51304_696# a_51134_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3960 a_46760_n6678# a_46168_n5789# a_44780_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X3961 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3962 a_48564_n10732# a_47946_n11559# a_48164_n11298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3963 a_10587_5953# a_11857_6408# a_12048_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3964 a_720_5708# a_747_6449# a_732_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3965 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3966 a_50666_1994# a_50307_1829# a_50305_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3967 VSS a_16145_n6869# a_25996_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3968 a_31335_773# a_32955_836# a_32779_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X3969 a_44341_n6843# a_44336_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3970 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3971 a_51098_6655# a_50223_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X3972 a_57360_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X3973 a_54214_n5622# a_53946_n5879# a_53775_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3974 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3975 a_4737_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3976 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3977 a_57871_5953# a_57157_6408# a_57775_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3978 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3979 VSS a_31249_n6869# a_31660_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3980 VSS a_31249_n6869# a_33548_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3981 a_35450_n10732# a_34736_n11559# a_35354_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X3982 VSS a_49210_6655# a_49160_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X3983 a_59761_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3984 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3985 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3986 VDD a_15232_6655# a_15182_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X3987 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3988 a_34698_5708# a_30830_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3989 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3990 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3991 a_36999_773# a_36731_836# a_36560_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3992 a_45663_n11370# a_44794_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X3993 a_53720_n5789# C[60] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X3994 a_35111_773# a_36505_690# a_36555_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3995 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3996 VSS a_818_1932# a_8246_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3997 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3998 a_12874_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3999 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4000 a_40775_773# a_40281_690# a_40336_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4001 a_37338_n10732# a_36624_n11559# a_37242_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4002 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4003 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4004 a_31433_1829# a_30841_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4005 VSS a_59988_n10732# a_59990_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4006 VDD a_46118_1932# a_56330_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4007 VDD a_1094_n5879# a_918_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4008 a_8121_n5795# a_7951_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4009 a_16343_7009# a_15627_6408# a_14363_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4010 a_17555_n5795# a_17385_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4011 a_47551_n11370# a_46676_n10732# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4012 VSS a_818_1932# a_4470_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4013 a_776_1994# a_689_1896# a_694_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4014 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4015 a_21895_773# a_23515_836# a_23339_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4016 a_29543_773# a_29179_836# a_29447_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X4017 a_47920_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4018 a_23219_n5795# a_23049_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4019 VSS a_3910_6655# a_3860_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4020 VSS a_35450_n10732# a_35452_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4021 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4022 a_8928_n10732# a_8258_n11533# a_8528_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4023 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4024 a_12571_5953# a_11805_6434# a_12475_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4025 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4026 a_50321_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4027 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4028 VDD a_12461_773# a_13386_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4029 a_51913_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4030 a_39226_n10732# a_38512_n11559# a_39130_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4031 a_54083_1829# a_53491_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4032 VDD C[75] a_38512_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4033 a_48646_n5622# a_48056_n5789# a_48550_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4034 a_31020_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4035 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4036 a_6384_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4037 a_36435_n5795# a_36265_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4038 a_23344_1994# a_23339_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4039 VDD a_32224_6655# a_32174_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4040 a_26766_696# a_26596_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4041 a_54310_n5622# a_53720_n5789# a_54214_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4042 a_8914_n5622# a_10308_n5789# a_10358_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4043 a_14363_5953# a_15627_6408# a_15818_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4044 a_42099_n5795# a_41929_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4045 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4046 a_43987_n5795# a_43817_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4047 a_29237_n6843# a_29232_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4048 VSS a_46347_n6869# a_48111_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4049 VSS a_37338_n10732# a_37340_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4050 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4051 a_40507_836# a_40281_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4052 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4053 VDD a_35111_773# a_36036_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4054 VDD a_48550_n5622# a_49475_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4055 a_53801_n10487# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4056 a_37111_7009# a_36395_6408# a_35125_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4057 a_12557_773# a_11967_690# a_12461_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4058 a_59990_n11788# a_59988_n10732# a_60291_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X4059 VSS a_16145_n6869# a_18444_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4060 a_24122_n10732# a_23408_n11559# a_24026_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4061 VSS a_46347_n6869# a_55663_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4062 a_14461_7009# a_14459_5953# a_14762_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4063 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4064 a_46662_n5622# a_46394_n5879# a_46223_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4065 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4066 a_29447_773# a_28953_690# a_29008_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4067 VSS a_38117_n11370# a_38067_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4068 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4069 a_27573_5953# a_26955_6408# a_27173_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4070 a_49416_696# a_49246_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4071 a_44379_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4072 VSS a_39226_n10732# a_39228_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4073 a_35452_n11788# a_35450_n10732# a_35753_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X4074 a_22220_n5622# a_22222_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4075 VSS a_13714_3465# a_36570_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4076 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4077 a_720_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4078 a_16644_5388# a_15726_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4079 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4080 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4081 VSS a_22234_n10732# a_22236_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4082 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4083 a_49796_5708# a_49823_6449# a_49808_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X4084 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4085 a_38887_773# a_40507_836# a_40331_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4086 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4087 VSS a_46118_1932# a_57322_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4088 a_35207_773# a_34617_690# a_35111_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4089 VSS a_31249_n6869# a_37324_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4090 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4091 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4092 VSS a_56762_6655# a_56712_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4093 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4094 a_42761_1829# a_42395_836# a_40775_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4095 a_31249_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4096 VDD a_22784_6655# a_22734_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4097 a_57496_n5789# C[62] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4098 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4099 a_37340_n11788# a_37338_n10732# a_37641_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4100 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4101 a_40336_1994# a_40331_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4102 a_41100_n5622# a_41102_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4103 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4104 a_54081_773# a_54083_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4105 VDD a_27291_836# a_27115_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X4106 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4107 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4108 a_16341_5953# a_15575_6434# a_16245_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4109 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4110 VSS a_24122_n10732# a_24124_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4111 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4112 a_12461_773# a_12193_836# a_12022_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4113 a_31349_5953# a_32619_6408# a_32810_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4114 a_30336_6655# a_29461_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4115 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4116 VDD a_6193_6408# a_6141_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4117 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4118 a_34843_836# a_34617_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4119 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4120 VSS a_36570_n7315# a_31249_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4121 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4122 a_10308_n5789# C[37] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4123 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4124 a_12690_n5622# a_12196_n5789# a_12251_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4125 a_57722_n5879# a_57496_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4126 a_37412_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4127 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4128 VSS a_27788_n5622# a_28713_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4129 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4130 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4131 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4132 a_39228_n11788# a_39226_n10732# a_39529_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4133 a_5021_7009# a_4305_6408# a_3035_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4134 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4135 a_49852_1994# a_49765_1896# a_49770_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4136 a_22124_n5622# a_23744_n5879# a_23568_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4137 a_39573_n6843# a_39214_n6678# a_39212_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4138 VDD a_2417_6408# a_2365_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4139 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4140 VSS a_26010_n10732# a_26012_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4141 a_22236_n11788# a_22234_n10732# a_22537_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4142 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4143 a_7124_n6678# a_6758_n5879# a_5138_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4144 a_44565_5953# a_43947_6408# a_44165_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4145 a_35111_773# a_34843_836# a_34672_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4146 a_9012_n6678# a_8646_n5879# a_7026_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4147 a_55873_773# a_57267_690# a_57317_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4148 a_2527_690# C[97] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4149 a_29676_n5622# a_31296_n5879# a_31120_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4150 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4151 a_4923_5953# a_6141_6434# a_6384_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4152 a_33636_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4153 a_10534_n5879# a_10308_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4154 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4155 a_31249_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4156 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4157 a_29774_n6678# a_29182_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4158 a_51533_n5795# a_51363_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4159 VSS a_53381_6408# a_53329_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4160 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4161 a_31662_n6678# a_31070_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4162 VDD a_35072_n5879# a_34896_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4163 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4164 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4165 a_46758_n5622# a_46394_n5879# a_46662_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4166 VDD a_2646_n11559# a_2864_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4167 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4168 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4169 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4170 a_55873_773# a_55379_690# a_55434_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4171 a_37242_n10732# a_38460_n11533# a_38703_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4172 VSS a_27898_n10732# a_27900_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4173 a_24124_n11788# a_24122_n10732# a_24425_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4174 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4175 a_21909_5953# a_23179_6408# a_23370_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4176 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4177 a_20896_6655# a_20021_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4178 a_39776_6655# a_38901_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4179 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4180 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4181 a_5138_n5622# a_6532_n5789# a_6582_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4182 a_2022_6655# a_1147_5953# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4183 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4184 VDD a_36570_n7315# a_31249_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4185 a_38985_1829# a_38393_690# a_36999_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4186 a_33333_5953# a_32567_6434# a_33237_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4187 a_14461_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4188 a_13855_690# C[103] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4189 a_857_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4190 a_46531_1829# a_46165_836# a_44551_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4191 VSS a_47946_n11559# a_47894_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4192 a_57551_n6843# a_57546_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4193 VDD a_4534_n11559# a_4752_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4194 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4195 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4196 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4197 a_20119_7009# a_20117_5953# a_20420_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4198 a_25996_n5622# a_25998_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4199 a_19823_n10487# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4200 a_38999_7009# a_38997_5953# a_39300_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4201 VDD a_27559_773# a_28484_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4202 a_26012_n11788# a_26010_n10732# a_26313_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4203 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4204 VSS C[17] a_26955_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4205 a_17555_n5795# a_17385_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4206 VDD a_53717_836# a_53541_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4207 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4208 a_33548_n5622# a_33550_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4209 VSS a_46347_n6869# a_52422_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4210 a_18446_n6678# a_17854_n5789# a_16460_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4211 VDD a_36341_2600# a_31020_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4212 a_10445_n6843# a_10358_n6611# a_10363_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4213 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4214 a_48335_5953# a_49553_6434# a_49796_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4215 a_36505_690# C[115] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4216 a_2756_n5789# C[33] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4217 a_23219_n5795# a_23049_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4218 VSS a_49834_n11559# a_49782_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4219 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4220 VDD a_55269_6408# a_55217_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4221 a_46347_n6869# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4222 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4223 a_24110_n6678# a_23518_n5789# a_22124_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4224 a_25998_n6678# a_25406_n5789# a_24012_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4225 a_38901_5953# a_38231_6434# a_38501_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4226 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4227 a_55605_836# a_55379_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4228 a_44876_n5622# a_44878_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4229 a_37242_n10732# a_36572_n11533# a_36842_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4230 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4231 a_1147_5953# a_477_6434# a_747_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4232 a_2893_n6843# a_2806_n6611# a_2811_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4233 a_27900_n11788# a_27898_n10732# a_28201_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4234 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4235 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4236 VDD a_6193_6408# a_6411_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4237 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4238 a_27655_773# a_27065_690# a_27559_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4239 a_818_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4240 a_36435_n5795# a_36265_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4241 VSS a_36570_n7315# a_46157_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4242 a_48335_5953# a_47717_6408# a_47935_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4243 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4244 a_23893_5953# a_23127_6434# a_23797_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4245 a_37326_n6678# a_36734_n5789# a_35340_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4246 VSS a_36570_n7315# a_46347_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4247 a_14578_n5622# a_16192_n5879# a_16016_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4248 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4249 a_1094_n5879# a_868_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4250 a_2982_n5879# a_2756_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4251 a_42099_n5795# a_41929_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4252 VSS a_36999_773# a_37924_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4253 a_41004_n5622# a_40736_n5879# a_40565_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4254 a_43987_n5795# a_43817_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4255 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4256 a_31431_773# a_31067_836# a_31335_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4257 VSS RESET a_13714_3465# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4258 a_16558_n6678# a_15966_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4259 VDD a_40400_n11559# a_40618_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4260 VSS a_9024_n10732# a_9026_n11788# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4261 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4262 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4263 a_44878_n6678# a_44286_n5789# a_42892_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4264 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4265 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4266 a_20464_1994# a_20105_1829# a_20103_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4267 a_39344_1994# a_38985_1829# a_38983_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4268 a_31662_n6678# a_31296_n5879# a_29676_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4269 VSS a_1243_5953# a_1245_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4270 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4271 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4272 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4273 VDD a_46118_1932# a_53628_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4274 a_39130_n10732# a_38460_n11533# a_38730_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4275 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4276 a_10305_836# a_10079_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4277 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4278 a_8914_n5622# a_8420_n5789# a_8475_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4279 a_54671_n6843# a_54312_n6678# a_54310_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X4280 a_6811_5953# a_6193_6408# a_6411_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4281 a_45928_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4282 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4283 a_27669_5953# a_26955_6408# a_27573_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4284 VSS a_19008_6655# a_18958_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4285 a_12800_n10732# a_12034_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4286 a_57775_5953# a_58993_6434# a_59236_5708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4287 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4288 a_33452_n5622# a_35072_n5879# a_34896_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4289 a_59990_n11788# a_59274_n11559# a_58004_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4290 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4291 VSS C[8] a_43947_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4292 VSS a_26789_n11370# a_26739_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4293 a_35438_n6678# a_34846_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4294 VDD a_42288_n11559# a_42506_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4295 a_46347_n6869# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4296 a_54081_773# a_53717_836# a_53985_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4297 a_50223_5953# a_49605_6408# a_49823_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4298 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4299 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4300 a_6758_n5879# a_6532_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4301 a_29034_5708# a_29061_6449# a_29046_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4302 VDD a_13714_3465# a_6139_2600# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4303 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4304 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4305 a_27559_773# a_27291_836# a_27120_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4306 VDD a_46347_n6869# a_57633_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4307 a_58174_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4308 a_55969_773# a_55605_836# a_55873_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4309 VSS a_31020_1932# a_37095_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4310 VDD a_53985_773# a_54910_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4311 VDD a_15916_1932# a_26128_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4312 VDD a_36570_n7315# a_46347_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4313 a_31059_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4314 VDD a_16145_n6869# a_26357_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4315 a_37109_5953# a_36343_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4316 a_31335_773# a_30841_690# a_30896_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4317 a_51304_696# a_51134_696# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4318 VDD RESET a_13714_3465# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4319 a_27884_n5622# a_27294_n5789# a_27788_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4320 VDD a_44176_n11559# a_44394_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4321 a_9026_n11788# a_9024_n10732# a_9327_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4322 a_29904_1994# a_29545_1829# a_29543_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4323 a_15673_n5795# a_15503_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4324 a_1474_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4325 VSS a_6368_n7315# a_16145_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4326 a_40885_5953# a_40119_6434# a_40789_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4327 a_2228_696# a_2058_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4328 a_2251_n11370# a_1376_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4329 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4330 VSS a_818_1932# a_8781_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4331 VSS a_16145_n6869# a_27349_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4332 VDD a_31249_n6869# a_39573_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4333 a_36570_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4334 VDD a_6139_2600# a_15726_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4335 VDD a_36341_2600# a_30830_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4336 a_48564_n10732# a_49782_n11533# a_50025_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4337 VSS a_38501_6449# a_38474_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4338 a_18348_n5622# a_18080_n5879# a_17909_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4339 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4340 a_44150_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4341 a_50223_5953# a_49553_6434# a_49823_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X4342 VDD a_27788_n5622# a_28713_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4343 a_50550_n11788# a_46157_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4344 VDD a_31249_n6869# a_45237_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4345 a_51327_n11370# a_50452_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4346 a_16145_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4347 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4348 a_44661_5953# a_43947_6408# a_44565_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4349 VSS a_36000_6655# a_35950_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4350 a_25900_n5622# a_25632_n5879# a_25461_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4351 a_3362_n11788# a_857_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4352 a_38999_7009# a_38231_6434# a_37013_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4353 a_628_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4354 a_16558_n6678# a_16192_n5879# a_14578_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4355 VSS a_25296_n11559# a_25244_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4356 a_1245_7009# a_477_6434# a_224_6410# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4357 a_31020_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4358 a_59747_1829# a_59155_690# a_57761_773# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4359 VDD a_59045_6408# a_59263_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X4360 a_20007_773# a_19513_690# a_19568_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X4361 a_6669_n6843# a_6582_n6611# a_6587_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4362 a_59974_n5622# a_59976_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4363 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4364 a_13714_3465# RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4365 a_26789_n11370# a_25914_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4366 a_46531_1829# a_45939_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4367 a_37228_n5622# a_36960_n5879# a_36789_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4368 VDD C[86] a_17744_n11559# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4369 VSS C[15] a_30731_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4370 a_51533_n5795# a_51363_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4371 VDD a_19632_n11559# a_19850_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4372 a_59988_n10732# a_59274_n11559# a_59878_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4373 a_28953_690# C[111] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4374 a_27669_5953# a_26903_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4375 a_29182_n5789# C[47] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4376 a_52424_n6678# a_51832_n5789# a_50438_n5622# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4377 VSS a_1047_n6869# a_14674_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4378 a_53215_n11370# a_52340_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4379 a_55887_5953# a_55269_6408# a_55487_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4380 a_48662_n11788# a_47946_n11559# a_46676_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4381 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4382 a_8795_5953# a_8029_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4383 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4384 VSS a_6139_2600# a_818_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4385 a_51658_1994# a_51653_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4386 a_31067_836# a_30841_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4387 a_44780_n5622# a_44512_n5879# a_44341_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4388 a_31564_n5622# a_31070_n5789# a_31125_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4389 VSS a_15461_n11370# a_15411_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4390 VSS C[77] a_34736_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4391 a_15955_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4392 VDD a_6368_n7315# a_16145_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4393 a_6909_7009# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4394 VDD a_31020_1932# a_43120_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4395 VDD a_30960_n11559# a_31178_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4396 a_21723_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4397 VSS a_54095_5953# a_54097_7009# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4398 VSS a_46662_n5622# a_47587_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4399 a_35438_n6678# a_35072_n5879# a_33452_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4400 VSS a_27184_n11559# a_27132_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4401 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4402 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4403 VSS a_36341_2600# a_30830_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4404 a_25914_n10732# a_27132_n11533# a_27375_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4405 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4406 a_58447_n6843# a_58088_n6678# a_58086_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4407 VDD a_6139_2600# a_15916_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4408 a_28677_n11370# a_27802_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4409 a_8685_773# a_10305_836# a_10129_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4410 VSS a_12461_773# a_13386_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4411 a_34710_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4412 VSS a_15916_1932# a_27120_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4413 VDD a_17851_836# a_17675_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4414 a_53985_773# a_53717_836# a_53546_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4415 a_59649_773# a_58993_6434# a_59263_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4416 a_628_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4417 VDD a_48282_n5879# a_48106_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4418 a_16145_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4419 a_48550_n5622# a_50170_n5879# a_49994_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4420 VSS a_26560_6655# a_26510_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4421 VSS a_36341_2600# a_46118_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4422 a_29408_n5879# a_29182_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4423 a_40005_n11370# a_39130_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4424 VSS a_17349_n11370# a_17299_n11535# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4425 VSS C[76] a_36624_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4426 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4427 a_50536_n6678# a_49944_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4428 VDD a_32848_n11559# a_33066_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4429 a_23611_n10237# a_15955_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4430 VDD a_55834_n5879# a_55658_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4431 VSS C[85] a_19632_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4432 VSS a_29072_n11559# a_29020_n11533# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4433 VDD a_49605_6408# a_49823_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4434 a_10134_1994# a_10129_1896# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4435 a_23879_773# a_23881_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4436 VDD a_1047_n6869# a_1005_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4437 a_30934_5388# a_30830_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4438 a_13714_3465# RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4439 VDD a_1047_n6869# a_2893_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4440 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4441 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4442 a_1047_n6869# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4443 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4444 VSS a_35111_773# a_36036_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4445 a_43758_696# a_43588_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4446 VSS C[30] a_2417_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4447 a_15916_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4448 a_46772_n10732# a_46058_n11559# a_46676_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4449 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4450 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4451 a_54097_7009# a_53329_6434# a_52111_5953# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4452 a_45928_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4453 a_42169_690# C[118] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4454 a_41116_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4455 a_48431_5953# a_47717_6408# a_48335_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X4456 a_8914_n5622# a_10534_n5879# a_10358_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4457 a_18444_n5622# a_18080_n5879# a_18348_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X4458 VDD a_34736_n11559# a_34954_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4459 VSS C[84] a_21520_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4460 a_44661_5953# a_43895_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4461 a_25403_836# a_25177_690# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4462 a_30771_n5795# a_30601_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4463 a_16021_n6843# a_16016_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4464 VSS a_40618_n11298# a_40591_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4465 a_818_1932# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4466 VDD a_36341_2600# a_46118_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4467 VDD a_29447_773# a_30372_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4468 a_17909_n6843# a_17904_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4469 VSS a_6368_n7315# a_1047_n6869# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4470 a_25258_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4471 a_30830_5620# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4472 a_19650_1994# a_19563_1896# a_19568_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4473 a_24108_n5622# a_23744_n5879# a_24012_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4474 a_55985_7009# a_55269_6408# a_53999_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4475 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4476 a_25996_n5622# a_25632_n5879# a_25900_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4477 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4478 VDD a_6368_n7315# a_857_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4479 VDD a_46347_n6869# a_54671_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4480 a_14363_5953# a_13745_6408# a_13963_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4481 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4482 VSS a_13714_3465# a_36341_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4483 a_16329_1829# a_15963_836# a_14349_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4484 a_25671_773# a_27065_690# a_27115_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4485 a_48660_n10732# a_47946_n11559# a_48564_n10732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4486 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4487 a_6907_5953# a_6193_6408# a_6811_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4488 a_43004_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4489 VDD a_46347_n6869# a_60335_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4490 VDD C[27] a_8081_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4491 a_36586_5708# a_36613_6449# a_36598_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4492 VSS a_31020_1932# a_44112_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4493 a_18215_773# a_17851_836# a_18119_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4494 VSS a_36341_2600# a_31020_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4495 VSS C[83] a_23408_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4496 VSS a_42506_n11298# a_42479_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4497 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4498 VDD a_52097_773# a_53022_696# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4499 a_36789_n6843# a_36784_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4500 VSS a_43552_6655# a_43502_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4501 a_14592_n10732# a_15804_n11533# a_16047_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4502 a_44876_n5622# a_44512_n5879# a_44780_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4503 VSS a_16145_n6869# a_24108_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4504 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4505 a_1047_n6869# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4506 a_6893_773# a_6529_836# a_6797_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4507 a_17349_n11370# a_16474_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4508 a_46157_n10335# a_36570_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4509 a_52326_n5622# a_52058_n5879# a_51887_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4510 a_40871_773# a_40873_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4511 a_46433_773# a_45939_690# a_45994_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4512 VSS a_16145_n6869# a_29772_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4513 a_44892_n11788# a_31059_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4514 a_15955_n10335# a_6368_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4515 VDD a_36341_2600# a_45928_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4516 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4517 VSS a_44394_n11298# a_44367_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4518 a_40591_n10487# a_40618_n11298# a_40603_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4519 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4520 a_15818_5708# a_15726_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4521 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4522 VDD a_6368_n7315# a_1047_n6869# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4523 a_50536_n6678# a_50170_n5879# a_48550_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4524 VSS C[2] a_55269_6408# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4525 VSS C[90] a_10198_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4526 a_16474_n10732# a_17692_n11533# a_17935_n10487# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4527 a_14688_n10732# a_13922_n11533# a_14592_n10732# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4528 VSS a_31249_n6869# a_42988_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4529 a_18460_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4530 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4531 VSS a_46118_1932# a_59745_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4532 a_9010_n5622# a_9012_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4533 a_19237_n11370# a_18362_n10732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4534 VDD a_6368_n7315# a_15955_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4535 VDD a_41893_n11370# a_41843_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4536 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4537 a_46118_1932# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4538 VDD a_6139_2600# a_818_1932# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4539 VDD a_818_1932# a_1590_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4540 a_36642_1994# a_36555_1896# a_36560_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4541 a_15673_n5795# a_15503_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4542 a_6625_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4543 VDD a_36570_n7315# a_31059_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4544 a_42663_773# a_44057_690# a_44107_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4545 VSS a_46118_1932# a_48417_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4546 a_18119_773# a_17625_690# a_17680_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4547 a_29788_n11788# a_15955_n10335# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4548 VDD a_25067_6408# a_25015_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4549 a_36341_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4550 VDD a_59610_n5879# a_59434_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4551 a_42479_n10487# a_42506_n11298# a_42491_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4552 a_48431_5953# a_47665_6434# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4553 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4554 a_21991_773# a_21627_836# a_21895_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4555 VSS C[89] a_12086_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4556 a_5798_6655# a_4923_5953# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4557 a_27065_690# C[110] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4558 VSS a_40171_6408# a_40119_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4559 a_10900_n6678# a_10534_n5879# a_8914_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4560 a_31059_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4561 a_8328_1994# a_8241_1896# a_8246_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4562 a_18133_5953# a_17515_6408# a_17733_6449# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4563 a_6797_773# a_6303_690# a_6358_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4564 a_31431_773# a_31433_1829# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4565 VDD a_43781_n11370# a_43731_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4566 VSS a_28843_6408# a_28791_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4567 a_8513_n10237# a_857_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4568 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4569 a_46165_836# a_45939_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4570 a_8699_5953# a_9969_6408# a_10160_5708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4571 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4572 VSS a_36570_n7315# a_31059_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4573 a_29447_773# a_31067_836# a_30891_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4574 a_18215_773# a_17625_690# a_18119_773# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4575 a_12690_n5622# a_14310_n5879# a_14134_n6611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4576 a_6368_n7315# a_13714_3465# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4577 VSS a_46118_1932# a_47882_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4578 a_55472_5388# a_45928_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4579 VSS a_6139_2600# a_15726_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4580 a_46758_n5622# a_46168_n5789# a_46662_n5622# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4581 a_44367_n10487# a_44394_n11298# a_44379_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4582 a_12788_n6678# a_12196_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4583 a_34547_n5795# a_34377_n5795# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X4584 a_16474_n10732# a_15804_n11533# a_16074_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4585 a_55983_5953# a_55269_6408# a_55887_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4586 a_15726_5620# a_6139_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4587 a_14676_n6678# a_14084_n5789# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4588 VSS C[88] a_13974_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4589 VSS a_31178_n11298# a_31151_n10487# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4590 VSS a_47322_6655# a_47272_6436# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4591 a_52097_773# a_51829_836# a_51658_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4592 VSS a_39116_n5622# a_40041_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4593 VSS a_41004_n5622# a_41929_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4594 VDD a_16145_n6869# a_29319_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4595 VSS a_6368_n7315# a_15955_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4596 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4597 VSS a_27559_773# a_28484_696# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4598 a_57589_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4599 a_15726_5620# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4600 VSS a_6139_2600# a_628_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4601 a_15916_1932# a_6139_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4602 VSS a_46347_n6869# a_46223_n6843# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4603 a_46545_7009# a_45928_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4604 a_46157_n10335# a_36570_n7315# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4605 VSS C[92] a_6422_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4606 VSS a_13714_3465# a_6368_n7315# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4607 VDD a_4641_836# a_4465_1896# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4608 VSS a_529_6408# a_477_6434# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4609 VDD a_46662_n5622# a_47587_n5795# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4610 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4611 VSS a_818_1932# a_6358_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4612 a_3250_n5622# a_4644_n5789# a_4694_n6611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4613 a_10986_5388# a_628_5620# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4614 VSS a_6139_2600# a_15916_1932# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4615 a_21895_773# a_21401_690# a_21456_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4616 a_31977_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4617 a_49999_n6843# a_49994_n6611# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4618 VDD a_46118_1932# a_54442_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4619 a_59878_n5622# a_59222_n11533# a_59492_n11298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4620 a_59477_n10237# a_46157_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4621 VDD a_42059_6408# a_42007_6434# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4622 VSS a_36341_2600# a_45928_5620# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4623 a_6529_836# a_6303_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4624 a_58856_696# a_58686_696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4625 VDD a_13714_3465# a_36570_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4626 a_30841_690# C[112] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4627 a_20332_n5622# a_20334_n6678# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4628 VSS a_818_1932# a_2582_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4629 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4630 a_57267_690# C[126] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4631 VDD a_30565_n11370# a_30515_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4632 VSS C[91] a_8310_n11559# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X4633 a_20007_773# a_21627_836# a_21451_1896# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X4634 a_18119_773# a_17851_836# a_17680_1994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4635 a_48056_n5789# C[57] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4636 a_6368_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4637 a_49944_n5789# C[58] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4638 a_6139_2600# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4639 VSS a_13714_3465# a_6139_2600# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4640 a_10683_5953# a_9917_6434# a_10587_5953# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X4641 VDD a_46118_1932# a_50666_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4642 a_50438_n5622# a_49944_n5789# a_49999_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4643 a_23881_1829# a_23515_836# a_21895_773# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4644 a_33865_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4645 a_31151_n10487# a_31178_n11298# a_31163_n10237# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4646 a_46118_1932# a_36341_2600# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4647 a_55608_n5789# C[61] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4648 a_48193_n6843# a_48106_n6611# a_48111_n6843# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4649 VDD a_36570_n7315# a_46157_n10335# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4650 a_857_n10335# a_6368_n7315# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4651 a_36570_n7315# a_13714_3465# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4652 a_57348_5708# a_57375_6449# a_57360_5388# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4653 VDD a_6139_2600# a_628_5620# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4654 a_4496_5708# a_628_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4655 VDD a_31020_1932# a_40418_1994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4656 a_53491_690# C[124] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4657 a_18805_n6843# a_18446_n6678# a_18444_n5622# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4658 VDD a_13714_3465# a_6368_n7315# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4659 a_20021_5953# a_19351_6434# a_19621_6449# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4660 VDD a_32453_n11370# a_32403_n11535# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4661 VDD a_30336_6655# a_30286_6436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X4662 a_35450_n10732# a_34684_n11533# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4663 a_30771_n5795# a_30601_n5795# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X4664 a_48282_n5879# a_48056_n5789# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X4665 a_14459_5953# a_13745_6408# a_14363_5953# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4666 VSS a_18348_n5622# a_19273_n5795# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X4667 a_30830_5620# a_36341_2600# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4668 VSS a_6368_n7315# a_857_n10335# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4669 VDD C[0] a_59045_6408# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X4670 a_21627_836# a_21401_690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X4671 a_35753_n10237# a_31059_n10335# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

