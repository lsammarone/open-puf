magic
tech sky130A
magscale 1 2
timestamp 1655262894
<< nwell >>
rect 33027 4847 33405 5966
rect 32760 4818 33405 4847
rect 32760 4526 33296 4818
rect 17040 4150 17422 4471
rect 47182 4310 47564 4631
<< nsubdiff >>
rect 47307 4483 47441 4502
rect 47307 4449 47379 4483
rect 47413 4449 47441 4483
rect 47307 4432 47441 4449
rect 17165 4323 17299 4342
rect 17165 4289 17237 4323
rect 17271 4289 17299 4323
rect 17165 4272 17299 4289
<< nsubdiffcont >>
rect 47379 4449 47413 4483
rect 17237 4289 17271 4323
<< locali >>
rect 32002 4524 32358 4530
rect 32002 4490 32049 4524
rect 32083 4490 32137 4524
rect 32171 4490 32358 4524
rect 32002 4480 32358 4490
rect 47104 4483 47647 4503
rect 47104 4449 47379 4483
rect 47413 4449 47647 4483
rect 47104 4431 47647 4449
rect 16962 4323 17505 4343
rect 16962 4289 17237 4323
rect 17271 4289 17505 4323
rect 16962 4271 17505 4289
<< viali >>
rect 32049 4490 32083 4524
rect 32137 4490 32171 4524
rect 32714 4522 32748 4556
rect 32985 4486 33019 4520
rect 33073 4486 33107 4520
rect 33161 4486 33195 4520
rect 33249 4486 33283 4520
rect 33337 4486 33371 4520
rect 33425 4486 33459 4520
rect 33513 4486 33547 4520
rect 33601 4486 33635 4520
rect 32714 4442 32748 4476
rect 33339 4384 33373 4418
rect 33505 4380 33539 4414
rect 33673 4386 33707 4420
rect 33840 4384 33874 4418
rect 34010 4385 34044 4419
rect 34174 4386 34208 4420
rect 45805 4363 45839 4408
rect 45973 4370 46007 4415
rect 46141 4360 46175 4405
rect 46309 4372 46343 4417
rect 46475 4370 46509 4415
rect 46641 4372 46675 4417
rect 46809 4372 46843 4417
rect 46983 4370 47017 4415
rect 47739 4364 47773 4409
rect 47901 4368 47935 4413
rect 48071 4372 48105 4417
rect 48235 4368 48269 4413
rect 48405 4368 48439 4413
rect 48573 4364 48607 4409
rect 48741 4368 48775 4413
rect 48915 4364 48949 4409
rect 46005 4272 46039 4306
rect 46105 4272 46139 4306
rect 46205 4272 46239 4306
rect 46305 4272 46339 4306
rect 46405 4272 46439 4306
rect 46505 4272 46539 4306
rect 46605 4272 46639 4306
rect 46705 4272 46739 4306
rect 47665 4272 47699 4306
rect 47765 4272 47799 4306
rect 47865 4272 47899 4306
rect 47965 4272 47999 4306
rect 48065 4272 48099 4306
rect 48165 4272 48199 4306
rect 48265 4272 48299 4306
rect 48365 4272 48399 4306
rect 15663 4203 15697 4248
rect 15831 4210 15865 4255
rect 15999 4200 16033 4245
rect 16167 4212 16201 4257
rect 16333 4210 16367 4255
rect 16499 4212 16533 4257
rect 16667 4212 16701 4257
rect 16841 4210 16875 4255
rect 17597 4204 17631 4249
rect 17759 4208 17793 4253
rect 17929 4212 17963 4257
rect 18093 4208 18127 4253
rect 18263 4208 18297 4253
rect 18431 4204 18465 4249
rect 18599 4208 18633 4253
rect 18773 4204 18807 4249
rect 15863 4112 15897 4146
rect 15963 4112 15997 4146
rect 16063 4112 16097 4146
rect 16163 4112 16197 4146
rect 16263 4112 16297 4146
rect 16363 4112 16397 4146
rect 16463 4112 16497 4146
rect 16563 4112 16597 4146
rect 17523 4112 17557 4146
rect 17623 4112 17657 4146
rect 17723 4112 17757 4146
rect 17823 4112 17857 4146
rect 17923 4112 17957 4146
rect 18023 4112 18057 4146
rect 18123 4112 18157 4146
rect 18223 4112 18257 4146
<< metal1 >>
rect 16714 5441 16969 5797
rect 32650 5464 32984 5788
rect 16714 5389 16734 5441
rect 16786 5389 16812 5441
rect 16864 5389 16905 5441
rect 16957 5389 16969 5441
rect 16714 5359 16969 5389
rect 32650 5412 32693 5464
rect 32745 5412 32806 5464
rect 32858 5412 32907 5464
rect 32959 5412 32984 5464
rect 32650 5368 32984 5412
rect 46854 5441 47081 5809
rect 46854 5389 46885 5441
rect 46937 5389 46968 5441
rect 47020 5389 47081 5441
rect 46854 5355 47081 5389
rect 9370 5224 9906 5308
rect 24404 5233 25012 5291
rect 39508 5241 40132 5299
rect 54514 5247 55247 5305
rect 32778 4844 32886 4857
rect 32778 4792 32808 4844
rect 32860 4792 32886 4844
rect 32778 4761 32886 4792
rect 34318 4761 34353 4857
rect 1 4690 19384 4691
rect 0 4626 19384 4690
rect 1 4625 19384 4626
rect 19318 4539 19384 4625
rect 47023 4617 47690 4626
rect 32699 4556 32778 4584
rect 47033 4568 47690 4617
rect 19318 4524 32265 4539
rect 19318 4490 32049 4524
rect 32083 4490 32137 4524
rect 32171 4490 32265 4524
rect 19318 4473 32265 4490
rect 32699 4522 32714 4556
rect 32748 4528 32778 4556
rect 32748 4522 33697 4528
rect 32699 4520 33697 4522
rect 32699 4486 32985 4520
rect 33019 4486 33073 4520
rect 33107 4486 33161 4520
rect 33195 4486 33249 4520
rect 33283 4486 33337 4520
rect 33371 4486 33425 4520
rect 33459 4486 33513 4520
rect 33547 4486 33601 4520
rect 33635 4486 33697 4520
rect 32699 4480 33697 4486
rect 32699 4476 32781 4480
rect 16933 4412 17582 4462
rect 32699 4442 32714 4476
rect 32748 4442 32781 4476
rect 32699 4424 32781 4442
rect 33270 4435 34215 4448
rect 16881 4404 17582 4412
rect 33270 4418 33486 4435
rect 33270 4384 33339 4418
rect 33373 4384 33486 4418
rect 33538 4414 33646 4435
rect 33698 4420 33779 4435
rect 33270 4383 33486 4384
rect 33539 4383 33646 4414
rect 33707 4386 33779 4420
rect 33698 4383 33779 4386
rect 33831 4418 33892 4435
rect 33831 4384 33840 4418
rect 33874 4384 33892 4418
rect 33831 4383 33892 4384
rect 33944 4420 34215 4435
rect 33944 4419 34174 4420
rect 33944 4385 34010 4419
rect 34044 4386 34174 4419
rect 34208 4386 34215 4420
rect 34044 4385 34215 4386
rect 33944 4383 34215 4385
rect 33270 4380 33505 4383
rect 33539 4380 34215 4383
rect 33270 4365 34215 4380
rect 39672 4417 55107 4427
rect 39672 4415 46309 4417
rect 39672 4408 45973 4415
rect 39672 4407 39854 4408
rect 39672 4355 39751 4407
rect 39803 4356 39854 4407
rect 39906 4363 45805 4408
rect 45839 4370 45973 4408
rect 46007 4405 46309 4415
rect 46007 4370 46141 4405
rect 45839 4363 46141 4370
rect 39906 4360 46141 4363
rect 46175 4372 46309 4405
rect 46343 4415 46641 4417
rect 46343 4372 46475 4415
rect 46175 4370 46475 4372
rect 46509 4372 46641 4415
rect 46675 4372 46809 4417
rect 46843 4415 48071 4417
rect 46843 4372 46983 4415
rect 46509 4370 46983 4372
rect 47017 4413 48071 4415
rect 47017 4409 47901 4413
rect 47017 4370 47739 4409
rect 46175 4364 47739 4370
rect 47773 4368 47901 4409
rect 47935 4372 48071 4413
rect 48105 4413 55107 4417
rect 48105 4372 48235 4413
rect 47935 4368 48235 4372
rect 48269 4368 48405 4413
rect 48439 4409 48741 4413
rect 48439 4368 48573 4409
rect 47773 4364 48573 4368
rect 48607 4368 48741 4409
rect 48775 4409 55107 4413
rect 48775 4368 48915 4409
rect 48607 4364 48915 4368
rect 48949 4408 55107 4409
rect 48949 4403 54955 4408
rect 48949 4364 54864 4403
rect 46175 4360 54864 4364
rect 39906 4356 54864 4360
rect 39803 4355 54864 4356
rect 39672 4351 54864 4355
rect 54916 4356 54955 4403
rect 55007 4356 55107 4408
rect 54916 4351 55107 4356
rect 39672 4346 55107 4351
rect 32778 4294 32881 4313
rect 32778 4291 32868 4294
rect 9515 4257 24881 4267
rect 9515 4255 16167 4257
rect 9515 4252 15831 4255
rect 9515 4200 9556 4252
rect 9608 4200 9652 4252
rect 9704 4248 15831 4252
rect 9704 4203 15663 4248
rect 15697 4210 15831 4248
rect 15865 4245 16167 4255
rect 15865 4210 15999 4245
rect 15697 4203 15999 4210
rect 9704 4200 15999 4203
rect 16033 4212 16167 4245
rect 16201 4255 16499 4257
rect 16201 4212 16333 4255
rect 16033 4210 16333 4212
rect 16367 4212 16499 4255
rect 16533 4212 16667 4257
rect 16701 4255 17929 4257
rect 16701 4212 16841 4255
rect 16367 4210 16841 4212
rect 16875 4253 17929 4255
rect 16875 4249 17759 4253
rect 16875 4210 17597 4249
rect 16033 4204 17597 4210
rect 17631 4208 17759 4249
rect 17793 4212 17929 4253
rect 17963 4253 24881 4257
rect 17963 4212 18093 4253
rect 17793 4208 18093 4212
rect 18127 4208 18263 4253
rect 18297 4249 18599 4253
rect 18297 4208 18431 4249
rect 17631 4204 18431 4208
rect 18465 4208 18599 4249
rect 18633 4250 24881 4253
rect 18633 4249 24766 4250
rect 18633 4208 18773 4249
rect 18465 4204 18773 4208
rect 18807 4243 24766 4249
rect 18807 4204 24667 4243
rect 16033 4200 24667 4204
rect 9515 4191 24667 4200
rect 24719 4198 24766 4243
rect 24818 4198 24881 4250
rect 32809 4242 32868 4291
rect 32809 4239 32881 4242
rect 32778 4217 32881 4239
rect 34318 4217 34353 4313
rect 45973 4306 48576 4312
rect 45973 4272 46005 4306
rect 46039 4272 46105 4306
rect 46139 4272 46205 4306
rect 46239 4272 46305 4306
rect 46339 4272 46405 4306
rect 46439 4272 46505 4306
rect 46539 4272 46605 4306
rect 46639 4272 46705 4306
rect 46739 4272 47665 4306
rect 47699 4272 47765 4306
rect 47799 4272 47865 4306
rect 47899 4272 47965 4306
rect 47999 4272 48065 4306
rect 48099 4272 48165 4306
rect 48199 4272 48265 4306
rect 48299 4272 48365 4306
rect 48399 4272 48576 4306
rect 45973 4267 48576 4272
rect 45973 4264 47419 4267
rect 47269 4263 47419 4264
rect 24719 4191 24881 4198
rect 9515 4186 24881 4191
rect 47269 4211 47314 4263
rect 47366 4215 47419 4263
rect 47471 4264 48576 4267
rect 47471 4215 47497 4264
rect 47366 4211 47497 4215
rect 47269 4172 47497 4211
rect 15831 4146 18434 4152
rect 15831 4112 15863 4146
rect 15897 4112 15963 4146
rect 15997 4112 16063 4146
rect 16097 4112 16163 4146
rect 16197 4112 16263 4146
rect 16297 4112 16363 4146
rect 16397 4112 16463 4146
rect 16497 4112 16563 4146
rect 16597 4112 17523 4146
rect 17557 4112 17623 4146
rect 17657 4112 17723 4146
rect 17757 4112 17823 4146
rect 17857 4112 17923 4146
rect 17957 4112 18023 4146
rect 18057 4112 18123 4146
rect 18157 4112 18223 4146
rect 18257 4112 18434 4146
rect 15831 4107 18434 4112
rect 15831 4104 17277 4107
rect 17127 4103 17277 4104
rect 17127 4051 17172 4103
rect 17224 4055 17277 4103
rect 17329 4104 18434 4107
rect 17329 4055 17355 4104
rect 17224 4051 17355 4055
rect 17127 4012 17355 4051
rect 47023 4020 47775 4078
rect 15493 3842 15544 3938
rect 16881 3866 17562 3924
rect 22012 3869 47523 3913
rect 22012 3867 47411 3869
rect 15493 3841 15543 3842
rect 22012 3815 33475 3867
rect 33527 3815 33619 3867
rect 33671 3815 33763 3867
rect 33815 3866 47411 3867
rect 33815 3815 47322 3866
rect 22012 3814 47322 3815
rect 47374 3817 47411 3866
rect 47463 3817 47523 3869
rect 47374 3814 47523 3817
rect 22012 3790 47523 3814
rect 22012 3783 47322 3790
rect 22012 3731 33474 3783
rect 33526 3731 33618 3783
rect 33670 3731 33762 3783
rect 33814 3738 47322 3783
rect 47374 3738 47415 3790
rect 47467 3738 47523 3790
rect 33814 3731 47523 3738
rect 17139 3707 47523 3731
rect 17139 3686 22218 3707
rect 17139 3634 17176 3686
rect 17228 3681 22218 3686
rect 17228 3634 17270 3681
rect 17139 3629 17270 3634
rect 17322 3629 22218 3681
rect 17139 3608 22218 3629
rect 17139 3606 17270 3608
rect 9306 3532 9969 3590
rect 17139 3554 17176 3606
rect 17228 3556 17270 3606
rect 17322 3556 22218 3608
rect 17228 3554 22218 3556
rect 17139 3525 22218 3554
rect 24404 3544 25032 3602
rect 39416 3544 40179 3602
rect 54606 3535 55257 3593
rect 62673 1474 62895 1552
<< via1 >>
rect 9555 5455 9607 5507
rect 9636 5454 9688 5506
rect 24671 5452 24723 5504
rect 24766 5452 24818 5504
rect 16734 5389 16786 5441
rect 16812 5389 16864 5441
rect 16905 5389 16957 5441
rect 32693 5412 32745 5464
rect 32806 5412 32858 5464
rect 32907 5412 32959 5464
rect 39748 5454 39800 5506
rect 39850 5454 39902 5506
rect 46885 5389 46937 5441
rect 46968 5389 47020 5441
rect 54866 5427 54918 5479
rect 54961 5427 55013 5479
rect 8563 5233 8615 5285
rect 8670 5235 8722 5287
rect 8772 5235 8824 5287
rect 8872 5236 8924 5288
rect 23593 5239 23645 5291
rect 23696 5239 23748 5291
rect 23779 5239 23831 5291
rect 23880 5239 23932 5291
rect 23967 5239 24019 5291
rect 38725 5235 38777 5287
rect 38813 5235 38865 5287
rect 38898 5240 38950 5292
rect 55641 5232 55693 5284
rect 55735 5232 55787 5284
rect 55812 5232 55864 5284
rect 55892 5231 55944 5283
rect 55966 5232 56018 5284
rect 32705 4789 32757 4841
rect 32808 4792 32860 4844
rect 32909 4792 32961 4844
rect 46891 4564 46943 4616
rect 46981 4565 47033 4617
rect 16758 4412 16810 4464
rect 16881 4412 16933 4464
rect 33486 4414 33538 4435
rect 33646 4420 33698 4435
rect 33486 4383 33505 4414
rect 33505 4383 33538 4414
rect 33646 4386 33673 4420
rect 33673 4386 33698 4420
rect 33646 4383 33698 4386
rect 33779 4383 33831 4435
rect 33892 4383 33944 4435
rect 39751 4355 39803 4407
rect 39854 4356 39906 4408
rect 54864 4351 54916 4403
rect 54955 4356 55007 4408
rect 9556 4200 9608 4252
rect 9652 4200 9704 4252
rect 24667 4191 24719 4243
rect 24766 4198 24818 4250
rect 32661 4237 32713 4289
rect 32757 4239 32809 4291
rect 32868 4242 32920 4294
rect 32960 4239 33012 4291
rect 47314 4211 47366 4263
rect 47419 4215 47471 4267
rect 17172 4051 17224 4103
rect 17277 4055 17329 4107
rect 48326 4024 48378 4076
rect 48418 4025 48470 4077
rect 48508 4024 48560 4076
rect 48596 4023 48648 4075
rect 15971 3863 16023 3915
rect 16055 3863 16107 3915
rect 16148 3864 16200 3916
rect 33475 3815 33527 3867
rect 33619 3815 33671 3867
rect 33763 3815 33815 3867
rect 47322 3814 47374 3866
rect 47411 3817 47463 3869
rect 33474 3731 33526 3783
rect 33618 3731 33670 3783
rect 33762 3731 33814 3783
rect 47322 3738 47374 3790
rect 47415 3738 47467 3790
rect 17176 3634 17228 3686
rect 17270 3629 17322 3681
rect 8557 3535 8609 3587
rect 8655 3535 8707 3587
rect 8750 3535 8802 3587
rect 8855 3535 8907 3587
rect 17176 3554 17228 3606
rect 17270 3556 17322 3608
rect 23607 3540 23659 3592
rect 23707 3540 23759 3592
rect 23806 3540 23858 3592
rect 23909 3540 23961 3592
rect 38715 3534 38767 3586
rect 38803 3534 38855 3586
rect 38901 3530 38953 3582
rect 55637 3531 55689 3583
rect 55725 3531 55777 3583
rect 55808 3531 55860 3583
rect 55895 3531 55947 3583
rect 9556 3317 9608 3369
rect 9636 3315 9688 3367
rect 24672 3332 24724 3384
rect 24755 3332 24807 3384
rect 39750 3322 39802 3374
rect 39841 3322 39893 3374
rect 54867 3307 54919 3359
rect 54950 3307 55002 3359
<< metal2 >>
rect 5569 7342 5613 8498
rect 7457 7342 7501 8498
rect 9345 7342 9389 8498
rect 11233 7342 11277 8498
rect 13121 7342 13165 8498
rect 15009 7342 15053 8498
rect 16897 7342 16941 8498
rect 18785 7342 18829 8498
rect 20673 7342 20717 8498
rect 22561 7342 22605 8498
rect 24449 7342 24493 8498
rect 26337 7342 26381 8498
rect 28225 7342 28269 8498
rect 30113 7342 30157 8498
rect 32001 7342 32045 8498
rect 33889 7342 33933 8498
rect 35777 7342 35821 8498
rect 37665 7342 37709 8498
rect 39553 7342 39597 8498
rect 41441 7342 41485 8498
rect 43329 7342 43373 8498
rect 45217 7342 45261 8498
rect 47105 7342 47149 8498
rect 48993 7342 49037 8498
rect 50881 7342 50925 8498
rect 52769 7342 52813 8498
rect 54657 7342 54701 8498
rect 56545 7342 56589 8498
rect 58433 7342 58477 8498
rect 60321 7342 60365 8498
rect 62209 7342 62253 8498
rect 208 6660 322 6695
rect 64230 6660 64344 6699
rect 208 6624 4285 6660
rect 62229 6624 64344 6660
rect 208 2204 322 6624
rect 9531 5507 9720 5537
rect 9531 5455 9555 5507
rect 9607 5506 9720 5507
rect 9607 5455 9636 5506
rect 9531 5454 9636 5455
rect 9688 5454 9720 5506
rect 8499 5288 8983 5413
rect 8499 5287 8872 5288
rect 8499 5285 8670 5287
rect 8499 5233 8563 5285
rect 8615 5235 8670 5285
rect 8722 5235 8772 5287
rect 8824 5236 8872 5287
rect 8924 5236 8983 5288
rect 8824 5235 8983 5236
rect 8615 5233 8983 5235
rect 8499 4066 8983 5233
rect 8499 4010 8566 4066
rect 8622 4010 8680 4066
rect 8736 4010 8794 4066
rect 8850 4010 8983 4066
rect 8499 3951 8983 4010
rect 8499 3895 8566 3951
rect 8622 3895 8680 3951
rect 8736 3895 8794 3951
rect 8850 3895 8983 3951
rect 8499 3836 8983 3895
rect 8499 3780 8566 3836
rect 8622 3780 8680 3836
rect 8736 3780 8794 3836
rect 8850 3780 8983 3836
rect 8499 3587 8983 3780
rect 8499 3535 8557 3587
rect 8609 3535 8655 3587
rect 8707 3535 8750 3587
rect 8802 3535 8855 3587
rect 8907 3535 8983 3587
rect 8499 3423 8983 3535
rect 9531 4252 9720 5454
rect 16714 5441 16974 5512
rect 16714 5389 16734 5441
rect 16786 5389 16812 5441
rect 16864 5389 16905 5441
rect 16957 5389 16974 5441
rect 24642 5504 24831 5527
rect 24642 5452 24671 5504
rect 24723 5452 24766 5504
rect 24818 5452 24831 5504
rect 16714 4464 16974 5389
rect 16714 4412 16758 4464
rect 16810 4412 16881 4464
rect 16933 4412 16974 4464
rect 16714 4368 16974 4412
rect 23555 5291 24022 5391
rect 23555 5239 23593 5291
rect 23645 5239 23696 5291
rect 23748 5239 23779 5291
rect 23831 5239 23880 5291
rect 23932 5239 23967 5291
rect 24019 5239 24022 5291
rect 9531 4200 9556 4252
rect 9608 4200 9652 4252
rect 9704 4200 9720 4252
rect 9531 3369 9720 4200
rect 17139 4107 17345 4152
rect 17139 4103 17277 4107
rect 17139 4051 17172 4103
rect 17224 4055 17277 4103
rect 17329 4055 17345 4107
rect 17224 4051 17345 4055
rect 9531 3317 9556 3369
rect 9608 3367 9720 3369
rect 9608 3317 9636 3367
rect 9531 3315 9636 3317
rect 9688 3315 9720 3367
rect 15920 3916 16273 3962
rect 15920 3915 16148 3916
rect 15920 3863 15971 3915
rect 16023 3863 16055 3915
rect 16107 3864 16148 3915
rect 16200 3864 16273 3916
rect 16107 3863 16273 3864
rect 15920 3505 16273 3863
rect 17139 3686 17345 4051
rect 17139 3634 17176 3686
rect 17228 3681 17345 3686
rect 17228 3634 17270 3681
rect 17139 3629 17270 3634
rect 17322 3629 17345 3681
rect 17139 3608 17345 3629
rect 17139 3606 17270 3608
rect 17139 3554 17176 3606
rect 17228 3556 17270 3606
rect 17322 3556 17345 3608
rect 17228 3554 17345 3556
rect 17139 3525 17345 3554
rect 23555 3976 24022 5239
rect 23555 3920 23605 3976
rect 23661 3920 23709 3976
rect 23765 3920 23813 3976
rect 23869 3920 23917 3976
rect 23973 3920 24022 3976
rect 23555 3860 24022 3920
rect 23555 3804 23605 3860
rect 23661 3804 23709 3860
rect 23765 3804 23813 3860
rect 23869 3804 23917 3860
rect 23973 3804 24022 3860
rect 23555 3744 24022 3804
rect 23555 3688 23605 3744
rect 23661 3688 23709 3744
rect 23765 3688 23813 3744
rect 23869 3688 23917 3744
rect 23973 3688 24022 3744
rect 23555 3592 24022 3688
rect 23555 3540 23607 3592
rect 23659 3540 23707 3592
rect 23759 3540 23806 3592
rect 23858 3540 23909 3592
rect 23961 3540 24022 3592
rect 15920 3449 15960 3505
rect 16016 3449 16068 3505
rect 16124 3449 16176 3505
rect 16232 3449 16273 3505
rect 15920 3411 16273 3449
rect 23555 3440 24022 3540
rect 24642 4250 24831 5452
rect 32647 5464 32982 5507
rect 32647 5412 32693 5464
rect 32745 5412 32806 5464
rect 32858 5412 32907 5464
rect 32959 5412 32982 5464
rect 32647 4844 32982 5412
rect 39733 5506 39920 5525
rect 39733 5454 39748 5506
rect 39800 5454 39850 5506
rect 39902 5454 39920 5506
rect 32647 4841 32808 4844
rect 32647 4789 32705 4841
rect 32757 4792 32808 4841
rect 32860 4792 32909 4844
rect 32961 4792 32982 4844
rect 32757 4789 32982 4792
rect 32647 4757 32982 4789
rect 38671 5292 38971 5389
rect 38671 5287 38898 5292
rect 38671 5235 38725 5287
rect 38777 5235 38813 5287
rect 38865 5240 38898 5287
rect 38950 5240 38971 5292
rect 38865 5235 38971 5240
rect 33418 4435 33957 4458
rect 33418 4383 33486 4435
rect 33538 4383 33646 4435
rect 33698 4383 33779 4435
rect 33831 4383 33892 4435
rect 33944 4383 33957 4435
rect 24642 4243 24766 4250
rect 24642 4191 24667 4243
rect 24719 4198 24766 4243
rect 24818 4198 24831 4250
rect 24719 4191 24831 4198
rect 15920 3355 15960 3411
rect 16016 3355 16068 3411
rect 16124 3355 16176 3411
rect 16232 3355 16273 3411
rect 15920 3329 16273 3355
rect 24642 3384 24831 4191
rect 32609 4294 33034 4312
rect 32609 4291 32868 4294
rect 32609 4289 32757 4291
rect 32609 4237 32661 4289
rect 32713 4239 32757 4289
rect 32809 4242 32868 4291
rect 32920 4291 33034 4294
rect 32920 4242 32960 4291
rect 32809 4239 32960 4242
rect 33012 4239 33034 4291
rect 32713 4237 33034 4239
rect 32609 3625 33034 4237
rect 33418 3867 33957 4383
rect 33418 3815 33475 3867
rect 33527 3815 33619 3867
rect 33671 3815 33763 3867
rect 33815 3815 33957 3867
rect 33418 3783 33957 3815
rect 33418 3731 33474 3783
rect 33526 3731 33618 3783
rect 33670 3731 33762 3783
rect 33814 3731 33957 3783
rect 33418 3657 33957 3731
rect 38671 4325 38971 5235
rect 38671 4269 38692 4325
rect 38748 4269 38786 4325
rect 38842 4269 38880 4325
rect 38936 4269 38971 4325
rect 38671 4237 38971 4269
rect 38671 4181 38692 4237
rect 38748 4181 38786 4237
rect 38842 4181 38880 4237
rect 38936 4181 38971 4237
rect 38671 4149 38971 4181
rect 38671 4093 38692 4149
rect 38748 4093 38786 4149
rect 38842 4093 38880 4149
rect 38936 4093 38971 4149
rect 32609 3569 32655 3625
rect 32711 3569 32780 3625
rect 32836 3569 32905 3625
rect 32961 3569 33034 3625
rect 32609 3529 33034 3569
rect 32609 3473 32655 3529
rect 32711 3473 32780 3529
rect 32836 3473 32905 3529
rect 32961 3473 33034 3529
rect 32609 3441 33034 3473
rect 38671 3586 38971 4093
rect 38671 3534 38715 3586
rect 38767 3534 38803 3586
rect 38855 3582 38971 3586
rect 38855 3534 38901 3582
rect 38671 3530 38901 3534
rect 38953 3530 38971 3582
rect 38671 3437 38971 3530
rect 39733 4408 39920 5454
rect 46862 5441 47081 5494
rect 46862 5389 46885 5441
rect 46937 5389 46968 5441
rect 47020 5389 47081 5441
rect 46862 4617 47081 5389
rect 46862 4616 46981 4617
rect 46862 4564 46891 4616
rect 46943 4565 46981 4616
rect 47033 4565 47081 4617
rect 46943 4564 47081 4565
rect 46862 4529 47081 4564
rect 54837 5479 55026 5502
rect 54837 5427 54866 5479
rect 54918 5427 54961 5479
rect 55013 5427 55026 5479
rect 39733 4407 39854 4408
rect 39733 4355 39751 4407
rect 39803 4356 39854 4407
rect 39906 4356 39920 4408
rect 39803 4355 39920 4356
rect 24642 3332 24672 3384
rect 24724 3332 24755 3384
rect 24807 3332 24831 3384
rect 24642 3319 24831 3332
rect 39733 3374 39920 4355
rect 54837 4408 55026 5427
rect 54837 4403 54955 4408
rect 54837 4351 54864 4403
rect 54916 4356 54955 4403
rect 55007 4356 55026 4408
rect 54916 4351 55026 4356
rect 47281 4267 47487 4312
rect 47281 4263 47419 4267
rect 47281 4211 47314 4263
rect 47366 4215 47419 4263
rect 47471 4215 47487 4267
rect 47366 4211 47487 4215
rect 47281 3869 47487 4211
rect 47281 3866 47411 3869
rect 47281 3814 47322 3866
rect 47374 3817 47411 3866
rect 47463 3817 47487 3869
rect 47374 3814 47487 3817
rect 47281 3790 47487 3814
rect 47281 3738 47322 3790
rect 47374 3738 47415 3790
rect 47467 3738 47487 3790
rect 47281 3695 47487 3738
rect 48289 4077 48703 4099
rect 48289 4076 48418 4077
rect 48289 4024 48326 4076
rect 48378 4025 48418 4076
rect 48470 4076 48703 4077
rect 48470 4025 48508 4076
rect 48378 4024 48508 4025
rect 48560 4075 48703 4076
rect 48560 4024 48596 4075
rect 48289 4023 48596 4024
rect 48648 4023 48703 4075
rect 39733 3322 39750 3374
rect 39802 3322 39841 3374
rect 39893 3322 39920 3374
rect 9531 3297 9720 3315
rect 39733 3314 39920 3322
rect 48289 3478 48703 4023
rect 48289 3422 48326 3478
rect 48382 3422 48419 3478
rect 48475 3422 48512 3478
rect 48568 3422 48605 3478
rect 48661 3422 48703 3478
rect 48289 3396 48703 3422
rect 48289 3340 48326 3396
rect 48382 3340 48419 3396
rect 48475 3340 48512 3396
rect 48568 3340 48605 3396
rect 48661 3340 48703 3396
rect 48289 3303 48703 3340
rect 54837 3359 55026 4351
rect 55602 5284 56023 5389
rect 55602 5232 55641 5284
rect 55693 5232 55735 5284
rect 55787 5232 55812 5284
rect 55864 5283 55966 5284
rect 55864 5232 55892 5283
rect 55602 5231 55892 5232
rect 55944 5232 55966 5283
rect 56018 5232 56023 5284
rect 55944 5231 56023 5232
rect 55602 3870 56023 5231
rect 55602 3814 55639 3870
rect 55695 3814 55743 3870
rect 55799 3814 55847 3870
rect 55903 3814 55951 3870
rect 56007 3814 56023 3870
rect 55602 3780 56023 3814
rect 55602 3724 55639 3780
rect 55695 3724 55743 3780
rect 55799 3724 55847 3780
rect 55903 3724 55951 3780
rect 56007 3724 56023 3780
rect 55602 3583 56023 3724
rect 55602 3531 55637 3583
rect 55689 3531 55725 3583
rect 55777 3531 55808 3583
rect 55860 3531 55895 3583
rect 55947 3531 56023 3583
rect 55602 3439 56023 3531
rect 54837 3307 54867 3359
rect 54919 3307 54950 3359
rect 55002 3307 55026 3359
rect 54837 3294 55026 3307
rect 932 3058 2360 3248
rect 932 2804 1818 3058
rect 932 2718 2340 2804
rect 932 2710 1818 2718
rect 64230 2204 64344 6624
rect 208 2168 603 2204
rect 1752 2168 2342 2204
rect 62578 2168 64344 2204
rect 208 2156 322 2168
rect 64230 2160 64344 2168
rect 2311 1168 2355 1486
rect 4199 1168 4243 1486
rect 6087 1168 6131 1486
rect 7975 1168 8019 1486
rect 9863 1168 9907 1486
rect 11751 1168 11795 1486
rect 13639 1168 13683 1486
rect 15527 1168 15571 1486
rect 17415 1168 17459 1486
rect 19303 1168 19347 1486
rect 21191 1168 21235 1486
rect 23079 1168 23123 1486
rect 24967 1168 25011 1486
rect 26855 1168 26899 1486
rect 28743 1168 28787 1486
rect 30631 1168 30675 1486
rect 32519 1168 32563 1486
rect 34407 1168 34451 1486
rect 36295 1168 36339 1486
rect 38183 1168 38227 1486
rect 40071 1168 40115 1486
rect 41959 1168 42003 1486
rect 43847 1168 43891 1486
rect 45735 1168 45779 1486
rect 47623 1168 47667 1486
rect 49511 1168 49555 1486
rect 51399 1168 51443 1486
rect 53287 1168 53331 1486
rect 55175 1168 55219 1486
rect 57063 1168 57107 1486
rect 58951 1366 58995 1486
rect 58951 1168 58997 1366
rect 422 22 467 1168
rect 2310 22 2355 1168
rect 4198 22 4243 1168
rect 6086 22 6131 1168
rect 7974 22 8019 1168
rect 9862 22 9907 1168
rect 11750 22 11795 1168
rect 13638 22 13683 1168
rect 15526 22 15571 1168
rect 17414 22 17459 1168
rect 19302 22 19347 1168
rect 21190 22 21235 1168
rect 23078 22 23123 1168
rect 24966 22 25011 1168
rect 26854 22 26899 1168
rect 28742 22 28787 1168
rect 30630 22 30675 1168
rect 32518 22 32563 1168
rect 34406 22 34451 1168
rect 36294 22 36339 1168
rect 38182 22 38227 1168
rect 40070 22 40115 1168
rect 41958 22 42003 1168
rect 43846 22 43891 1168
rect 45734 22 45779 1168
rect 47622 22 47667 1168
rect 49510 22 49555 1168
rect 51398 22 51443 1168
rect 53286 22 53331 1168
rect 55174 22 55219 1168
rect 57062 22 57107 1168
rect 58950 468 58997 1168
rect 58950 22 58995 468
rect 60827 0 60883 1486
<< via2 >>
rect 8566 4010 8622 4066
rect 8680 4010 8736 4066
rect 8794 4010 8850 4066
rect 8566 3895 8622 3951
rect 8680 3895 8736 3951
rect 8794 3895 8850 3951
rect 8566 3780 8622 3836
rect 8680 3780 8736 3836
rect 8794 3780 8850 3836
rect 23605 3920 23661 3976
rect 23709 3920 23765 3976
rect 23813 3920 23869 3976
rect 23917 3920 23973 3976
rect 23605 3804 23661 3860
rect 23709 3804 23765 3860
rect 23813 3804 23869 3860
rect 23917 3804 23973 3860
rect 23605 3688 23661 3744
rect 23709 3688 23765 3744
rect 23813 3688 23869 3744
rect 23917 3688 23973 3744
rect 15960 3449 16016 3505
rect 16068 3449 16124 3505
rect 16176 3449 16232 3505
rect 15960 3355 16016 3411
rect 16068 3355 16124 3411
rect 16176 3355 16232 3411
rect 38692 4269 38748 4325
rect 38786 4269 38842 4325
rect 38880 4269 38936 4325
rect 38692 4181 38748 4237
rect 38786 4181 38842 4237
rect 38880 4181 38936 4237
rect 38692 4093 38748 4149
rect 38786 4093 38842 4149
rect 38880 4093 38936 4149
rect 32655 3569 32711 3625
rect 32780 3569 32836 3625
rect 32905 3569 32961 3625
rect 32655 3473 32711 3529
rect 32780 3473 32836 3529
rect 32905 3473 32961 3529
rect 48326 3422 48382 3478
rect 48419 3422 48475 3478
rect 48512 3422 48568 3478
rect 48605 3422 48661 3478
rect 48326 3340 48382 3396
rect 48419 3340 48475 3396
rect 48512 3340 48568 3396
rect 48605 3340 48661 3396
rect 55639 3814 55695 3870
rect 55743 3814 55799 3870
rect 55847 3814 55903 3870
rect 55951 3814 56007 3870
rect 55639 3724 55695 3780
rect 55743 3724 55799 3780
rect 55847 3724 55903 3780
rect 55951 3724 56007 3780
<< metal3 >>
rect 3463 5966 4358 6012
rect 3463 5965 3747 5966
rect 3463 5787 3575 5965
rect 3681 5788 3747 5965
rect 3853 5965 4358 5966
rect 3853 5788 3921 5965
rect 3681 5787 3921 5788
rect 4027 5787 4358 5965
rect 3463 5758 4358 5787
rect 38669 4325 38973 4339
rect 38669 4269 38692 4325
rect 38748 4269 38786 4325
rect 38842 4269 38880 4325
rect 38936 4269 38973 4325
rect 38669 4237 38973 4269
rect 38669 4181 38692 4237
rect 38748 4226 38786 4237
rect 38842 4227 38880 4237
rect 38936 4227 38973 4237
rect 38842 4181 38859 4227
rect 38669 4149 38705 4181
rect 38792 4149 38859 4181
rect 8565 4092 8907 4125
rect 38669 4093 38692 4149
rect 38842 4115 38859 4149
rect 38946 4115 38973 4227
rect 38748 4093 38786 4114
rect 38842 4093 38880 4115
rect 38936 4093 38973 4115
rect 8497 4066 8986 4092
rect 38669 4073 38973 4093
rect 8497 4010 8566 4066
rect 8622 4010 8680 4066
rect 8736 4010 8794 4066
rect 8850 4010 8986 4066
rect 8497 3951 8986 4010
rect 8497 3923 8566 3951
rect 8622 3923 8680 3951
rect 8736 3929 8794 3951
rect 8850 3929 8986 3951
rect 8497 3832 8563 3923
rect 8649 3895 8680 3923
rect 8850 3895 8859 3929
rect 8649 3838 8714 3895
rect 8800 3838 8859 3895
rect 8945 3838 8986 3929
rect 8649 3836 8986 3838
rect 8649 3832 8680 3836
rect 8497 3780 8566 3832
rect 8622 3780 8680 3832
rect 8736 3780 8794 3836
rect 8850 3780 8986 3836
rect 8497 3725 8986 3780
rect 23555 3976 24022 4030
rect 23555 3933 23605 3976
rect 23661 3933 23709 3976
rect 23555 3849 23603 3933
rect 23696 3920 23709 3933
rect 23765 3933 23813 3976
rect 23765 3920 23770 3933
rect 23869 3920 23917 3976
rect 23973 3920 24022 3976
rect 23696 3860 23770 3920
rect 23863 3860 24022 3920
rect 23696 3849 23709 3860
rect 23555 3804 23605 3849
rect 23661 3804 23709 3849
rect 23765 3849 23770 3860
rect 23765 3804 23813 3849
rect 23869 3804 23917 3860
rect 23973 3804 24022 3860
rect 23555 3772 24022 3804
rect 23555 3688 23603 3772
rect 23696 3744 23770 3772
rect 23863 3744 24022 3772
rect 23696 3688 23709 3744
rect 23765 3688 23770 3744
rect 23869 3688 23917 3744
rect 23973 3688 24022 3744
rect 55602 3877 56024 3898
rect 55602 3870 55646 3877
rect 55730 3870 55767 3877
rect 55851 3870 55905 3877
rect 55989 3870 56024 3877
rect 55602 3814 55639 3870
rect 55730 3814 55743 3870
rect 55903 3814 55905 3870
rect 56007 3814 56024 3870
rect 55602 3780 55646 3814
rect 55730 3780 55767 3814
rect 55851 3780 55905 3814
rect 55989 3780 56024 3814
rect 55602 3724 55639 3780
rect 55730 3724 55743 3780
rect 55903 3724 55905 3780
rect 56007 3724 56024 3780
rect 55602 3719 55646 3724
rect 55730 3719 55767 3724
rect 55851 3719 55905 3724
rect 55989 3719 56024 3724
rect 55602 3690 56024 3719
rect 23555 3644 24022 3688
rect 32607 3625 33032 3663
rect 32607 3586 32655 3625
rect 32711 3586 32780 3625
rect 32836 3586 32905 3625
rect 32961 3586 33032 3625
rect 15920 3505 16273 3528
rect 15920 3457 15960 3505
rect 16016 3457 16068 3505
rect 16124 3457 16176 3505
rect 15920 3388 15944 3457
rect 16021 3388 16047 3457
rect 16124 3388 16150 3457
rect 16232 3449 16273 3505
rect 16227 3411 16273 3449
rect 32607 3474 32653 3586
rect 32740 3474 32772 3586
rect 32859 3474 32891 3586
rect 32978 3474 33032 3586
rect 32607 3473 32655 3474
rect 32711 3473 32780 3474
rect 32836 3473 32905 3474
rect 32961 3473 33032 3474
rect 32607 3436 33032 3473
rect 48289 3502 48704 3545
rect 48289 3501 48467 3502
rect 48289 3478 48327 3501
rect 48411 3478 48467 3501
rect 48551 3478 48595 3502
rect 15920 3355 15960 3388
rect 16016 3355 16068 3388
rect 16124 3355 16176 3388
rect 16232 3355 16273 3411
rect 15920 3329 16273 3355
rect 48289 3422 48326 3478
rect 48411 3422 48419 3478
rect 48568 3422 48595 3478
rect 48289 3396 48327 3422
rect 48411 3396 48467 3422
rect 48551 3396 48595 3422
rect 48289 3340 48326 3396
rect 48411 3343 48419 3396
rect 48568 3344 48595 3396
rect 48679 3344 48704 3502
rect 48382 3340 48419 3343
rect 48475 3340 48512 3344
rect 48568 3340 48605 3344
rect 48661 3340 48704 3344
rect 48289 3304 48704 3340
<< via3 >>
rect 4809 7905 4915 8083
rect 5018 7904 5124 8082
rect 5184 7904 5290 8082
rect 5364 7906 5470 8084
rect 21438 7922 21544 8100
rect 21654 7922 21760 8100
rect 21870 7922 21976 8100
rect 29930 7921 30036 8099
rect 30146 7921 30252 8099
rect 30362 7921 30468 8099
rect 43458 7927 43564 8105
rect 43674 7927 43780 8105
rect 43890 7927 43996 8105
rect 59943 7920 60049 8098
rect 60159 7920 60265 8098
rect 60375 7920 60481 8098
rect 3575 5787 3681 5965
rect 3747 5788 3853 5966
rect 3921 5787 4027 5965
rect 19903 5808 20009 5986
rect 20119 5808 20225 5986
rect 20335 5808 20441 5986
rect 28411 5800 28517 5978
rect 28627 5800 28733 5978
rect 28843 5800 28949 5978
rect 41883 5795 41989 5973
rect 42099 5795 42205 5973
rect 42315 5795 42421 5973
rect 58434 5787 58540 5965
rect 58650 5787 58756 5965
rect 58866 5787 58972 5965
rect 38705 4181 38748 4226
rect 38748 4181 38786 4226
rect 38786 4181 38792 4226
rect 38859 4181 38880 4227
rect 38880 4181 38936 4227
rect 38936 4181 38946 4227
rect 38705 4149 38792 4181
rect 38859 4149 38946 4181
rect 38705 4114 38748 4149
rect 38748 4114 38786 4149
rect 38786 4114 38792 4149
rect 38859 4115 38880 4149
rect 38880 4115 38936 4149
rect 38936 4115 38946 4149
rect 8563 3895 8566 3923
rect 8566 3895 8622 3923
rect 8622 3895 8649 3923
rect 8714 3895 8736 3929
rect 8736 3895 8794 3929
rect 8794 3895 8800 3929
rect 8563 3836 8649 3895
rect 8714 3838 8800 3895
rect 8859 3838 8945 3929
rect 8563 3832 8566 3836
rect 8566 3832 8622 3836
rect 8622 3832 8649 3836
rect 23603 3920 23605 3933
rect 23605 3920 23661 3933
rect 23661 3920 23696 3933
rect 23770 3920 23813 3933
rect 23813 3920 23863 3933
rect 23603 3860 23696 3920
rect 23770 3860 23863 3920
rect 23603 3849 23605 3860
rect 23605 3849 23661 3860
rect 23661 3849 23696 3860
rect 23770 3849 23813 3860
rect 23813 3849 23863 3860
rect 23603 3744 23696 3772
rect 23770 3744 23863 3772
rect 23603 3688 23605 3744
rect 23605 3688 23661 3744
rect 23661 3688 23696 3744
rect 23770 3688 23813 3744
rect 23813 3688 23863 3744
rect 55646 3870 55730 3877
rect 55767 3870 55851 3877
rect 55905 3870 55989 3877
rect 55646 3814 55695 3870
rect 55695 3814 55730 3870
rect 55767 3814 55799 3870
rect 55799 3814 55847 3870
rect 55847 3814 55851 3870
rect 55905 3814 55951 3870
rect 55951 3814 55989 3870
rect 55646 3780 55730 3814
rect 55767 3780 55851 3814
rect 55905 3780 55989 3814
rect 55646 3724 55695 3780
rect 55695 3724 55730 3780
rect 55767 3724 55799 3780
rect 55799 3724 55847 3780
rect 55847 3724 55851 3780
rect 55905 3724 55951 3780
rect 55951 3724 55989 3780
rect 55646 3719 55730 3724
rect 55767 3719 55851 3724
rect 55905 3719 55989 3724
rect 15944 3449 15960 3457
rect 15960 3449 16016 3457
rect 16016 3449 16021 3457
rect 15944 3411 16021 3449
rect 15944 3388 15960 3411
rect 15960 3388 16016 3411
rect 16016 3388 16021 3411
rect 16047 3449 16068 3457
rect 16068 3449 16124 3457
rect 16047 3411 16124 3449
rect 16047 3388 16068 3411
rect 16068 3388 16124 3411
rect 16150 3449 16176 3457
rect 16176 3449 16227 3457
rect 16150 3411 16227 3449
rect 32653 3569 32655 3586
rect 32655 3569 32711 3586
rect 32711 3569 32740 3586
rect 32653 3529 32740 3569
rect 32653 3474 32655 3529
rect 32655 3474 32711 3529
rect 32711 3474 32740 3529
rect 32772 3569 32780 3586
rect 32780 3569 32836 3586
rect 32836 3569 32859 3586
rect 32772 3529 32859 3569
rect 32772 3474 32780 3529
rect 32780 3474 32836 3529
rect 32836 3474 32859 3529
rect 32891 3569 32905 3586
rect 32905 3569 32961 3586
rect 32961 3569 32978 3586
rect 32891 3529 32978 3569
rect 32891 3474 32905 3529
rect 32905 3474 32961 3529
rect 32961 3474 32978 3529
rect 48327 3478 48411 3501
rect 48467 3478 48551 3502
rect 48595 3478 48679 3502
rect 16150 3388 16176 3411
rect 16176 3388 16227 3411
rect 48327 3422 48382 3478
rect 48382 3422 48411 3478
rect 48467 3422 48475 3478
rect 48475 3422 48512 3478
rect 48512 3422 48551 3478
rect 48595 3422 48605 3478
rect 48605 3422 48661 3478
rect 48661 3422 48679 3478
rect 48327 3396 48411 3422
rect 48467 3396 48551 3422
rect 48595 3396 48679 3422
rect 48327 3343 48382 3396
rect 48382 3343 48411 3396
rect 48467 3344 48475 3396
rect 48475 3344 48512 3396
rect 48512 3344 48551 3396
rect 48595 3344 48605 3396
rect 48605 3344 48661 3396
rect 48661 3344 48679 3396
rect 3577 2839 3683 3017
rect 3782 2841 3888 3019
rect 3981 2841 4087 3019
rect 19894 2857 20000 3035
rect 20110 2857 20216 3035
rect 20326 2857 20432 3035
rect 28416 2852 28522 3030
rect 28632 2852 28738 3030
rect 28848 2852 28954 3030
rect 41919 2854 42025 3032
rect 42135 2854 42241 3032
rect 42351 2854 42457 3032
rect 58414 2865 58520 3043
rect 58630 2865 58736 3043
rect 58846 2865 58952 3043
rect 4823 728 4929 906
rect 5044 728 5150 906
rect 5253 728 5359 906
rect 5427 728 5533 906
rect 8551 760 8637 851
rect 8699 760 8785 851
rect 8847 760 8933 851
rect 16070 834 16147 903
rect 16093 715 16170 784
rect 21456 727 21562 905
rect 21672 727 21778 905
rect 21888 727 21994 905
rect 23608 755 23704 863
rect 23741 755 23837 863
rect 23874 755 23970 863
rect 29885 732 29991 910
rect 30101 732 30207 910
rect 30317 732 30423 910
rect 32674 742 32761 854
rect 32797 742 32884 854
rect 32929 742 33016 854
rect 38703 739 38790 851
rect 38872 739 38959 851
rect 43403 722 43509 900
rect 43619 722 43725 900
rect 43835 722 43941 900
rect 48329 726 48413 884
rect 48442 726 48526 884
rect 48557 726 48641 884
rect 55652 736 55736 894
rect 55771 736 55855 894
rect 55900 736 55984 894
rect 59915 717 60021 895
rect 60131 717 60237 895
rect 60347 717 60453 895
<< metal4 >>
rect 3431 5966 4237 8265
rect 3431 5965 3747 5966
rect 3431 5787 3575 5965
rect 3681 5788 3747 5965
rect 3853 5965 4237 5966
rect 3853 5788 3921 5965
rect 3681 5787 3921 5788
rect 4027 5787 4237 5965
rect 3431 3019 4237 5787
rect 3431 3017 3782 3019
rect 3431 2839 3577 3017
rect 3683 2841 3782 3017
rect 3888 2841 3981 3019
rect 4087 2841 4237 3019
rect 3683 2839 4237 2841
rect 3431 559 4237 2839
rect 4774 8084 5580 8266
rect 4774 8083 5364 8084
rect 4774 7905 4809 8083
rect 4915 8082 5364 8083
rect 4915 7905 5018 8082
rect 4774 7904 5018 7905
rect 5124 7904 5184 8082
rect 5290 7906 5364 8082
rect 5470 7906 5580 8084
rect 5290 7904 5580 7906
rect 4774 906 5580 7904
rect 19774 5986 20580 8266
rect 19774 5808 19903 5986
rect 20009 5808 20119 5986
rect 20225 5808 20335 5986
rect 20441 5808 20580 5986
rect 4774 728 4823 906
rect 4929 728 5044 906
rect 5150 728 5253 906
rect 5359 728 5427 906
rect 5533 728 5580 906
rect 4774 560 5580 728
rect 8505 3929 8974 4044
rect 8505 3923 8714 3929
rect 8505 3832 8563 3923
rect 8649 3838 8714 3923
rect 8800 3838 8859 3929
rect 8945 3838 8974 3929
rect 8649 3832 8974 3838
rect 8505 851 8974 3832
rect 15920 3457 16274 3529
rect 15920 3388 15944 3457
rect 16021 3388 16047 3457
rect 16124 3388 16150 3457
rect 16227 3388 16274 3457
rect 15920 3328 16274 3388
rect 8505 760 8551 851
rect 8637 760 8699 851
rect 8785 760 8847 851
rect 8933 760 8974 851
rect 8505 661 8974 760
rect 15996 903 16197 3328
rect 15996 834 16070 903
rect 16147 834 16197 903
rect 15996 784 16197 834
rect 15996 715 16093 784
rect 16170 715 16197 784
rect 15996 636 16197 715
rect 19774 3035 20580 5808
rect 19774 2857 19894 3035
rect 20000 2857 20110 3035
rect 20216 2857 20326 3035
rect 20432 2857 20580 3035
rect 19774 560 20580 2857
rect 21274 8100 22080 8266
rect 21274 7922 21438 8100
rect 21544 7922 21654 8100
rect 21760 7922 21870 8100
rect 21976 7922 22080 8100
rect 21274 905 22080 7922
rect 28274 5978 29080 8266
rect 28274 5800 28411 5978
rect 28517 5800 28627 5978
rect 28733 5800 28843 5978
rect 28949 5800 29080 5978
rect 21274 727 21456 905
rect 21562 727 21672 905
rect 21778 727 21888 905
rect 21994 727 22080 905
rect 21274 560 22080 727
rect 23555 3933 24022 4058
rect 23555 3849 23603 3933
rect 23696 3849 23770 3933
rect 23863 3849 24022 3933
rect 23555 3772 24022 3849
rect 23555 3688 23603 3772
rect 23696 3688 23770 3772
rect 23863 3688 24022 3772
rect 23555 863 24022 3688
rect 23555 755 23608 863
rect 23704 755 23741 863
rect 23837 755 23874 863
rect 23970 755 24022 863
rect 23555 686 24022 755
rect 28274 3030 29080 5800
rect 28274 2852 28416 3030
rect 28522 2852 28632 3030
rect 28738 2852 28848 3030
rect 28954 2852 29080 3030
rect 28274 560 29080 2852
rect 29774 8099 30580 8266
rect 29774 7921 29930 8099
rect 30036 7921 30146 8099
rect 30252 7921 30362 8099
rect 30468 7921 30580 8099
rect 29774 910 30580 7921
rect 41774 5973 42580 8266
rect 41774 5795 41883 5973
rect 41989 5795 42099 5973
rect 42205 5795 42315 5973
rect 42421 5795 42580 5973
rect 38669 4227 38974 4384
rect 38669 4226 38859 4227
rect 38669 4114 38705 4226
rect 38792 4115 38859 4226
rect 38946 4115 38974 4227
rect 38792 4114 38974 4115
rect 29774 732 29885 910
rect 29991 732 30101 910
rect 30207 732 30317 910
rect 30423 732 30580 910
rect 29774 560 30580 732
rect 32607 3586 33032 3665
rect 32607 3474 32653 3586
rect 32740 3474 32772 3586
rect 32859 3474 32891 3586
rect 32978 3474 33032 3586
rect 32607 854 33032 3474
rect 32607 742 32674 854
rect 32761 742 32797 854
rect 32884 742 32929 854
rect 33016 742 33032 854
rect 32607 700 33032 742
rect 38669 851 38974 4114
rect 38669 739 38703 851
rect 38790 739 38872 851
rect 38959 739 38974 851
rect 38669 691 38974 739
rect 41774 3032 42580 5795
rect 41774 2854 41919 3032
rect 42025 2854 42135 3032
rect 42241 2854 42351 3032
rect 42457 2854 42580 3032
rect 41774 560 42580 2854
rect 43274 8105 44080 8266
rect 43274 7927 43458 8105
rect 43564 7927 43674 8105
rect 43780 7927 43890 8105
rect 43996 7927 44080 8105
rect 43274 900 44080 7927
rect 58274 5965 59080 8266
rect 58274 5787 58434 5965
rect 58540 5787 58650 5965
rect 58756 5787 58866 5965
rect 58972 5787 59080 5965
rect 55602 3877 56027 3900
rect 55602 3719 55646 3877
rect 55730 3719 55767 3877
rect 55851 3719 55905 3877
rect 55989 3719 56027 3877
rect 43274 722 43403 900
rect 43509 722 43619 900
rect 43725 722 43835 900
rect 43941 722 44080 900
rect 43274 560 44080 722
rect 48289 3502 48703 3591
rect 48289 3501 48467 3502
rect 48289 3343 48327 3501
rect 48411 3344 48467 3501
rect 48551 3344 48595 3502
rect 48679 3344 48703 3502
rect 48411 3343 48703 3344
rect 48289 884 48703 3343
rect 48289 726 48329 884
rect 48413 726 48442 884
rect 48526 726 48557 884
rect 48641 726 48703 884
rect 48289 638 48703 726
rect 55602 894 56027 3719
rect 55602 736 55652 894
rect 55736 736 55771 894
rect 55855 736 55900 894
rect 55984 736 56027 894
rect 55602 650 56027 736
rect 58274 3043 59080 5787
rect 58274 2865 58414 3043
rect 58520 2865 58630 3043
rect 58736 2865 58846 3043
rect 58952 2865 59080 3043
rect 58274 560 59080 2865
rect 59774 8098 60580 8266
rect 59774 7920 59943 8098
rect 60049 7920 60159 8098
rect 60265 7920 60375 8098
rect 60481 7920 60580 8098
rect 59774 895 60580 7920
rect 59774 717 59915 895
rect 60021 717 60131 895
rect 60237 717 60347 895
rect 60453 717 60580 895
rect 59774 560 60580 717
use brbufhalf  brbufhalf_0
timestamp 1654663570
transform 1 0 5843 0 1 -1834
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_1
timestamp 1654663570
transform 1 0 36045 0 1 -1834
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_2
timestamp 1654663570
transform -1 0 58721 0 -1 10662
box -3552 2527 26658 5446
use brbufhalf_64  brbufhalf_64_0
timestamp 1655064284
transform -1 0 28519 0 -1 10662
box -3552 2527 26308 5446
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1653697408
transform 1 0 32318 0 1 4265
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654402208
transform 1 0 17460 0 1 3889
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654402208
transform 1 0 15530 0 1 3889
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1654402208
transform 1 0 32866 0 1 4265
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1654402208
transform 1 0 47602 0 1 4049
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1654402208
transform 1 0 45672 0 1 4049
box -38 -48 1510 592
use unitcell2buf  unitcell2buf_13
timestamp 1654643405
transform 1 0 977 0 1 1878
box -574 -1185 1322 1192
<< labels >>
flabel metal1 62673 1474 62895 1552 1 FreeSans 1600 0 0 0 OUT
port 3 n
flabel metal4 3431 559 4237 8265 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 4774 560 5580 8266 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 19774 560 20580 8266 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 21274 560 22080 8266 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 28274 560 29080 8266 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 29774 560 30580 8266 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 41774 560 42580 8266 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 43274 560 44080 8266 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 58274 560 59080 8266 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 59774 560 60580 8266 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal1 0 4626 534 4690 1 FreeSans 1600 0 0 0 RESET
port 71 n
flabel metal2 62209 7342 62253 8498 1 FreeSans 1600 0 0 0 C[0]
port 72 n
flabel metal2 60321 7342 60365 8498 1 FreeSans 1600 0 0 0 C[1]
port 73 n
flabel metal2 58433 7342 58477 8498 1 FreeSans 1600 0 0 0 C[2]
port 74 n
flabel metal2 56545 7342 56589 8498 1 FreeSans 1600 0 0 0 C[3]
port 75 n
flabel metal2 54657 7342 54701 8498 1 FreeSans 1600 0 0 0 C[4]
port 76 n
flabel metal2 52769 7342 52813 8498 1 FreeSans 1600 0 0 0 C[5]
port 77 n
flabel metal2 50881 7342 50925 8498 1 FreeSans 1600 0 0 0 C[6]
port 78 n
flabel metal2 48993 7342 49037 8498 1 FreeSans 1600 0 0 0 C[7]
port 79 n
flabel metal2 47105 7342 47149 8498 1 FreeSans 1600 0 0 0 C[8]
port 80 n
flabel metal2 45217 7342 45261 8498 1 FreeSans 1600 0 0 0 C[9]
port 81 n
flabel metal2 43329 7342 43373 8498 1 FreeSans 1600 0 0 0 C[10]
port 82 n
flabel metal2 41441 7342 41485 8498 1 FreeSans 1600 0 0 0 C[11]
port 83 n
flabel metal2 39553 7342 39597 8498 1 FreeSans 1600 0 0 0 C[12]
port 84 n
flabel metal2 37665 7342 37709 8498 1 FreeSans 1600 0 0 0 C[13]
port 85 n
flabel metal2 35777 7342 35821 8498 1 FreeSans 1600 0 0 0 C[14]
port 86 n
flabel metal2 33889 7342 33933 8498 1 FreeSans 1600 0 0 0 C[15]
port 87 n
flabel metal2 32001 7342 32045 8498 1 FreeSans 1600 0 0 0 C[16]
port 88 n
flabel metal2 30113 7342 30157 8498 1 FreeSans 1600 0 0 0 C[17]
port 89 n
flabel metal2 28225 7342 28269 8498 1 FreeSans 1600 0 0 0 C[18]
port 90 n
flabel metal2 26337 7342 26381 8498 1 FreeSans 1600 0 0 0 C[19]
port 91 n
flabel metal2 24449 7342 24493 8498 1 FreeSans 1600 0 0 0 C[20]
port 92 n
flabel metal2 22561 7342 22605 8498 1 FreeSans 1600 0 0 0 C[21]
port 93 n
flabel metal2 20673 7342 20717 8498 1 FreeSans 1600 0 0 0 C[22]
port 94 n
flabel metal2 18785 7342 18829 8498 1 FreeSans 1600 0 0 0 C[23]
port 95 n
flabel metal2 16897 7342 16941 8498 1 FreeSans 1600 0 0 0 C[24]
port 96 n
flabel metal2 15009 7342 15053 8498 1 FreeSans 1600 0 0 0 C[25]
port 97 n
flabel metal2 13121 7342 13165 8498 1 FreeSans 1600 0 0 0 C[26]
port 98 n
flabel metal2 11233 7342 11277 8498 1 FreeSans 1600 0 0 0 C[27]
port 99 n
flabel metal2 9345 7342 9389 8498 1 FreeSans 1600 0 0 0 C[28]
port 100 n
flabel metal2 7457 7342 7501 8498 1 FreeSans 1600 0 0 0 C[29]
port 101 n
flabel metal2 5569 7342 5613 8498 1 FreeSans 1600 0 0 0 C[30]
port 102 n
flabel metal2 422 22 467 1168 1 FreeSans 1600 0 0 0 C[31]
port 103 n
flabel metal2 2310 22 2355 1168 1 FreeSans 1600 0 0 0 C[32]
port 104 n
flabel metal2 4198 22 4243 1168 1 FreeSans 1600 0 0 0 C[33]
port 105 n
flabel metal2 6086 22 6131 1168 1 FreeSans 1600 0 0 0 C[34]
port 106 n
flabel metal2 7974 22 8019 1168 1 FreeSans 1600 0 0 0 C[35]
port 107 n
flabel metal2 9862 22 9907 1168 1 FreeSans 1600 0 0 0 C[36]
port 108 n
flabel metal2 11750 22 11795 1168 1 FreeSans 1600 0 0 0 C[37]
port 109 n
flabel metal2 13638 22 13683 1168 1 FreeSans 1600 0 0 0 C[38]
port 110 n
flabel metal2 15526 22 15571 1168 1 FreeSans 1600 0 0 0 C[39]
port 111 n
flabel metal2 17414 22 17459 1168 1 FreeSans 1600 0 0 0 C[40]
port 112 n
flabel metal2 19302 22 19347 1168 1 FreeSans 1600 0 0 0 C[41]
port 113 n
flabel metal2 21190 22 21235 1168 1 FreeSans 1600 0 0 0 C[42]
port 114 n
flabel metal2 23078 22 23123 1168 1 FreeSans 1600 0 0 0 C[43]
port 115 n
flabel metal2 24966 22 25011 1168 1 FreeSans 1600 0 0 0 C[44]
port 116 n
flabel metal2 26854 22 26899 1168 1 FreeSans 1600 0 0 0 C[45]
port 117 n
flabel metal2 28742 22 28787 1168 1 FreeSans 1600 0 0 0 C[46]
port 118 n
flabel metal2 30630 22 30675 1168 1 FreeSans 1600 0 0 0 C[47]
port 119 n
flabel metal2 32518 22 32563 1168 1 FreeSans 1600 0 0 0 C[48]
port 120 n
flabel metal2 34406 22 34451 1168 1 FreeSans 1600 0 0 0 C[49]
port 121 n
flabel metal2 36294 22 36339 1168 1 FreeSans 1600 0 0 0 C[50]
port 122 n
flabel metal2 38182 22 38227 1168 1 FreeSans 1600 0 0 0 C[51]
port 123 n
flabel metal2 40070 22 40115 1168 1 FreeSans 1600 0 0 0 C[52]
port 124 n
flabel metal2 41958 22 42003 1168 1 FreeSans 1600 0 0 0 C[53]
port 125 n
flabel metal2 43846 22 43891 1168 1 FreeSans 1600 0 0 0 C[54]
port 126 n
flabel metal2 45734 22 45779 1168 1 FreeSans 1600 0 0 0 C[55]
port 127 n
flabel metal2 47622 22 47667 1168 1 FreeSans 1600 0 0 0 C[56]
port 128 n
flabel metal2 49510 22 49555 1168 1 FreeSans 1600 0 0 0 C[57]
port 129 n
flabel metal2 51398 22 51443 1168 1 FreeSans 1600 0 0 0 C[58]
port 130 n
flabel metal2 53286 22 53331 1168 1 FreeSans 1600 0 0 0 C[59]
port 131 n
flabel metal2 55174 22 55219 1168 1 FreeSans 1600 0 0 0 C[60]
port 132 n
flabel metal2 57062 22 57107 1168 1 FreeSans 1600 0 0 0 C[61]
port 133 n
flabel metal2 58950 22 58995 1168 1 FreeSans 1600 0 0 0 C[62]
port 134 n
flabel metal2 60827 0 60883 1486 1 FreeSans 1600 0 0 0 C[63]
port 135 n
<< end >>
