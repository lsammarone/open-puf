/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/parameters/fast.spice