magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< locali >>
rect 207 1140 243 1174
rect 277 1140 315 1174
rect 349 1140 387 1174
rect 421 1140 459 1174
rect 493 1140 531 1174
rect 565 1140 603 1174
rect 637 1140 675 1174
rect 709 1140 747 1174
rect 781 1140 817 1174
rect 207 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 531 54
rect 565 20 603 54
rect 637 20 675 54
rect 709 20 747 54
rect 781 20 817 54
<< viali >>
rect 243 1140 277 1174
rect 315 1140 349 1174
rect 387 1140 421 1174
rect 459 1140 493 1174
rect 531 1140 565 1174
rect 603 1140 637 1174
rect 675 1140 709 1174
rect 747 1140 781 1174
rect 243 20 277 54
rect 315 20 349 54
rect 387 20 421 54
rect 459 20 493 54
rect 531 20 565 54
rect 603 20 637 54
rect 675 20 709 54
rect 747 20 781 54
<< obsli1 >>
rect 48 1010 82 1048
rect 48 938 82 976
rect 48 866 82 904
rect 48 794 82 832
rect 48 722 82 760
rect 48 650 82 688
rect 48 578 82 616
rect 48 506 82 544
rect 48 434 82 472
rect 48 362 82 400
rect 48 290 82 328
rect 48 218 82 256
rect 48 112 82 184
rect 183 88 217 1106
rect 339 88 373 1106
rect 495 88 529 1106
rect 651 88 685 1106
rect 807 88 841 1106
rect 942 1010 976 1048
rect 942 938 976 976
rect 942 866 976 904
rect 942 794 976 832
rect 942 722 976 760
rect 942 650 976 688
rect 942 578 976 616
rect 942 506 976 544
rect 942 434 976 472
rect 942 362 976 400
rect 942 290 976 328
rect 942 218 976 256
rect 942 112 976 184
<< obsli1c >>
rect 48 1048 82 1082
rect 48 976 82 1010
rect 48 904 82 938
rect 48 832 82 866
rect 48 760 82 794
rect 48 688 82 722
rect 48 616 82 650
rect 48 544 82 578
rect 48 472 82 506
rect 48 400 82 434
rect 48 328 82 362
rect 48 256 82 290
rect 48 184 82 218
rect 942 1048 976 1082
rect 942 976 976 1010
rect 942 904 976 938
rect 942 832 976 866
rect 942 760 976 794
rect 942 688 976 722
rect 942 616 976 650
rect 942 544 976 578
rect 942 472 976 506
rect 942 400 976 434
rect 942 328 976 362
rect 942 256 976 290
rect 942 184 976 218
<< metal1 >>
rect 231 1174 793 1194
rect 231 1140 243 1174
rect 277 1140 315 1174
rect 349 1140 387 1174
rect 421 1140 459 1174
rect 493 1140 531 1174
rect 565 1140 603 1174
rect 637 1140 675 1174
rect 709 1140 747 1174
rect 781 1140 793 1174
rect 231 1128 793 1140
rect 36 1082 95 1094
rect 36 1048 48 1082
rect 82 1048 95 1082
rect 36 1010 95 1048
rect 36 976 48 1010
rect 82 976 95 1010
rect 36 938 95 976
rect 36 904 48 938
rect 82 904 95 938
rect 36 866 95 904
rect 36 832 48 866
rect 82 832 95 866
rect 36 794 95 832
rect 36 760 48 794
rect 82 760 95 794
rect 36 722 95 760
rect 36 688 48 722
rect 82 688 95 722
rect 36 650 95 688
rect 36 616 48 650
rect 82 616 95 650
rect 36 578 95 616
rect 36 544 48 578
rect 82 544 95 578
rect 36 506 95 544
rect 36 472 48 506
rect 82 472 95 506
rect 36 434 95 472
rect 36 400 48 434
rect 82 400 95 434
rect 36 362 95 400
rect 36 328 48 362
rect 82 328 95 362
rect 36 290 95 328
rect 36 256 48 290
rect 82 256 95 290
rect 36 218 95 256
rect 36 184 48 218
rect 82 184 95 218
rect 36 100 95 184
rect 930 1082 989 1094
rect 930 1048 942 1082
rect 976 1048 989 1082
rect 930 1010 989 1048
rect 930 976 942 1010
rect 976 976 989 1010
rect 930 938 989 976
rect 930 904 942 938
rect 976 904 989 938
rect 930 866 989 904
rect 930 832 942 866
rect 976 832 989 866
rect 930 794 989 832
rect 930 760 942 794
rect 976 760 989 794
rect 930 722 989 760
rect 930 688 942 722
rect 976 688 989 722
rect 930 650 989 688
rect 930 616 942 650
rect 976 616 989 650
rect 930 578 989 616
rect 930 544 942 578
rect 976 544 989 578
rect 930 506 989 544
rect 930 472 942 506
rect 976 472 989 506
rect 930 434 989 472
rect 930 400 942 434
rect 976 400 989 434
rect 930 362 989 400
rect 930 328 942 362
rect 976 328 989 362
rect 930 290 989 328
rect 930 256 942 290
rect 976 256 989 290
rect 930 218 989 256
rect 930 184 942 218
rect 976 184 989 218
rect 930 100 989 184
rect 231 54 793 66
rect 231 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 531 54
rect 565 20 603 54
rect 637 20 675 54
rect 709 20 747 54
rect 781 20 793 54
rect 231 0 793 20
<< obsm1 >>
rect 174 100 226 1094
rect 330 100 382 1094
rect 486 100 538 1094
rect 642 100 694 1094
rect 798 100 850 1094
<< metal2 >>
rect 10 622 1014 1094
rect 10 100 1014 572
<< labels >>
rlabel metal2 s 10 622 1014 1094 6 DRAIN
port 1 nsew
rlabel viali s 747 1140 781 1174 6 GATE
port 2 nsew
rlabel viali s 747 20 781 54 6 GATE
port 2 nsew
rlabel viali s 675 1140 709 1174 6 GATE
port 2 nsew
rlabel viali s 675 20 709 54 6 GATE
port 2 nsew
rlabel viali s 603 1140 637 1174 6 GATE
port 2 nsew
rlabel viali s 603 20 637 54 6 GATE
port 2 nsew
rlabel viali s 531 1140 565 1174 6 GATE
port 2 nsew
rlabel viali s 531 20 565 54 6 GATE
port 2 nsew
rlabel viali s 459 1140 493 1174 6 GATE
port 2 nsew
rlabel viali s 459 20 493 54 6 GATE
port 2 nsew
rlabel viali s 387 1140 421 1174 6 GATE
port 2 nsew
rlabel viali s 387 20 421 54 6 GATE
port 2 nsew
rlabel viali s 315 1140 349 1174 6 GATE
port 2 nsew
rlabel viali s 315 20 349 54 6 GATE
port 2 nsew
rlabel viali s 243 1140 277 1174 6 GATE
port 2 nsew
rlabel viali s 243 20 277 54 6 GATE
port 2 nsew
rlabel locali s 207 1140 817 1174 6 GATE
port 2 nsew
rlabel locali s 207 20 817 54 6 GATE
port 2 nsew
rlabel metal1 s 231 1128 793 1194 6 GATE
port 2 nsew
rlabel metal1 s 231 0 793 66 6 GATE
port 2 nsew
rlabel metal2 s 10 100 1014 572 6 SOURCE
port 3 nsew
rlabel metal1 s 36 100 95 1094 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 930 100 989 1094 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 10 0 1014 1194
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7314062
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7291100
<< end >>
