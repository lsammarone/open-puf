/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8__leak_discrete.corner.spice