VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 32BR
  CLASS BLOCK ;
  FOREIGN 32BR ;
  ORIGIN 0.750 0.000 ;
  SIZE 126.720 BY 33.460 ;
  PIN VDD
    ANTENNADIFFAREA 81.137398 ;
    PORT
      LAYER nwell ;
        RECT 3.520 31.000 4.650 31.190 ;
        RECT 11.230 31.000 12.360 31.190 ;
        RECT 18.940 31.000 20.070 31.190 ;
        RECT 26.650 31.000 27.780 31.190 ;
        RECT 34.360 31.000 35.490 31.190 ;
        RECT 42.070 31.000 43.200 31.190 ;
        RECT 49.780 31.000 50.910 31.190 ;
        RECT 57.490 31.000 58.620 31.190 ;
        RECT 65.200 31.000 66.330 31.190 ;
        RECT 72.910 31.000 74.040 31.190 ;
        RECT 80.620 31.000 81.750 31.190 ;
        RECT 88.330 31.000 89.460 31.190 ;
        RECT 96.040 31.000 97.170 31.190 ;
        RECT 103.750 31.000 104.880 31.190 ;
        RECT 111.460 31.000 112.590 31.190 ;
        RECT 119.170 31.000 120.300 31.190 ;
        RECT 3.040 30.390 4.650 31.000 ;
        RECT 10.750 30.390 12.360 31.000 ;
        RECT 18.460 30.390 20.070 31.000 ;
        RECT 26.170 30.390 27.780 31.000 ;
        RECT 33.880 30.390 35.490 31.000 ;
        RECT 41.590 30.390 43.200 31.000 ;
        RECT 49.300 30.390 50.910 31.000 ;
        RECT 57.010 30.390 58.620 31.000 ;
        RECT 64.720 30.390 66.330 31.000 ;
        RECT 72.430 30.390 74.040 31.000 ;
        RECT 80.140 30.390 81.750 31.000 ;
        RECT 87.850 30.390 89.460 31.000 ;
        RECT 95.560 30.390 97.170 31.000 ;
        RECT 103.270 30.390 104.880 31.000 ;
        RECT 110.980 30.390 112.590 31.000 ;
        RECT 118.690 30.390 120.300 31.000 ;
        RECT 1.410 30.005 5.730 30.390 ;
        RECT 9.120 30.005 13.440 30.390 ;
        RECT 16.830 30.005 21.150 30.390 ;
        RECT 24.540 30.005 28.860 30.390 ;
        RECT 32.250 30.005 36.570 30.390 ;
        RECT 39.960 30.005 44.280 30.390 ;
        RECT 47.670 30.005 51.990 30.390 ;
        RECT 55.380 30.005 59.700 30.390 ;
        RECT 63.090 30.005 67.410 30.390 ;
        RECT 70.800 30.005 75.120 30.390 ;
        RECT 78.510 30.005 82.830 30.390 ;
        RECT 86.220 30.005 90.540 30.390 ;
        RECT 93.930 30.005 98.250 30.390 ;
        RECT 101.640 30.005 105.960 30.390 ;
        RECT 109.350 30.005 113.670 30.390 ;
        RECT 117.060 30.005 121.380 30.390 ;
        RECT 1.410 29.995 7.390 30.005 ;
        RECT 9.120 29.995 15.100 30.005 ;
        RECT 16.830 29.995 22.810 30.005 ;
        RECT 24.540 29.995 30.520 30.005 ;
        RECT 32.250 29.995 38.230 30.005 ;
        RECT 39.960 29.995 45.940 30.005 ;
        RECT 47.670 29.995 53.650 30.005 ;
        RECT 55.380 29.995 61.360 30.005 ;
        RECT 63.090 29.995 69.070 30.005 ;
        RECT 70.800 29.995 76.780 30.005 ;
        RECT 78.510 29.995 84.490 30.005 ;
        RECT 86.220 29.995 92.200 30.005 ;
        RECT 93.930 29.995 99.910 30.005 ;
        RECT 101.640 29.995 107.620 30.005 ;
        RECT 109.350 29.995 115.330 30.005 ;
        RECT 117.060 29.995 123.040 30.005 ;
        RECT -0.320 28.400 123.040 29.995 ;
        RECT -0.320 28.390 5.730 28.400 ;
        RECT 7.390 28.390 13.440 28.400 ;
        RECT 15.100 28.390 21.150 28.400 ;
        RECT 22.810 28.390 28.860 28.400 ;
        RECT 30.520 28.390 36.570 28.400 ;
        RECT 38.230 28.390 44.280 28.400 ;
        RECT 45.940 28.390 51.990 28.400 ;
        RECT 53.650 28.390 59.700 28.400 ;
        RECT 61.360 28.390 67.410 28.400 ;
        RECT 69.070 28.390 75.120 28.400 ;
        RECT 76.780 28.390 82.830 28.400 ;
        RECT 84.490 28.390 90.540 28.400 ;
        RECT 92.200 28.390 98.250 28.400 ;
        RECT 99.910 28.390 105.960 28.400 ;
        RECT 107.620 28.390 113.670 28.400 ;
        RECT 115.330 28.390 121.380 28.400 ;
        RECT 3.510 25.720 4.640 25.910 ;
        RECT 11.220 25.720 12.350 25.910 ;
        RECT 18.930 25.720 20.060 25.910 ;
        RECT 26.640 25.720 27.770 25.910 ;
        RECT 34.350 25.720 35.480 25.910 ;
        RECT 42.060 25.720 43.190 25.910 ;
        RECT 49.770 25.720 50.900 25.910 ;
        RECT 57.480 25.720 58.610 25.910 ;
        RECT 65.190 25.720 66.320 25.910 ;
        RECT 72.900 25.720 74.030 25.910 ;
        RECT 80.610 25.720 81.740 25.910 ;
        RECT 88.320 25.720 89.450 25.910 ;
        RECT 96.030 25.720 97.160 25.910 ;
        RECT 103.740 25.720 104.870 25.910 ;
        RECT 111.450 25.720 112.580 25.910 ;
        RECT 119.160 25.720 120.290 25.910 ;
        RECT 3.030 24.780 4.640 25.720 ;
        RECT 10.740 24.780 12.350 25.720 ;
        RECT 18.450 24.780 20.060 25.720 ;
        RECT 26.160 24.780 27.770 25.720 ;
        RECT 33.870 24.780 35.480 25.720 ;
        RECT 41.580 24.780 43.190 25.720 ;
        RECT 49.290 24.780 50.900 25.720 ;
        RECT 57.000 24.780 58.610 25.720 ;
        RECT 64.710 24.780 66.320 25.720 ;
        RECT 72.420 24.780 74.030 25.720 ;
        RECT 80.130 24.780 81.740 25.720 ;
        RECT 87.840 24.780 89.450 25.720 ;
        RECT 95.550 24.780 97.160 25.720 ;
        RECT 103.260 24.780 104.870 25.720 ;
        RECT 110.970 24.780 112.580 25.720 ;
        RECT 118.680 24.780 120.290 25.720 ;
        RECT 0.700 23.110 6.540 24.780 ;
        RECT 8.410 23.110 14.250 24.780 ;
        RECT 16.120 23.110 21.960 24.780 ;
        RECT 23.830 23.110 29.670 24.780 ;
        RECT 31.540 23.110 37.380 24.780 ;
        RECT 39.250 23.110 45.090 24.780 ;
        RECT 46.960 23.110 52.800 24.780 ;
        RECT 54.670 23.110 60.510 24.780 ;
        RECT 62.380 23.110 68.220 24.780 ;
        RECT 70.090 23.110 75.930 24.780 ;
        RECT 77.800 23.110 83.640 24.780 ;
        RECT 85.510 23.110 91.350 24.780 ;
        RECT 93.220 23.110 99.060 24.780 ;
        RECT 100.930 23.110 106.770 24.780 ;
        RECT 108.640 23.110 114.480 24.780 ;
        RECT 116.350 23.110 122.190 24.780 ;
        RECT 22.010 19.010 29.750 20.615 ;
        RECT 22.010 18.570 24.830 19.010 ;
        RECT 55.220 18.270 59.740 19.875 ;
        RECT 83.670 19.040 91.410 20.645 ;
        RECT 55.260 16.685 59.600 18.270 ;
        RECT 56.920 16.675 59.600 16.685 ;
        RECT 22.150 13.990 25.890 14.190 ;
        RECT 22.140 13.860 25.890 13.990 ;
        RECT 22.140 12.255 29.880 13.860 ;
        RECT 83.670 13.830 85.275 19.040 ;
        RECT 124.365 17.720 125.970 18.780 ;
        RECT 124.210 16.115 125.970 17.720 ;
        RECT 55.200 12.060 59.720 13.665 ;
        RECT 83.670 12.230 91.540 13.830 ;
        RECT 83.800 12.225 91.540 12.230 ;
        RECT 55.200 11.625 57.880 12.060 ;
        RECT 55.190 10.350 57.880 11.625 ;
        RECT 0.850 8.680 6.690 10.350 ;
        RECT 8.560 8.680 14.400 10.350 ;
        RECT 16.270 8.680 22.110 10.350 ;
        RECT 23.980 8.680 29.820 10.350 ;
        RECT 31.690 8.680 37.530 10.350 ;
        RECT 39.400 8.680 45.240 10.350 ;
        RECT 47.110 8.680 52.950 10.350 ;
        RECT 54.820 8.680 60.660 10.350 ;
        RECT 62.530 8.680 68.370 10.350 ;
        RECT 70.240 8.680 76.080 10.350 ;
        RECT 77.950 8.680 83.790 10.350 ;
        RECT 85.660 8.680 91.500 10.350 ;
        RECT 93.370 8.680 99.210 10.350 ;
        RECT 101.080 8.680 106.920 10.350 ;
        RECT 108.790 8.680 114.630 10.350 ;
        RECT 116.500 8.680 122.340 10.350 ;
        RECT 2.750 7.740 4.360 8.680 ;
        RECT 10.460 7.740 12.070 8.680 ;
        RECT 18.170 7.740 19.780 8.680 ;
        RECT 25.880 7.740 27.490 8.680 ;
        RECT 33.590 7.740 35.200 8.680 ;
        RECT 41.300 7.740 42.910 8.680 ;
        RECT 49.010 7.740 50.620 8.680 ;
        RECT 56.720 7.740 58.330 8.680 ;
        RECT 64.430 7.740 66.040 8.680 ;
        RECT 72.140 7.740 73.750 8.680 ;
        RECT 79.850 7.740 81.460 8.680 ;
        RECT 87.560 7.740 89.170 8.680 ;
        RECT 95.270 7.740 96.880 8.680 ;
        RECT 102.980 7.740 104.590 8.680 ;
        RECT 110.690 7.740 112.300 8.680 ;
        RECT 118.400 7.740 120.010 8.680 ;
        RECT 2.750 7.550 3.880 7.740 ;
        RECT 10.460 7.550 11.590 7.740 ;
        RECT 18.170 7.550 19.300 7.740 ;
        RECT 25.880 7.550 27.010 7.740 ;
        RECT 33.590 7.550 34.720 7.740 ;
        RECT 41.300 7.550 42.430 7.740 ;
        RECT 49.010 7.550 50.140 7.740 ;
        RECT 56.720 7.550 57.850 7.740 ;
        RECT 64.430 7.550 65.560 7.740 ;
        RECT 72.140 7.550 73.270 7.740 ;
        RECT 79.850 7.550 80.980 7.740 ;
        RECT 87.560 7.550 88.690 7.740 ;
        RECT 95.270 7.550 96.400 7.740 ;
        RECT 102.980 7.550 104.110 7.740 ;
        RECT 110.690 7.550 111.820 7.740 ;
        RECT 118.400 7.550 119.530 7.740 ;
        RECT 1.660 5.060 7.710 5.070 ;
        RECT 9.370 5.060 15.420 5.070 ;
        RECT 17.080 5.060 23.130 5.070 ;
        RECT 24.790 5.060 30.840 5.070 ;
        RECT 32.500 5.060 38.550 5.070 ;
        RECT 40.210 5.060 46.260 5.070 ;
        RECT 47.920 5.060 53.970 5.070 ;
        RECT 55.630 5.060 61.680 5.070 ;
        RECT 63.340 5.060 69.390 5.070 ;
        RECT 71.050 5.060 77.100 5.070 ;
        RECT 78.760 5.060 84.810 5.070 ;
        RECT 86.470 5.060 92.520 5.070 ;
        RECT 94.180 5.060 100.230 5.070 ;
        RECT 101.890 5.060 107.940 5.070 ;
        RECT 109.600 5.060 115.650 5.070 ;
        RECT 117.310 5.060 123.360 5.070 ;
        RECT 0.000 3.465 123.360 5.060 ;
        RECT 0.000 3.455 5.980 3.465 ;
        RECT 7.710 3.455 13.690 3.465 ;
        RECT 15.420 3.455 21.400 3.465 ;
        RECT 23.130 3.455 29.110 3.465 ;
        RECT 30.840 3.455 36.820 3.465 ;
        RECT 38.550 3.455 44.530 3.465 ;
        RECT 46.260 3.455 52.240 3.465 ;
        RECT 53.970 3.455 59.950 3.465 ;
        RECT 61.680 3.455 67.660 3.465 ;
        RECT 69.390 3.455 75.370 3.465 ;
        RECT 77.100 3.455 83.080 3.465 ;
        RECT 84.810 3.455 90.790 3.465 ;
        RECT 92.520 3.455 98.500 3.465 ;
        RECT 100.230 3.455 106.210 3.465 ;
        RECT 107.940 3.455 113.920 3.465 ;
        RECT 115.650 3.455 121.630 3.465 ;
        RECT 1.660 3.070 5.980 3.455 ;
        RECT 9.370 3.070 13.690 3.455 ;
        RECT 17.080 3.070 21.400 3.455 ;
        RECT 24.790 3.070 29.110 3.455 ;
        RECT 32.500 3.070 36.820 3.455 ;
        RECT 40.210 3.070 44.530 3.455 ;
        RECT 47.920 3.070 52.240 3.455 ;
        RECT 55.630 3.070 59.950 3.455 ;
        RECT 63.340 3.070 67.660 3.455 ;
        RECT 71.050 3.070 75.370 3.455 ;
        RECT 78.760 3.070 83.080 3.455 ;
        RECT 86.470 3.070 90.790 3.455 ;
        RECT 94.180 3.070 98.500 3.455 ;
        RECT 101.890 3.070 106.210 3.455 ;
        RECT 109.600 3.070 113.920 3.455 ;
        RECT 117.310 3.070 121.630 3.455 ;
        RECT 2.740 2.460 4.350 3.070 ;
        RECT 10.450 2.460 12.060 3.070 ;
        RECT 18.160 2.460 19.770 3.070 ;
        RECT 25.870 2.460 27.480 3.070 ;
        RECT 33.580 2.460 35.190 3.070 ;
        RECT 41.290 2.460 42.900 3.070 ;
        RECT 49.000 2.460 50.610 3.070 ;
        RECT 56.710 2.460 58.320 3.070 ;
        RECT 64.420 2.460 66.030 3.070 ;
        RECT 72.130 2.460 73.740 3.070 ;
        RECT 79.840 2.460 81.450 3.070 ;
        RECT 87.550 2.460 89.160 3.070 ;
        RECT 95.260 2.460 96.870 3.070 ;
        RECT 102.970 2.460 104.580 3.070 ;
        RECT 110.680 2.460 112.290 3.070 ;
        RECT 118.390 2.460 120.000 3.070 ;
        RECT 2.740 2.270 3.870 2.460 ;
        RECT 10.450 2.270 11.580 2.460 ;
        RECT 18.160 2.270 19.290 2.460 ;
        RECT 25.870 2.270 27.000 2.460 ;
        RECT 33.580 2.270 34.710 2.460 ;
        RECT 41.290 2.270 42.420 2.460 ;
        RECT 49.000 2.270 50.130 2.460 ;
        RECT 56.710 2.270 57.840 2.460 ;
        RECT 64.420 2.270 65.550 2.460 ;
        RECT 72.130 2.270 73.260 2.460 ;
        RECT 79.840 2.270 80.970 2.460 ;
        RECT 87.550 2.270 88.680 2.460 ;
        RECT 95.260 2.270 96.390 2.460 ;
        RECT 102.970 2.270 104.100 2.460 ;
        RECT 110.680 2.270 111.810 2.460 ;
        RECT 118.390 2.270 119.520 2.460 ;
      LAYER li1 ;
        RECT 0.700 28.665 0.910 29.805 ;
        RECT 2.090 29.090 2.260 29.910 ;
        RECT 4.880 29.090 5.050 29.910 ;
        RECT 2.090 28.870 5.060 29.090 ;
        RECT -0.130 28.495 1.250 28.665 ;
        RECT 2.820 28.550 4.230 28.870 ;
        RECT 6.650 28.675 6.860 29.815 ;
        RECT 3.660 28.540 4.230 28.550 ;
        RECT 5.820 28.505 7.200 28.675 ;
        RECT 8.410 28.665 8.620 29.805 ;
        RECT 9.800 29.090 9.970 29.910 ;
        RECT 12.590 29.090 12.760 29.910 ;
        RECT 9.800 28.870 12.770 29.090 ;
        RECT 0.985 23.435 1.315 24.575 ;
        RECT 2.810 23.435 4.220 23.810 ;
        RECT 5.055 23.435 5.385 24.575 ;
        RECT 0.890 23.430 6.340 23.435 ;
        RECT 6.685 23.430 6.855 28.505 ;
        RECT 7.580 28.495 8.960 28.665 ;
        RECT 10.530 28.550 11.940 28.870 ;
        RECT 14.360 28.675 14.570 29.815 ;
        RECT 11.370 28.540 11.940 28.550 ;
        RECT 13.530 28.505 14.910 28.675 ;
        RECT 16.120 28.665 16.330 29.805 ;
        RECT 17.510 29.090 17.680 29.910 ;
        RECT 20.300 29.090 20.470 29.910 ;
        RECT 17.510 28.870 20.480 29.090 ;
        RECT 8.695 23.435 9.025 24.575 ;
        RECT 10.520 23.435 11.930 23.810 ;
        RECT 12.765 23.435 13.095 24.575 ;
        RECT 0.890 23.265 6.855 23.430 ;
        RECT 8.600 23.430 14.050 23.435 ;
        RECT 14.395 23.430 14.565 28.505 ;
        RECT 15.290 28.495 16.670 28.665 ;
        RECT 18.240 28.550 19.650 28.870 ;
        RECT 22.070 28.675 22.280 29.815 ;
        RECT 19.080 28.540 19.650 28.550 ;
        RECT 21.240 28.505 22.620 28.675 ;
        RECT 23.830 28.665 24.040 29.805 ;
        RECT 25.220 29.090 25.390 29.910 ;
        RECT 28.010 29.090 28.180 29.910 ;
        RECT 25.220 28.870 28.190 29.090 ;
        RECT 16.405 23.435 16.735 24.575 ;
        RECT 18.230 23.435 19.640 23.810 ;
        RECT 20.475 23.435 20.805 24.575 ;
        RECT 8.600 23.265 14.565 23.430 ;
        RECT 16.310 23.430 21.760 23.435 ;
        RECT 22.105 23.430 22.275 28.505 ;
        RECT 23.000 28.495 24.380 28.665 ;
        RECT 25.950 28.550 27.360 28.870 ;
        RECT 29.780 28.675 29.990 29.815 ;
        RECT 26.790 28.540 27.360 28.550 ;
        RECT 28.950 28.505 30.330 28.675 ;
        RECT 31.540 28.665 31.750 29.805 ;
        RECT 32.930 29.090 33.100 29.910 ;
        RECT 35.720 29.090 35.890 29.910 ;
        RECT 32.930 28.870 35.900 29.090 ;
        RECT 24.115 23.435 24.445 24.575 ;
        RECT 25.940 23.435 27.350 23.810 ;
        RECT 28.185 23.435 28.515 24.575 ;
        RECT 16.310 23.265 22.275 23.430 ;
        RECT 24.020 23.430 29.470 23.435 ;
        RECT 29.815 23.430 29.985 28.505 ;
        RECT 30.710 28.495 32.090 28.665 ;
        RECT 33.660 28.550 35.070 28.870 ;
        RECT 37.490 28.675 37.700 29.815 ;
        RECT 34.500 28.540 35.070 28.550 ;
        RECT 36.660 28.505 38.040 28.675 ;
        RECT 39.250 28.665 39.460 29.805 ;
        RECT 40.640 29.090 40.810 29.910 ;
        RECT 43.430 29.090 43.600 29.910 ;
        RECT 40.640 28.870 43.610 29.090 ;
        RECT 31.825 23.435 32.155 24.575 ;
        RECT 33.650 23.435 35.060 23.810 ;
        RECT 35.895 23.435 36.225 24.575 ;
        RECT 24.020 23.265 29.985 23.430 ;
        RECT 31.730 23.430 37.180 23.435 ;
        RECT 37.525 23.430 37.695 28.505 ;
        RECT 38.420 28.495 39.800 28.665 ;
        RECT 41.370 28.550 42.780 28.870 ;
        RECT 45.200 28.675 45.410 29.815 ;
        RECT 42.210 28.540 42.780 28.550 ;
        RECT 44.370 28.505 45.750 28.675 ;
        RECT 46.960 28.665 47.170 29.805 ;
        RECT 48.350 29.090 48.520 29.910 ;
        RECT 51.140 29.090 51.310 29.910 ;
        RECT 48.350 28.870 51.320 29.090 ;
        RECT 39.535 23.435 39.865 24.575 ;
        RECT 41.360 23.435 42.770 23.810 ;
        RECT 43.605 23.435 43.935 24.575 ;
        RECT 31.730 23.265 37.695 23.430 ;
        RECT 39.440 23.430 44.890 23.435 ;
        RECT 45.235 23.430 45.405 28.505 ;
        RECT 46.130 28.495 47.510 28.665 ;
        RECT 49.080 28.550 50.490 28.870 ;
        RECT 52.910 28.675 53.120 29.815 ;
        RECT 49.920 28.540 50.490 28.550 ;
        RECT 52.080 28.505 53.460 28.675 ;
        RECT 54.670 28.665 54.880 29.805 ;
        RECT 56.060 29.090 56.230 29.910 ;
        RECT 58.850 29.090 59.020 29.910 ;
        RECT 56.060 28.870 59.030 29.090 ;
        RECT 47.245 23.435 47.575 24.575 ;
        RECT 49.070 23.435 50.480 23.810 ;
        RECT 51.315 23.435 51.645 24.575 ;
        RECT 39.440 23.265 45.405 23.430 ;
        RECT 47.150 23.430 52.600 23.435 ;
        RECT 52.945 23.430 53.115 28.505 ;
        RECT 53.840 28.495 55.220 28.665 ;
        RECT 56.790 28.550 58.200 28.870 ;
        RECT 60.620 28.675 60.830 29.815 ;
        RECT 57.630 28.540 58.200 28.550 ;
        RECT 59.790 28.505 61.170 28.675 ;
        RECT 62.380 28.665 62.590 29.805 ;
        RECT 63.770 29.090 63.940 29.910 ;
        RECT 66.560 29.090 66.730 29.910 ;
        RECT 63.770 28.870 66.740 29.090 ;
        RECT 54.955 23.435 55.285 24.575 ;
        RECT 56.780 23.435 58.190 23.810 ;
        RECT 59.025 23.435 59.355 24.575 ;
        RECT 47.150 23.265 53.115 23.430 ;
        RECT 54.860 23.430 60.310 23.435 ;
        RECT 60.655 23.430 60.825 28.505 ;
        RECT 61.550 28.495 62.930 28.665 ;
        RECT 64.500 28.550 65.910 28.870 ;
        RECT 68.330 28.675 68.540 29.815 ;
        RECT 65.340 28.540 65.910 28.550 ;
        RECT 67.500 28.505 68.880 28.675 ;
        RECT 70.090 28.665 70.300 29.805 ;
        RECT 71.480 29.090 71.650 29.910 ;
        RECT 74.270 29.090 74.440 29.910 ;
        RECT 71.480 28.870 74.450 29.090 ;
        RECT 62.665 23.435 62.995 24.575 ;
        RECT 64.490 23.435 65.900 23.810 ;
        RECT 66.735 23.435 67.065 24.575 ;
        RECT 54.860 23.265 60.825 23.430 ;
        RECT 62.570 23.430 68.020 23.435 ;
        RECT 68.365 23.430 68.535 28.505 ;
        RECT 69.260 28.495 70.640 28.665 ;
        RECT 72.210 28.550 73.620 28.870 ;
        RECT 76.040 28.675 76.250 29.815 ;
        RECT 73.050 28.540 73.620 28.550 ;
        RECT 75.210 28.505 76.590 28.675 ;
        RECT 77.800 28.665 78.010 29.805 ;
        RECT 79.190 29.090 79.360 29.910 ;
        RECT 81.980 29.090 82.150 29.910 ;
        RECT 79.190 28.870 82.160 29.090 ;
        RECT 70.375 23.435 70.705 24.575 ;
        RECT 72.200 23.435 73.610 23.810 ;
        RECT 74.445 23.435 74.775 24.575 ;
        RECT 62.570 23.265 68.535 23.430 ;
        RECT 70.280 23.430 75.730 23.435 ;
        RECT 76.075 23.430 76.245 28.505 ;
        RECT 76.970 28.495 78.350 28.665 ;
        RECT 79.920 28.550 81.330 28.870 ;
        RECT 83.750 28.675 83.960 29.815 ;
        RECT 80.760 28.540 81.330 28.550 ;
        RECT 82.920 28.505 84.300 28.675 ;
        RECT 85.510 28.665 85.720 29.805 ;
        RECT 86.900 29.090 87.070 29.910 ;
        RECT 89.690 29.090 89.860 29.910 ;
        RECT 86.900 28.870 89.870 29.090 ;
        RECT 78.085 23.435 78.415 24.575 ;
        RECT 79.910 23.435 81.320 23.810 ;
        RECT 82.155 23.435 82.485 24.575 ;
        RECT 70.280 23.265 76.245 23.430 ;
        RECT 77.990 23.430 83.440 23.435 ;
        RECT 83.785 23.430 83.955 28.505 ;
        RECT 84.680 28.495 86.060 28.665 ;
        RECT 87.630 28.550 89.040 28.870 ;
        RECT 91.460 28.675 91.670 29.815 ;
        RECT 88.470 28.540 89.040 28.550 ;
        RECT 90.630 28.505 92.010 28.675 ;
        RECT 93.220 28.665 93.430 29.805 ;
        RECT 94.610 29.090 94.780 29.910 ;
        RECT 97.400 29.090 97.570 29.910 ;
        RECT 94.610 28.870 97.580 29.090 ;
        RECT 85.795 23.435 86.125 24.575 ;
        RECT 87.620 23.435 89.030 23.810 ;
        RECT 89.865 23.435 90.195 24.575 ;
        RECT 77.990 23.265 83.955 23.430 ;
        RECT 85.700 23.430 91.150 23.435 ;
        RECT 91.495 23.430 91.665 28.505 ;
        RECT 92.390 28.495 93.770 28.665 ;
        RECT 95.340 28.550 96.750 28.870 ;
        RECT 99.170 28.675 99.380 29.815 ;
        RECT 96.180 28.540 96.750 28.550 ;
        RECT 98.340 28.505 99.720 28.675 ;
        RECT 100.930 28.665 101.140 29.805 ;
        RECT 102.320 29.090 102.490 29.910 ;
        RECT 105.110 29.090 105.280 29.910 ;
        RECT 102.320 28.870 105.290 29.090 ;
        RECT 93.505 23.435 93.835 24.575 ;
        RECT 95.330 23.435 96.740 23.810 ;
        RECT 97.575 23.435 97.905 24.575 ;
        RECT 85.700 23.265 91.665 23.430 ;
        RECT 93.410 23.430 98.860 23.435 ;
        RECT 99.205 23.430 99.375 28.505 ;
        RECT 100.100 28.495 101.480 28.665 ;
        RECT 103.050 28.550 104.460 28.870 ;
        RECT 106.880 28.675 107.090 29.815 ;
        RECT 103.890 28.540 104.460 28.550 ;
        RECT 106.050 28.505 107.430 28.675 ;
        RECT 108.640 28.665 108.850 29.805 ;
        RECT 110.030 29.090 110.200 29.910 ;
        RECT 112.820 29.090 112.990 29.910 ;
        RECT 110.030 28.870 113.000 29.090 ;
        RECT 101.215 23.435 101.545 24.575 ;
        RECT 103.040 23.435 104.450 23.810 ;
        RECT 105.285 23.435 105.615 24.575 ;
        RECT 93.410 23.265 99.375 23.430 ;
        RECT 101.120 23.430 106.570 23.435 ;
        RECT 106.915 23.430 107.085 28.505 ;
        RECT 107.810 28.495 109.190 28.665 ;
        RECT 110.760 28.550 112.170 28.870 ;
        RECT 114.590 28.675 114.800 29.815 ;
        RECT 111.600 28.540 112.170 28.550 ;
        RECT 113.760 28.505 115.140 28.675 ;
        RECT 116.350 28.665 116.560 29.805 ;
        RECT 117.740 29.090 117.910 29.910 ;
        RECT 120.530 29.090 120.700 29.910 ;
        RECT 117.740 28.870 120.710 29.090 ;
        RECT 108.925 23.435 109.255 24.575 ;
        RECT 110.750 23.435 112.160 23.810 ;
        RECT 112.995 23.435 113.325 24.575 ;
        RECT 101.120 23.265 107.085 23.430 ;
        RECT 108.830 23.430 114.280 23.435 ;
        RECT 114.625 23.430 114.795 28.505 ;
        RECT 115.520 28.495 116.900 28.665 ;
        RECT 118.470 28.550 119.880 28.870 ;
        RECT 122.300 28.675 122.510 29.815 ;
        RECT 119.310 28.540 119.880 28.550 ;
        RECT 121.470 28.505 122.850 28.675 ;
        RECT 116.635 23.435 116.965 24.575 ;
        RECT 118.460 23.435 119.870 23.810 ;
        RECT 120.705 23.435 121.035 24.575 ;
        RECT 108.830 23.265 114.795 23.430 ;
        RECT 116.540 23.430 121.990 23.435 ;
        RECT 122.335 23.430 122.505 28.505 ;
        RECT 116.540 23.265 122.505 23.430 ;
        RECT 2.270 23.260 4.220 23.265 ;
        RECT 6.240 23.260 6.855 23.265 ;
        RECT 9.980 23.260 11.930 23.265 ;
        RECT 13.950 23.260 14.565 23.265 ;
        RECT 17.690 23.260 19.640 23.265 ;
        RECT 21.660 23.260 22.275 23.265 ;
        RECT 25.400 23.260 27.350 23.265 ;
        RECT 29.370 23.260 29.985 23.265 ;
        RECT 33.110 23.260 35.060 23.265 ;
        RECT 37.080 23.260 37.695 23.265 ;
        RECT 40.820 23.260 42.770 23.265 ;
        RECT 44.790 23.260 45.405 23.265 ;
        RECT 48.530 23.260 50.480 23.265 ;
        RECT 52.500 23.260 53.115 23.265 ;
        RECT 56.240 23.260 58.190 23.265 ;
        RECT 60.210 23.260 60.825 23.265 ;
        RECT 63.950 23.260 65.900 23.265 ;
        RECT 67.920 23.260 68.535 23.265 ;
        RECT 71.660 23.260 73.610 23.265 ;
        RECT 75.630 23.260 76.245 23.265 ;
        RECT 79.370 23.260 81.320 23.265 ;
        RECT 83.340 23.260 83.955 23.265 ;
        RECT 87.080 23.260 89.030 23.265 ;
        RECT 91.050 23.260 91.665 23.265 ;
        RECT 94.790 23.260 96.740 23.265 ;
        RECT 98.760 23.260 99.375 23.265 ;
        RECT 102.500 23.260 104.450 23.265 ;
        RECT 106.470 23.260 107.085 23.265 ;
        RECT 110.210 23.260 112.160 23.265 ;
        RECT 114.180 23.260 114.795 23.265 ;
        RECT 117.920 23.260 119.870 23.265 ;
        RECT 121.890 23.260 122.505 23.265 ;
        RECT 22.400 19.285 22.610 20.435 ;
        RECT 23.280 19.285 23.450 20.085 ;
        RECT 24.120 19.285 24.290 20.085 ;
        RECT 24.960 19.285 25.130 20.085 ;
        RECT 25.800 19.285 25.970 20.085 ;
        RECT 26.640 19.285 26.810 20.085 ;
        RECT 27.480 19.285 27.650 20.085 ;
        RECT 28.320 19.285 28.490 20.085 ;
        RECT 29.160 19.285 29.370 20.085 ;
        RECT 22.200 19.115 29.560 19.285 ;
        RECT 23.040 18.880 23.550 19.115 ;
        RECT 55.665 18.545 55.920 19.345 ;
        RECT 56.590 18.545 56.760 19.345 ;
        RECT 57.430 18.545 57.600 19.345 ;
        RECT 58.270 18.545 58.440 19.345 ;
        RECT 59.110 18.545 59.410 19.345 ;
        RECT 84.060 19.315 84.270 20.465 ;
        RECT 84.940 19.315 85.110 20.115 ;
        RECT 85.780 19.315 85.950 20.115 ;
        RECT 86.620 19.315 86.790 20.115 ;
        RECT 87.460 19.315 87.630 20.115 ;
        RECT 88.300 19.315 88.470 20.115 ;
        RECT 89.140 19.315 89.310 20.115 ;
        RECT 89.980 19.315 90.150 20.115 ;
        RECT 90.820 19.315 91.030 20.115 ;
        RECT 83.860 19.145 91.220 19.315 ;
        RECT 55.410 18.375 59.550 18.545 ;
        RECT 55.450 18.015 56.830 18.185 ;
        RECT 55.790 16.875 56.000 18.015 ;
        RECT 57.110 18.005 59.410 18.175 ;
        RECT 125.280 18.020 125.620 18.270 ;
        RECT 57.240 17.580 57.505 18.005 ;
        RECT 56.670 16.880 57.505 17.580 ;
        RECT 58.175 17.205 58.345 18.005 ;
        RECT 59.015 17.545 59.225 18.005 ;
        RECT 125.280 17.615 125.450 18.020 ;
        RECT 124.400 17.445 125.780 17.615 ;
        RECT 56.770 16.870 57.505 16.880 ;
        RECT 57.240 16.865 57.505 16.870 ;
        RECT 124.925 16.685 125.255 17.445 ;
        RECT 23.240 13.755 23.750 13.940 ;
        RECT 22.330 13.585 29.690 13.755 ;
        RECT 84.190 13.725 84.770 14.190 ;
        RECT 22.530 12.435 22.740 13.585 ;
        RECT 23.410 12.785 23.580 13.585 ;
        RECT 24.250 12.785 24.420 13.585 ;
        RECT 25.090 12.785 25.260 13.585 ;
        RECT 25.930 12.785 26.100 13.585 ;
        RECT 26.770 12.785 26.940 13.585 ;
        RECT 27.610 12.785 27.780 13.585 ;
        RECT 28.450 12.785 28.620 13.585 ;
        RECT 29.290 12.785 29.500 13.585 ;
        RECT 83.990 13.555 91.350 13.725 ;
        RECT 55.645 12.335 55.900 13.135 ;
        RECT 56.570 12.335 56.740 13.135 ;
        RECT 57.410 12.335 57.580 13.135 ;
        RECT 58.250 12.335 58.420 13.135 ;
        RECT 59.090 12.335 59.390 13.135 ;
        RECT 84.190 12.405 84.400 13.555 ;
        RECT 85.070 12.755 85.240 13.555 ;
        RECT 85.910 12.755 86.080 13.555 ;
        RECT 86.750 12.755 86.920 13.555 ;
        RECT 87.590 12.755 87.760 13.555 ;
        RECT 88.430 12.755 88.600 13.555 ;
        RECT 89.270 12.755 89.440 13.555 ;
        RECT 90.110 12.755 90.280 13.555 ;
        RECT 90.950 12.755 91.160 13.555 ;
        RECT 55.390 12.165 59.530 12.335 ;
        RECT 0.535 10.195 1.150 10.200 ;
        RECT 3.170 10.195 5.120 10.200 ;
        RECT 8.245 10.195 8.860 10.200 ;
        RECT 10.880 10.195 12.830 10.200 ;
        RECT 15.955 10.195 16.570 10.200 ;
        RECT 18.590 10.195 20.540 10.200 ;
        RECT 23.665 10.195 24.280 10.200 ;
        RECT 26.300 10.195 28.250 10.200 ;
        RECT 31.375 10.195 31.990 10.200 ;
        RECT 34.010 10.195 35.960 10.200 ;
        RECT 39.085 10.195 39.700 10.200 ;
        RECT 41.720 10.195 43.670 10.200 ;
        RECT 46.795 10.195 47.410 10.200 ;
        RECT 49.430 10.195 51.380 10.200 ;
        RECT 54.505 10.195 55.120 10.200 ;
        RECT 57.140 10.195 59.090 10.200 ;
        RECT 62.215 10.195 62.830 10.200 ;
        RECT 64.850 10.195 66.800 10.200 ;
        RECT 69.925 10.195 70.540 10.200 ;
        RECT 72.560 10.195 74.510 10.200 ;
        RECT 77.635 10.195 78.250 10.200 ;
        RECT 80.270 10.195 82.220 10.200 ;
        RECT 85.345 10.195 85.960 10.200 ;
        RECT 87.980 10.195 89.930 10.200 ;
        RECT 93.055 10.195 93.670 10.200 ;
        RECT 95.690 10.195 97.640 10.200 ;
        RECT 100.765 10.195 101.380 10.200 ;
        RECT 103.400 10.195 105.350 10.200 ;
        RECT 108.475 10.195 109.090 10.200 ;
        RECT 111.110 10.195 113.060 10.200 ;
        RECT 116.185 10.195 116.800 10.200 ;
        RECT 118.820 10.195 120.770 10.200 ;
        RECT 0.535 10.030 6.500 10.195 ;
        RECT 0.535 4.955 0.705 10.030 ;
        RECT 1.050 10.025 6.500 10.030 ;
        RECT 8.245 10.030 14.210 10.195 ;
        RECT 2.005 8.885 2.335 10.025 ;
        RECT 3.170 9.650 4.580 10.025 ;
        RECT 6.075 8.885 6.405 10.025 ;
        RECT 0.190 4.785 1.570 4.955 ;
        RECT 3.160 4.910 3.730 4.920 ;
        RECT 0.530 3.645 0.740 4.785 ;
        RECT 3.160 4.590 4.570 4.910 ;
        RECT 6.140 4.795 7.520 4.965 ;
        RECT 8.245 4.955 8.415 10.030 ;
        RECT 8.760 10.025 14.210 10.030 ;
        RECT 15.955 10.030 21.920 10.195 ;
        RECT 9.715 8.885 10.045 10.025 ;
        RECT 10.880 9.650 12.290 10.025 ;
        RECT 13.785 8.885 14.115 10.025 ;
        RECT 2.330 4.370 5.300 4.590 ;
        RECT 2.340 3.550 2.510 4.370 ;
        RECT 5.130 3.550 5.300 4.370 ;
        RECT 6.480 3.655 6.690 4.795 ;
        RECT 7.900 4.785 9.280 4.955 ;
        RECT 10.870 4.910 11.440 4.920 ;
        RECT 8.240 3.645 8.450 4.785 ;
        RECT 10.870 4.590 12.280 4.910 ;
        RECT 13.850 4.795 15.230 4.965 ;
        RECT 15.955 4.955 16.125 10.030 ;
        RECT 16.470 10.025 21.920 10.030 ;
        RECT 23.665 10.030 29.630 10.195 ;
        RECT 17.425 8.885 17.755 10.025 ;
        RECT 18.590 9.650 20.000 10.025 ;
        RECT 21.495 8.885 21.825 10.025 ;
        RECT 10.040 4.370 13.010 4.590 ;
        RECT 10.050 3.550 10.220 4.370 ;
        RECT 12.840 3.550 13.010 4.370 ;
        RECT 14.190 3.655 14.400 4.795 ;
        RECT 15.610 4.785 16.990 4.955 ;
        RECT 18.580 4.910 19.150 4.920 ;
        RECT 15.950 3.645 16.160 4.785 ;
        RECT 18.580 4.590 19.990 4.910 ;
        RECT 21.560 4.795 22.940 4.965 ;
        RECT 23.665 4.955 23.835 10.030 ;
        RECT 24.180 10.025 29.630 10.030 ;
        RECT 31.375 10.030 37.340 10.195 ;
        RECT 25.135 8.885 25.465 10.025 ;
        RECT 26.300 9.650 27.710 10.025 ;
        RECT 29.205 8.885 29.535 10.025 ;
        RECT 17.750 4.370 20.720 4.590 ;
        RECT 17.760 3.550 17.930 4.370 ;
        RECT 20.550 3.550 20.720 4.370 ;
        RECT 21.900 3.655 22.110 4.795 ;
        RECT 23.320 4.785 24.700 4.955 ;
        RECT 26.290 4.910 26.860 4.920 ;
        RECT 23.660 3.645 23.870 4.785 ;
        RECT 26.290 4.590 27.700 4.910 ;
        RECT 29.270 4.795 30.650 4.965 ;
        RECT 31.375 4.955 31.545 10.030 ;
        RECT 31.890 10.025 37.340 10.030 ;
        RECT 39.085 10.030 45.050 10.195 ;
        RECT 32.845 8.885 33.175 10.025 ;
        RECT 34.010 9.650 35.420 10.025 ;
        RECT 36.915 8.885 37.245 10.025 ;
        RECT 25.460 4.370 28.430 4.590 ;
        RECT 25.470 3.550 25.640 4.370 ;
        RECT 28.260 3.550 28.430 4.370 ;
        RECT 29.610 3.655 29.820 4.795 ;
        RECT 31.030 4.785 32.410 4.955 ;
        RECT 34.000 4.910 34.570 4.920 ;
        RECT 31.370 3.645 31.580 4.785 ;
        RECT 34.000 4.590 35.410 4.910 ;
        RECT 36.980 4.795 38.360 4.965 ;
        RECT 39.085 4.955 39.255 10.030 ;
        RECT 39.600 10.025 45.050 10.030 ;
        RECT 46.795 10.030 52.760 10.195 ;
        RECT 40.555 8.885 40.885 10.025 ;
        RECT 41.720 9.650 43.130 10.025 ;
        RECT 44.625 8.885 44.955 10.025 ;
        RECT 33.170 4.370 36.140 4.590 ;
        RECT 33.180 3.550 33.350 4.370 ;
        RECT 35.970 3.550 36.140 4.370 ;
        RECT 37.320 3.655 37.530 4.795 ;
        RECT 38.740 4.785 40.120 4.955 ;
        RECT 41.710 4.910 42.280 4.920 ;
        RECT 39.080 3.645 39.290 4.785 ;
        RECT 41.710 4.590 43.120 4.910 ;
        RECT 44.690 4.795 46.070 4.965 ;
        RECT 46.795 4.955 46.965 10.030 ;
        RECT 47.310 10.025 52.760 10.030 ;
        RECT 54.505 10.030 60.470 10.195 ;
        RECT 48.265 8.885 48.595 10.025 ;
        RECT 49.430 9.650 50.840 10.025 ;
        RECT 52.335 8.885 52.665 10.025 ;
        RECT 40.880 4.370 43.850 4.590 ;
        RECT 40.890 3.550 41.060 4.370 ;
        RECT 43.680 3.550 43.850 4.370 ;
        RECT 45.030 3.655 45.240 4.795 ;
        RECT 46.450 4.785 47.830 4.955 ;
        RECT 49.420 4.910 49.990 4.920 ;
        RECT 46.790 3.645 47.000 4.785 ;
        RECT 49.420 4.590 50.830 4.910 ;
        RECT 52.400 4.795 53.780 4.965 ;
        RECT 54.505 4.955 54.675 10.030 ;
        RECT 55.020 10.025 60.470 10.030 ;
        RECT 62.215 10.030 68.180 10.195 ;
        RECT 55.975 8.885 56.305 10.025 ;
        RECT 57.140 9.650 58.550 10.025 ;
        RECT 60.045 8.885 60.375 10.025 ;
        RECT 48.590 4.370 51.560 4.590 ;
        RECT 48.600 3.550 48.770 4.370 ;
        RECT 51.390 3.550 51.560 4.370 ;
        RECT 52.740 3.655 52.950 4.795 ;
        RECT 54.160 4.785 55.540 4.955 ;
        RECT 57.130 4.910 57.700 4.920 ;
        RECT 54.500 3.645 54.710 4.785 ;
        RECT 57.130 4.590 58.540 4.910 ;
        RECT 60.110 4.795 61.490 4.965 ;
        RECT 62.215 4.955 62.385 10.030 ;
        RECT 62.730 10.025 68.180 10.030 ;
        RECT 69.925 10.030 75.890 10.195 ;
        RECT 63.685 8.885 64.015 10.025 ;
        RECT 64.850 9.650 66.260 10.025 ;
        RECT 67.755 8.885 68.085 10.025 ;
        RECT 56.300 4.370 59.270 4.590 ;
        RECT 56.310 3.550 56.480 4.370 ;
        RECT 59.100 3.550 59.270 4.370 ;
        RECT 60.450 3.655 60.660 4.795 ;
        RECT 61.870 4.785 63.250 4.955 ;
        RECT 64.840 4.910 65.410 4.920 ;
        RECT 62.210 3.645 62.420 4.785 ;
        RECT 64.840 4.590 66.250 4.910 ;
        RECT 67.820 4.795 69.200 4.965 ;
        RECT 69.925 4.955 70.095 10.030 ;
        RECT 70.440 10.025 75.890 10.030 ;
        RECT 77.635 10.030 83.600 10.195 ;
        RECT 71.395 8.885 71.725 10.025 ;
        RECT 72.560 9.650 73.970 10.025 ;
        RECT 75.465 8.885 75.795 10.025 ;
        RECT 64.010 4.370 66.980 4.590 ;
        RECT 64.020 3.550 64.190 4.370 ;
        RECT 66.810 3.550 66.980 4.370 ;
        RECT 68.160 3.655 68.370 4.795 ;
        RECT 69.580 4.785 70.960 4.955 ;
        RECT 72.550 4.910 73.120 4.920 ;
        RECT 69.920 3.645 70.130 4.785 ;
        RECT 72.550 4.590 73.960 4.910 ;
        RECT 75.530 4.795 76.910 4.965 ;
        RECT 77.635 4.955 77.805 10.030 ;
        RECT 78.150 10.025 83.600 10.030 ;
        RECT 85.345 10.030 91.310 10.195 ;
        RECT 79.105 8.885 79.435 10.025 ;
        RECT 80.270 9.650 81.680 10.025 ;
        RECT 83.175 8.885 83.505 10.025 ;
        RECT 71.720 4.370 74.690 4.590 ;
        RECT 71.730 3.550 71.900 4.370 ;
        RECT 74.520 3.550 74.690 4.370 ;
        RECT 75.870 3.655 76.080 4.795 ;
        RECT 77.290 4.785 78.670 4.955 ;
        RECT 80.260 4.910 80.830 4.920 ;
        RECT 77.630 3.645 77.840 4.785 ;
        RECT 80.260 4.590 81.670 4.910 ;
        RECT 83.240 4.795 84.620 4.965 ;
        RECT 85.345 4.955 85.515 10.030 ;
        RECT 85.860 10.025 91.310 10.030 ;
        RECT 93.055 10.030 99.020 10.195 ;
        RECT 86.815 8.885 87.145 10.025 ;
        RECT 87.980 9.650 89.390 10.025 ;
        RECT 90.885 8.885 91.215 10.025 ;
        RECT 79.430 4.370 82.400 4.590 ;
        RECT 79.440 3.550 79.610 4.370 ;
        RECT 82.230 3.550 82.400 4.370 ;
        RECT 83.580 3.655 83.790 4.795 ;
        RECT 85.000 4.785 86.380 4.955 ;
        RECT 87.970 4.910 88.540 4.920 ;
        RECT 85.340 3.645 85.550 4.785 ;
        RECT 87.970 4.590 89.380 4.910 ;
        RECT 90.950 4.795 92.330 4.965 ;
        RECT 93.055 4.955 93.225 10.030 ;
        RECT 93.570 10.025 99.020 10.030 ;
        RECT 100.765 10.030 106.730 10.195 ;
        RECT 94.525 8.885 94.855 10.025 ;
        RECT 95.690 9.650 97.100 10.025 ;
        RECT 98.595 8.885 98.925 10.025 ;
        RECT 87.140 4.370 90.110 4.590 ;
        RECT 87.150 3.550 87.320 4.370 ;
        RECT 89.940 3.550 90.110 4.370 ;
        RECT 91.290 3.655 91.500 4.795 ;
        RECT 92.710 4.785 94.090 4.955 ;
        RECT 95.680 4.910 96.250 4.920 ;
        RECT 93.050 3.645 93.260 4.785 ;
        RECT 95.680 4.590 97.090 4.910 ;
        RECT 98.660 4.795 100.040 4.965 ;
        RECT 100.765 4.955 100.935 10.030 ;
        RECT 101.280 10.025 106.730 10.030 ;
        RECT 108.475 10.030 114.440 10.195 ;
        RECT 102.235 8.885 102.565 10.025 ;
        RECT 103.400 9.650 104.810 10.025 ;
        RECT 106.305 8.885 106.635 10.025 ;
        RECT 94.850 4.370 97.820 4.590 ;
        RECT 94.860 3.550 95.030 4.370 ;
        RECT 97.650 3.550 97.820 4.370 ;
        RECT 99.000 3.655 99.210 4.795 ;
        RECT 100.420 4.785 101.800 4.955 ;
        RECT 103.390 4.910 103.960 4.920 ;
        RECT 100.760 3.645 100.970 4.785 ;
        RECT 103.390 4.590 104.800 4.910 ;
        RECT 106.370 4.795 107.750 4.965 ;
        RECT 108.475 4.955 108.645 10.030 ;
        RECT 108.990 10.025 114.440 10.030 ;
        RECT 116.185 10.030 122.150 10.195 ;
        RECT 109.945 8.885 110.275 10.025 ;
        RECT 111.110 9.650 112.520 10.025 ;
        RECT 114.015 8.885 114.345 10.025 ;
        RECT 102.560 4.370 105.530 4.590 ;
        RECT 102.570 3.550 102.740 4.370 ;
        RECT 105.360 3.550 105.530 4.370 ;
        RECT 106.710 3.655 106.920 4.795 ;
        RECT 108.130 4.785 109.510 4.955 ;
        RECT 111.100 4.910 111.670 4.920 ;
        RECT 108.470 3.645 108.680 4.785 ;
        RECT 111.100 4.590 112.510 4.910 ;
        RECT 114.080 4.795 115.460 4.965 ;
        RECT 116.185 4.955 116.355 10.030 ;
        RECT 116.700 10.025 122.150 10.030 ;
        RECT 117.655 8.885 117.985 10.025 ;
        RECT 118.820 9.650 120.230 10.025 ;
        RECT 121.725 8.885 122.055 10.025 ;
        RECT 110.270 4.370 113.240 4.590 ;
        RECT 110.280 3.550 110.450 4.370 ;
        RECT 113.070 3.550 113.240 4.370 ;
        RECT 114.420 3.655 114.630 4.795 ;
        RECT 115.840 4.785 117.220 4.955 ;
        RECT 118.810 4.910 119.380 4.920 ;
        RECT 116.180 3.645 116.390 4.785 ;
        RECT 118.810 4.590 120.220 4.910 ;
        RECT 121.790 4.795 123.170 4.965 ;
        RECT 117.980 4.370 120.950 4.590 ;
        RECT 117.990 3.550 118.160 4.370 ;
        RECT 120.780 3.550 120.950 4.370 ;
        RECT 122.130 3.655 122.340 4.795 ;
      LAYER mcon ;
        RECT 2.090 28.950 2.260 29.830 ;
        RECT 4.880 28.950 5.050 29.830 ;
        RECT 3.840 28.710 4.060 28.950 ;
        RECT 0.015 28.495 0.185 28.665 ;
        RECT 0.475 28.495 0.645 28.665 ;
        RECT 0.935 28.495 1.105 28.665 ;
        RECT 5.965 28.505 6.135 28.675 ;
        RECT 6.425 28.505 6.595 28.675 ;
        RECT 6.885 28.505 7.055 28.675 ;
        RECT 9.800 28.950 9.970 29.830 ;
        RECT 12.590 28.950 12.760 29.830 ;
        RECT 11.550 28.710 11.770 28.950 ;
        RECT 1.035 23.265 1.205 23.435 ;
        RECT 1.495 23.265 1.665 23.435 ;
        RECT 1.955 23.265 2.125 23.435 ;
        RECT 3.830 23.430 4.050 23.670 ;
        RECT 5.105 23.265 5.275 23.435 ;
        RECT 5.565 23.265 5.735 23.435 ;
        RECT 6.025 23.265 6.195 23.435 ;
        RECT 7.725 28.495 7.895 28.665 ;
        RECT 8.185 28.495 8.355 28.665 ;
        RECT 8.645 28.495 8.815 28.665 ;
        RECT 13.675 28.505 13.845 28.675 ;
        RECT 14.135 28.505 14.305 28.675 ;
        RECT 14.595 28.505 14.765 28.675 ;
        RECT 17.510 28.950 17.680 29.830 ;
        RECT 20.300 28.950 20.470 29.830 ;
        RECT 19.260 28.710 19.480 28.950 ;
        RECT 8.745 23.265 8.915 23.435 ;
        RECT 9.205 23.265 9.375 23.435 ;
        RECT 9.665 23.265 9.835 23.435 ;
        RECT 11.540 23.430 11.760 23.670 ;
        RECT 12.815 23.265 12.985 23.435 ;
        RECT 13.275 23.265 13.445 23.435 ;
        RECT 13.735 23.265 13.905 23.435 ;
        RECT 15.435 28.495 15.605 28.665 ;
        RECT 15.895 28.495 16.065 28.665 ;
        RECT 16.355 28.495 16.525 28.665 ;
        RECT 21.385 28.505 21.555 28.675 ;
        RECT 21.845 28.505 22.015 28.675 ;
        RECT 22.305 28.505 22.475 28.675 ;
        RECT 25.220 28.950 25.390 29.830 ;
        RECT 28.010 28.950 28.180 29.830 ;
        RECT 26.970 28.710 27.190 28.950 ;
        RECT 16.455 23.265 16.625 23.435 ;
        RECT 16.915 23.265 17.085 23.435 ;
        RECT 17.375 23.265 17.545 23.435 ;
        RECT 19.250 23.430 19.470 23.670 ;
        RECT 20.525 23.265 20.695 23.435 ;
        RECT 20.985 23.265 21.155 23.435 ;
        RECT 21.445 23.265 21.615 23.435 ;
        RECT 23.145 28.495 23.315 28.665 ;
        RECT 23.605 28.495 23.775 28.665 ;
        RECT 24.065 28.495 24.235 28.665 ;
        RECT 29.095 28.505 29.265 28.675 ;
        RECT 29.555 28.505 29.725 28.675 ;
        RECT 30.015 28.505 30.185 28.675 ;
        RECT 32.930 28.950 33.100 29.830 ;
        RECT 35.720 28.950 35.890 29.830 ;
        RECT 34.680 28.710 34.900 28.950 ;
        RECT 24.165 23.265 24.335 23.435 ;
        RECT 24.625 23.265 24.795 23.435 ;
        RECT 25.085 23.265 25.255 23.435 ;
        RECT 26.960 23.430 27.180 23.670 ;
        RECT 28.235 23.265 28.405 23.435 ;
        RECT 28.695 23.265 28.865 23.435 ;
        RECT 29.155 23.265 29.325 23.435 ;
        RECT 30.855 28.495 31.025 28.665 ;
        RECT 31.315 28.495 31.485 28.665 ;
        RECT 31.775 28.495 31.945 28.665 ;
        RECT 36.805 28.505 36.975 28.675 ;
        RECT 37.265 28.505 37.435 28.675 ;
        RECT 37.725 28.505 37.895 28.675 ;
        RECT 40.640 28.950 40.810 29.830 ;
        RECT 43.430 28.950 43.600 29.830 ;
        RECT 42.390 28.710 42.610 28.950 ;
        RECT 31.875 23.265 32.045 23.435 ;
        RECT 32.335 23.265 32.505 23.435 ;
        RECT 32.795 23.265 32.965 23.435 ;
        RECT 34.670 23.430 34.890 23.670 ;
        RECT 35.945 23.265 36.115 23.435 ;
        RECT 36.405 23.265 36.575 23.435 ;
        RECT 36.865 23.265 37.035 23.435 ;
        RECT 38.565 28.495 38.735 28.665 ;
        RECT 39.025 28.495 39.195 28.665 ;
        RECT 39.485 28.495 39.655 28.665 ;
        RECT 44.515 28.505 44.685 28.675 ;
        RECT 44.975 28.505 45.145 28.675 ;
        RECT 45.435 28.505 45.605 28.675 ;
        RECT 48.350 28.950 48.520 29.830 ;
        RECT 51.140 28.950 51.310 29.830 ;
        RECT 50.100 28.710 50.320 28.950 ;
        RECT 39.585 23.265 39.755 23.435 ;
        RECT 40.045 23.265 40.215 23.435 ;
        RECT 40.505 23.265 40.675 23.435 ;
        RECT 42.380 23.430 42.600 23.670 ;
        RECT 43.655 23.265 43.825 23.435 ;
        RECT 44.115 23.265 44.285 23.435 ;
        RECT 44.575 23.265 44.745 23.435 ;
        RECT 46.275 28.495 46.445 28.665 ;
        RECT 46.735 28.495 46.905 28.665 ;
        RECT 47.195 28.495 47.365 28.665 ;
        RECT 52.225 28.505 52.395 28.675 ;
        RECT 52.685 28.505 52.855 28.675 ;
        RECT 53.145 28.505 53.315 28.675 ;
        RECT 56.060 28.950 56.230 29.830 ;
        RECT 58.850 28.950 59.020 29.830 ;
        RECT 57.810 28.710 58.030 28.950 ;
        RECT 47.295 23.265 47.465 23.435 ;
        RECT 47.755 23.265 47.925 23.435 ;
        RECT 48.215 23.265 48.385 23.435 ;
        RECT 50.090 23.430 50.310 23.670 ;
        RECT 51.365 23.265 51.535 23.435 ;
        RECT 51.825 23.265 51.995 23.435 ;
        RECT 52.285 23.265 52.455 23.435 ;
        RECT 53.985 28.495 54.155 28.665 ;
        RECT 54.445 28.495 54.615 28.665 ;
        RECT 54.905 28.495 55.075 28.665 ;
        RECT 59.935 28.505 60.105 28.675 ;
        RECT 60.395 28.505 60.565 28.675 ;
        RECT 60.855 28.505 61.025 28.675 ;
        RECT 63.770 28.950 63.940 29.830 ;
        RECT 66.560 28.950 66.730 29.830 ;
        RECT 65.520 28.710 65.740 28.950 ;
        RECT 55.005 23.265 55.175 23.435 ;
        RECT 55.465 23.265 55.635 23.435 ;
        RECT 55.925 23.265 56.095 23.435 ;
        RECT 57.800 23.430 58.020 23.670 ;
        RECT 59.075 23.265 59.245 23.435 ;
        RECT 59.535 23.265 59.705 23.435 ;
        RECT 59.995 23.265 60.165 23.435 ;
        RECT 61.695 28.495 61.865 28.665 ;
        RECT 62.155 28.495 62.325 28.665 ;
        RECT 62.615 28.495 62.785 28.665 ;
        RECT 67.645 28.505 67.815 28.675 ;
        RECT 68.105 28.505 68.275 28.675 ;
        RECT 68.565 28.505 68.735 28.675 ;
        RECT 71.480 28.950 71.650 29.830 ;
        RECT 74.270 28.950 74.440 29.830 ;
        RECT 73.230 28.710 73.450 28.950 ;
        RECT 62.715 23.265 62.885 23.435 ;
        RECT 63.175 23.265 63.345 23.435 ;
        RECT 63.635 23.265 63.805 23.435 ;
        RECT 65.510 23.430 65.730 23.670 ;
        RECT 66.785 23.265 66.955 23.435 ;
        RECT 67.245 23.265 67.415 23.435 ;
        RECT 67.705 23.265 67.875 23.435 ;
        RECT 69.405 28.495 69.575 28.665 ;
        RECT 69.865 28.495 70.035 28.665 ;
        RECT 70.325 28.495 70.495 28.665 ;
        RECT 75.355 28.505 75.525 28.675 ;
        RECT 75.815 28.505 75.985 28.675 ;
        RECT 76.275 28.505 76.445 28.675 ;
        RECT 79.190 28.950 79.360 29.830 ;
        RECT 81.980 28.950 82.150 29.830 ;
        RECT 80.940 28.710 81.160 28.950 ;
        RECT 70.425 23.265 70.595 23.435 ;
        RECT 70.885 23.265 71.055 23.435 ;
        RECT 71.345 23.265 71.515 23.435 ;
        RECT 73.220 23.430 73.440 23.670 ;
        RECT 74.495 23.265 74.665 23.435 ;
        RECT 74.955 23.265 75.125 23.435 ;
        RECT 75.415 23.265 75.585 23.435 ;
        RECT 77.115 28.495 77.285 28.665 ;
        RECT 77.575 28.495 77.745 28.665 ;
        RECT 78.035 28.495 78.205 28.665 ;
        RECT 83.065 28.505 83.235 28.675 ;
        RECT 83.525 28.505 83.695 28.675 ;
        RECT 83.985 28.505 84.155 28.675 ;
        RECT 86.900 28.950 87.070 29.830 ;
        RECT 89.690 28.950 89.860 29.830 ;
        RECT 88.650 28.710 88.870 28.950 ;
        RECT 78.135 23.265 78.305 23.435 ;
        RECT 78.595 23.265 78.765 23.435 ;
        RECT 79.055 23.265 79.225 23.435 ;
        RECT 80.930 23.430 81.150 23.670 ;
        RECT 82.205 23.265 82.375 23.435 ;
        RECT 82.665 23.265 82.835 23.435 ;
        RECT 83.125 23.265 83.295 23.435 ;
        RECT 84.825 28.495 84.995 28.665 ;
        RECT 85.285 28.495 85.455 28.665 ;
        RECT 85.745 28.495 85.915 28.665 ;
        RECT 90.775 28.505 90.945 28.675 ;
        RECT 91.235 28.505 91.405 28.675 ;
        RECT 91.695 28.505 91.865 28.675 ;
        RECT 94.610 28.950 94.780 29.830 ;
        RECT 97.400 28.950 97.570 29.830 ;
        RECT 96.360 28.710 96.580 28.950 ;
        RECT 85.845 23.265 86.015 23.435 ;
        RECT 86.305 23.265 86.475 23.435 ;
        RECT 86.765 23.265 86.935 23.435 ;
        RECT 88.640 23.430 88.860 23.670 ;
        RECT 89.915 23.265 90.085 23.435 ;
        RECT 90.375 23.265 90.545 23.435 ;
        RECT 90.835 23.265 91.005 23.435 ;
        RECT 92.535 28.495 92.705 28.665 ;
        RECT 92.995 28.495 93.165 28.665 ;
        RECT 93.455 28.495 93.625 28.665 ;
        RECT 98.485 28.505 98.655 28.675 ;
        RECT 98.945 28.505 99.115 28.675 ;
        RECT 99.405 28.505 99.575 28.675 ;
        RECT 102.320 28.950 102.490 29.830 ;
        RECT 105.110 28.950 105.280 29.830 ;
        RECT 104.070 28.710 104.290 28.950 ;
        RECT 93.555 23.265 93.725 23.435 ;
        RECT 94.015 23.265 94.185 23.435 ;
        RECT 94.475 23.265 94.645 23.435 ;
        RECT 96.350 23.430 96.570 23.670 ;
        RECT 97.625 23.265 97.795 23.435 ;
        RECT 98.085 23.265 98.255 23.435 ;
        RECT 98.545 23.265 98.715 23.435 ;
        RECT 100.245 28.495 100.415 28.665 ;
        RECT 100.705 28.495 100.875 28.665 ;
        RECT 101.165 28.495 101.335 28.665 ;
        RECT 106.195 28.505 106.365 28.675 ;
        RECT 106.655 28.505 106.825 28.675 ;
        RECT 107.115 28.505 107.285 28.675 ;
        RECT 110.030 28.950 110.200 29.830 ;
        RECT 112.820 28.950 112.990 29.830 ;
        RECT 111.780 28.710 112.000 28.950 ;
        RECT 101.265 23.265 101.435 23.435 ;
        RECT 101.725 23.265 101.895 23.435 ;
        RECT 102.185 23.265 102.355 23.435 ;
        RECT 104.060 23.430 104.280 23.670 ;
        RECT 105.335 23.265 105.505 23.435 ;
        RECT 105.795 23.265 105.965 23.435 ;
        RECT 106.255 23.265 106.425 23.435 ;
        RECT 107.955 28.495 108.125 28.665 ;
        RECT 108.415 28.495 108.585 28.665 ;
        RECT 108.875 28.495 109.045 28.665 ;
        RECT 113.905 28.505 114.075 28.675 ;
        RECT 114.365 28.505 114.535 28.675 ;
        RECT 114.825 28.505 114.995 28.675 ;
        RECT 117.740 28.950 117.910 29.830 ;
        RECT 120.530 28.950 120.700 29.830 ;
        RECT 119.490 28.710 119.710 28.950 ;
        RECT 108.975 23.265 109.145 23.435 ;
        RECT 109.435 23.265 109.605 23.435 ;
        RECT 109.895 23.265 110.065 23.435 ;
        RECT 111.770 23.430 111.990 23.670 ;
        RECT 113.045 23.265 113.215 23.435 ;
        RECT 113.505 23.265 113.675 23.435 ;
        RECT 113.965 23.265 114.135 23.435 ;
        RECT 115.665 28.495 115.835 28.665 ;
        RECT 116.125 28.495 116.295 28.665 ;
        RECT 116.585 28.495 116.755 28.665 ;
        RECT 121.615 28.505 121.785 28.675 ;
        RECT 122.075 28.505 122.245 28.675 ;
        RECT 122.535 28.505 122.705 28.675 ;
        RECT 116.685 23.265 116.855 23.435 ;
        RECT 117.145 23.265 117.315 23.435 ;
        RECT 117.605 23.265 117.775 23.435 ;
        RECT 119.480 23.430 119.700 23.670 ;
        RECT 120.755 23.265 120.925 23.435 ;
        RECT 121.215 23.265 121.385 23.435 ;
        RECT 121.675 23.265 121.845 23.435 ;
        RECT 22.345 19.115 22.515 19.285 ;
        RECT 22.805 19.115 22.975 19.285 ;
        RECT 23.265 19.115 23.435 19.285 ;
        RECT 23.725 19.115 23.895 19.285 ;
        RECT 24.185 19.115 24.355 19.285 ;
        RECT 24.645 19.115 24.815 19.285 ;
        RECT 25.105 19.115 25.275 19.285 ;
        RECT 25.565 19.115 25.735 19.285 ;
        RECT 26.025 19.115 26.195 19.285 ;
        RECT 26.485 19.115 26.655 19.285 ;
        RECT 26.945 19.115 27.115 19.285 ;
        RECT 27.405 19.115 27.575 19.285 ;
        RECT 27.865 19.115 28.035 19.285 ;
        RECT 28.325 19.115 28.495 19.285 ;
        RECT 28.785 19.115 28.955 19.285 ;
        RECT 29.245 19.115 29.415 19.285 ;
        RECT 84.005 19.145 84.175 19.315 ;
        RECT 84.465 19.145 84.635 19.315 ;
        RECT 84.925 19.145 85.095 19.315 ;
        RECT 85.385 19.145 85.555 19.315 ;
        RECT 85.845 19.145 86.015 19.315 ;
        RECT 86.305 19.145 86.475 19.315 ;
        RECT 86.765 19.145 86.935 19.315 ;
        RECT 87.225 19.145 87.395 19.315 ;
        RECT 87.685 19.145 87.855 19.315 ;
        RECT 88.145 19.145 88.315 19.315 ;
        RECT 88.605 19.145 88.775 19.315 ;
        RECT 89.065 19.145 89.235 19.315 ;
        RECT 89.525 19.145 89.695 19.315 ;
        RECT 89.985 19.145 90.155 19.315 ;
        RECT 90.445 19.145 90.615 19.315 ;
        RECT 90.905 19.145 91.075 19.315 ;
        RECT 55.555 18.375 55.725 18.545 ;
        RECT 56.015 18.375 56.185 18.545 ;
        RECT 56.475 18.375 56.645 18.545 ;
        RECT 56.935 18.375 57.105 18.545 ;
        RECT 57.395 18.375 57.565 18.545 ;
        RECT 57.855 18.375 58.025 18.545 ;
        RECT 58.315 18.375 58.485 18.545 ;
        RECT 58.775 18.375 58.945 18.545 ;
        RECT 59.235 18.375 59.405 18.545 ;
        RECT 55.595 18.015 55.765 18.185 ;
        RECT 56.055 18.015 56.225 18.185 ;
        RECT 56.515 18.015 56.685 18.185 ;
        RECT 57.255 18.005 57.425 18.175 ;
        RECT 57.715 18.005 57.885 18.175 ;
        RECT 58.175 18.005 58.345 18.175 ;
        RECT 58.635 18.005 58.805 18.175 ;
        RECT 59.095 18.005 59.265 18.175 ;
        RECT 124.545 17.445 124.715 17.615 ;
        RECT 125.005 17.445 125.175 17.615 ;
        RECT 125.465 17.445 125.635 17.615 ;
        RECT 22.475 13.585 22.645 13.755 ;
        RECT 22.935 13.585 23.105 13.755 ;
        RECT 23.395 13.585 23.565 13.755 ;
        RECT 23.855 13.585 24.025 13.755 ;
        RECT 24.315 13.585 24.485 13.755 ;
        RECT 24.775 13.585 24.945 13.755 ;
        RECT 25.235 13.585 25.405 13.755 ;
        RECT 25.695 13.585 25.865 13.755 ;
        RECT 26.155 13.585 26.325 13.755 ;
        RECT 26.615 13.585 26.785 13.755 ;
        RECT 27.075 13.585 27.245 13.755 ;
        RECT 27.535 13.585 27.705 13.755 ;
        RECT 27.995 13.585 28.165 13.755 ;
        RECT 28.455 13.585 28.625 13.755 ;
        RECT 28.915 13.585 29.085 13.755 ;
        RECT 29.375 13.585 29.545 13.755 ;
        RECT 84.135 13.555 84.305 13.725 ;
        RECT 84.595 13.555 84.765 13.725 ;
        RECT 85.055 13.555 85.225 13.725 ;
        RECT 85.515 13.555 85.685 13.725 ;
        RECT 85.975 13.555 86.145 13.725 ;
        RECT 86.435 13.555 86.605 13.725 ;
        RECT 86.895 13.555 87.065 13.725 ;
        RECT 87.355 13.555 87.525 13.725 ;
        RECT 87.815 13.555 87.985 13.725 ;
        RECT 88.275 13.555 88.445 13.725 ;
        RECT 88.735 13.555 88.905 13.725 ;
        RECT 89.195 13.555 89.365 13.725 ;
        RECT 89.655 13.555 89.825 13.725 ;
        RECT 90.115 13.555 90.285 13.725 ;
        RECT 90.575 13.555 90.745 13.725 ;
        RECT 91.035 13.555 91.205 13.725 ;
        RECT 55.535 12.165 55.705 12.335 ;
        RECT 55.995 12.165 56.165 12.335 ;
        RECT 56.455 12.165 56.625 12.335 ;
        RECT 56.915 12.165 57.085 12.335 ;
        RECT 57.375 12.165 57.545 12.335 ;
        RECT 57.835 12.165 58.005 12.335 ;
        RECT 58.295 12.165 58.465 12.335 ;
        RECT 58.755 12.165 58.925 12.335 ;
        RECT 59.215 12.165 59.385 12.335 ;
        RECT 1.195 10.025 1.365 10.195 ;
        RECT 1.655 10.025 1.825 10.195 ;
        RECT 2.115 10.025 2.285 10.195 ;
        RECT 3.340 9.790 3.560 10.030 ;
        RECT 5.265 10.025 5.435 10.195 ;
        RECT 5.725 10.025 5.895 10.195 ;
        RECT 6.185 10.025 6.355 10.195 ;
        RECT 0.335 4.785 0.505 4.955 ;
        RECT 0.795 4.785 0.965 4.955 ;
        RECT 1.255 4.785 1.425 4.955 ;
        RECT 6.285 4.795 6.455 4.965 ;
        RECT 6.745 4.795 6.915 4.965 ;
        RECT 7.205 4.795 7.375 4.965 ;
        RECT 8.905 10.025 9.075 10.195 ;
        RECT 9.365 10.025 9.535 10.195 ;
        RECT 9.825 10.025 9.995 10.195 ;
        RECT 11.050 9.790 11.270 10.030 ;
        RECT 12.975 10.025 13.145 10.195 ;
        RECT 13.435 10.025 13.605 10.195 ;
        RECT 13.895 10.025 14.065 10.195 ;
        RECT 3.330 4.510 3.550 4.750 ;
        RECT 2.340 3.630 2.510 4.510 ;
        RECT 5.130 3.630 5.300 4.510 ;
        RECT 8.045 4.785 8.215 4.955 ;
        RECT 8.505 4.785 8.675 4.955 ;
        RECT 8.965 4.785 9.135 4.955 ;
        RECT 13.995 4.795 14.165 4.965 ;
        RECT 14.455 4.795 14.625 4.965 ;
        RECT 14.915 4.795 15.085 4.965 ;
        RECT 16.615 10.025 16.785 10.195 ;
        RECT 17.075 10.025 17.245 10.195 ;
        RECT 17.535 10.025 17.705 10.195 ;
        RECT 18.760 9.790 18.980 10.030 ;
        RECT 20.685 10.025 20.855 10.195 ;
        RECT 21.145 10.025 21.315 10.195 ;
        RECT 21.605 10.025 21.775 10.195 ;
        RECT 11.040 4.510 11.260 4.750 ;
        RECT 10.050 3.630 10.220 4.510 ;
        RECT 12.840 3.630 13.010 4.510 ;
        RECT 15.755 4.785 15.925 4.955 ;
        RECT 16.215 4.785 16.385 4.955 ;
        RECT 16.675 4.785 16.845 4.955 ;
        RECT 21.705 4.795 21.875 4.965 ;
        RECT 22.165 4.795 22.335 4.965 ;
        RECT 22.625 4.795 22.795 4.965 ;
        RECT 24.325 10.025 24.495 10.195 ;
        RECT 24.785 10.025 24.955 10.195 ;
        RECT 25.245 10.025 25.415 10.195 ;
        RECT 26.470 9.790 26.690 10.030 ;
        RECT 28.395 10.025 28.565 10.195 ;
        RECT 28.855 10.025 29.025 10.195 ;
        RECT 29.315 10.025 29.485 10.195 ;
        RECT 18.750 4.510 18.970 4.750 ;
        RECT 17.760 3.630 17.930 4.510 ;
        RECT 20.550 3.630 20.720 4.510 ;
        RECT 23.465 4.785 23.635 4.955 ;
        RECT 23.925 4.785 24.095 4.955 ;
        RECT 24.385 4.785 24.555 4.955 ;
        RECT 29.415 4.795 29.585 4.965 ;
        RECT 29.875 4.795 30.045 4.965 ;
        RECT 30.335 4.795 30.505 4.965 ;
        RECT 32.035 10.025 32.205 10.195 ;
        RECT 32.495 10.025 32.665 10.195 ;
        RECT 32.955 10.025 33.125 10.195 ;
        RECT 34.180 9.790 34.400 10.030 ;
        RECT 36.105 10.025 36.275 10.195 ;
        RECT 36.565 10.025 36.735 10.195 ;
        RECT 37.025 10.025 37.195 10.195 ;
        RECT 26.460 4.510 26.680 4.750 ;
        RECT 25.470 3.630 25.640 4.510 ;
        RECT 28.260 3.630 28.430 4.510 ;
        RECT 31.175 4.785 31.345 4.955 ;
        RECT 31.635 4.785 31.805 4.955 ;
        RECT 32.095 4.785 32.265 4.955 ;
        RECT 37.125 4.795 37.295 4.965 ;
        RECT 37.585 4.795 37.755 4.965 ;
        RECT 38.045 4.795 38.215 4.965 ;
        RECT 39.745 10.025 39.915 10.195 ;
        RECT 40.205 10.025 40.375 10.195 ;
        RECT 40.665 10.025 40.835 10.195 ;
        RECT 41.890 9.790 42.110 10.030 ;
        RECT 43.815 10.025 43.985 10.195 ;
        RECT 44.275 10.025 44.445 10.195 ;
        RECT 44.735 10.025 44.905 10.195 ;
        RECT 34.170 4.510 34.390 4.750 ;
        RECT 33.180 3.630 33.350 4.510 ;
        RECT 35.970 3.630 36.140 4.510 ;
        RECT 38.885 4.785 39.055 4.955 ;
        RECT 39.345 4.785 39.515 4.955 ;
        RECT 39.805 4.785 39.975 4.955 ;
        RECT 44.835 4.795 45.005 4.965 ;
        RECT 45.295 4.795 45.465 4.965 ;
        RECT 45.755 4.795 45.925 4.965 ;
        RECT 47.455 10.025 47.625 10.195 ;
        RECT 47.915 10.025 48.085 10.195 ;
        RECT 48.375 10.025 48.545 10.195 ;
        RECT 49.600 9.790 49.820 10.030 ;
        RECT 51.525 10.025 51.695 10.195 ;
        RECT 51.985 10.025 52.155 10.195 ;
        RECT 52.445 10.025 52.615 10.195 ;
        RECT 41.880 4.510 42.100 4.750 ;
        RECT 40.890 3.630 41.060 4.510 ;
        RECT 43.680 3.630 43.850 4.510 ;
        RECT 46.595 4.785 46.765 4.955 ;
        RECT 47.055 4.785 47.225 4.955 ;
        RECT 47.515 4.785 47.685 4.955 ;
        RECT 52.545 4.795 52.715 4.965 ;
        RECT 53.005 4.795 53.175 4.965 ;
        RECT 53.465 4.795 53.635 4.965 ;
        RECT 55.165 10.025 55.335 10.195 ;
        RECT 55.625 10.025 55.795 10.195 ;
        RECT 56.085 10.025 56.255 10.195 ;
        RECT 57.310 9.790 57.530 10.030 ;
        RECT 59.235 10.025 59.405 10.195 ;
        RECT 59.695 10.025 59.865 10.195 ;
        RECT 60.155 10.025 60.325 10.195 ;
        RECT 49.590 4.510 49.810 4.750 ;
        RECT 48.600 3.630 48.770 4.510 ;
        RECT 51.390 3.630 51.560 4.510 ;
        RECT 54.305 4.785 54.475 4.955 ;
        RECT 54.765 4.785 54.935 4.955 ;
        RECT 55.225 4.785 55.395 4.955 ;
        RECT 60.255 4.795 60.425 4.965 ;
        RECT 60.715 4.795 60.885 4.965 ;
        RECT 61.175 4.795 61.345 4.965 ;
        RECT 62.875 10.025 63.045 10.195 ;
        RECT 63.335 10.025 63.505 10.195 ;
        RECT 63.795 10.025 63.965 10.195 ;
        RECT 65.020 9.790 65.240 10.030 ;
        RECT 66.945 10.025 67.115 10.195 ;
        RECT 67.405 10.025 67.575 10.195 ;
        RECT 67.865 10.025 68.035 10.195 ;
        RECT 57.300 4.510 57.520 4.750 ;
        RECT 56.310 3.630 56.480 4.510 ;
        RECT 59.100 3.630 59.270 4.510 ;
        RECT 62.015 4.785 62.185 4.955 ;
        RECT 62.475 4.785 62.645 4.955 ;
        RECT 62.935 4.785 63.105 4.955 ;
        RECT 67.965 4.795 68.135 4.965 ;
        RECT 68.425 4.795 68.595 4.965 ;
        RECT 68.885 4.795 69.055 4.965 ;
        RECT 70.585 10.025 70.755 10.195 ;
        RECT 71.045 10.025 71.215 10.195 ;
        RECT 71.505 10.025 71.675 10.195 ;
        RECT 72.730 9.790 72.950 10.030 ;
        RECT 74.655 10.025 74.825 10.195 ;
        RECT 75.115 10.025 75.285 10.195 ;
        RECT 75.575 10.025 75.745 10.195 ;
        RECT 65.010 4.510 65.230 4.750 ;
        RECT 64.020 3.630 64.190 4.510 ;
        RECT 66.810 3.630 66.980 4.510 ;
        RECT 69.725 4.785 69.895 4.955 ;
        RECT 70.185 4.785 70.355 4.955 ;
        RECT 70.645 4.785 70.815 4.955 ;
        RECT 75.675 4.795 75.845 4.965 ;
        RECT 76.135 4.795 76.305 4.965 ;
        RECT 76.595 4.795 76.765 4.965 ;
        RECT 78.295 10.025 78.465 10.195 ;
        RECT 78.755 10.025 78.925 10.195 ;
        RECT 79.215 10.025 79.385 10.195 ;
        RECT 80.440 9.790 80.660 10.030 ;
        RECT 82.365 10.025 82.535 10.195 ;
        RECT 82.825 10.025 82.995 10.195 ;
        RECT 83.285 10.025 83.455 10.195 ;
        RECT 72.720 4.510 72.940 4.750 ;
        RECT 71.730 3.630 71.900 4.510 ;
        RECT 74.520 3.630 74.690 4.510 ;
        RECT 77.435 4.785 77.605 4.955 ;
        RECT 77.895 4.785 78.065 4.955 ;
        RECT 78.355 4.785 78.525 4.955 ;
        RECT 83.385 4.795 83.555 4.965 ;
        RECT 83.845 4.795 84.015 4.965 ;
        RECT 84.305 4.795 84.475 4.965 ;
        RECT 86.005 10.025 86.175 10.195 ;
        RECT 86.465 10.025 86.635 10.195 ;
        RECT 86.925 10.025 87.095 10.195 ;
        RECT 88.150 9.790 88.370 10.030 ;
        RECT 90.075 10.025 90.245 10.195 ;
        RECT 90.535 10.025 90.705 10.195 ;
        RECT 90.995 10.025 91.165 10.195 ;
        RECT 80.430 4.510 80.650 4.750 ;
        RECT 79.440 3.630 79.610 4.510 ;
        RECT 82.230 3.630 82.400 4.510 ;
        RECT 85.145 4.785 85.315 4.955 ;
        RECT 85.605 4.785 85.775 4.955 ;
        RECT 86.065 4.785 86.235 4.955 ;
        RECT 91.095 4.795 91.265 4.965 ;
        RECT 91.555 4.795 91.725 4.965 ;
        RECT 92.015 4.795 92.185 4.965 ;
        RECT 93.715 10.025 93.885 10.195 ;
        RECT 94.175 10.025 94.345 10.195 ;
        RECT 94.635 10.025 94.805 10.195 ;
        RECT 95.860 9.790 96.080 10.030 ;
        RECT 97.785 10.025 97.955 10.195 ;
        RECT 98.245 10.025 98.415 10.195 ;
        RECT 98.705 10.025 98.875 10.195 ;
        RECT 88.140 4.510 88.360 4.750 ;
        RECT 87.150 3.630 87.320 4.510 ;
        RECT 89.940 3.630 90.110 4.510 ;
        RECT 92.855 4.785 93.025 4.955 ;
        RECT 93.315 4.785 93.485 4.955 ;
        RECT 93.775 4.785 93.945 4.955 ;
        RECT 98.805 4.795 98.975 4.965 ;
        RECT 99.265 4.795 99.435 4.965 ;
        RECT 99.725 4.795 99.895 4.965 ;
        RECT 101.425 10.025 101.595 10.195 ;
        RECT 101.885 10.025 102.055 10.195 ;
        RECT 102.345 10.025 102.515 10.195 ;
        RECT 103.570 9.790 103.790 10.030 ;
        RECT 105.495 10.025 105.665 10.195 ;
        RECT 105.955 10.025 106.125 10.195 ;
        RECT 106.415 10.025 106.585 10.195 ;
        RECT 95.850 4.510 96.070 4.750 ;
        RECT 94.860 3.630 95.030 4.510 ;
        RECT 97.650 3.630 97.820 4.510 ;
        RECT 100.565 4.785 100.735 4.955 ;
        RECT 101.025 4.785 101.195 4.955 ;
        RECT 101.485 4.785 101.655 4.955 ;
        RECT 106.515 4.795 106.685 4.965 ;
        RECT 106.975 4.795 107.145 4.965 ;
        RECT 107.435 4.795 107.605 4.965 ;
        RECT 109.135 10.025 109.305 10.195 ;
        RECT 109.595 10.025 109.765 10.195 ;
        RECT 110.055 10.025 110.225 10.195 ;
        RECT 111.280 9.790 111.500 10.030 ;
        RECT 113.205 10.025 113.375 10.195 ;
        RECT 113.665 10.025 113.835 10.195 ;
        RECT 114.125 10.025 114.295 10.195 ;
        RECT 103.560 4.510 103.780 4.750 ;
        RECT 102.570 3.630 102.740 4.510 ;
        RECT 105.360 3.630 105.530 4.510 ;
        RECT 108.275 4.785 108.445 4.955 ;
        RECT 108.735 4.785 108.905 4.955 ;
        RECT 109.195 4.785 109.365 4.955 ;
        RECT 114.225 4.795 114.395 4.965 ;
        RECT 114.685 4.795 114.855 4.965 ;
        RECT 115.145 4.795 115.315 4.965 ;
        RECT 116.845 10.025 117.015 10.195 ;
        RECT 117.305 10.025 117.475 10.195 ;
        RECT 117.765 10.025 117.935 10.195 ;
        RECT 118.990 9.790 119.210 10.030 ;
        RECT 120.915 10.025 121.085 10.195 ;
        RECT 121.375 10.025 121.545 10.195 ;
        RECT 121.835 10.025 122.005 10.195 ;
        RECT 111.270 4.510 111.490 4.750 ;
        RECT 110.280 3.630 110.450 4.510 ;
        RECT 113.070 3.630 113.240 4.510 ;
        RECT 115.985 4.785 116.155 4.955 ;
        RECT 116.445 4.785 116.615 4.955 ;
        RECT 116.905 4.785 117.075 4.955 ;
        RECT 121.935 4.795 122.105 4.965 ;
        RECT 122.395 4.795 122.565 4.965 ;
        RECT 122.855 4.795 123.025 4.965 ;
        RECT 118.980 4.510 119.200 4.750 ;
        RECT 117.990 3.630 118.160 4.510 ;
        RECT 120.780 3.630 120.950 4.510 ;
      LAYER met1 ;
        RECT 2.060 29.210 2.290 29.890 ;
        RECT 4.850 29.320 5.080 29.890 ;
        RECT 2.000 28.890 2.330 29.210 ;
        RECT -0.130 28.340 1.250 28.820 ;
        RECT 3.730 28.640 4.180 29.020 ;
        RECT 4.740 28.990 5.080 29.320 ;
        RECT 9.770 29.210 10.000 29.890 ;
        RECT 12.560 29.320 12.790 29.890 ;
        RECT 4.850 28.890 5.080 28.990 ;
        RECT 9.710 28.890 10.040 29.210 ;
        RECT 5.820 28.350 7.200 28.830 ;
        RECT 7.580 28.340 8.960 28.820 ;
        RECT 11.440 28.640 11.890 29.020 ;
        RECT 12.450 28.990 12.790 29.320 ;
        RECT 17.480 29.210 17.710 29.890 ;
        RECT 20.270 29.320 20.500 29.890 ;
        RECT 12.560 28.890 12.790 28.990 ;
        RECT 17.420 28.890 17.750 29.210 ;
        RECT 13.530 28.350 14.910 28.830 ;
        RECT 15.290 28.340 16.670 28.820 ;
        RECT 19.150 28.640 19.600 29.020 ;
        RECT 20.160 28.990 20.500 29.320 ;
        RECT 25.190 29.210 25.420 29.890 ;
        RECT 27.980 29.320 28.210 29.890 ;
        RECT 20.270 28.890 20.500 28.990 ;
        RECT 25.130 28.890 25.460 29.210 ;
        RECT 21.240 28.350 22.620 28.830 ;
        RECT 23.000 28.340 24.380 28.820 ;
        RECT 26.860 28.640 27.310 29.020 ;
        RECT 27.870 28.990 28.210 29.320 ;
        RECT 32.900 29.210 33.130 29.890 ;
        RECT 35.690 29.320 35.920 29.890 ;
        RECT 27.980 28.890 28.210 28.990 ;
        RECT 32.840 28.890 33.170 29.210 ;
        RECT 28.950 28.350 30.330 28.830 ;
        RECT 30.710 28.340 32.090 28.820 ;
        RECT 34.570 28.640 35.020 29.020 ;
        RECT 35.580 28.990 35.920 29.320 ;
        RECT 40.610 29.210 40.840 29.890 ;
        RECT 43.400 29.320 43.630 29.890 ;
        RECT 35.690 28.890 35.920 28.990 ;
        RECT 40.550 28.890 40.880 29.210 ;
        RECT 36.660 28.350 38.040 28.830 ;
        RECT 38.420 28.340 39.800 28.820 ;
        RECT 42.280 28.640 42.730 29.020 ;
        RECT 43.290 28.990 43.630 29.320 ;
        RECT 48.320 29.210 48.550 29.890 ;
        RECT 51.110 29.320 51.340 29.890 ;
        RECT 43.400 28.890 43.630 28.990 ;
        RECT 48.260 28.890 48.590 29.210 ;
        RECT 44.370 28.350 45.750 28.830 ;
        RECT 46.130 28.340 47.510 28.820 ;
        RECT 49.990 28.640 50.440 29.020 ;
        RECT 51.000 28.990 51.340 29.320 ;
        RECT 56.030 29.210 56.260 29.890 ;
        RECT 58.820 29.320 59.050 29.890 ;
        RECT 51.110 28.890 51.340 28.990 ;
        RECT 55.970 28.890 56.300 29.210 ;
        RECT 52.080 28.350 53.460 28.830 ;
        RECT 53.840 28.340 55.220 28.820 ;
        RECT 57.700 28.640 58.150 29.020 ;
        RECT 58.710 28.990 59.050 29.320 ;
        RECT 63.740 29.210 63.970 29.890 ;
        RECT 66.530 29.320 66.760 29.890 ;
        RECT 58.820 28.890 59.050 28.990 ;
        RECT 63.680 28.890 64.010 29.210 ;
        RECT 59.790 28.350 61.170 28.830 ;
        RECT 61.550 28.340 62.930 28.820 ;
        RECT 65.410 28.640 65.860 29.020 ;
        RECT 66.420 28.990 66.760 29.320 ;
        RECT 71.450 29.210 71.680 29.890 ;
        RECT 74.240 29.320 74.470 29.890 ;
        RECT 66.530 28.890 66.760 28.990 ;
        RECT 71.390 28.890 71.720 29.210 ;
        RECT 67.500 28.350 68.880 28.830 ;
        RECT 69.260 28.340 70.640 28.820 ;
        RECT 73.120 28.640 73.570 29.020 ;
        RECT 74.130 28.990 74.470 29.320 ;
        RECT 79.160 29.210 79.390 29.890 ;
        RECT 81.950 29.320 82.180 29.890 ;
        RECT 74.240 28.890 74.470 28.990 ;
        RECT 79.100 28.890 79.430 29.210 ;
        RECT 75.210 28.350 76.590 28.830 ;
        RECT 76.970 28.340 78.350 28.820 ;
        RECT 80.830 28.640 81.280 29.020 ;
        RECT 81.840 28.990 82.180 29.320 ;
        RECT 86.870 29.210 87.100 29.890 ;
        RECT 89.660 29.320 89.890 29.890 ;
        RECT 81.950 28.890 82.180 28.990 ;
        RECT 86.810 28.890 87.140 29.210 ;
        RECT 82.920 28.350 84.300 28.830 ;
        RECT 84.680 28.340 86.060 28.820 ;
        RECT 88.540 28.640 88.990 29.020 ;
        RECT 89.550 28.990 89.890 29.320 ;
        RECT 94.580 29.210 94.810 29.890 ;
        RECT 97.370 29.320 97.600 29.890 ;
        RECT 89.660 28.890 89.890 28.990 ;
        RECT 94.520 28.890 94.850 29.210 ;
        RECT 90.630 28.350 92.010 28.830 ;
        RECT 92.390 28.340 93.770 28.820 ;
        RECT 96.250 28.640 96.700 29.020 ;
        RECT 97.260 28.990 97.600 29.320 ;
        RECT 102.290 29.210 102.520 29.890 ;
        RECT 105.080 29.320 105.310 29.890 ;
        RECT 97.370 28.890 97.600 28.990 ;
        RECT 102.230 28.890 102.560 29.210 ;
        RECT 98.340 28.350 99.720 28.830 ;
        RECT 100.100 28.340 101.480 28.820 ;
        RECT 103.960 28.640 104.410 29.020 ;
        RECT 104.970 28.990 105.310 29.320 ;
        RECT 110.000 29.210 110.230 29.890 ;
        RECT 112.790 29.320 113.020 29.890 ;
        RECT 105.080 28.890 105.310 28.990 ;
        RECT 109.940 28.890 110.270 29.210 ;
        RECT 106.050 28.350 107.430 28.830 ;
        RECT 107.810 28.340 109.190 28.820 ;
        RECT 111.670 28.640 112.120 29.020 ;
        RECT 112.680 28.990 113.020 29.320 ;
        RECT 117.710 29.210 117.940 29.890 ;
        RECT 120.500 29.320 120.730 29.890 ;
        RECT 112.790 28.890 113.020 28.990 ;
        RECT 117.650 28.890 117.980 29.210 ;
        RECT 113.760 28.350 115.140 28.830 ;
        RECT 115.520 28.340 116.900 28.820 ;
        RECT 119.380 28.640 119.830 29.020 ;
        RECT 120.390 28.990 120.730 29.320 ;
        RECT 120.500 28.890 120.730 28.990 ;
        RECT 121.470 28.350 122.850 28.830 ;
        RECT 3.720 23.590 4.170 23.740 ;
        RECT 11.430 23.590 11.880 23.740 ;
        RECT 19.140 23.590 19.590 23.740 ;
        RECT 26.850 23.590 27.300 23.740 ;
        RECT 34.560 23.590 35.010 23.740 ;
        RECT 42.270 23.590 42.720 23.740 ;
        RECT 49.980 23.590 50.430 23.740 ;
        RECT 57.690 23.590 58.140 23.740 ;
        RECT 65.400 23.590 65.850 23.740 ;
        RECT 73.110 23.590 73.560 23.740 ;
        RECT 80.820 23.590 81.270 23.740 ;
        RECT 88.530 23.590 88.980 23.740 ;
        RECT 96.240 23.590 96.690 23.740 ;
        RECT 103.950 23.590 104.400 23.740 ;
        RECT 111.660 23.590 112.110 23.740 ;
        RECT 119.370 23.590 119.820 23.740 ;
        RECT -0.320 23.110 124.760 23.590 ;
        RECT 22.200 19.420 29.560 19.440 ;
        RECT 29.870 19.420 30.280 23.110 ;
        RECT 22.200 19.015 30.280 19.420 ;
        RECT 83.135 19.390 83.505 23.110 ;
        RECT 124.280 22.470 124.760 23.110 ;
        RECT 124.260 22.260 124.760 22.470 ;
        RECT 83.860 19.390 91.340 19.470 ;
        RECT 83.135 19.020 91.340 19.390 ;
        RECT 22.200 18.960 29.560 19.015 ;
        RECT 29.870 19.010 30.280 19.015 ;
        RECT 83.860 18.990 91.340 19.020 ;
        RECT 22.200 13.910 22.720 18.960 ;
        RECT 55.410 18.470 59.550 18.700 ;
        RECT 54.435 18.220 59.550 18.470 ;
        RECT 54.435 18.000 56.830 18.220 ;
        RECT 22.200 13.810 29.690 13.910 ;
        RECT 22.200 13.435 30.275 13.810 ;
        RECT 22.200 13.430 29.690 13.435 ;
        RECT 29.900 10.350 30.270 13.435 ;
        RECT 54.435 12.515 54.905 18.000 ;
        RECT 55.450 17.860 56.830 18.000 ;
        RECT 57.110 17.850 59.410 18.220 ;
        RECT 90.830 13.880 91.340 18.990 ;
        RECT 124.260 17.770 124.740 22.260 ;
        RECT 124.260 17.310 125.780 17.770 ;
        RECT 124.400 17.290 125.780 17.310 ;
        RECT 83.990 13.830 91.350 13.880 ;
        RECT 83.345 13.455 91.350 13.830 ;
        RECT 54.435 12.490 55.875 12.515 ;
        RECT 54.435 12.045 59.530 12.490 ;
        RECT 54.435 10.350 54.905 12.045 ;
        RECT 55.390 12.010 59.530 12.045 ;
        RECT 83.345 10.350 83.720 13.455 ;
        RECT 83.990 13.400 91.350 13.455 ;
        RECT 0.000 9.870 123.360 10.350 ;
        RECT 3.220 9.720 3.670 9.870 ;
        RECT 10.930 9.720 11.380 9.870 ;
        RECT 18.640 9.720 19.090 9.870 ;
        RECT 26.350 9.720 26.800 9.870 ;
        RECT 34.060 9.720 34.510 9.870 ;
        RECT 41.770 9.720 42.220 9.870 ;
        RECT 49.480 9.720 49.930 9.870 ;
        RECT 54.435 9.865 55.165 9.870 ;
        RECT 57.190 9.720 57.640 9.870 ;
        RECT 64.900 9.720 65.350 9.870 ;
        RECT 72.610 9.720 73.060 9.870 ;
        RECT 80.320 9.720 80.770 9.870 ;
        RECT 88.030 9.720 88.480 9.870 ;
        RECT 95.740 9.720 96.190 9.870 ;
        RECT 103.450 9.720 103.900 9.870 ;
        RECT 111.160 9.720 111.610 9.870 ;
        RECT 118.870 9.720 119.320 9.870 ;
        RECT 0.190 4.630 1.570 5.110 ;
        RECT 2.310 4.470 2.540 4.570 ;
        RECT 2.310 4.140 2.650 4.470 ;
        RECT 3.210 4.440 3.660 4.820 ;
        RECT 6.140 4.640 7.520 5.120 ;
        RECT 7.900 4.630 9.280 5.110 ;
        RECT 5.060 4.250 5.390 4.570 ;
        RECT 10.020 4.470 10.250 4.570 ;
        RECT 2.310 3.570 2.540 4.140 ;
        RECT 5.100 3.570 5.330 4.250 ;
        RECT 10.020 4.140 10.360 4.470 ;
        RECT 10.920 4.440 11.370 4.820 ;
        RECT 13.850 4.640 15.230 5.120 ;
        RECT 15.610 4.630 16.990 5.110 ;
        RECT 12.770 4.250 13.100 4.570 ;
        RECT 17.730 4.470 17.960 4.570 ;
        RECT 10.020 3.570 10.250 4.140 ;
        RECT 12.810 3.570 13.040 4.250 ;
        RECT 17.730 4.140 18.070 4.470 ;
        RECT 18.630 4.440 19.080 4.820 ;
        RECT 21.560 4.640 22.940 5.120 ;
        RECT 23.320 4.630 24.700 5.110 ;
        RECT 20.480 4.250 20.810 4.570 ;
        RECT 25.440 4.470 25.670 4.570 ;
        RECT 17.730 3.570 17.960 4.140 ;
        RECT 20.520 3.570 20.750 4.250 ;
        RECT 25.440 4.140 25.780 4.470 ;
        RECT 26.340 4.440 26.790 4.820 ;
        RECT 29.270 4.640 30.650 5.120 ;
        RECT 31.030 4.630 32.410 5.110 ;
        RECT 28.190 4.250 28.520 4.570 ;
        RECT 33.150 4.470 33.380 4.570 ;
        RECT 25.440 3.570 25.670 4.140 ;
        RECT 28.230 3.570 28.460 4.250 ;
        RECT 33.150 4.140 33.490 4.470 ;
        RECT 34.050 4.440 34.500 4.820 ;
        RECT 36.980 4.640 38.360 5.120 ;
        RECT 38.740 4.630 40.120 5.110 ;
        RECT 35.900 4.250 36.230 4.570 ;
        RECT 40.860 4.470 41.090 4.570 ;
        RECT 33.150 3.570 33.380 4.140 ;
        RECT 35.940 3.570 36.170 4.250 ;
        RECT 40.860 4.140 41.200 4.470 ;
        RECT 41.760 4.440 42.210 4.820 ;
        RECT 44.690 4.640 46.070 5.120 ;
        RECT 46.450 4.630 47.830 5.110 ;
        RECT 43.610 4.250 43.940 4.570 ;
        RECT 48.570 4.470 48.800 4.570 ;
        RECT 40.860 3.570 41.090 4.140 ;
        RECT 43.650 3.570 43.880 4.250 ;
        RECT 48.570 4.140 48.910 4.470 ;
        RECT 49.470 4.440 49.920 4.820 ;
        RECT 52.400 4.640 53.780 5.120 ;
        RECT 54.160 4.630 55.540 5.110 ;
        RECT 51.320 4.250 51.650 4.570 ;
        RECT 56.280 4.470 56.510 4.570 ;
        RECT 48.570 3.570 48.800 4.140 ;
        RECT 51.360 3.570 51.590 4.250 ;
        RECT 56.280 4.140 56.620 4.470 ;
        RECT 57.180 4.440 57.630 4.820 ;
        RECT 60.110 4.640 61.490 5.120 ;
        RECT 61.870 4.630 63.250 5.110 ;
        RECT 59.030 4.250 59.360 4.570 ;
        RECT 63.990 4.470 64.220 4.570 ;
        RECT 56.280 3.570 56.510 4.140 ;
        RECT 59.070 3.570 59.300 4.250 ;
        RECT 63.990 4.140 64.330 4.470 ;
        RECT 64.890 4.440 65.340 4.820 ;
        RECT 67.820 4.640 69.200 5.120 ;
        RECT 69.580 4.630 70.960 5.110 ;
        RECT 66.740 4.250 67.070 4.570 ;
        RECT 71.700 4.470 71.930 4.570 ;
        RECT 63.990 3.570 64.220 4.140 ;
        RECT 66.780 3.570 67.010 4.250 ;
        RECT 71.700 4.140 72.040 4.470 ;
        RECT 72.600 4.440 73.050 4.820 ;
        RECT 75.530 4.640 76.910 5.120 ;
        RECT 77.290 4.630 78.670 5.110 ;
        RECT 74.450 4.250 74.780 4.570 ;
        RECT 79.410 4.470 79.640 4.570 ;
        RECT 71.700 3.570 71.930 4.140 ;
        RECT 74.490 3.570 74.720 4.250 ;
        RECT 79.410 4.140 79.750 4.470 ;
        RECT 80.310 4.440 80.760 4.820 ;
        RECT 83.240 4.640 84.620 5.120 ;
        RECT 85.000 4.630 86.380 5.110 ;
        RECT 82.160 4.250 82.490 4.570 ;
        RECT 87.120 4.470 87.350 4.570 ;
        RECT 79.410 3.570 79.640 4.140 ;
        RECT 82.200 3.570 82.430 4.250 ;
        RECT 87.120 4.140 87.460 4.470 ;
        RECT 88.020 4.440 88.470 4.820 ;
        RECT 90.950 4.640 92.330 5.120 ;
        RECT 92.710 4.630 94.090 5.110 ;
        RECT 89.870 4.250 90.200 4.570 ;
        RECT 94.830 4.470 95.060 4.570 ;
        RECT 87.120 3.570 87.350 4.140 ;
        RECT 89.910 3.570 90.140 4.250 ;
        RECT 94.830 4.140 95.170 4.470 ;
        RECT 95.730 4.440 96.180 4.820 ;
        RECT 98.660 4.640 100.040 5.120 ;
        RECT 100.420 4.630 101.800 5.110 ;
        RECT 97.580 4.250 97.910 4.570 ;
        RECT 102.540 4.470 102.770 4.570 ;
        RECT 94.830 3.570 95.060 4.140 ;
        RECT 97.620 3.570 97.850 4.250 ;
        RECT 102.540 4.140 102.880 4.470 ;
        RECT 103.440 4.440 103.890 4.820 ;
        RECT 106.370 4.640 107.750 5.120 ;
        RECT 108.130 4.630 109.510 5.110 ;
        RECT 105.290 4.250 105.620 4.570 ;
        RECT 110.250 4.470 110.480 4.570 ;
        RECT 102.540 3.570 102.770 4.140 ;
        RECT 105.330 3.570 105.560 4.250 ;
        RECT 110.250 4.140 110.590 4.470 ;
        RECT 111.150 4.440 111.600 4.820 ;
        RECT 114.080 4.640 115.460 5.120 ;
        RECT 115.840 4.630 117.220 5.110 ;
        RECT 113.000 4.250 113.330 4.570 ;
        RECT 117.960 4.470 118.190 4.570 ;
        RECT 110.250 3.570 110.480 4.140 ;
        RECT 113.040 3.570 113.270 4.250 ;
        RECT 117.960 4.140 118.300 4.470 ;
        RECT 118.860 4.440 119.310 4.820 ;
        RECT 121.790 4.640 123.170 5.120 ;
        RECT 120.710 4.250 121.040 4.570 ;
        RECT 117.960 3.570 118.190 4.140 ;
        RECT 120.750 3.570 120.980 4.250 ;
      LAYER via ;
        RECT 2.030 28.920 2.290 29.180 ;
        RECT 4.780 29.020 5.040 29.280 ;
        RECT 0.840 28.470 1.100 28.750 ;
        RECT 9.740 28.920 10.000 29.180 ;
        RECT 12.490 29.020 12.750 29.280 ;
        RECT 6.010 28.450 6.270 28.710 ;
        RECT 8.550 28.470 8.810 28.750 ;
        RECT 17.450 28.920 17.710 29.180 ;
        RECT 20.200 29.020 20.460 29.280 ;
        RECT 13.720 28.450 13.980 28.710 ;
        RECT 16.260 28.470 16.520 28.750 ;
        RECT 25.160 28.920 25.420 29.180 ;
        RECT 27.910 29.020 28.170 29.280 ;
        RECT 21.430 28.450 21.690 28.710 ;
        RECT 23.970 28.470 24.230 28.750 ;
        RECT 32.870 28.920 33.130 29.180 ;
        RECT 35.620 29.020 35.880 29.280 ;
        RECT 29.140 28.450 29.400 28.710 ;
        RECT 31.680 28.470 31.940 28.750 ;
        RECT 40.580 28.920 40.840 29.180 ;
        RECT 43.330 29.020 43.590 29.280 ;
        RECT 36.850 28.450 37.110 28.710 ;
        RECT 39.390 28.470 39.650 28.750 ;
        RECT 48.290 28.920 48.550 29.180 ;
        RECT 51.040 29.020 51.300 29.280 ;
        RECT 44.560 28.450 44.820 28.710 ;
        RECT 47.100 28.470 47.360 28.750 ;
        RECT 56.000 28.920 56.260 29.180 ;
        RECT 58.750 29.020 59.010 29.280 ;
        RECT 52.270 28.450 52.530 28.710 ;
        RECT 54.810 28.470 55.070 28.750 ;
        RECT 63.710 28.920 63.970 29.180 ;
        RECT 66.460 29.020 66.720 29.280 ;
        RECT 59.980 28.450 60.240 28.710 ;
        RECT 62.520 28.470 62.780 28.750 ;
        RECT 71.420 28.920 71.680 29.180 ;
        RECT 74.170 29.020 74.430 29.280 ;
        RECT 67.690 28.450 67.950 28.710 ;
        RECT 70.230 28.470 70.490 28.750 ;
        RECT 79.130 28.920 79.390 29.180 ;
        RECT 81.880 29.020 82.140 29.280 ;
        RECT 75.400 28.450 75.660 28.710 ;
        RECT 77.940 28.470 78.200 28.750 ;
        RECT 86.840 28.920 87.100 29.180 ;
        RECT 89.590 29.020 89.850 29.280 ;
        RECT 83.110 28.450 83.370 28.710 ;
        RECT 85.650 28.470 85.910 28.750 ;
        RECT 94.550 28.920 94.810 29.180 ;
        RECT 97.300 29.020 97.560 29.280 ;
        RECT 90.820 28.450 91.080 28.710 ;
        RECT 93.360 28.470 93.620 28.750 ;
        RECT 102.260 28.920 102.520 29.180 ;
        RECT 105.010 29.020 105.270 29.280 ;
        RECT 98.530 28.450 98.790 28.710 ;
        RECT 101.070 28.470 101.330 28.750 ;
        RECT 109.970 28.920 110.230 29.180 ;
        RECT 112.720 29.020 112.980 29.280 ;
        RECT 106.240 28.450 106.500 28.710 ;
        RECT 108.780 28.470 109.040 28.750 ;
        RECT 117.680 28.920 117.940 29.180 ;
        RECT 120.430 29.020 120.690 29.280 ;
        RECT 113.950 28.450 114.210 28.710 ;
        RECT 116.490 28.470 116.750 28.750 ;
        RECT 121.660 28.450 121.920 28.710 ;
        RECT 1.120 4.750 1.380 5.010 ;
        RECT 6.290 4.710 6.550 4.990 ;
        RECT 8.830 4.750 9.090 5.010 ;
        RECT 2.350 4.180 2.610 4.440 ;
        RECT 5.100 4.280 5.360 4.540 ;
        RECT 14.000 4.710 14.260 4.990 ;
        RECT 16.540 4.750 16.800 5.010 ;
        RECT 10.060 4.180 10.320 4.440 ;
        RECT 12.810 4.280 13.070 4.540 ;
        RECT 21.710 4.710 21.970 4.990 ;
        RECT 24.250 4.750 24.510 5.010 ;
        RECT 17.770 4.180 18.030 4.440 ;
        RECT 20.520 4.280 20.780 4.540 ;
        RECT 29.420 4.710 29.680 4.990 ;
        RECT 31.960 4.750 32.220 5.010 ;
        RECT 25.480 4.180 25.740 4.440 ;
        RECT 28.230 4.280 28.490 4.540 ;
        RECT 37.130 4.710 37.390 4.990 ;
        RECT 39.670 4.750 39.930 5.010 ;
        RECT 33.190 4.180 33.450 4.440 ;
        RECT 35.940 4.280 36.200 4.540 ;
        RECT 44.840 4.710 45.100 4.990 ;
        RECT 47.380 4.750 47.640 5.010 ;
        RECT 40.900 4.180 41.160 4.440 ;
        RECT 43.650 4.280 43.910 4.540 ;
        RECT 52.550 4.710 52.810 4.990 ;
        RECT 55.090 4.750 55.350 5.010 ;
        RECT 48.610 4.180 48.870 4.440 ;
        RECT 51.360 4.280 51.620 4.540 ;
        RECT 60.260 4.710 60.520 4.990 ;
        RECT 62.800 4.750 63.060 5.010 ;
        RECT 56.320 4.180 56.580 4.440 ;
        RECT 59.070 4.280 59.330 4.540 ;
        RECT 67.970 4.710 68.230 4.990 ;
        RECT 70.510 4.750 70.770 5.010 ;
        RECT 64.030 4.180 64.290 4.440 ;
        RECT 66.780 4.280 67.040 4.540 ;
        RECT 75.680 4.710 75.940 4.990 ;
        RECT 78.220 4.750 78.480 5.010 ;
        RECT 71.740 4.180 72.000 4.440 ;
        RECT 74.490 4.280 74.750 4.540 ;
        RECT 83.390 4.710 83.650 4.990 ;
        RECT 85.930 4.750 86.190 5.010 ;
        RECT 79.450 4.180 79.710 4.440 ;
        RECT 82.200 4.280 82.460 4.540 ;
        RECT 91.100 4.710 91.360 4.990 ;
        RECT 93.640 4.750 93.900 5.010 ;
        RECT 87.160 4.180 87.420 4.440 ;
        RECT 89.910 4.280 90.170 4.540 ;
        RECT 98.810 4.710 99.070 4.990 ;
        RECT 101.350 4.750 101.610 5.010 ;
        RECT 94.870 4.180 95.130 4.440 ;
        RECT 97.620 4.280 97.880 4.540 ;
        RECT 106.520 4.710 106.780 4.990 ;
        RECT 109.060 4.750 109.320 5.010 ;
        RECT 102.580 4.180 102.840 4.440 ;
        RECT 105.330 4.280 105.590 4.540 ;
        RECT 114.230 4.710 114.490 4.990 ;
        RECT 116.770 4.750 117.030 5.010 ;
        RECT 110.290 4.180 110.550 4.440 ;
        RECT 113.040 4.280 113.300 4.540 ;
        RECT 121.940 4.710 122.200 4.990 ;
        RECT 118.000 4.180 118.260 4.440 ;
        RECT 120.750 4.280 121.010 4.540 ;
      LAYER met2 ;
        RECT 0.990 29.070 2.330 29.210 ;
        RECT 0.990 28.780 1.130 29.070 ;
        RECT 2.000 28.890 2.330 29.070 ;
        RECT 4.740 29.110 5.070 29.320 ;
        RECT 4.740 28.990 6.150 29.110 ;
        RECT 4.930 28.970 6.150 28.990 ;
        RECT 0.810 28.440 1.130 28.780 ;
        RECT 6.010 28.740 6.150 28.970 ;
        RECT 8.700 29.070 10.040 29.210 ;
        RECT 8.700 28.780 8.840 29.070 ;
        RECT 9.710 28.890 10.040 29.070 ;
        RECT 12.450 29.110 12.780 29.320 ;
        RECT 12.450 28.990 13.860 29.110 ;
        RECT 12.640 28.970 13.860 28.990 ;
        RECT 6.010 28.420 6.320 28.740 ;
        RECT 8.520 28.440 8.840 28.780 ;
        RECT 13.720 28.740 13.860 28.970 ;
        RECT 16.410 29.070 17.750 29.210 ;
        RECT 16.410 28.780 16.550 29.070 ;
        RECT 17.420 28.890 17.750 29.070 ;
        RECT 20.160 29.110 20.490 29.320 ;
        RECT 20.160 28.990 21.570 29.110 ;
        RECT 20.350 28.970 21.570 28.990 ;
        RECT 13.720 28.420 14.030 28.740 ;
        RECT 16.230 28.440 16.550 28.780 ;
        RECT 21.430 28.740 21.570 28.970 ;
        RECT 24.120 29.070 25.460 29.210 ;
        RECT 24.120 28.780 24.260 29.070 ;
        RECT 25.130 28.890 25.460 29.070 ;
        RECT 27.870 29.110 28.200 29.320 ;
        RECT 27.870 28.990 29.280 29.110 ;
        RECT 28.060 28.970 29.280 28.990 ;
        RECT 21.430 28.420 21.740 28.740 ;
        RECT 23.940 28.440 24.260 28.780 ;
        RECT 29.140 28.740 29.280 28.970 ;
        RECT 31.830 29.070 33.170 29.210 ;
        RECT 31.830 28.780 31.970 29.070 ;
        RECT 32.840 28.890 33.170 29.070 ;
        RECT 35.580 29.110 35.910 29.320 ;
        RECT 35.580 28.990 36.990 29.110 ;
        RECT 35.770 28.970 36.990 28.990 ;
        RECT 29.140 28.420 29.450 28.740 ;
        RECT 31.650 28.440 31.970 28.780 ;
        RECT 36.850 28.740 36.990 28.970 ;
        RECT 39.540 29.070 40.880 29.210 ;
        RECT 39.540 28.780 39.680 29.070 ;
        RECT 40.550 28.890 40.880 29.070 ;
        RECT 43.290 29.110 43.620 29.320 ;
        RECT 43.290 28.990 44.700 29.110 ;
        RECT 43.480 28.970 44.700 28.990 ;
        RECT 36.850 28.420 37.160 28.740 ;
        RECT 39.360 28.440 39.680 28.780 ;
        RECT 44.560 28.740 44.700 28.970 ;
        RECT 47.250 29.070 48.590 29.210 ;
        RECT 47.250 28.780 47.390 29.070 ;
        RECT 48.260 28.890 48.590 29.070 ;
        RECT 51.000 29.110 51.330 29.320 ;
        RECT 51.000 28.990 52.410 29.110 ;
        RECT 51.190 28.970 52.410 28.990 ;
        RECT 44.560 28.420 44.870 28.740 ;
        RECT 47.070 28.440 47.390 28.780 ;
        RECT 52.270 28.740 52.410 28.970 ;
        RECT 54.960 29.070 56.300 29.210 ;
        RECT 54.960 28.780 55.100 29.070 ;
        RECT 55.970 28.890 56.300 29.070 ;
        RECT 58.710 29.110 59.040 29.320 ;
        RECT 58.710 28.990 60.120 29.110 ;
        RECT 58.900 28.970 60.120 28.990 ;
        RECT 52.270 28.420 52.580 28.740 ;
        RECT 54.780 28.440 55.100 28.780 ;
        RECT 59.980 28.740 60.120 28.970 ;
        RECT 62.670 29.070 64.010 29.210 ;
        RECT 62.670 28.780 62.810 29.070 ;
        RECT 63.680 28.890 64.010 29.070 ;
        RECT 66.420 29.110 66.750 29.320 ;
        RECT 66.420 28.990 67.830 29.110 ;
        RECT 66.610 28.970 67.830 28.990 ;
        RECT 59.980 28.420 60.290 28.740 ;
        RECT 62.490 28.440 62.810 28.780 ;
        RECT 67.690 28.740 67.830 28.970 ;
        RECT 70.380 29.070 71.720 29.210 ;
        RECT 70.380 28.780 70.520 29.070 ;
        RECT 71.390 28.890 71.720 29.070 ;
        RECT 74.130 29.110 74.460 29.320 ;
        RECT 74.130 28.990 75.540 29.110 ;
        RECT 74.320 28.970 75.540 28.990 ;
        RECT 67.690 28.420 68.000 28.740 ;
        RECT 70.200 28.440 70.520 28.780 ;
        RECT 75.400 28.740 75.540 28.970 ;
        RECT 78.090 29.070 79.430 29.210 ;
        RECT 78.090 28.780 78.230 29.070 ;
        RECT 79.100 28.890 79.430 29.070 ;
        RECT 81.840 29.110 82.170 29.320 ;
        RECT 81.840 28.990 83.250 29.110 ;
        RECT 82.030 28.970 83.250 28.990 ;
        RECT 75.400 28.420 75.710 28.740 ;
        RECT 77.910 28.440 78.230 28.780 ;
        RECT 83.110 28.740 83.250 28.970 ;
        RECT 85.800 29.070 87.140 29.210 ;
        RECT 85.800 28.780 85.940 29.070 ;
        RECT 86.810 28.890 87.140 29.070 ;
        RECT 89.550 29.110 89.880 29.320 ;
        RECT 89.550 28.990 90.960 29.110 ;
        RECT 89.740 28.970 90.960 28.990 ;
        RECT 83.110 28.420 83.420 28.740 ;
        RECT 85.620 28.440 85.940 28.780 ;
        RECT 90.820 28.740 90.960 28.970 ;
        RECT 93.510 29.070 94.850 29.210 ;
        RECT 93.510 28.780 93.650 29.070 ;
        RECT 94.520 28.890 94.850 29.070 ;
        RECT 97.260 29.110 97.590 29.320 ;
        RECT 97.260 28.990 98.670 29.110 ;
        RECT 97.450 28.970 98.670 28.990 ;
        RECT 90.820 28.420 91.130 28.740 ;
        RECT 93.330 28.440 93.650 28.780 ;
        RECT 98.530 28.740 98.670 28.970 ;
        RECT 101.220 29.070 102.560 29.210 ;
        RECT 101.220 28.780 101.360 29.070 ;
        RECT 102.230 28.890 102.560 29.070 ;
        RECT 104.970 29.110 105.300 29.320 ;
        RECT 104.970 28.990 106.380 29.110 ;
        RECT 105.160 28.970 106.380 28.990 ;
        RECT 98.530 28.420 98.840 28.740 ;
        RECT 101.040 28.440 101.360 28.780 ;
        RECT 106.240 28.740 106.380 28.970 ;
        RECT 108.930 29.070 110.270 29.210 ;
        RECT 108.930 28.780 109.070 29.070 ;
        RECT 109.940 28.890 110.270 29.070 ;
        RECT 112.680 29.110 113.010 29.320 ;
        RECT 112.680 28.990 114.090 29.110 ;
        RECT 112.870 28.970 114.090 28.990 ;
        RECT 106.240 28.420 106.550 28.740 ;
        RECT 108.750 28.440 109.070 28.780 ;
        RECT 113.950 28.740 114.090 28.970 ;
        RECT 116.640 29.070 117.980 29.210 ;
        RECT 116.640 28.780 116.780 29.070 ;
        RECT 117.650 28.890 117.980 29.070 ;
        RECT 120.390 29.110 120.720 29.320 ;
        RECT 120.390 28.990 121.800 29.110 ;
        RECT 120.580 28.970 121.800 28.990 ;
        RECT 113.950 28.420 114.260 28.740 ;
        RECT 116.460 28.440 116.780 28.780 ;
        RECT 121.660 28.740 121.800 28.970 ;
        RECT 121.660 28.420 121.970 28.740 ;
        RECT 1.070 4.720 1.380 5.040 ;
        RECT 1.240 4.490 1.380 4.720 ;
        RECT 6.260 4.680 6.580 5.020 ;
        RECT 8.780 4.720 9.090 5.040 ;
        RECT 1.240 4.470 2.460 4.490 ;
        RECT 1.240 4.350 2.650 4.470 ;
        RECT 2.320 4.140 2.650 4.350 ;
        RECT 5.060 4.390 5.390 4.570 ;
        RECT 6.260 4.390 6.400 4.680 ;
        RECT 5.060 4.250 6.400 4.390 ;
        RECT 8.950 4.490 9.090 4.720 ;
        RECT 13.970 4.680 14.290 5.020 ;
        RECT 16.490 4.720 16.800 5.040 ;
        RECT 8.950 4.470 10.170 4.490 ;
        RECT 8.950 4.350 10.360 4.470 ;
        RECT 10.030 4.140 10.360 4.350 ;
        RECT 12.770 4.390 13.100 4.570 ;
        RECT 13.970 4.390 14.110 4.680 ;
        RECT 12.770 4.250 14.110 4.390 ;
        RECT 16.660 4.490 16.800 4.720 ;
        RECT 21.680 4.680 22.000 5.020 ;
        RECT 24.200 4.720 24.510 5.040 ;
        RECT 16.660 4.470 17.880 4.490 ;
        RECT 16.660 4.350 18.070 4.470 ;
        RECT 17.740 4.140 18.070 4.350 ;
        RECT 20.480 4.390 20.810 4.570 ;
        RECT 21.680 4.390 21.820 4.680 ;
        RECT 20.480 4.250 21.820 4.390 ;
        RECT 24.370 4.490 24.510 4.720 ;
        RECT 29.390 4.680 29.710 5.020 ;
        RECT 31.910 4.720 32.220 5.040 ;
        RECT 24.370 4.470 25.590 4.490 ;
        RECT 24.370 4.350 25.780 4.470 ;
        RECT 25.450 4.140 25.780 4.350 ;
        RECT 28.190 4.390 28.520 4.570 ;
        RECT 29.390 4.390 29.530 4.680 ;
        RECT 28.190 4.250 29.530 4.390 ;
        RECT 32.080 4.490 32.220 4.720 ;
        RECT 37.100 4.680 37.420 5.020 ;
        RECT 39.620 4.720 39.930 5.040 ;
        RECT 32.080 4.470 33.300 4.490 ;
        RECT 32.080 4.350 33.490 4.470 ;
        RECT 33.160 4.140 33.490 4.350 ;
        RECT 35.900 4.390 36.230 4.570 ;
        RECT 37.100 4.390 37.240 4.680 ;
        RECT 35.900 4.250 37.240 4.390 ;
        RECT 39.790 4.490 39.930 4.720 ;
        RECT 44.810 4.680 45.130 5.020 ;
        RECT 47.330 4.720 47.640 5.040 ;
        RECT 39.790 4.470 41.010 4.490 ;
        RECT 39.790 4.350 41.200 4.470 ;
        RECT 40.870 4.140 41.200 4.350 ;
        RECT 43.610 4.390 43.940 4.570 ;
        RECT 44.810 4.390 44.950 4.680 ;
        RECT 43.610 4.250 44.950 4.390 ;
        RECT 47.500 4.490 47.640 4.720 ;
        RECT 52.520 4.680 52.840 5.020 ;
        RECT 55.040 4.720 55.350 5.040 ;
        RECT 47.500 4.470 48.720 4.490 ;
        RECT 47.500 4.350 48.910 4.470 ;
        RECT 48.580 4.140 48.910 4.350 ;
        RECT 51.320 4.390 51.650 4.570 ;
        RECT 52.520 4.390 52.660 4.680 ;
        RECT 51.320 4.250 52.660 4.390 ;
        RECT 55.210 4.490 55.350 4.720 ;
        RECT 60.230 4.680 60.550 5.020 ;
        RECT 62.750 4.720 63.060 5.040 ;
        RECT 55.210 4.470 56.430 4.490 ;
        RECT 55.210 4.350 56.620 4.470 ;
        RECT 56.290 4.140 56.620 4.350 ;
        RECT 59.030 4.390 59.360 4.570 ;
        RECT 60.230 4.390 60.370 4.680 ;
        RECT 59.030 4.250 60.370 4.390 ;
        RECT 62.920 4.490 63.060 4.720 ;
        RECT 67.940 4.680 68.260 5.020 ;
        RECT 70.460 4.720 70.770 5.040 ;
        RECT 62.920 4.470 64.140 4.490 ;
        RECT 62.920 4.350 64.330 4.470 ;
        RECT 64.000 4.140 64.330 4.350 ;
        RECT 66.740 4.390 67.070 4.570 ;
        RECT 67.940 4.390 68.080 4.680 ;
        RECT 66.740 4.250 68.080 4.390 ;
        RECT 70.630 4.490 70.770 4.720 ;
        RECT 75.650 4.680 75.970 5.020 ;
        RECT 78.170 4.720 78.480 5.040 ;
        RECT 70.630 4.470 71.850 4.490 ;
        RECT 70.630 4.350 72.040 4.470 ;
        RECT 71.710 4.140 72.040 4.350 ;
        RECT 74.450 4.390 74.780 4.570 ;
        RECT 75.650 4.390 75.790 4.680 ;
        RECT 74.450 4.250 75.790 4.390 ;
        RECT 78.340 4.490 78.480 4.720 ;
        RECT 83.360 4.680 83.680 5.020 ;
        RECT 85.880 4.720 86.190 5.040 ;
        RECT 78.340 4.470 79.560 4.490 ;
        RECT 78.340 4.350 79.750 4.470 ;
        RECT 79.420 4.140 79.750 4.350 ;
        RECT 82.160 4.390 82.490 4.570 ;
        RECT 83.360 4.390 83.500 4.680 ;
        RECT 82.160 4.250 83.500 4.390 ;
        RECT 86.050 4.490 86.190 4.720 ;
        RECT 91.070 4.680 91.390 5.020 ;
        RECT 93.590 4.720 93.900 5.040 ;
        RECT 86.050 4.470 87.270 4.490 ;
        RECT 86.050 4.350 87.460 4.470 ;
        RECT 87.130 4.140 87.460 4.350 ;
        RECT 89.870 4.390 90.200 4.570 ;
        RECT 91.070 4.390 91.210 4.680 ;
        RECT 89.870 4.250 91.210 4.390 ;
        RECT 93.760 4.490 93.900 4.720 ;
        RECT 98.780 4.680 99.100 5.020 ;
        RECT 101.300 4.720 101.610 5.040 ;
        RECT 93.760 4.470 94.980 4.490 ;
        RECT 93.760 4.350 95.170 4.470 ;
        RECT 94.840 4.140 95.170 4.350 ;
        RECT 97.580 4.390 97.910 4.570 ;
        RECT 98.780 4.390 98.920 4.680 ;
        RECT 97.580 4.250 98.920 4.390 ;
        RECT 101.470 4.490 101.610 4.720 ;
        RECT 106.490 4.680 106.810 5.020 ;
        RECT 109.010 4.720 109.320 5.040 ;
        RECT 101.470 4.470 102.690 4.490 ;
        RECT 101.470 4.350 102.880 4.470 ;
        RECT 102.550 4.140 102.880 4.350 ;
        RECT 105.290 4.390 105.620 4.570 ;
        RECT 106.490 4.390 106.630 4.680 ;
        RECT 105.290 4.250 106.630 4.390 ;
        RECT 109.180 4.490 109.320 4.720 ;
        RECT 114.200 4.680 114.520 5.020 ;
        RECT 116.720 4.720 117.030 5.040 ;
        RECT 109.180 4.470 110.400 4.490 ;
        RECT 109.180 4.350 110.590 4.470 ;
        RECT 110.260 4.140 110.590 4.350 ;
        RECT 113.000 4.390 113.330 4.570 ;
        RECT 114.200 4.390 114.340 4.680 ;
        RECT 113.000 4.250 114.340 4.390 ;
        RECT 116.890 4.490 117.030 4.720 ;
        RECT 121.910 4.680 122.230 5.020 ;
        RECT 116.890 4.470 118.110 4.490 ;
        RECT 116.890 4.350 118.300 4.470 ;
        RECT 117.970 4.140 118.300 4.350 ;
        RECT 120.710 4.390 121.040 4.570 ;
        RECT 121.910 4.390 122.050 4.680 ;
        RECT 120.710 4.250 122.050 4.390 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 53.765900 ;
    PORT
      LAYER pwell ;
        RECT 3.000 31.660 4.660 33.460 ;
        RECT 10.710 31.660 12.370 33.460 ;
        RECT 18.420 31.660 20.080 33.460 ;
        RECT 26.130 31.660 27.790 33.460 ;
        RECT 33.840 31.660 35.500 33.460 ;
        RECT 41.550 31.660 43.210 33.460 ;
        RECT 49.260 31.660 50.920 33.460 ;
        RECT 56.970 31.660 58.630 33.460 ;
        RECT 64.680 31.660 66.340 33.460 ;
        RECT 72.390 31.660 74.050 33.460 ;
        RECT 80.100 31.660 81.760 33.460 ;
        RECT 87.810 31.660 89.470 33.460 ;
        RECT 95.520 31.660 97.180 33.460 ;
        RECT 103.230 31.660 104.890 33.460 ;
        RECT 110.940 31.660 112.600 33.460 ;
        RECT 118.650 31.660 120.310 33.460 ;
        RECT 2.990 26.380 4.650 28.180 ;
        RECT 10.700 26.380 12.360 28.180 ;
        RECT 18.410 26.380 20.070 28.180 ;
        RECT 26.120 26.380 27.780 28.180 ;
        RECT 33.830 26.380 35.490 28.180 ;
        RECT 41.540 26.380 43.200 28.180 ;
        RECT 49.250 26.380 50.910 28.180 ;
        RECT 56.960 26.380 58.620 28.180 ;
        RECT 64.670 26.380 66.330 28.180 ;
        RECT 72.380 26.380 74.040 28.180 ;
        RECT 80.090 26.380 81.750 28.180 ;
        RECT 87.800 26.380 89.460 28.180 ;
        RECT 95.510 26.380 97.170 28.180 ;
        RECT 103.220 26.380 104.880 28.180 ;
        RECT 110.930 26.380 112.590 28.180 ;
        RECT 118.640 26.380 120.300 28.180 ;
        RECT 22.270 21.815 23.180 22.805 ;
        RECT 22.270 20.905 29.500 21.815 ;
        RECT 2.740 5.280 4.400 7.080 ;
        RECT 10.450 5.280 12.110 7.080 ;
        RECT 18.160 5.280 19.820 7.080 ;
        RECT 25.870 5.280 27.530 7.080 ;
        RECT 33.580 5.280 35.240 7.080 ;
        RECT 41.290 5.280 42.950 7.080 ;
        RECT 49.000 5.280 50.660 7.080 ;
        RECT 56.710 5.280 58.370 7.080 ;
        RECT 64.420 5.280 66.080 7.080 ;
        RECT 72.130 5.280 73.790 7.080 ;
        RECT 79.840 5.280 81.500 7.080 ;
        RECT 87.550 5.280 89.210 7.080 ;
        RECT 95.260 5.280 96.920 7.080 ;
        RECT 102.970 5.280 104.630 7.080 ;
        RECT 110.680 5.280 112.340 7.080 ;
        RECT 118.390 5.280 120.050 7.080 ;
        RECT 2.730 0.000 4.390 1.800 ;
        RECT 10.440 0.000 12.100 1.800 ;
        RECT 18.150 0.000 19.810 1.800 ;
        RECT 25.860 0.000 27.520 1.800 ;
        RECT 33.570 0.000 35.230 1.800 ;
        RECT 41.280 0.000 42.940 1.800 ;
        RECT 48.990 0.000 50.650 1.800 ;
        RECT 56.700 0.000 58.360 1.800 ;
        RECT 64.410 0.000 66.070 1.800 ;
        RECT 72.120 0.000 73.780 1.800 ;
        RECT 79.830 0.000 81.490 1.800 ;
        RECT 87.540 0.000 89.200 1.800 ;
        RECT 95.250 0.000 96.910 1.800 ;
        RECT 102.960 0.000 104.620 1.800 ;
        RECT 110.670 0.000 112.330 1.800 ;
        RECT 118.380 0.000 120.040 1.800 ;
      LAYER li1 ;
        RECT 3.220 33.170 4.570 33.340 ;
        RECT 10.930 33.170 12.280 33.340 ;
        RECT 18.640 33.170 19.990 33.340 ;
        RECT 26.350 33.170 27.700 33.340 ;
        RECT 34.060 33.170 35.410 33.340 ;
        RECT 41.770 33.170 43.120 33.340 ;
        RECT 49.480 33.170 50.830 33.340 ;
        RECT 57.190 33.170 58.540 33.340 ;
        RECT 64.900 33.170 66.250 33.340 ;
        RECT 72.610 33.170 73.960 33.340 ;
        RECT 80.320 33.170 81.670 33.340 ;
        RECT 88.030 33.170 89.380 33.340 ;
        RECT 95.740 33.170 97.090 33.340 ;
        RECT 103.450 33.170 104.800 33.340 ;
        RECT 111.160 33.170 112.510 33.340 ;
        RECT 118.870 33.170 120.220 33.340 ;
        RECT 1.475 32.960 4.570 33.170 ;
        RECT 1.475 31.425 1.685 32.960 ;
        RECT 3.220 32.950 4.570 32.960 ;
        RECT 9.185 32.960 12.280 33.170 ;
        RECT 9.185 31.425 9.395 32.960 ;
        RECT 10.930 32.950 12.280 32.960 ;
        RECT 16.895 32.960 19.990 33.170 ;
        RECT 16.895 31.425 17.105 32.960 ;
        RECT 18.640 32.950 19.990 32.960 ;
        RECT 24.605 32.960 27.700 33.170 ;
        RECT 24.605 31.425 24.815 32.960 ;
        RECT 26.350 32.950 27.700 32.960 ;
        RECT 32.315 32.960 35.410 33.170 ;
        RECT 32.315 31.425 32.525 32.960 ;
        RECT 34.060 32.950 35.410 32.960 ;
        RECT 40.025 32.960 43.120 33.170 ;
        RECT 40.025 31.425 40.235 32.960 ;
        RECT 41.770 32.950 43.120 32.960 ;
        RECT 47.735 32.960 50.830 33.170 ;
        RECT 47.735 31.425 47.945 32.960 ;
        RECT 49.480 32.950 50.830 32.960 ;
        RECT 55.445 32.960 58.540 33.170 ;
        RECT 55.445 31.425 55.655 32.960 ;
        RECT 57.190 32.950 58.540 32.960 ;
        RECT 63.155 32.960 66.250 33.170 ;
        RECT 63.155 31.425 63.365 32.960 ;
        RECT 64.900 32.950 66.250 32.960 ;
        RECT 70.865 32.960 73.960 33.170 ;
        RECT 70.865 31.425 71.075 32.960 ;
        RECT 72.610 32.950 73.960 32.960 ;
        RECT 78.575 32.960 81.670 33.170 ;
        RECT 78.575 31.425 78.785 32.960 ;
        RECT 80.320 32.950 81.670 32.960 ;
        RECT 86.285 32.960 89.380 33.170 ;
        RECT 86.285 31.425 86.495 32.960 ;
        RECT 88.030 32.950 89.380 32.960 ;
        RECT 93.995 32.960 97.090 33.170 ;
        RECT 93.995 31.425 94.205 32.960 ;
        RECT 95.740 32.950 97.090 32.960 ;
        RECT 101.705 32.960 104.800 33.170 ;
        RECT 101.705 31.425 101.915 32.960 ;
        RECT 103.450 32.950 104.800 32.960 ;
        RECT 109.415 32.960 112.510 33.170 ;
        RECT 109.415 31.425 109.625 32.960 ;
        RECT 111.160 32.950 112.510 32.960 ;
        RECT 117.125 32.960 120.220 33.170 ;
        RECT 117.125 31.425 117.335 32.960 ;
        RECT 118.870 32.950 120.220 32.960 ;
        RECT 0.965 31.385 1.685 31.425 ;
        RECT -0.130 31.215 1.685 31.385 ;
        RECT 5.820 31.225 7.200 31.395 ;
        RECT 8.675 31.385 9.395 31.425 ;
        RECT 0.700 30.395 0.930 31.215 ;
        RECT 6.650 30.405 6.880 31.225 ;
        RECT 7.580 31.215 9.395 31.385 ;
        RECT 13.530 31.225 14.910 31.395 ;
        RECT 16.385 31.385 17.105 31.425 ;
        RECT 8.410 30.395 8.640 31.215 ;
        RECT 14.360 30.405 14.590 31.225 ;
        RECT 15.290 31.215 17.105 31.385 ;
        RECT 21.240 31.225 22.620 31.395 ;
        RECT 24.095 31.385 24.815 31.425 ;
        RECT 16.120 30.395 16.350 31.215 ;
        RECT 22.070 30.405 22.300 31.225 ;
        RECT 23.000 31.215 24.815 31.385 ;
        RECT 28.950 31.225 30.330 31.395 ;
        RECT 31.805 31.385 32.525 31.425 ;
        RECT 23.830 30.395 24.060 31.215 ;
        RECT 29.780 30.405 30.010 31.225 ;
        RECT 30.710 31.215 32.525 31.385 ;
        RECT 36.660 31.225 38.040 31.395 ;
        RECT 39.515 31.385 40.235 31.425 ;
        RECT 31.540 30.395 31.770 31.215 ;
        RECT 37.490 30.405 37.720 31.225 ;
        RECT 38.420 31.215 40.235 31.385 ;
        RECT 44.370 31.225 45.750 31.395 ;
        RECT 47.225 31.385 47.945 31.425 ;
        RECT 39.250 30.395 39.480 31.215 ;
        RECT 45.200 30.405 45.430 31.225 ;
        RECT 46.130 31.215 47.945 31.385 ;
        RECT 52.080 31.225 53.460 31.395 ;
        RECT 54.935 31.385 55.655 31.425 ;
        RECT 46.960 30.395 47.190 31.215 ;
        RECT 52.910 30.405 53.140 31.225 ;
        RECT 53.840 31.215 55.655 31.385 ;
        RECT 59.790 31.225 61.170 31.395 ;
        RECT 62.645 31.385 63.365 31.425 ;
        RECT 54.670 30.395 54.900 31.215 ;
        RECT 60.620 30.405 60.850 31.225 ;
        RECT 61.550 31.215 63.365 31.385 ;
        RECT 67.500 31.225 68.880 31.395 ;
        RECT 70.355 31.385 71.075 31.425 ;
        RECT 62.380 30.395 62.610 31.215 ;
        RECT 68.330 30.405 68.560 31.225 ;
        RECT 69.260 31.215 71.075 31.385 ;
        RECT 75.210 31.225 76.590 31.395 ;
        RECT 78.065 31.385 78.785 31.425 ;
        RECT 70.090 30.395 70.320 31.215 ;
        RECT 76.040 30.405 76.270 31.225 ;
        RECT 76.970 31.215 78.785 31.385 ;
        RECT 82.920 31.225 84.300 31.395 ;
        RECT 85.775 31.385 86.495 31.425 ;
        RECT 77.800 30.395 78.030 31.215 ;
        RECT 83.750 30.405 83.980 31.225 ;
        RECT 84.680 31.215 86.495 31.385 ;
        RECT 90.630 31.225 92.010 31.395 ;
        RECT 93.485 31.385 94.205 31.425 ;
        RECT 85.510 30.395 85.740 31.215 ;
        RECT 91.460 30.405 91.690 31.225 ;
        RECT 92.390 31.215 94.205 31.385 ;
        RECT 98.340 31.225 99.720 31.395 ;
        RECT 101.195 31.385 101.915 31.425 ;
        RECT 93.220 30.395 93.450 31.215 ;
        RECT 99.170 30.405 99.400 31.225 ;
        RECT 100.100 31.215 101.915 31.385 ;
        RECT 106.050 31.225 107.430 31.395 ;
        RECT 108.905 31.385 109.625 31.425 ;
        RECT 100.930 30.395 101.160 31.215 ;
        RECT 106.880 30.405 107.110 31.225 ;
        RECT 107.810 31.215 109.625 31.385 ;
        RECT 113.760 31.225 115.140 31.395 ;
        RECT 116.615 31.385 117.335 31.425 ;
        RECT 108.640 30.395 108.870 31.215 ;
        RECT 114.590 30.405 114.820 31.225 ;
        RECT 115.520 31.215 117.335 31.385 ;
        RECT 121.470 31.225 122.850 31.395 ;
        RECT 116.350 30.395 116.580 31.215 ;
        RECT 122.300 30.405 122.530 31.225 ;
        RECT 2.120 28.060 2.350 28.090 ;
        RECT 9.830 28.060 10.060 28.090 ;
        RECT 17.540 28.060 17.770 28.090 ;
        RECT 25.250 28.060 25.480 28.090 ;
        RECT 32.960 28.060 33.190 28.090 ;
        RECT 40.670 28.060 40.900 28.090 ;
        RECT 48.380 28.060 48.610 28.090 ;
        RECT 56.090 28.060 56.320 28.090 ;
        RECT 63.800 28.060 64.030 28.090 ;
        RECT 71.510 28.060 71.740 28.090 ;
        RECT 79.220 28.060 79.450 28.090 ;
        RECT 86.930 28.060 87.160 28.090 ;
        RECT 94.640 28.060 94.870 28.090 ;
        RECT 102.350 28.060 102.580 28.090 ;
        RECT 110.060 28.060 110.290 28.090 ;
        RECT 117.770 28.060 118.000 28.090 ;
        RECT 2.120 27.890 4.560 28.060 ;
        RECT 2.120 27.870 2.350 27.890 ;
        RECT 3.210 27.840 4.560 27.890 ;
        RECT 9.830 27.890 12.270 28.060 ;
        RECT 9.830 27.870 10.060 27.890 ;
        RECT 10.920 27.840 12.270 27.890 ;
        RECT 17.540 27.890 19.980 28.060 ;
        RECT 17.540 27.870 17.770 27.890 ;
        RECT 18.630 27.840 19.980 27.890 ;
        RECT 25.250 27.890 27.690 28.060 ;
        RECT 25.250 27.870 25.480 27.890 ;
        RECT 26.340 27.840 27.690 27.890 ;
        RECT 32.960 27.890 35.400 28.060 ;
        RECT 32.960 27.870 33.190 27.890 ;
        RECT 34.050 27.840 35.400 27.890 ;
        RECT 40.670 27.890 43.110 28.060 ;
        RECT 40.670 27.870 40.900 27.890 ;
        RECT 41.760 27.840 43.110 27.890 ;
        RECT 48.380 27.890 50.820 28.060 ;
        RECT 48.380 27.870 48.610 27.890 ;
        RECT 49.470 27.840 50.820 27.890 ;
        RECT 56.090 27.890 58.530 28.060 ;
        RECT 56.090 27.870 56.320 27.890 ;
        RECT 57.180 27.840 58.530 27.890 ;
        RECT 63.800 27.890 66.240 28.060 ;
        RECT 63.800 27.870 64.030 27.890 ;
        RECT 64.890 27.840 66.240 27.890 ;
        RECT 71.510 27.890 73.950 28.060 ;
        RECT 71.510 27.870 71.740 27.890 ;
        RECT 72.600 27.840 73.950 27.890 ;
        RECT 79.220 27.890 81.660 28.060 ;
        RECT 79.220 27.870 79.450 27.890 ;
        RECT 80.310 27.840 81.660 27.890 ;
        RECT 86.930 27.890 89.370 28.060 ;
        RECT 86.930 27.870 87.160 27.890 ;
        RECT 88.020 27.840 89.370 27.890 ;
        RECT 94.640 27.890 97.080 28.060 ;
        RECT 94.640 27.870 94.870 27.890 ;
        RECT 95.730 27.840 97.080 27.890 ;
        RECT 102.350 27.890 104.790 28.060 ;
        RECT 102.350 27.870 102.580 27.890 ;
        RECT 103.440 27.840 104.790 27.890 ;
        RECT 110.060 27.890 112.500 28.060 ;
        RECT 110.060 27.870 110.290 27.890 ;
        RECT 111.150 27.840 112.500 27.890 ;
        RECT 117.770 27.890 120.210 28.060 ;
        RECT 117.770 27.870 118.000 27.890 ;
        RECT 118.860 27.840 120.210 27.890 ;
        RECT 3.210 27.670 5.060 27.840 ;
        RECT 10.920 27.670 12.770 27.840 ;
        RECT 18.630 27.670 20.480 27.840 ;
        RECT 26.340 27.670 28.190 27.840 ;
        RECT 34.050 27.670 35.900 27.840 ;
        RECT 41.760 27.670 43.610 27.840 ;
        RECT 49.470 27.670 51.320 27.840 ;
        RECT 57.180 27.670 59.030 27.840 ;
        RECT 64.890 27.670 66.740 27.840 ;
        RECT 72.600 27.670 74.450 27.840 ;
        RECT 80.310 27.670 82.160 27.840 ;
        RECT 88.020 27.670 89.870 27.840 ;
        RECT 95.730 27.670 97.580 27.840 ;
        RECT 103.440 27.670 105.290 27.840 ;
        RECT 111.150 27.670 113.000 27.840 ;
        RECT 118.860 27.670 120.710 27.840 ;
        RECT 4.890 26.155 5.060 27.670 ;
        RECT 6.170 26.155 6.340 27.380 ;
        RECT 12.600 26.155 12.770 27.670 ;
        RECT 13.880 26.155 14.050 27.380 ;
        RECT 20.310 26.155 20.480 27.670 ;
        RECT 21.590 26.155 21.760 27.380 ;
        RECT 28.020 26.155 28.190 27.670 ;
        RECT 29.300 26.155 29.470 27.380 ;
        RECT 35.730 26.155 35.900 27.670 ;
        RECT 37.010 26.155 37.180 27.380 ;
        RECT 43.440 26.155 43.610 27.670 ;
        RECT 44.720 26.155 44.890 27.380 ;
        RECT 51.150 26.155 51.320 27.670 ;
        RECT 52.430 26.155 52.600 27.380 ;
        RECT 58.860 26.155 59.030 27.670 ;
        RECT 60.140 26.155 60.310 27.380 ;
        RECT 0.890 25.985 2.270 26.155 ;
        RECT 4.890 25.985 6.340 26.155 ;
        RECT 8.600 25.985 9.980 26.155 ;
        RECT 12.600 25.985 14.050 26.155 ;
        RECT 16.310 25.985 17.690 26.155 ;
        RECT 20.310 25.985 21.760 26.155 ;
        RECT 24.020 25.985 25.400 26.155 ;
        RECT 28.020 25.985 29.470 26.155 ;
        RECT 31.730 25.985 33.110 26.155 ;
        RECT 35.730 25.985 37.180 26.155 ;
        RECT 39.440 25.985 40.820 26.155 ;
        RECT 43.440 25.985 44.890 26.155 ;
        RECT 47.150 25.985 48.530 26.155 ;
        RECT 51.150 25.985 52.600 26.155 ;
        RECT 54.860 25.985 56.240 26.155 ;
        RECT 58.860 25.985 60.310 26.155 ;
        RECT 61.370 26.180 61.710 26.210 ;
        RECT 61.370 26.155 62.820 26.180 ;
        RECT 66.570 26.155 66.740 27.670 ;
        RECT 67.850 26.155 68.020 27.380 ;
        RECT 74.280 26.155 74.450 27.670 ;
        RECT 75.560 26.155 75.730 27.380 ;
        RECT 81.990 26.155 82.160 27.670 ;
        RECT 83.270 26.155 83.440 27.380 ;
        RECT 89.700 26.155 89.870 27.670 ;
        RECT 90.980 26.155 91.150 27.380 ;
        RECT 61.370 25.985 63.950 26.155 ;
        RECT 66.570 25.985 68.020 26.155 ;
        RECT 70.280 25.985 71.660 26.155 ;
        RECT 74.280 25.985 75.730 26.155 ;
        RECT 77.990 25.985 79.370 26.155 ;
        RECT 81.990 25.985 83.440 26.155 ;
        RECT 85.700 25.985 87.080 26.155 ;
        RECT 89.700 25.985 91.150 26.155 ;
        RECT 92.325 26.155 93.755 26.275 ;
        RECT 97.410 26.155 97.580 27.670 ;
        RECT 98.690 26.155 98.860 27.380 ;
        RECT 105.120 26.155 105.290 27.670 ;
        RECT 106.400 26.155 106.570 27.380 ;
        RECT 112.830 26.155 113.000 27.670 ;
        RECT 114.110 26.155 114.280 27.380 ;
        RECT 120.540 26.155 120.710 27.670 ;
        RECT 121.820 26.155 121.990 27.380 ;
        RECT 92.325 25.985 94.790 26.155 ;
        RECT 97.410 25.985 98.860 26.155 ;
        RECT 101.120 25.985 102.500 26.155 ;
        RECT 105.120 25.985 106.570 26.155 ;
        RECT 108.830 25.985 110.210 26.155 ;
        RECT 112.830 25.985 114.280 26.155 ;
        RECT 116.540 25.985 117.920 26.155 ;
        RECT 120.540 25.985 121.990 26.155 ;
        RECT 0.985 25.175 1.255 25.985 ;
        RECT 1.925 25.175 2.165 25.985 ;
        RECT 4.890 25.980 5.325 25.985 ;
        RECT 5.055 25.175 5.325 25.980 ;
        RECT 5.995 25.175 6.235 25.985 ;
        RECT 8.695 25.175 8.965 25.985 ;
        RECT 9.635 25.175 9.875 25.985 ;
        RECT 12.600 25.980 13.035 25.985 ;
        RECT 12.765 25.175 13.035 25.980 ;
        RECT 13.705 25.175 13.945 25.985 ;
        RECT 16.405 25.175 16.675 25.985 ;
        RECT 17.345 25.175 17.585 25.985 ;
        RECT 20.310 25.980 20.745 25.985 ;
        RECT 20.475 25.175 20.745 25.980 ;
        RECT 21.415 25.175 21.655 25.985 ;
        RECT 24.115 25.175 24.385 25.985 ;
        RECT 25.055 25.175 25.295 25.985 ;
        RECT 28.020 25.980 28.455 25.985 ;
        RECT 28.185 25.175 28.455 25.980 ;
        RECT 29.125 25.175 29.365 25.985 ;
        RECT 31.825 25.175 32.095 25.985 ;
        RECT 32.765 25.175 33.005 25.985 ;
        RECT 35.730 25.980 36.165 25.985 ;
        RECT 35.895 25.175 36.165 25.980 ;
        RECT 36.835 25.175 37.075 25.985 ;
        RECT 39.535 25.175 39.805 25.985 ;
        RECT 40.475 25.175 40.715 25.985 ;
        RECT 43.440 25.980 43.875 25.985 ;
        RECT 43.605 25.175 43.875 25.980 ;
        RECT 44.545 25.175 44.785 25.985 ;
        RECT 47.245 25.175 47.515 25.985 ;
        RECT 48.185 25.175 48.425 25.985 ;
        RECT 51.150 25.980 51.585 25.985 ;
        RECT 51.315 25.175 51.585 25.980 ;
        RECT 52.255 25.175 52.495 25.985 ;
        RECT 54.955 25.175 55.225 25.985 ;
        RECT 55.895 25.175 56.135 25.985 ;
        RECT 58.860 25.980 59.295 25.985 ;
        RECT 59.025 25.175 59.295 25.980 ;
        RECT 59.965 25.175 60.205 25.985 ;
        RECT 61.370 25.840 62.935 25.985 ;
        RECT 61.370 22.790 61.710 25.840 ;
        RECT 62.665 25.175 62.935 25.840 ;
        RECT 63.605 25.175 63.845 25.985 ;
        RECT 66.570 25.980 67.005 25.985 ;
        RECT 66.735 25.175 67.005 25.980 ;
        RECT 67.675 25.175 67.915 25.985 ;
        RECT 70.375 25.175 70.645 25.985 ;
        RECT 71.315 25.175 71.555 25.985 ;
        RECT 74.280 25.980 74.715 25.985 ;
        RECT 74.445 25.175 74.715 25.980 ;
        RECT 75.385 25.175 75.625 25.985 ;
        RECT 78.085 25.175 78.355 25.985 ;
        RECT 79.025 25.175 79.265 25.985 ;
        RECT 81.990 25.980 82.425 25.985 ;
        RECT 82.155 25.175 82.425 25.980 ;
        RECT 83.095 25.175 83.335 25.985 ;
        RECT 85.795 25.175 86.065 25.985 ;
        RECT 86.735 25.175 86.975 25.985 ;
        RECT 89.700 25.980 90.135 25.985 ;
        RECT 89.865 25.175 90.135 25.980 ;
        RECT 90.805 25.175 91.045 25.985 ;
        RECT 92.325 25.965 93.775 25.985 ;
        RECT 22.670 22.170 23.170 22.610 ;
        RECT 22.200 22.165 23.170 22.170 ;
        RECT 20.445 22.005 23.170 22.165 ;
        RECT 60.840 22.450 61.710 22.790 ;
        RECT 20.445 21.835 29.560 22.005 ;
        RECT 20.445 21.775 22.610 21.835 ;
        RECT 20.445 17.715 20.835 21.775 ;
        RECT 22.380 21.035 22.610 21.775 ;
        RECT 23.280 21.375 23.450 21.835 ;
        RECT 24.120 21.375 24.290 21.835 ;
        RECT 24.960 21.375 25.130 21.835 ;
        RECT 25.800 21.375 25.970 21.835 ;
        RECT 26.640 21.375 26.810 21.835 ;
        RECT 27.480 21.375 27.650 21.835 ;
        RECT 28.320 21.375 28.490 21.835 ;
        RECT 29.160 21.035 29.370 21.835 ;
        RECT 60.840 21.450 61.180 22.450 ;
        RECT 92.325 22.425 92.635 25.965 ;
        RECT 93.505 25.175 93.775 25.965 ;
        RECT 94.445 25.175 94.685 25.985 ;
        RECT 97.410 25.980 97.845 25.985 ;
        RECT 97.575 25.175 97.845 25.980 ;
        RECT 98.515 25.175 98.755 25.985 ;
        RECT 101.215 25.175 101.485 25.985 ;
        RECT 102.155 25.175 102.395 25.985 ;
        RECT 105.120 25.980 105.555 25.985 ;
        RECT 105.285 25.175 105.555 25.980 ;
        RECT 106.225 25.175 106.465 25.985 ;
        RECT 108.925 25.175 109.195 25.985 ;
        RECT 109.865 25.175 110.105 25.985 ;
        RECT 112.830 25.980 113.265 25.985 ;
        RECT 112.995 25.175 113.265 25.980 ;
        RECT 113.935 25.175 114.175 25.985 ;
        RECT 116.635 25.175 116.905 25.985 ;
        RECT 117.575 25.175 117.815 25.985 ;
        RECT 120.540 25.980 120.975 25.985 ;
        RECT 120.705 25.175 120.975 25.980 ;
        RECT 121.645 25.175 121.885 25.985 ;
        RECT 91.775 22.115 92.635 22.425 ;
        RECT 83.860 22.025 91.220 22.035 ;
        RECT 83.860 22.020 91.340 22.025 ;
        RECT 91.775 22.020 92.085 22.115 ;
        RECT 83.860 21.865 92.085 22.020 ;
        RECT 59.110 21.265 61.180 21.450 ;
        RECT 55.410 21.110 61.180 21.265 ;
        RECT 55.410 21.095 59.550 21.110 ;
        RECT 55.665 20.635 55.920 21.095 ;
        RECT 56.590 20.635 56.760 21.095 ;
        RECT 57.430 20.635 57.600 21.095 ;
        RECT 58.270 20.635 58.440 21.095 ;
        RECT 59.110 20.635 59.415 21.095 ;
        RECT 84.040 21.065 84.270 21.865 ;
        RECT 84.940 21.405 85.110 21.865 ;
        RECT 85.780 21.405 85.950 21.865 ;
        RECT 86.620 21.405 86.790 21.865 ;
        RECT 87.460 21.405 87.630 21.865 ;
        RECT 88.300 21.405 88.470 21.865 ;
        RECT 89.140 21.405 89.310 21.865 ;
        RECT 89.980 21.405 90.150 21.865 ;
        RECT 90.820 21.715 92.085 21.865 ;
        RECT 90.820 21.065 91.030 21.715 ;
        RECT 20.445 17.325 21.375 17.715 ;
        RECT 20.985 11.100 21.375 17.325 ;
        RECT 55.770 15.465 56.000 16.285 ;
        RECT 55.450 15.295 56.830 15.465 ;
        RECT 57.240 15.455 57.505 15.915 ;
        RECT 58.175 15.455 58.345 15.915 ;
        RECT 59.015 15.455 59.265 15.920 ;
        RECT 57.110 15.285 59.410 15.455 ;
        RECT 55.390 14.885 59.530 15.055 ;
        RECT 55.645 14.425 55.900 14.885 ;
        RECT 56.570 14.425 56.740 14.885 ;
        RECT 57.410 14.425 57.580 14.885 ;
        RECT 58.250 14.425 58.420 14.885 ;
        RECT 59.090 14.425 59.395 14.885 ;
        RECT 22.510 11.100 22.740 11.835 ;
        RECT 20.985 11.035 22.740 11.100 ;
        RECT 23.410 11.035 23.580 11.495 ;
        RECT 24.250 11.035 24.420 11.495 ;
        RECT 25.090 11.035 25.260 11.495 ;
        RECT 25.930 11.035 26.100 11.495 ;
        RECT 26.770 11.035 26.940 11.495 ;
        RECT 27.610 11.035 27.780 11.495 ;
        RECT 28.450 11.035 28.620 11.495 ;
        RECT 29.290 11.035 29.500 11.835 ;
        RECT 20.985 10.865 29.690 11.035 ;
        RECT 84.170 11.005 84.400 11.805 ;
        RECT 85.070 11.005 85.240 11.465 ;
        RECT 85.910 11.005 86.080 11.465 ;
        RECT 86.750 11.005 86.920 11.465 ;
        RECT 87.590 11.005 87.760 11.465 ;
        RECT 88.430 11.005 88.600 11.465 ;
        RECT 89.270 11.005 89.440 11.465 ;
        RECT 90.110 11.005 90.280 11.465 ;
        RECT 90.950 11.010 91.160 11.805 ;
        RECT 91.775 11.010 92.085 21.715 ;
        RECT 124.925 14.895 125.255 15.275 ;
        RECT 124.400 14.725 125.780 14.895 ;
        RECT 90.950 11.005 92.110 11.010 ;
        RECT 20.985 10.710 22.740 10.865 ;
        RECT 83.990 10.835 92.110 11.005 ;
        RECT 1.155 7.475 1.395 8.285 ;
        RECT 2.065 7.480 2.335 8.285 ;
        RECT 2.065 7.475 2.500 7.480 ;
        RECT 5.225 7.475 5.465 8.285 ;
        RECT 6.135 7.475 6.405 8.285 ;
        RECT 8.865 7.475 9.105 8.285 ;
        RECT 9.775 7.480 10.045 8.285 ;
        RECT 9.775 7.475 10.210 7.480 ;
        RECT 12.935 7.475 13.175 8.285 ;
        RECT 13.845 7.475 14.115 8.285 ;
        RECT 16.575 7.475 16.815 8.285 ;
        RECT 17.485 7.480 17.755 8.285 ;
        RECT 17.485 7.475 17.920 7.480 ;
        RECT 20.645 7.475 20.885 8.285 ;
        RECT 21.555 7.555 21.825 8.285 ;
        RECT 22.335 7.555 22.725 10.710 ;
        RECT 90.960 10.700 92.110 10.835 ;
        RECT 21.545 7.475 22.725 7.555 ;
        RECT 24.285 7.475 24.525 8.285 ;
        RECT 25.195 7.480 25.465 8.285 ;
        RECT 25.195 7.475 25.630 7.480 ;
        RECT 28.355 7.475 28.595 8.285 ;
        RECT 29.265 7.475 29.535 8.285 ;
        RECT 31.995 7.475 32.235 8.285 ;
        RECT 32.905 7.480 33.175 8.285 ;
        RECT 32.905 7.475 33.340 7.480 ;
        RECT 36.065 7.475 36.305 8.285 ;
        RECT 36.975 7.475 37.245 8.285 ;
        RECT 39.705 7.475 39.945 8.285 ;
        RECT 40.615 7.480 40.885 8.285 ;
        RECT 40.615 7.475 41.050 7.480 ;
        RECT 43.775 7.475 44.015 8.285 ;
        RECT 44.685 7.475 44.955 8.285 ;
        RECT 47.415 7.475 47.655 8.285 ;
        RECT 48.325 7.480 48.595 8.285 ;
        RECT 48.325 7.475 48.760 7.480 ;
        RECT 51.485 7.475 51.725 8.285 ;
        RECT 52.395 7.475 52.665 8.285 ;
        RECT 55.125 7.475 55.365 8.285 ;
        RECT 56.035 7.480 56.305 8.285 ;
        RECT 56.035 7.475 56.470 7.480 ;
        RECT 59.195 7.475 59.435 8.285 ;
        RECT 60.105 7.475 60.375 8.285 ;
        RECT 62.835 7.475 63.075 8.285 ;
        RECT 63.745 7.480 64.015 8.285 ;
        RECT 63.745 7.475 64.180 7.480 ;
        RECT 66.905 7.475 67.145 8.285 ;
        RECT 67.815 7.475 68.085 8.285 ;
        RECT 70.545 7.475 70.785 8.285 ;
        RECT 71.455 7.480 71.725 8.285 ;
        RECT 71.455 7.475 71.890 7.480 ;
        RECT 74.615 7.475 74.855 8.285 ;
        RECT 75.525 7.475 75.795 8.285 ;
        RECT 78.255 7.475 78.495 8.285 ;
        RECT 79.165 7.480 79.435 8.285 ;
        RECT 79.165 7.475 79.600 7.480 ;
        RECT 82.325 7.475 82.565 8.285 ;
        RECT 83.235 7.475 83.505 8.285 ;
        RECT 85.965 7.475 86.205 8.285 ;
        RECT 86.875 7.480 87.145 8.285 ;
        RECT 86.875 7.475 87.310 7.480 ;
        RECT 90.035 7.475 90.275 8.285 ;
        RECT 90.945 7.605 91.215 8.285 ;
        RECT 91.755 7.605 92.065 10.700 ;
        RECT 90.945 7.475 92.065 7.605 ;
        RECT 93.675 7.475 93.915 8.285 ;
        RECT 94.585 7.480 94.855 8.285 ;
        RECT 94.585 7.475 95.020 7.480 ;
        RECT 97.745 7.475 97.985 8.285 ;
        RECT 98.655 7.475 98.925 8.285 ;
        RECT 101.385 7.475 101.625 8.285 ;
        RECT 102.295 7.480 102.565 8.285 ;
        RECT 102.295 7.475 102.730 7.480 ;
        RECT 105.455 7.475 105.695 8.285 ;
        RECT 106.365 7.475 106.635 8.285 ;
        RECT 109.095 7.475 109.335 8.285 ;
        RECT 110.005 7.480 110.275 8.285 ;
        RECT 110.005 7.475 110.440 7.480 ;
        RECT 113.165 7.475 113.405 8.285 ;
        RECT 114.075 7.475 114.345 8.285 ;
        RECT 116.805 7.475 117.045 8.285 ;
        RECT 117.715 7.480 117.985 8.285 ;
        RECT 117.715 7.475 118.150 7.480 ;
        RECT 120.875 7.475 121.115 8.285 ;
        RECT 121.785 7.475 122.055 8.285 ;
        RECT 1.050 7.305 2.500 7.475 ;
        RECT 5.120 7.305 6.500 7.475 ;
        RECT 8.760 7.305 10.210 7.475 ;
        RECT 12.830 7.305 14.210 7.475 ;
        RECT 16.470 7.305 17.920 7.475 ;
        RECT 20.540 7.305 22.725 7.475 ;
        RECT 1.050 6.080 1.220 7.305 ;
        RECT 2.330 5.790 2.500 7.305 ;
        RECT 8.760 6.080 8.930 7.305 ;
        RECT 10.040 5.790 10.210 7.305 ;
        RECT 16.470 6.080 16.640 7.305 ;
        RECT 17.750 5.790 17.920 7.305 ;
        RECT 21.545 7.165 22.725 7.305 ;
        RECT 24.180 7.305 25.630 7.475 ;
        RECT 28.250 7.305 29.630 7.475 ;
        RECT 31.890 7.305 33.340 7.475 ;
        RECT 35.960 7.305 37.340 7.475 ;
        RECT 39.600 7.305 41.050 7.475 ;
        RECT 43.670 7.305 45.050 7.475 ;
        RECT 47.310 7.305 48.760 7.475 ;
        RECT 51.380 7.305 52.760 7.475 ;
        RECT 55.020 7.305 56.470 7.475 ;
        RECT 59.090 7.305 60.470 7.475 ;
        RECT 62.730 7.305 64.180 7.475 ;
        RECT 66.800 7.305 68.180 7.475 ;
        RECT 70.440 7.305 71.890 7.475 ;
        RECT 74.510 7.305 75.890 7.475 ;
        RECT 78.150 7.305 79.600 7.475 ;
        RECT 82.220 7.305 83.600 7.475 ;
        RECT 85.860 7.305 87.310 7.475 ;
        RECT 89.930 7.305 92.065 7.475 ;
        RECT 24.180 6.080 24.350 7.305 ;
        RECT 25.460 5.790 25.630 7.305 ;
        RECT 31.890 6.080 32.060 7.305 ;
        RECT 33.170 5.790 33.340 7.305 ;
        RECT 39.600 6.080 39.770 7.305 ;
        RECT 40.880 5.790 41.050 7.305 ;
        RECT 47.310 6.080 47.480 7.305 ;
        RECT 48.590 5.790 48.760 7.305 ;
        RECT 55.020 6.080 55.190 7.305 ;
        RECT 56.300 5.790 56.470 7.305 ;
        RECT 62.730 6.080 62.900 7.305 ;
        RECT 64.010 5.790 64.180 7.305 ;
        RECT 70.440 6.080 70.610 7.305 ;
        RECT 71.720 5.790 71.890 7.305 ;
        RECT 78.150 6.080 78.320 7.305 ;
        RECT 79.430 5.790 79.600 7.305 ;
        RECT 85.860 6.080 86.030 7.305 ;
        RECT 87.140 5.790 87.310 7.305 ;
        RECT 90.995 7.295 92.065 7.305 ;
        RECT 93.570 7.305 95.020 7.475 ;
        RECT 97.640 7.305 99.020 7.475 ;
        RECT 101.280 7.305 102.730 7.475 ;
        RECT 105.350 7.305 106.730 7.475 ;
        RECT 108.990 7.305 110.440 7.475 ;
        RECT 113.060 7.305 114.440 7.475 ;
        RECT 116.700 7.305 118.150 7.475 ;
        RECT 120.770 7.305 122.150 7.475 ;
        RECT 93.570 6.080 93.740 7.305 ;
        RECT 94.850 5.790 95.020 7.305 ;
        RECT 101.280 6.080 101.450 7.305 ;
        RECT 102.560 5.790 102.730 7.305 ;
        RECT 108.990 6.080 109.160 7.305 ;
        RECT 110.270 5.790 110.440 7.305 ;
        RECT 116.700 6.080 116.870 7.305 ;
        RECT 117.980 5.790 118.150 7.305 ;
        RECT 2.330 5.620 4.180 5.790 ;
        RECT 10.040 5.620 11.890 5.790 ;
        RECT 17.750 5.620 19.600 5.790 ;
        RECT 25.460 5.620 27.310 5.790 ;
        RECT 33.170 5.620 35.020 5.790 ;
        RECT 40.880 5.620 42.730 5.790 ;
        RECT 48.590 5.620 50.440 5.790 ;
        RECT 56.300 5.620 58.150 5.790 ;
        RECT 64.010 5.620 65.860 5.790 ;
        RECT 71.720 5.620 73.570 5.790 ;
        RECT 79.430 5.620 81.280 5.790 ;
        RECT 87.140 5.620 88.990 5.790 ;
        RECT 94.850 5.620 96.700 5.790 ;
        RECT 102.560 5.620 104.410 5.790 ;
        RECT 110.270 5.620 112.120 5.790 ;
        RECT 117.980 5.620 119.830 5.790 ;
        RECT 2.830 5.570 4.180 5.620 ;
        RECT 5.040 5.570 5.270 5.590 ;
        RECT 2.830 5.400 5.270 5.570 ;
        RECT 10.540 5.570 11.890 5.620 ;
        RECT 12.750 5.570 12.980 5.590 ;
        RECT 10.540 5.400 12.980 5.570 ;
        RECT 18.250 5.570 19.600 5.620 ;
        RECT 20.460 5.570 20.690 5.590 ;
        RECT 18.250 5.400 20.690 5.570 ;
        RECT 25.960 5.570 27.310 5.620 ;
        RECT 28.170 5.570 28.400 5.590 ;
        RECT 25.960 5.400 28.400 5.570 ;
        RECT 33.670 5.570 35.020 5.620 ;
        RECT 35.880 5.570 36.110 5.590 ;
        RECT 33.670 5.400 36.110 5.570 ;
        RECT 41.380 5.570 42.730 5.620 ;
        RECT 43.590 5.570 43.820 5.590 ;
        RECT 41.380 5.400 43.820 5.570 ;
        RECT 49.090 5.570 50.440 5.620 ;
        RECT 51.300 5.570 51.530 5.590 ;
        RECT 49.090 5.400 51.530 5.570 ;
        RECT 56.800 5.570 58.150 5.620 ;
        RECT 59.010 5.570 59.240 5.590 ;
        RECT 56.800 5.400 59.240 5.570 ;
        RECT 64.510 5.570 65.860 5.620 ;
        RECT 66.720 5.570 66.950 5.590 ;
        RECT 64.510 5.400 66.950 5.570 ;
        RECT 72.220 5.570 73.570 5.620 ;
        RECT 74.430 5.570 74.660 5.590 ;
        RECT 72.220 5.400 74.660 5.570 ;
        RECT 79.930 5.570 81.280 5.620 ;
        RECT 82.140 5.570 82.370 5.590 ;
        RECT 79.930 5.400 82.370 5.570 ;
        RECT 87.640 5.570 88.990 5.620 ;
        RECT 89.850 5.570 90.080 5.590 ;
        RECT 87.640 5.400 90.080 5.570 ;
        RECT 95.350 5.570 96.700 5.620 ;
        RECT 97.560 5.570 97.790 5.590 ;
        RECT 95.350 5.400 97.790 5.570 ;
        RECT 103.060 5.570 104.410 5.620 ;
        RECT 105.270 5.570 105.500 5.590 ;
        RECT 103.060 5.400 105.500 5.570 ;
        RECT 110.770 5.570 112.120 5.620 ;
        RECT 112.980 5.570 113.210 5.590 ;
        RECT 110.770 5.400 113.210 5.570 ;
        RECT 118.480 5.570 119.830 5.620 ;
        RECT 120.690 5.570 120.920 5.590 ;
        RECT 118.480 5.400 120.920 5.570 ;
        RECT 5.040 5.370 5.270 5.400 ;
        RECT 12.750 5.370 12.980 5.400 ;
        RECT 20.460 5.370 20.690 5.400 ;
        RECT 28.170 5.370 28.400 5.400 ;
        RECT 35.880 5.370 36.110 5.400 ;
        RECT 43.590 5.370 43.820 5.400 ;
        RECT 51.300 5.370 51.530 5.400 ;
        RECT 59.010 5.370 59.240 5.400 ;
        RECT 66.720 5.370 66.950 5.400 ;
        RECT 74.430 5.370 74.660 5.400 ;
        RECT 82.140 5.370 82.370 5.400 ;
        RECT 89.850 5.370 90.080 5.400 ;
        RECT 97.560 5.370 97.790 5.400 ;
        RECT 105.270 5.370 105.500 5.400 ;
        RECT 112.980 5.370 113.210 5.400 ;
        RECT 120.690 5.370 120.920 5.400 ;
        RECT 0.510 2.235 0.740 3.055 ;
        RECT 6.460 2.245 6.690 3.065 ;
        RECT 0.190 2.065 1.570 2.235 ;
        RECT 5.705 2.075 7.520 2.245 ;
        RECT 8.220 2.235 8.450 3.055 ;
        RECT 14.170 2.245 14.400 3.065 ;
        RECT 5.705 2.035 6.425 2.075 ;
        RECT 7.900 2.065 9.280 2.235 ;
        RECT 13.415 2.075 15.230 2.245 ;
        RECT 15.930 2.235 16.160 3.055 ;
        RECT 21.880 2.245 22.110 3.065 ;
        RECT 13.415 2.035 14.135 2.075 ;
        RECT 15.610 2.065 16.990 2.235 ;
        RECT 21.125 2.075 22.940 2.245 ;
        RECT 23.640 2.235 23.870 3.055 ;
        RECT 29.590 2.245 29.820 3.065 ;
        RECT 21.125 2.035 21.845 2.075 ;
        RECT 23.320 2.065 24.700 2.235 ;
        RECT 28.835 2.075 30.650 2.245 ;
        RECT 31.350 2.235 31.580 3.055 ;
        RECT 37.300 2.245 37.530 3.065 ;
        RECT 28.835 2.035 29.555 2.075 ;
        RECT 31.030 2.065 32.410 2.235 ;
        RECT 36.545 2.075 38.360 2.245 ;
        RECT 39.060 2.235 39.290 3.055 ;
        RECT 45.010 2.245 45.240 3.065 ;
        RECT 36.545 2.035 37.265 2.075 ;
        RECT 38.740 2.065 40.120 2.235 ;
        RECT 44.255 2.075 46.070 2.245 ;
        RECT 46.770 2.235 47.000 3.055 ;
        RECT 52.720 2.245 52.950 3.065 ;
        RECT 44.255 2.035 44.975 2.075 ;
        RECT 46.450 2.065 47.830 2.235 ;
        RECT 51.965 2.075 53.780 2.245 ;
        RECT 54.480 2.235 54.710 3.055 ;
        RECT 60.430 2.245 60.660 3.065 ;
        RECT 51.965 2.035 52.685 2.075 ;
        RECT 54.160 2.065 55.540 2.235 ;
        RECT 59.675 2.075 61.490 2.245 ;
        RECT 62.190 2.235 62.420 3.055 ;
        RECT 68.140 2.245 68.370 3.065 ;
        RECT 59.675 2.035 60.395 2.075 ;
        RECT 61.870 2.065 63.250 2.235 ;
        RECT 67.385 2.075 69.200 2.245 ;
        RECT 69.900 2.235 70.130 3.055 ;
        RECT 75.850 2.245 76.080 3.065 ;
        RECT 67.385 2.035 68.105 2.075 ;
        RECT 69.580 2.065 70.960 2.235 ;
        RECT 75.095 2.075 76.910 2.245 ;
        RECT 77.610 2.235 77.840 3.055 ;
        RECT 83.560 2.245 83.790 3.065 ;
        RECT 75.095 2.035 75.815 2.075 ;
        RECT 77.290 2.065 78.670 2.235 ;
        RECT 82.805 2.075 84.620 2.245 ;
        RECT 85.320 2.235 85.550 3.055 ;
        RECT 91.270 2.245 91.500 3.065 ;
        RECT 82.805 2.035 83.525 2.075 ;
        RECT 85.000 2.065 86.380 2.235 ;
        RECT 90.515 2.075 92.330 2.245 ;
        RECT 93.030 2.235 93.260 3.055 ;
        RECT 98.980 2.245 99.210 3.065 ;
        RECT 90.515 2.035 91.235 2.075 ;
        RECT 92.710 2.065 94.090 2.235 ;
        RECT 98.225 2.075 100.040 2.245 ;
        RECT 100.740 2.235 100.970 3.055 ;
        RECT 106.690 2.245 106.920 3.065 ;
        RECT 98.225 2.035 98.945 2.075 ;
        RECT 100.420 2.065 101.800 2.235 ;
        RECT 105.935 2.075 107.750 2.245 ;
        RECT 108.450 2.235 108.680 3.055 ;
        RECT 114.400 2.245 114.630 3.065 ;
        RECT 105.935 2.035 106.655 2.075 ;
        RECT 108.130 2.065 109.510 2.235 ;
        RECT 113.645 2.075 115.460 2.245 ;
        RECT 116.160 2.235 116.390 3.055 ;
        RECT 122.110 2.245 122.340 3.065 ;
        RECT 113.645 2.035 114.365 2.075 ;
        RECT 115.840 2.065 117.220 2.235 ;
        RECT 121.355 2.075 123.170 2.245 ;
        RECT 121.355 2.035 122.075 2.075 ;
        RECT 2.820 0.500 4.170 0.510 ;
        RECT 5.705 0.500 5.915 2.035 ;
        RECT 2.820 0.290 5.915 0.500 ;
        RECT 10.530 0.500 11.880 0.510 ;
        RECT 13.415 0.500 13.625 2.035 ;
        RECT 10.530 0.290 13.625 0.500 ;
        RECT 18.240 0.500 19.590 0.510 ;
        RECT 21.125 0.500 21.335 2.035 ;
        RECT 18.240 0.290 21.335 0.500 ;
        RECT 25.950 0.500 27.300 0.510 ;
        RECT 28.835 0.500 29.045 2.035 ;
        RECT 25.950 0.290 29.045 0.500 ;
        RECT 33.660 0.500 35.010 0.510 ;
        RECT 36.545 0.500 36.755 2.035 ;
        RECT 33.660 0.290 36.755 0.500 ;
        RECT 41.370 0.500 42.720 0.510 ;
        RECT 44.255 0.500 44.465 2.035 ;
        RECT 41.370 0.290 44.465 0.500 ;
        RECT 49.080 0.500 50.430 0.510 ;
        RECT 51.965 0.500 52.175 2.035 ;
        RECT 49.080 0.290 52.175 0.500 ;
        RECT 56.790 0.500 58.140 0.510 ;
        RECT 59.675 0.500 59.885 2.035 ;
        RECT 56.790 0.290 59.885 0.500 ;
        RECT 64.500 0.500 65.850 0.510 ;
        RECT 67.385 0.500 67.595 2.035 ;
        RECT 64.500 0.290 67.595 0.500 ;
        RECT 72.210 0.500 73.560 0.510 ;
        RECT 75.095 0.500 75.305 2.035 ;
        RECT 72.210 0.290 75.305 0.500 ;
        RECT 79.920 0.500 81.270 0.510 ;
        RECT 82.805 0.500 83.015 2.035 ;
        RECT 79.920 0.290 83.015 0.500 ;
        RECT 87.630 0.500 88.980 0.510 ;
        RECT 90.515 0.500 90.725 2.035 ;
        RECT 87.630 0.290 90.725 0.500 ;
        RECT 95.340 0.500 96.690 0.510 ;
        RECT 98.225 0.500 98.435 2.035 ;
        RECT 95.340 0.290 98.435 0.500 ;
        RECT 103.050 0.500 104.400 0.510 ;
        RECT 105.935 0.500 106.145 2.035 ;
        RECT 103.050 0.290 106.145 0.500 ;
        RECT 110.760 0.500 112.110 0.510 ;
        RECT 113.645 0.500 113.855 2.035 ;
        RECT 110.760 0.290 113.855 0.500 ;
        RECT 118.470 0.500 119.820 0.510 ;
        RECT 121.355 0.500 121.565 2.035 ;
        RECT 118.470 0.290 121.565 0.500 ;
        RECT 2.820 0.120 4.170 0.290 ;
        RECT 10.530 0.120 11.880 0.290 ;
        RECT 18.240 0.120 19.590 0.290 ;
        RECT 25.950 0.120 27.300 0.290 ;
        RECT 33.660 0.120 35.010 0.290 ;
        RECT 41.370 0.120 42.720 0.290 ;
        RECT 49.080 0.120 50.430 0.290 ;
        RECT 56.790 0.120 58.140 0.290 ;
        RECT 64.500 0.120 65.850 0.290 ;
        RECT 72.210 0.120 73.560 0.290 ;
        RECT 79.920 0.120 81.270 0.290 ;
        RECT 87.630 0.120 88.980 0.290 ;
        RECT 95.340 0.120 96.690 0.290 ;
        RECT 103.050 0.120 104.400 0.290 ;
        RECT 110.760 0.120 112.110 0.290 ;
        RECT 118.470 0.120 119.820 0.290 ;
      LAYER mcon ;
        RECT 4.290 33.060 4.520 33.260 ;
        RECT 12.000 33.060 12.230 33.260 ;
        RECT 19.710 33.060 19.940 33.260 ;
        RECT 27.420 33.060 27.650 33.260 ;
        RECT 35.130 33.060 35.360 33.260 ;
        RECT 42.840 33.060 43.070 33.260 ;
        RECT 50.550 33.060 50.780 33.260 ;
        RECT 58.260 33.060 58.490 33.260 ;
        RECT 65.970 33.060 66.200 33.260 ;
        RECT 73.680 33.060 73.910 33.260 ;
        RECT 81.390 33.060 81.620 33.260 ;
        RECT 89.100 33.060 89.330 33.260 ;
        RECT 96.810 33.060 97.040 33.260 ;
        RECT 104.520 33.060 104.750 33.260 ;
        RECT 112.230 33.060 112.460 33.260 ;
        RECT 119.940 33.060 120.170 33.260 ;
        RECT 0.015 31.215 0.185 31.385 ;
        RECT 0.475 31.215 0.645 31.385 ;
        RECT 0.935 31.215 1.105 31.385 ;
        RECT 5.965 31.225 6.135 31.395 ;
        RECT 6.425 31.225 6.595 31.395 ;
        RECT 6.885 31.225 7.055 31.395 ;
        RECT 7.725 31.215 7.895 31.385 ;
        RECT 8.185 31.215 8.355 31.385 ;
        RECT 8.645 31.215 8.815 31.385 ;
        RECT 13.675 31.225 13.845 31.395 ;
        RECT 14.135 31.225 14.305 31.395 ;
        RECT 14.595 31.225 14.765 31.395 ;
        RECT 15.435 31.215 15.605 31.385 ;
        RECT 15.895 31.215 16.065 31.385 ;
        RECT 16.355 31.215 16.525 31.385 ;
        RECT 21.385 31.225 21.555 31.395 ;
        RECT 21.845 31.225 22.015 31.395 ;
        RECT 22.305 31.225 22.475 31.395 ;
        RECT 23.145 31.215 23.315 31.385 ;
        RECT 23.605 31.215 23.775 31.385 ;
        RECT 24.065 31.215 24.235 31.385 ;
        RECT 29.095 31.225 29.265 31.395 ;
        RECT 29.555 31.225 29.725 31.395 ;
        RECT 30.015 31.225 30.185 31.395 ;
        RECT 30.855 31.215 31.025 31.385 ;
        RECT 31.315 31.215 31.485 31.385 ;
        RECT 31.775 31.215 31.945 31.385 ;
        RECT 36.805 31.225 36.975 31.395 ;
        RECT 37.265 31.225 37.435 31.395 ;
        RECT 37.725 31.225 37.895 31.395 ;
        RECT 38.565 31.215 38.735 31.385 ;
        RECT 39.025 31.215 39.195 31.385 ;
        RECT 39.485 31.215 39.655 31.385 ;
        RECT 44.515 31.225 44.685 31.395 ;
        RECT 44.975 31.225 45.145 31.395 ;
        RECT 45.435 31.225 45.605 31.395 ;
        RECT 46.275 31.215 46.445 31.385 ;
        RECT 46.735 31.215 46.905 31.385 ;
        RECT 47.195 31.215 47.365 31.385 ;
        RECT 52.225 31.225 52.395 31.395 ;
        RECT 52.685 31.225 52.855 31.395 ;
        RECT 53.145 31.225 53.315 31.395 ;
        RECT 53.985 31.215 54.155 31.385 ;
        RECT 54.445 31.215 54.615 31.385 ;
        RECT 54.905 31.215 55.075 31.385 ;
        RECT 59.935 31.225 60.105 31.395 ;
        RECT 60.395 31.225 60.565 31.395 ;
        RECT 60.855 31.225 61.025 31.395 ;
        RECT 61.695 31.215 61.865 31.385 ;
        RECT 62.155 31.215 62.325 31.385 ;
        RECT 62.615 31.215 62.785 31.385 ;
        RECT 67.645 31.225 67.815 31.395 ;
        RECT 68.105 31.225 68.275 31.395 ;
        RECT 68.565 31.225 68.735 31.395 ;
        RECT 69.405 31.215 69.575 31.385 ;
        RECT 69.865 31.215 70.035 31.385 ;
        RECT 70.325 31.215 70.495 31.385 ;
        RECT 75.355 31.225 75.525 31.395 ;
        RECT 75.815 31.225 75.985 31.395 ;
        RECT 76.275 31.225 76.445 31.395 ;
        RECT 77.115 31.215 77.285 31.385 ;
        RECT 77.575 31.215 77.745 31.385 ;
        RECT 78.035 31.215 78.205 31.385 ;
        RECT 83.065 31.225 83.235 31.395 ;
        RECT 83.525 31.225 83.695 31.395 ;
        RECT 83.985 31.225 84.155 31.395 ;
        RECT 84.825 31.215 84.995 31.385 ;
        RECT 85.285 31.215 85.455 31.385 ;
        RECT 85.745 31.215 85.915 31.385 ;
        RECT 90.775 31.225 90.945 31.395 ;
        RECT 91.235 31.225 91.405 31.395 ;
        RECT 91.695 31.225 91.865 31.395 ;
        RECT 92.535 31.215 92.705 31.385 ;
        RECT 92.995 31.215 93.165 31.385 ;
        RECT 93.455 31.215 93.625 31.385 ;
        RECT 98.485 31.225 98.655 31.395 ;
        RECT 98.945 31.225 99.115 31.395 ;
        RECT 99.405 31.225 99.575 31.395 ;
        RECT 100.245 31.215 100.415 31.385 ;
        RECT 100.705 31.215 100.875 31.385 ;
        RECT 101.165 31.215 101.335 31.385 ;
        RECT 106.195 31.225 106.365 31.395 ;
        RECT 106.655 31.225 106.825 31.395 ;
        RECT 107.115 31.225 107.285 31.395 ;
        RECT 107.955 31.215 108.125 31.385 ;
        RECT 108.415 31.215 108.585 31.385 ;
        RECT 108.875 31.215 109.045 31.385 ;
        RECT 113.905 31.225 114.075 31.395 ;
        RECT 114.365 31.225 114.535 31.395 ;
        RECT 114.825 31.225 114.995 31.395 ;
        RECT 115.665 31.215 115.835 31.385 ;
        RECT 116.125 31.215 116.295 31.385 ;
        RECT 116.585 31.215 116.755 31.385 ;
        RECT 121.615 31.225 121.785 31.395 ;
        RECT 122.075 31.225 122.245 31.395 ;
        RECT 122.535 31.225 122.705 31.395 ;
        RECT 2.140 27.880 2.350 28.050 ;
        RECT 4.280 27.780 4.510 27.980 ;
        RECT 9.850 27.880 10.060 28.050 ;
        RECT 11.990 27.780 12.220 27.980 ;
        RECT 17.560 27.880 17.770 28.050 ;
        RECT 19.700 27.780 19.930 27.980 ;
        RECT 25.270 27.880 25.480 28.050 ;
        RECT 27.410 27.780 27.640 27.980 ;
        RECT 32.980 27.880 33.190 28.050 ;
        RECT 35.120 27.780 35.350 27.980 ;
        RECT 40.690 27.880 40.900 28.050 ;
        RECT 42.830 27.780 43.060 27.980 ;
        RECT 48.400 27.880 48.610 28.050 ;
        RECT 50.540 27.780 50.770 27.980 ;
        RECT 56.110 27.880 56.320 28.050 ;
        RECT 58.250 27.780 58.480 27.980 ;
        RECT 63.820 27.880 64.030 28.050 ;
        RECT 65.960 27.780 66.190 27.980 ;
        RECT 71.530 27.880 71.740 28.050 ;
        RECT 73.670 27.780 73.900 27.980 ;
        RECT 79.240 27.880 79.450 28.050 ;
        RECT 81.380 27.780 81.610 27.980 ;
        RECT 86.950 27.880 87.160 28.050 ;
        RECT 89.090 27.780 89.320 27.980 ;
        RECT 94.660 27.880 94.870 28.050 ;
        RECT 96.800 27.780 97.030 27.980 ;
        RECT 102.370 27.880 102.580 28.050 ;
        RECT 104.510 27.780 104.740 27.980 ;
        RECT 110.080 27.880 110.290 28.050 ;
        RECT 112.220 27.780 112.450 27.980 ;
        RECT 117.790 27.880 118.000 28.050 ;
        RECT 119.930 27.780 120.160 27.980 ;
        RECT 6.170 27.210 6.340 27.380 ;
        RECT 13.880 27.210 14.050 27.380 ;
        RECT 21.590 27.210 21.760 27.380 ;
        RECT 29.300 27.210 29.470 27.380 ;
        RECT 37.010 27.210 37.180 27.380 ;
        RECT 44.720 27.210 44.890 27.380 ;
        RECT 52.430 27.210 52.600 27.380 ;
        RECT 60.140 27.210 60.310 27.380 ;
        RECT 1.035 25.985 1.205 26.155 ;
        RECT 1.495 25.985 1.665 26.155 ;
        RECT 1.955 25.985 2.125 26.155 ;
        RECT 5.105 25.985 5.275 26.155 ;
        RECT 5.565 25.985 5.735 26.155 ;
        RECT 6.025 25.985 6.195 26.155 ;
        RECT 8.745 25.985 8.915 26.155 ;
        RECT 9.205 25.985 9.375 26.155 ;
        RECT 9.665 25.985 9.835 26.155 ;
        RECT 12.815 25.985 12.985 26.155 ;
        RECT 13.275 25.985 13.445 26.155 ;
        RECT 13.735 25.985 13.905 26.155 ;
        RECT 16.455 25.985 16.625 26.155 ;
        RECT 16.915 25.985 17.085 26.155 ;
        RECT 17.375 25.985 17.545 26.155 ;
        RECT 20.525 25.985 20.695 26.155 ;
        RECT 20.985 25.985 21.155 26.155 ;
        RECT 21.445 25.985 21.615 26.155 ;
        RECT 24.165 25.985 24.335 26.155 ;
        RECT 24.625 25.985 24.795 26.155 ;
        RECT 25.085 25.985 25.255 26.155 ;
        RECT 28.235 25.985 28.405 26.155 ;
        RECT 28.695 25.985 28.865 26.155 ;
        RECT 29.155 25.985 29.325 26.155 ;
        RECT 31.875 25.985 32.045 26.155 ;
        RECT 32.335 25.985 32.505 26.155 ;
        RECT 32.795 25.985 32.965 26.155 ;
        RECT 35.945 25.985 36.115 26.155 ;
        RECT 36.405 25.985 36.575 26.155 ;
        RECT 36.865 25.985 37.035 26.155 ;
        RECT 39.585 25.985 39.755 26.155 ;
        RECT 40.045 25.985 40.215 26.155 ;
        RECT 40.505 25.985 40.675 26.155 ;
        RECT 43.655 25.985 43.825 26.155 ;
        RECT 44.115 25.985 44.285 26.155 ;
        RECT 44.575 25.985 44.745 26.155 ;
        RECT 47.295 25.985 47.465 26.155 ;
        RECT 47.755 25.985 47.925 26.155 ;
        RECT 48.215 25.985 48.385 26.155 ;
        RECT 51.365 25.985 51.535 26.155 ;
        RECT 51.825 25.985 51.995 26.155 ;
        RECT 52.285 25.985 52.455 26.155 ;
        RECT 55.005 25.985 55.175 26.155 ;
        RECT 55.465 25.985 55.635 26.155 ;
        RECT 55.925 25.985 56.095 26.155 ;
        RECT 59.075 25.985 59.245 26.155 ;
        RECT 59.535 25.985 59.705 26.155 ;
        RECT 59.995 25.985 60.165 26.155 ;
        RECT 67.850 27.210 68.020 27.380 ;
        RECT 75.560 27.210 75.730 27.380 ;
        RECT 83.270 27.210 83.440 27.380 ;
        RECT 90.980 27.210 91.150 27.380 ;
        RECT 62.715 25.985 62.885 26.155 ;
        RECT 63.175 25.985 63.345 26.155 ;
        RECT 63.635 25.985 63.805 26.155 ;
        RECT 66.785 25.985 66.955 26.155 ;
        RECT 67.245 25.985 67.415 26.155 ;
        RECT 67.705 25.985 67.875 26.155 ;
        RECT 70.425 25.985 70.595 26.155 ;
        RECT 70.885 25.985 71.055 26.155 ;
        RECT 71.345 25.985 71.515 26.155 ;
        RECT 74.495 25.985 74.665 26.155 ;
        RECT 74.955 25.985 75.125 26.155 ;
        RECT 75.415 25.985 75.585 26.155 ;
        RECT 78.135 25.985 78.305 26.155 ;
        RECT 78.595 25.985 78.765 26.155 ;
        RECT 79.055 25.985 79.225 26.155 ;
        RECT 82.205 25.985 82.375 26.155 ;
        RECT 82.665 25.985 82.835 26.155 ;
        RECT 83.125 25.985 83.295 26.155 ;
        RECT 85.845 25.985 86.015 26.155 ;
        RECT 86.305 25.985 86.475 26.155 ;
        RECT 86.765 25.985 86.935 26.155 ;
        RECT 89.915 25.985 90.085 26.155 ;
        RECT 90.375 25.985 90.545 26.155 ;
        RECT 90.835 25.985 91.005 26.155 ;
        RECT 98.690 27.210 98.860 27.380 ;
        RECT 106.400 27.210 106.570 27.380 ;
        RECT 114.110 27.210 114.280 27.380 ;
        RECT 121.820 27.210 121.990 27.380 ;
        RECT 93.555 25.985 93.725 26.155 ;
        RECT 94.015 25.985 94.185 26.155 ;
        RECT 94.475 25.985 94.645 26.155 ;
        RECT 97.625 25.985 97.795 26.155 ;
        RECT 98.085 25.985 98.255 26.155 ;
        RECT 98.545 25.985 98.715 26.155 ;
        RECT 101.265 25.985 101.435 26.155 ;
        RECT 101.725 25.985 101.895 26.155 ;
        RECT 102.185 25.985 102.355 26.155 ;
        RECT 105.335 25.985 105.505 26.155 ;
        RECT 105.795 25.985 105.965 26.155 ;
        RECT 106.255 25.985 106.425 26.155 ;
        RECT 108.975 25.985 109.145 26.155 ;
        RECT 109.435 25.985 109.605 26.155 ;
        RECT 109.895 25.985 110.065 26.155 ;
        RECT 113.045 25.985 113.215 26.155 ;
        RECT 113.505 25.985 113.675 26.155 ;
        RECT 113.965 25.985 114.135 26.155 ;
        RECT 116.685 25.985 116.855 26.155 ;
        RECT 117.145 25.985 117.315 26.155 ;
        RECT 117.605 25.985 117.775 26.155 ;
        RECT 120.755 25.985 120.925 26.155 ;
        RECT 121.215 25.985 121.385 26.155 ;
        RECT 121.675 25.985 121.845 26.155 ;
        RECT 22.345 21.835 22.515 22.005 ;
        RECT 22.805 21.835 22.975 22.005 ;
        RECT 23.265 21.835 23.435 22.005 ;
        RECT 23.725 21.835 23.895 22.005 ;
        RECT 24.185 21.835 24.355 22.005 ;
        RECT 24.645 21.835 24.815 22.005 ;
        RECT 25.105 21.835 25.275 22.005 ;
        RECT 25.565 21.835 25.735 22.005 ;
        RECT 26.025 21.835 26.195 22.005 ;
        RECT 26.485 21.835 26.655 22.005 ;
        RECT 26.945 21.835 27.115 22.005 ;
        RECT 27.405 21.835 27.575 22.005 ;
        RECT 27.865 21.835 28.035 22.005 ;
        RECT 28.325 21.835 28.495 22.005 ;
        RECT 28.785 21.835 28.955 22.005 ;
        RECT 29.245 21.835 29.415 22.005 ;
        RECT 84.005 21.865 84.175 22.035 ;
        RECT 84.465 21.865 84.635 22.035 ;
        RECT 84.925 21.865 85.095 22.035 ;
        RECT 85.385 21.865 85.555 22.035 ;
        RECT 85.845 21.865 86.015 22.035 ;
        RECT 86.305 21.865 86.475 22.035 ;
        RECT 86.765 21.865 86.935 22.035 ;
        RECT 87.225 21.865 87.395 22.035 ;
        RECT 87.685 21.865 87.855 22.035 ;
        RECT 88.145 21.865 88.315 22.035 ;
        RECT 88.605 21.865 88.775 22.035 ;
        RECT 89.065 21.865 89.235 22.035 ;
        RECT 89.525 21.865 89.695 22.035 ;
        RECT 89.985 21.865 90.155 22.035 ;
        RECT 90.445 21.865 90.615 22.035 ;
        RECT 90.905 21.865 91.075 22.035 ;
        RECT 55.555 21.095 55.725 21.265 ;
        RECT 56.015 21.095 56.185 21.265 ;
        RECT 56.475 21.095 56.645 21.265 ;
        RECT 56.935 21.095 57.105 21.265 ;
        RECT 57.395 21.095 57.565 21.265 ;
        RECT 57.855 21.095 58.025 21.265 ;
        RECT 58.315 21.095 58.485 21.265 ;
        RECT 58.775 21.095 58.945 21.265 ;
        RECT 59.235 21.095 59.405 21.265 ;
        RECT 55.595 15.295 55.765 15.465 ;
        RECT 56.055 15.295 56.225 15.465 ;
        RECT 56.515 15.295 56.685 15.465 ;
        RECT 57.255 15.285 57.425 15.455 ;
        RECT 57.715 15.285 57.885 15.455 ;
        RECT 58.175 15.285 58.345 15.455 ;
        RECT 58.635 15.285 58.805 15.455 ;
        RECT 59.095 15.285 59.265 15.455 ;
        RECT 55.535 14.885 55.705 15.055 ;
        RECT 55.995 14.885 56.165 15.055 ;
        RECT 56.455 14.885 56.625 15.055 ;
        RECT 56.915 14.885 57.085 15.055 ;
        RECT 57.375 14.885 57.545 15.055 ;
        RECT 57.835 14.885 58.005 15.055 ;
        RECT 58.295 14.885 58.465 15.055 ;
        RECT 58.755 14.885 58.925 15.055 ;
        RECT 59.215 14.885 59.385 15.055 ;
        RECT 22.475 10.865 22.645 11.035 ;
        RECT 22.935 10.865 23.105 11.035 ;
        RECT 23.395 10.865 23.565 11.035 ;
        RECT 23.855 10.865 24.025 11.035 ;
        RECT 24.315 10.865 24.485 11.035 ;
        RECT 24.775 10.865 24.945 11.035 ;
        RECT 25.235 10.865 25.405 11.035 ;
        RECT 25.695 10.865 25.865 11.035 ;
        RECT 26.155 10.865 26.325 11.035 ;
        RECT 26.615 10.865 26.785 11.035 ;
        RECT 27.075 10.865 27.245 11.035 ;
        RECT 27.535 10.865 27.705 11.035 ;
        RECT 27.995 10.865 28.165 11.035 ;
        RECT 28.455 10.865 28.625 11.035 ;
        RECT 28.915 10.865 29.085 11.035 ;
        RECT 29.375 10.865 29.545 11.035 ;
        RECT 124.545 14.725 124.715 14.895 ;
        RECT 125.005 14.725 125.175 14.895 ;
        RECT 125.465 14.725 125.635 14.895 ;
        RECT 84.135 10.835 84.305 11.005 ;
        RECT 84.595 10.835 84.765 11.005 ;
        RECT 85.055 10.835 85.225 11.005 ;
        RECT 85.515 10.835 85.685 11.005 ;
        RECT 85.975 10.835 86.145 11.005 ;
        RECT 86.435 10.835 86.605 11.005 ;
        RECT 86.895 10.835 87.065 11.005 ;
        RECT 87.355 10.835 87.525 11.005 ;
        RECT 87.815 10.835 87.985 11.005 ;
        RECT 88.275 10.835 88.445 11.005 ;
        RECT 88.735 10.835 88.905 11.005 ;
        RECT 89.195 10.835 89.365 11.005 ;
        RECT 89.655 10.835 89.825 11.005 ;
        RECT 90.115 10.835 90.285 11.005 ;
        RECT 90.575 10.835 90.745 11.005 ;
        RECT 91.035 10.835 91.205 11.005 ;
        RECT 1.195 7.305 1.365 7.475 ;
        RECT 1.655 7.305 1.825 7.475 ;
        RECT 2.115 7.305 2.285 7.475 ;
        RECT 5.265 7.305 5.435 7.475 ;
        RECT 5.725 7.305 5.895 7.475 ;
        RECT 6.185 7.305 6.355 7.475 ;
        RECT 8.905 7.305 9.075 7.475 ;
        RECT 9.365 7.305 9.535 7.475 ;
        RECT 9.825 7.305 9.995 7.475 ;
        RECT 12.975 7.305 13.145 7.475 ;
        RECT 13.435 7.305 13.605 7.475 ;
        RECT 13.895 7.305 14.065 7.475 ;
        RECT 16.615 7.305 16.785 7.475 ;
        RECT 17.075 7.305 17.245 7.475 ;
        RECT 17.535 7.305 17.705 7.475 ;
        RECT 20.685 7.305 20.855 7.475 ;
        RECT 21.145 7.305 21.315 7.475 ;
        RECT 21.605 7.305 21.775 7.475 ;
        RECT 24.325 7.305 24.495 7.475 ;
        RECT 24.785 7.305 24.955 7.475 ;
        RECT 25.245 7.305 25.415 7.475 ;
        RECT 28.395 7.305 28.565 7.475 ;
        RECT 28.855 7.305 29.025 7.475 ;
        RECT 29.315 7.305 29.485 7.475 ;
        RECT 32.035 7.305 32.205 7.475 ;
        RECT 32.495 7.305 32.665 7.475 ;
        RECT 32.955 7.305 33.125 7.475 ;
        RECT 36.105 7.305 36.275 7.475 ;
        RECT 36.565 7.305 36.735 7.475 ;
        RECT 37.025 7.305 37.195 7.475 ;
        RECT 39.745 7.305 39.915 7.475 ;
        RECT 40.205 7.305 40.375 7.475 ;
        RECT 40.665 7.305 40.835 7.475 ;
        RECT 43.815 7.305 43.985 7.475 ;
        RECT 44.275 7.305 44.445 7.475 ;
        RECT 44.735 7.305 44.905 7.475 ;
        RECT 47.455 7.305 47.625 7.475 ;
        RECT 47.915 7.305 48.085 7.475 ;
        RECT 48.375 7.305 48.545 7.475 ;
        RECT 51.525 7.305 51.695 7.475 ;
        RECT 51.985 7.305 52.155 7.475 ;
        RECT 52.445 7.305 52.615 7.475 ;
        RECT 55.165 7.305 55.335 7.475 ;
        RECT 55.625 7.305 55.795 7.475 ;
        RECT 56.085 7.305 56.255 7.475 ;
        RECT 59.235 7.305 59.405 7.475 ;
        RECT 59.695 7.305 59.865 7.475 ;
        RECT 60.155 7.305 60.325 7.475 ;
        RECT 62.875 7.305 63.045 7.475 ;
        RECT 63.335 7.305 63.505 7.475 ;
        RECT 63.795 7.305 63.965 7.475 ;
        RECT 66.945 7.305 67.115 7.475 ;
        RECT 67.405 7.305 67.575 7.475 ;
        RECT 67.865 7.305 68.035 7.475 ;
        RECT 70.585 7.305 70.755 7.475 ;
        RECT 71.045 7.305 71.215 7.475 ;
        RECT 71.505 7.305 71.675 7.475 ;
        RECT 74.655 7.305 74.825 7.475 ;
        RECT 75.115 7.305 75.285 7.475 ;
        RECT 75.575 7.305 75.745 7.475 ;
        RECT 78.295 7.305 78.465 7.475 ;
        RECT 78.755 7.305 78.925 7.475 ;
        RECT 79.215 7.305 79.385 7.475 ;
        RECT 82.365 7.305 82.535 7.475 ;
        RECT 82.825 7.305 82.995 7.475 ;
        RECT 83.285 7.305 83.455 7.475 ;
        RECT 86.005 7.305 86.175 7.475 ;
        RECT 86.465 7.305 86.635 7.475 ;
        RECT 86.925 7.305 87.095 7.475 ;
        RECT 90.075 7.305 90.245 7.475 ;
        RECT 90.535 7.305 90.705 7.475 ;
        RECT 90.995 7.305 91.165 7.475 ;
        RECT 93.715 7.305 93.885 7.475 ;
        RECT 94.175 7.305 94.345 7.475 ;
        RECT 94.635 7.305 94.805 7.475 ;
        RECT 97.785 7.305 97.955 7.475 ;
        RECT 98.245 7.305 98.415 7.475 ;
        RECT 98.705 7.305 98.875 7.475 ;
        RECT 101.425 7.305 101.595 7.475 ;
        RECT 101.885 7.305 102.055 7.475 ;
        RECT 102.345 7.305 102.515 7.475 ;
        RECT 105.495 7.305 105.665 7.475 ;
        RECT 105.955 7.305 106.125 7.475 ;
        RECT 106.415 7.305 106.585 7.475 ;
        RECT 109.135 7.305 109.305 7.475 ;
        RECT 109.595 7.305 109.765 7.475 ;
        RECT 110.055 7.305 110.225 7.475 ;
        RECT 113.205 7.305 113.375 7.475 ;
        RECT 113.665 7.305 113.835 7.475 ;
        RECT 114.125 7.305 114.295 7.475 ;
        RECT 116.845 7.305 117.015 7.475 ;
        RECT 117.305 7.305 117.475 7.475 ;
        RECT 117.765 7.305 117.935 7.475 ;
        RECT 120.915 7.305 121.085 7.475 ;
        RECT 121.375 7.305 121.545 7.475 ;
        RECT 121.835 7.305 122.005 7.475 ;
        RECT 2.880 5.480 3.110 5.680 ;
        RECT 5.040 5.410 5.250 5.580 ;
        RECT 10.590 5.480 10.820 5.680 ;
        RECT 12.750 5.410 12.960 5.580 ;
        RECT 18.300 5.480 18.530 5.680 ;
        RECT 20.460 5.410 20.670 5.580 ;
        RECT 26.010 5.480 26.240 5.680 ;
        RECT 28.170 5.410 28.380 5.580 ;
        RECT 33.720 5.480 33.950 5.680 ;
        RECT 35.880 5.410 36.090 5.580 ;
        RECT 41.430 5.480 41.660 5.680 ;
        RECT 43.590 5.410 43.800 5.580 ;
        RECT 49.140 5.480 49.370 5.680 ;
        RECT 51.300 5.410 51.510 5.580 ;
        RECT 56.850 5.480 57.080 5.680 ;
        RECT 59.010 5.410 59.220 5.580 ;
        RECT 64.560 5.480 64.790 5.680 ;
        RECT 66.720 5.410 66.930 5.580 ;
        RECT 72.270 5.480 72.500 5.680 ;
        RECT 74.430 5.410 74.640 5.580 ;
        RECT 79.980 5.480 80.210 5.680 ;
        RECT 82.140 5.410 82.350 5.580 ;
        RECT 87.690 5.480 87.920 5.680 ;
        RECT 89.850 5.410 90.060 5.580 ;
        RECT 95.400 5.480 95.630 5.680 ;
        RECT 97.560 5.410 97.770 5.580 ;
        RECT 103.110 5.480 103.340 5.680 ;
        RECT 105.270 5.410 105.480 5.580 ;
        RECT 110.820 5.480 111.050 5.680 ;
        RECT 112.980 5.410 113.190 5.580 ;
        RECT 118.530 5.480 118.760 5.680 ;
        RECT 120.690 5.410 120.900 5.580 ;
        RECT 0.335 2.065 0.505 2.235 ;
        RECT 0.795 2.065 0.965 2.235 ;
        RECT 1.255 2.065 1.425 2.235 ;
        RECT 6.285 2.075 6.455 2.245 ;
        RECT 6.745 2.075 6.915 2.245 ;
        RECT 7.205 2.075 7.375 2.245 ;
        RECT 8.045 2.065 8.215 2.235 ;
        RECT 8.505 2.065 8.675 2.235 ;
        RECT 8.965 2.065 9.135 2.235 ;
        RECT 13.995 2.075 14.165 2.245 ;
        RECT 14.455 2.075 14.625 2.245 ;
        RECT 14.915 2.075 15.085 2.245 ;
        RECT 15.755 2.065 15.925 2.235 ;
        RECT 16.215 2.065 16.385 2.235 ;
        RECT 16.675 2.065 16.845 2.235 ;
        RECT 21.705 2.075 21.875 2.245 ;
        RECT 22.165 2.075 22.335 2.245 ;
        RECT 22.625 2.075 22.795 2.245 ;
        RECT 23.465 2.065 23.635 2.235 ;
        RECT 23.925 2.065 24.095 2.235 ;
        RECT 24.385 2.065 24.555 2.235 ;
        RECT 29.415 2.075 29.585 2.245 ;
        RECT 29.875 2.075 30.045 2.245 ;
        RECT 30.335 2.075 30.505 2.245 ;
        RECT 31.175 2.065 31.345 2.235 ;
        RECT 31.635 2.065 31.805 2.235 ;
        RECT 32.095 2.065 32.265 2.235 ;
        RECT 37.125 2.075 37.295 2.245 ;
        RECT 37.585 2.075 37.755 2.245 ;
        RECT 38.045 2.075 38.215 2.245 ;
        RECT 38.885 2.065 39.055 2.235 ;
        RECT 39.345 2.065 39.515 2.235 ;
        RECT 39.805 2.065 39.975 2.235 ;
        RECT 44.835 2.075 45.005 2.245 ;
        RECT 45.295 2.075 45.465 2.245 ;
        RECT 45.755 2.075 45.925 2.245 ;
        RECT 46.595 2.065 46.765 2.235 ;
        RECT 47.055 2.065 47.225 2.235 ;
        RECT 47.515 2.065 47.685 2.235 ;
        RECT 52.545 2.075 52.715 2.245 ;
        RECT 53.005 2.075 53.175 2.245 ;
        RECT 53.465 2.075 53.635 2.245 ;
        RECT 54.305 2.065 54.475 2.235 ;
        RECT 54.765 2.065 54.935 2.235 ;
        RECT 55.225 2.065 55.395 2.235 ;
        RECT 60.255 2.075 60.425 2.245 ;
        RECT 60.715 2.075 60.885 2.245 ;
        RECT 61.175 2.075 61.345 2.245 ;
        RECT 62.015 2.065 62.185 2.235 ;
        RECT 62.475 2.065 62.645 2.235 ;
        RECT 62.935 2.065 63.105 2.235 ;
        RECT 67.965 2.075 68.135 2.245 ;
        RECT 68.425 2.075 68.595 2.245 ;
        RECT 68.885 2.075 69.055 2.245 ;
        RECT 69.725 2.065 69.895 2.235 ;
        RECT 70.185 2.065 70.355 2.235 ;
        RECT 70.645 2.065 70.815 2.235 ;
        RECT 75.675 2.075 75.845 2.245 ;
        RECT 76.135 2.075 76.305 2.245 ;
        RECT 76.595 2.075 76.765 2.245 ;
        RECT 77.435 2.065 77.605 2.235 ;
        RECT 77.895 2.065 78.065 2.235 ;
        RECT 78.355 2.065 78.525 2.235 ;
        RECT 83.385 2.075 83.555 2.245 ;
        RECT 83.845 2.075 84.015 2.245 ;
        RECT 84.305 2.075 84.475 2.245 ;
        RECT 85.145 2.065 85.315 2.235 ;
        RECT 85.605 2.065 85.775 2.235 ;
        RECT 86.065 2.065 86.235 2.235 ;
        RECT 91.095 2.075 91.265 2.245 ;
        RECT 91.555 2.075 91.725 2.245 ;
        RECT 92.015 2.075 92.185 2.245 ;
        RECT 92.855 2.065 93.025 2.235 ;
        RECT 93.315 2.065 93.485 2.235 ;
        RECT 93.775 2.065 93.945 2.235 ;
        RECT 98.805 2.075 98.975 2.245 ;
        RECT 99.265 2.075 99.435 2.245 ;
        RECT 99.725 2.075 99.895 2.245 ;
        RECT 100.565 2.065 100.735 2.235 ;
        RECT 101.025 2.065 101.195 2.235 ;
        RECT 101.485 2.065 101.655 2.235 ;
        RECT 106.515 2.075 106.685 2.245 ;
        RECT 106.975 2.075 107.145 2.245 ;
        RECT 107.435 2.075 107.605 2.245 ;
        RECT 108.275 2.065 108.445 2.235 ;
        RECT 108.735 2.065 108.905 2.235 ;
        RECT 109.195 2.065 109.365 2.235 ;
        RECT 114.225 2.075 114.395 2.245 ;
        RECT 114.685 2.075 114.855 2.245 ;
        RECT 115.145 2.075 115.315 2.245 ;
        RECT 115.985 2.065 116.155 2.235 ;
        RECT 116.445 2.065 116.615 2.235 ;
        RECT 116.905 2.065 117.075 2.235 ;
        RECT 121.935 2.075 122.105 2.245 ;
        RECT 122.395 2.075 122.565 2.245 ;
        RECT 122.855 2.075 123.025 2.245 ;
        RECT 2.870 0.200 3.100 0.400 ;
        RECT 10.580 0.200 10.810 0.400 ;
        RECT 18.290 0.200 18.520 0.400 ;
        RECT 26.000 0.200 26.230 0.400 ;
        RECT 33.710 0.200 33.940 0.400 ;
        RECT 41.420 0.200 41.650 0.400 ;
        RECT 49.130 0.200 49.360 0.400 ;
        RECT 56.840 0.200 57.070 0.400 ;
        RECT 64.550 0.200 64.780 0.400 ;
        RECT 72.260 0.200 72.490 0.400 ;
        RECT 79.970 0.200 80.200 0.400 ;
        RECT 87.680 0.200 87.910 0.400 ;
        RECT 95.390 0.200 95.620 0.400 ;
        RECT 103.100 0.200 103.330 0.400 ;
        RECT 110.810 0.200 111.040 0.400 ;
        RECT 118.520 0.200 118.750 0.400 ;
      LAYER met1 ;
        RECT -0.320 32.930 123.040 33.340 ;
        RECT 5.005 31.550 5.175 32.930 ;
        RECT 12.715 31.550 12.885 32.930 ;
        RECT 20.425 31.550 20.595 32.930 ;
        RECT 28.135 31.550 28.305 32.930 ;
        RECT 35.845 31.550 36.015 32.930 ;
        RECT 43.555 31.550 43.725 32.930 ;
        RECT 51.265 31.550 51.435 32.930 ;
        RECT 58.975 31.550 59.145 32.930 ;
        RECT 66.685 31.550 66.855 32.930 ;
        RECT 74.395 31.550 74.565 32.930 ;
        RECT 82.105 31.550 82.275 32.930 ;
        RECT 89.815 31.550 89.985 32.930 ;
        RECT 97.525 31.550 97.695 32.930 ;
        RECT 105.235 31.550 105.405 32.930 ;
        RECT 112.945 31.550 113.115 32.930 ;
        RECT 120.655 31.550 120.825 32.930 ;
        RECT -0.130 31.060 1.250 31.540 ;
        RECT 5.005 31.380 7.200 31.550 ;
        RECT 5.820 31.070 7.200 31.380 ;
        RECT 7.580 31.060 8.960 31.540 ;
        RECT 12.715 31.380 14.910 31.550 ;
        RECT 13.530 31.070 14.910 31.380 ;
        RECT 15.290 31.060 16.670 31.540 ;
        RECT 20.425 31.380 22.620 31.550 ;
        RECT 21.240 31.070 22.620 31.380 ;
        RECT 23.000 31.060 24.380 31.540 ;
        RECT 28.135 31.380 30.330 31.550 ;
        RECT 28.950 31.070 30.330 31.380 ;
        RECT 30.710 31.060 32.090 31.540 ;
        RECT 35.845 31.380 38.040 31.550 ;
        RECT 36.660 31.070 38.040 31.380 ;
        RECT 38.420 31.060 39.800 31.540 ;
        RECT 43.555 31.380 45.750 31.550 ;
        RECT 44.370 31.070 45.750 31.380 ;
        RECT 46.130 31.060 47.510 31.540 ;
        RECT 51.265 31.380 53.460 31.550 ;
        RECT 52.080 31.070 53.460 31.380 ;
        RECT 53.840 31.060 55.220 31.540 ;
        RECT 58.975 31.380 61.170 31.550 ;
        RECT 59.790 31.070 61.170 31.380 ;
        RECT 61.550 31.060 62.930 31.540 ;
        RECT 66.685 31.380 68.880 31.550 ;
        RECT 67.500 31.070 68.880 31.380 ;
        RECT 69.260 31.060 70.640 31.540 ;
        RECT 74.395 31.380 76.590 31.550 ;
        RECT 75.210 31.070 76.590 31.380 ;
        RECT 76.970 31.060 78.350 31.540 ;
        RECT 82.105 31.380 84.300 31.550 ;
        RECT 82.920 31.070 84.300 31.380 ;
        RECT 84.680 31.060 86.060 31.540 ;
        RECT 89.815 31.380 92.010 31.550 ;
        RECT 90.630 31.070 92.010 31.380 ;
        RECT 92.390 31.060 93.770 31.540 ;
        RECT 97.525 31.380 99.720 31.550 ;
        RECT 98.340 31.070 99.720 31.380 ;
        RECT 100.100 31.060 101.480 31.540 ;
        RECT 105.235 31.380 107.430 31.550 ;
        RECT 106.050 31.070 107.430 31.380 ;
        RECT 107.810 31.060 109.190 31.540 ;
        RECT 112.945 31.380 115.140 31.550 ;
        RECT 113.760 31.070 115.140 31.380 ;
        RECT 115.520 31.060 116.900 31.540 ;
        RECT 120.655 31.380 122.850 31.550 ;
        RECT 121.470 31.070 122.850 31.380 ;
        RECT 2.070 27.830 2.410 28.120 ;
        RECT 2.270 26.310 2.410 27.830 ;
        RECT 4.210 27.680 4.570 28.060 ;
        RECT 9.780 27.830 10.120 28.120 ;
        RECT 6.100 27.130 6.430 27.450 ;
        RECT 9.980 26.310 10.120 27.830 ;
        RECT 11.920 27.680 12.280 28.060 ;
        RECT 17.490 27.830 17.830 28.120 ;
        RECT 13.810 27.130 14.140 27.450 ;
        RECT 17.690 26.310 17.830 27.830 ;
        RECT 19.630 27.680 19.990 28.060 ;
        RECT 25.200 27.830 25.540 28.120 ;
        RECT 21.520 27.130 21.850 27.450 ;
        RECT 25.400 26.310 25.540 27.830 ;
        RECT 27.340 27.680 27.700 28.060 ;
        RECT 32.910 27.830 33.250 28.120 ;
        RECT 29.230 27.130 29.560 27.450 ;
        RECT 33.110 26.310 33.250 27.830 ;
        RECT 35.050 27.680 35.410 28.060 ;
        RECT 40.620 27.830 40.960 28.120 ;
        RECT 36.940 27.130 37.270 27.450 ;
        RECT 40.820 26.310 40.960 27.830 ;
        RECT 42.760 27.680 43.120 28.060 ;
        RECT 48.330 27.830 48.670 28.120 ;
        RECT 44.650 27.130 44.980 27.450 ;
        RECT 48.530 26.310 48.670 27.830 ;
        RECT 50.470 27.680 50.830 28.060 ;
        RECT 56.040 27.830 56.380 28.120 ;
        RECT 52.360 27.130 52.690 27.450 ;
        RECT 56.240 26.310 56.380 27.830 ;
        RECT 58.180 27.680 58.540 28.060 ;
        RECT 63.750 27.830 64.090 28.120 ;
        RECT 60.070 27.130 60.400 27.450 ;
        RECT 63.950 26.310 64.090 27.830 ;
        RECT 65.890 27.680 66.250 28.060 ;
        RECT 71.460 27.830 71.800 28.120 ;
        RECT 67.780 27.130 68.110 27.450 ;
        RECT 71.660 26.310 71.800 27.830 ;
        RECT 73.600 27.680 73.960 28.060 ;
        RECT 79.170 27.830 79.510 28.120 ;
        RECT 75.490 27.130 75.820 27.450 ;
        RECT 79.370 26.310 79.510 27.830 ;
        RECT 81.310 27.680 81.670 28.060 ;
        RECT 86.880 27.830 87.220 28.120 ;
        RECT 83.200 27.130 83.530 27.450 ;
        RECT 87.080 26.310 87.220 27.830 ;
        RECT 89.020 27.680 89.380 28.060 ;
        RECT 94.590 27.830 94.930 28.120 ;
        RECT 90.910 27.130 91.240 27.450 ;
        RECT 94.790 26.310 94.930 27.830 ;
        RECT 96.730 27.680 97.090 28.060 ;
        RECT 102.300 27.830 102.640 28.120 ;
        RECT 98.620 27.130 98.950 27.450 ;
        RECT 102.500 26.310 102.640 27.830 ;
        RECT 104.440 27.680 104.800 28.060 ;
        RECT 110.010 27.830 110.350 28.120 ;
        RECT 106.330 27.130 106.660 27.450 ;
        RECT 110.210 26.310 110.350 27.830 ;
        RECT 112.150 27.680 112.510 28.060 ;
        RECT 117.720 27.830 118.060 28.120 ;
        RECT 114.040 27.130 114.370 27.450 ;
        RECT 117.920 26.310 118.060 27.830 ;
        RECT 119.860 27.680 120.220 28.060 ;
        RECT 121.750 27.130 122.080 27.450 ;
        RECT 0.890 26.170 2.410 26.310 ;
        RECT 0.890 25.830 2.270 26.170 ;
        RECT 4.960 25.830 6.340 26.310 ;
        RECT 8.600 26.170 10.120 26.310 ;
        RECT 8.600 25.830 9.980 26.170 ;
        RECT 12.670 25.830 14.050 26.310 ;
        RECT 16.310 26.170 17.830 26.310 ;
        RECT 16.310 25.830 17.690 26.170 ;
        RECT 20.380 25.830 21.760 26.310 ;
        RECT 24.020 26.170 25.540 26.310 ;
        RECT 24.020 25.830 25.400 26.170 ;
        RECT 28.090 25.830 29.470 26.310 ;
        RECT 31.730 26.170 33.250 26.310 ;
        RECT 31.730 25.830 33.110 26.170 ;
        RECT 35.800 25.830 37.180 26.310 ;
        RECT 39.440 26.170 40.960 26.310 ;
        RECT 39.440 25.830 40.820 26.170 ;
        RECT 43.510 25.830 44.890 26.310 ;
        RECT 47.150 26.170 48.670 26.310 ;
        RECT 47.150 25.830 48.530 26.170 ;
        RECT 51.220 25.830 52.600 26.310 ;
        RECT 54.860 26.170 56.380 26.310 ;
        RECT 54.860 25.830 56.240 26.170 ;
        RECT 58.930 25.830 60.310 26.310 ;
        RECT 62.570 26.170 64.090 26.310 ;
        RECT 62.570 25.830 63.950 26.170 ;
        RECT 66.640 25.830 68.020 26.310 ;
        RECT 70.280 26.170 71.800 26.310 ;
        RECT 70.280 25.830 71.660 26.170 ;
        RECT 74.350 25.830 75.730 26.310 ;
        RECT 77.990 26.170 79.510 26.310 ;
        RECT 77.990 25.830 79.370 26.170 ;
        RECT 82.060 25.830 83.440 26.310 ;
        RECT 85.700 26.170 87.220 26.310 ;
        RECT 85.700 25.830 87.080 26.170 ;
        RECT 89.770 25.830 91.150 26.310 ;
        RECT 93.410 26.170 94.930 26.310 ;
        RECT 93.410 25.830 94.790 26.170 ;
        RECT 97.480 25.830 98.860 26.310 ;
        RECT 101.120 26.170 102.640 26.310 ;
        RECT 101.120 25.830 102.500 26.170 ;
        RECT 105.190 25.830 106.570 26.310 ;
        RECT 108.830 26.170 110.350 26.310 ;
        RECT 108.830 25.830 110.210 26.170 ;
        RECT 112.900 25.830 114.280 26.310 ;
        RECT 116.540 26.170 118.060 26.310 ;
        RECT 116.540 25.830 117.920 26.170 ;
        RECT 120.610 25.830 121.990 26.310 ;
        RECT 83.860 22.165 91.220 22.190 ;
        RECT 22.200 21.680 29.560 22.160 ;
        RECT 83.860 21.850 91.270 22.165 ;
        RECT 83.860 21.710 91.220 21.850 ;
        RECT 55.410 21.415 59.550 21.420 ;
        RECT 55.410 20.940 60.425 21.415 ;
        RECT 58.985 20.925 60.425 20.940 ;
        RECT 55.450 15.210 56.830 15.620 ;
        RECT 57.110 15.430 59.410 15.610 ;
        RECT 59.935 15.430 60.425 20.925 ;
        RECT 57.110 15.210 60.425 15.430 ;
        RECT 55.390 14.940 60.425 15.210 ;
        RECT 124.400 15.015 125.780 15.050 ;
        RECT 55.390 14.730 59.530 14.940 ;
        RECT 124.325 14.570 125.780 15.015 ;
        RECT 22.330 11.180 29.690 11.190 ;
        RECT 22.080 11.145 29.690 11.180 ;
        RECT 22.010 10.750 29.690 11.145 ;
        RECT 22.080 10.710 29.690 10.750 ;
        RECT 83.990 11.115 91.520 11.160 ;
        RECT 83.990 10.800 91.540 11.115 ;
        RECT 83.990 10.690 91.520 10.800 ;
        RECT 83.990 10.680 91.350 10.690 ;
        RECT 1.050 7.150 2.430 7.630 ;
        RECT 5.120 7.290 6.500 7.630 ;
        RECT 4.980 7.150 6.500 7.290 ;
        RECT 8.760 7.150 10.140 7.630 ;
        RECT 12.830 7.290 14.210 7.630 ;
        RECT 12.690 7.150 14.210 7.290 ;
        RECT 16.470 7.150 17.850 7.630 ;
        RECT 20.540 7.290 21.920 7.630 ;
        RECT 20.400 7.150 21.920 7.290 ;
        RECT 24.180 7.150 25.560 7.630 ;
        RECT 28.250 7.290 29.630 7.630 ;
        RECT 28.110 7.150 29.630 7.290 ;
        RECT 31.890 7.150 33.270 7.630 ;
        RECT 35.960 7.290 37.340 7.630 ;
        RECT 35.820 7.150 37.340 7.290 ;
        RECT 39.600 7.150 40.980 7.630 ;
        RECT 43.670 7.290 45.050 7.630 ;
        RECT 43.530 7.150 45.050 7.290 ;
        RECT 47.310 7.150 48.690 7.630 ;
        RECT 51.380 7.290 52.760 7.630 ;
        RECT 51.240 7.150 52.760 7.290 ;
        RECT 55.020 7.150 56.400 7.630 ;
        RECT 59.090 7.290 60.470 7.630 ;
        RECT 58.950 7.150 60.470 7.290 ;
        RECT 62.730 7.150 64.110 7.630 ;
        RECT 66.800 7.290 68.180 7.630 ;
        RECT 66.660 7.150 68.180 7.290 ;
        RECT 70.440 7.150 71.820 7.630 ;
        RECT 74.510 7.290 75.890 7.630 ;
        RECT 74.370 7.150 75.890 7.290 ;
        RECT 78.150 7.150 79.530 7.630 ;
        RECT 82.220 7.290 83.600 7.630 ;
        RECT 82.080 7.150 83.600 7.290 ;
        RECT 85.860 7.150 87.240 7.630 ;
        RECT 89.930 7.290 91.310 7.630 ;
        RECT 89.790 7.150 91.310 7.290 ;
        RECT 93.570 7.150 94.950 7.630 ;
        RECT 97.640 7.290 99.020 7.630 ;
        RECT 97.500 7.150 99.020 7.290 ;
        RECT 101.280 7.150 102.660 7.630 ;
        RECT 105.350 7.290 106.730 7.630 ;
        RECT 105.210 7.150 106.730 7.290 ;
        RECT 108.990 7.150 110.370 7.630 ;
        RECT 113.060 7.290 114.440 7.630 ;
        RECT 112.920 7.150 114.440 7.290 ;
        RECT 116.700 7.150 118.080 7.630 ;
        RECT 120.770 7.290 122.150 7.630 ;
        RECT 120.630 7.150 122.150 7.290 ;
        RECT 0.960 6.010 1.290 6.330 ;
        RECT 2.820 5.400 3.180 5.780 ;
        RECT 4.980 5.630 5.120 7.150 ;
        RECT 8.670 6.010 9.000 6.330 ;
        RECT 4.980 5.340 5.320 5.630 ;
        RECT 10.530 5.400 10.890 5.780 ;
        RECT 12.690 5.630 12.830 7.150 ;
        RECT 16.380 6.010 16.710 6.330 ;
        RECT 12.690 5.340 13.030 5.630 ;
        RECT 18.240 5.400 18.600 5.780 ;
        RECT 20.400 5.630 20.540 7.150 ;
        RECT 24.090 6.010 24.420 6.330 ;
        RECT 20.400 5.340 20.740 5.630 ;
        RECT 25.950 5.400 26.310 5.780 ;
        RECT 28.110 5.630 28.250 7.150 ;
        RECT 31.800 6.010 32.130 6.330 ;
        RECT 28.110 5.340 28.450 5.630 ;
        RECT 33.660 5.400 34.020 5.780 ;
        RECT 35.820 5.630 35.960 7.150 ;
        RECT 39.510 6.010 39.840 6.330 ;
        RECT 35.820 5.340 36.160 5.630 ;
        RECT 41.370 5.400 41.730 5.780 ;
        RECT 43.530 5.630 43.670 7.150 ;
        RECT 47.220 6.010 47.550 6.330 ;
        RECT 43.530 5.340 43.870 5.630 ;
        RECT 49.080 5.400 49.440 5.780 ;
        RECT 51.240 5.630 51.380 7.150 ;
        RECT 54.930 6.010 55.260 6.330 ;
        RECT 51.240 5.340 51.580 5.630 ;
        RECT 56.790 5.400 57.150 5.780 ;
        RECT 58.950 5.630 59.090 7.150 ;
        RECT 62.640 6.010 62.970 6.330 ;
        RECT 58.950 5.340 59.290 5.630 ;
        RECT 64.500 5.400 64.860 5.780 ;
        RECT 66.660 5.630 66.800 7.150 ;
        RECT 70.350 6.010 70.680 6.330 ;
        RECT 66.660 5.340 67.000 5.630 ;
        RECT 72.210 5.400 72.570 5.780 ;
        RECT 74.370 5.630 74.510 7.150 ;
        RECT 78.060 6.010 78.390 6.330 ;
        RECT 74.370 5.340 74.710 5.630 ;
        RECT 79.920 5.400 80.280 5.780 ;
        RECT 82.080 5.630 82.220 7.150 ;
        RECT 85.770 6.010 86.100 6.330 ;
        RECT 82.080 5.340 82.420 5.630 ;
        RECT 87.630 5.400 87.990 5.780 ;
        RECT 89.790 5.630 89.930 7.150 ;
        RECT 93.480 6.010 93.810 6.330 ;
        RECT 89.790 5.340 90.130 5.630 ;
        RECT 95.340 5.400 95.700 5.780 ;
        RECT 97.500 5.630 97.640 7.150 ;
        RECT 101.190 6.010 101.520 6.330 ;
        RECT 97.500 5.340 97.840 5.630 ;
        RECT 103.050 5.400 103.410 5.780 ;
        RECT 105.210 5.630 105.350 7.150 ;
        RECT 108.900 6.010 109.230 6.330 ;
        RECT 105.210 5.340 105.550 5.630 ;
        RECT 110.760 5.400 111.120 5.780 ;
        RECT 112.920 5.630 113.060 7.150 ;
        RECT 116.610 6.010 116.940 6.330 ;
        RECT 112.920 5.340 113.260 5.630 ;
        RECT 118.470 5.400 118.830 5.780 ;
        RECT 120.630 5.630 120.770 7.150 ;
        RECT 120.630 5.340 120.970 5.630 ;
        RECT 0.190 2.080 1.570 2.390 ;
        RECT 0.190 1.910 2.385 2.080 ;
        RECT 6.140 1.920 7.520 2.400 ;
        RECT 7.900 2.080 9.280 2.390 ;
        RECT 7.900 1.910 10.095 2.080 ;
        RECT 13.850 1.920 15.230 2.400 ;
        RECT 15.610 2.080 16.990 2.390 ;
        RECT 15.610 1.910 17.805 2.080 ;
        RECT 21.560 1.920 22.940 2.400 ;
        RECT 23.320 2.080 24.700 2.390 ;
        RECT 23.320 1.910 25.515 2.080 ;
        RECT 29.270 1.920 30.650 2.400 ;
        RECT 31.030 2.080 32.410 2.390 ;
        RECT 31.030 1.910 33.225 2.080 ;
        RECT 36.980 1.920 38.360 2.400 ;
        RECT 38.740 2.080 40.120 2.390 ;
        RECT 38.740 1.910 40.935 2.080 ;
        RECT 44.690 1.920 46.070 2.400 ;
        RECT 46.450 2.080 47.830 2.390 ;
        RECT 46.450 1.910 48.645 2.080 ;
        RECT 52.400 1.920 53.780 2.400 ;
        RECT 54.160 2.080 55.540 2.390 ;
        RECT 54.160 1.910 56.355 2.080 ;
        RECT 60.110 1.920 61.490 2.400 ;
        RECT 61.870 2.080 63.250 2.390 ;
        RECT 61.870 1.910 64.065 2.080 ;
        RECT 67.820 1.920 69.200 2.400 ;
        RECT 69.580 2.080 70.960 2.390 ;
        RECT 69.580 1.910 71.775 2.080 ;
        RECT 75.530 1.920 76.910 2.400 ;
        RECT 77.290 2.080 78.670 2.390 ;
        RECT 77.290 1.910 79.485 2.080 ;
        RECT 83.240 1.920 84.620 2.400 ;
        RECT 85.000 2.080 86.380 2.390 ;
        RECT 85.000 1.910 87.195 2.080 ;
        RECT 90.950 1.920 92.330 2.400 ;
        RECT 92.710 2.080 94.090 2.390 ;
        RECT 92.710 1.910 94.905 2.080 ;
        RECT 98.660 1.920 100.040 2.400 ;
        RECT 100.420 2.080 101.800 2.390 ;
        RECT 100.420 1.910 102.615 2.080 ;
        RECT 106.370 1.920 107.750 2.400 ;
        RECT 108.130 2.080 109.510 2.390 ;
        RECT 108.130 1.910 110.325 2.080 ;
        RECT 114.080 1.920 115.460 2.400 ;
        RECT 115.840 2.080 117.220 2.390 ;
        RECT 115.840 1.910 118.035 2.080 ;
        RECT 121.790 1.920 123.170 2.400 ;
        RECT 2.215 0.530 2.385 1.910 ;
        RECT 9.925 0.530 10.095 1.910 ;
        RECT 17.635 0.530 17.805 1.910 ;
        RECT 25.345 0.530 25.515 1.910 ;
        RECT 33.055 0.530 33.225 1.910 ;
        RECT 40.765 0.530 40.935 1.910 ;
        RECT 48.475 0.530 48.645 1.910 ;
        RECT 56.185 0.530 56.355 1.910 ;
        RECT 63.895 0.530 64.065 1.910 ;
        RECT 71.605 0.530 71.775 1.910 ;
        RECT 79.315 0.530 79.485 1.910 ;
        RECT 87.025 0.530 87.195 1.910 ;
        RECT 94.735 0.530 94.905 1.910 ;
        RECT 102.445 0.530 102.615 1.910 ;
        RECT 110.155 0.530 110.325 1.910 ;
        RECT 117.865 0.530 118.035 1.910 ;
        RECT 124.325 0.530 124.735 14.570 ;
        RECT 0.000 0.120 124.735 0.530 ;
      LAYER via ;
        RECT 6.340 31.160 6.630 31.480 ;
        RECT 14.050 31.160 14.340 31.480 ;
        RECT 21.760 31.160 22.050 31.480 ;
        RECT 29.470 31.160 29.760 31.480 ;
        RECT 37.180 31.160 37.470 31.480 ;
        RECT 44.890 31.160 45.180 31.480 ;
        RECT 52.600 31.160 52.890 31.480 ;
        RECT 60.310 31.160 60.600 31.480 ;
        RECT 68.020 31.160 68.310 31.480 ;
        RECT 75.730 31.160 76.020 31.480 ;
        RECT 83.440 31.160 83.730 31.480 ;
        RECT 91.150 31.160 91.440 31.480 ;
        RECT 98.860 31.160 99.150 31.480 ;
        RECT 106.570 31.160 106.860 31.480 ;
        RECT 114.280 31.160 114.570 31.480 ;
        RECT 121.990 31.160 122.280 31.480 ;
        RECT 4.240 27.720 4.540 28.020 ;
        RECT 6.130 27.160 6.390 27.420 ;
        RECT 11.950 27.720 12.250 28.020 ;
        RECT 13.840 27.160 14.100 27.420 ;
        RECT 19.660 27.720 19.960 28.020 ;
        RECT 21.550 27.160 21.810 27.420 ;
        RECT 27.370 27.720 27.670 28.020 ;
        RECT 29.260 27.160 29.520 27.420 ;
        RECT 35.080 27.720 35.380 28.020 ;
        RECT 36.970 27.160 37.230 27.420 ;
        RECT 42.790 27.720 43.090 28.020 ;
        RECT 44.680 27.160 44.940 27.420 ;
        RECT 50.500 27.720 50.800 28.020 ;
        RECT 52.390 27.160 52.650 27.420 ;
        RECT 58.210 27.720 58.510 28.020 ;
        RECT 60.100 27.160 60.360 27.420 ;
        RECT 65.920 27.720 66.220 28.020 ;
        RECT 67.810 27.160 68.070 27.420 ;
        RECT 73.630 27.720 73.930 28.020 ;
        RECT 75.520 27.160 75.780 27.420 ;
        RECT 81.340 27.720 81.640 28.020 ;
        RECT 83.230 27.160 83.490 27.420 ;
        RECT 89.050 27.720 89.350 28.020 ;
        RECT 90.940 27.160 91.200 27.420 ;
        RECT 96.760 27.720 97.060 28.020 ;
        RECT 98.650 27.160 98.910 27.420 ;
        RECT 104.470 27.720 104.770 28.020 ;
        RECT 106.360 27.160 106.620 27.420 ;
        RECT 112.180 27.720 112.480 28.020 ;
        RECT 114.070 27.160 114.330 27.420 ;
        RECT 119.890 27.720 120.190 28.020 ;
        RECT 121.780 27.160 122.040 27.420 ;
        RECT 1.000 6.040 1.260 6.300 ;
        RECT 2.850 5.440 3.150 5.740 ;
        RECT 8.710 6.040 8.970 6.300 ;
        RECT 10.560 5.440 10.860 5.740 ;
        RECT 16.420 6.040 16.680 6.300 ;
        RECT 18.270 5.440 18.570 5.740 ;
        RECT 24.130 6.040 24.390 6.300 ;
        RECT 25.980 5.440 26.280 5.740 ;
        RECT 31.840 6.040 32.100 6.300 ;
        RECT 33.690 5.440 33.990 5.740 ;
        RECT 39.550 6.040 39.810 6.300 ;
        RECT 41.400 5.440 41.700 5.740 ;
        RECT 47.260 6.040 47.520 6.300 ;
        RECT 49.110 5.440 49.410 5.740 ;
        RECT 54.970 6.040 55.230 6.300 ;
        RECT 56.820 5.440 57.120 5.740 ;
        RECT 62.680 6.040 62.940 6.300 ;
        RECT 64.530 5.440 64.830 5.740 ;
        RECT 70.390 6.040 70.650 6.300 ;
        RECT 72.240 5.440 72.540 5.740 ;
        RECT 78.100 6.040 78.360 6.300 ;
        RECT 79.950 5.440 80.250 5.740 ;
        RECT 85.810 6.040 86.070 6.300 ;
        RECT 87.660 5.440 87.960 5.740 ;
        RECT 93.520 6.040 93.780 6.300 ;
        RECT 95.370 5.440 95.670 5.740 ;
        RECT 101.230 6.040 101.490 6.300 ;
        RECT 103.080 5.440 103.380 5.740 ;
        RECT 108.940 6.040 109.200 6.300 ;
        RECT 110.790 5.440 111.090 5.740 ;
        RECT 116.650 6.040 116.910 6.300 ;
        RECT 118.500 5.440 118.800 5.740 ;
        RECT 0.760 1.980 1.050 2.300 ;
        RECT 8.470 1.980 8.760 2.300 ;
        RECT 16.180 1.980 16.470 2.300 ;
        RECT 23.890 1.980 24.180 2.300 ;
        RECT 31.600 1.980 31.890 2.300 ;
        RECT 39.310 1.980 39.600 2.300 ;
        RECT 47.020 1.980 47.310 2.300 ;
        RECT 54.730 1.980 55.020 2.300 ;
        RECT 62.440 1.980 62.730 2.300 ;
        RECT 70.150 1.980 70.440 2.300 ;
        RECT 77.860 1.980 78.150 2.300 ;
        RECT 85.570 1.980 85.860 2.300 ;
        RECT 93.280 1.980 93.570 2.300 ;
        RECT 100.990 1.980 101.280 2.300 ;
        RECT 108.700 1.980 108.990 2.300 ;
        RECT 116.410 1.980 116.700 2.300 ;
      LAYER met2 ;
        RECT 6.310 31.120 6.630 31.530 ;
        RECT 14.020 31.120 14.340 31.530 ;
        RECT 21.730 31.120 22.050 31.530 ;
        RECT 29.440 31.120 29.760 31.530 ;
        RECT 37.150 31.120 37.470 31.530 ;
        RECT 44.860 31.120 45.180 31.530 ;
        RECT 52.570 31.120 52.890 31.530 ;
        RECT 60.280 31.120 60.600 31.530 ;
        RECT 67.990 31.120 68.310 31.530 ;
        RECT 75.700 31.120 76.020 31.530 ;
        RECT 83.410 31.120 83.730 31.530 ;
        RECT 91.120 31.120 91.440 31.530 ;
        RECT 98.830 31.120 99.150 31.530 ;
        RECT 106.540 31.120 106.860 31.530 ;
        RECT 114.250 31.120 114.570 31.530 ;
        RECT 121.960 31.120 122.280 31.530 ;
        RECT 6.490 28.200 6.630 31.120 ;
        RECT 14.200 28.200 14.340 31.120 ;
        RECT 21.910 28.200 22.050 31.120 ;
        RECT 29.620 28.200 29.760 31.120 ;
        RECT 37.330 28.200 37.470 31.120 ;
        RECT 45.040 28.200 45.180 31.120 ;
        RECT 52.750 28.200 52.890 31.120 ;
        RECT 60.460 28.200 60.600 31.120 ;
        RECT 68.170 28.200 68.310 31.120 ;
        RECT 75.880 28.200 76.020 31.120 ;
        RECT 83.590 28.200 83.730 31.120 ;
        RECT 91.300 28.200 91.440 31.120 ;
        RECT 99.010 28.200 99.150 31.120 ;
        RECT 106.720 28.200 106.860 31.120 ;
        RECT 114.430 28.200 114.570 31.120 ;
        RECT 122.140 28.200 122.280 31.120 ;
        RECT 4.210 28.060 4.390 28.070 ;
        RECT 6.290 28.060 6.630 28.200 ;
        RECT 11.920 28.060 12.100 28.070 ;
        RECT 14.000 28.060 14.340 28.200 ;
        RECT 19.630 28.060 19.810 28.070 ;
        RECT 21.710 28.060 22.050 28.200 ;
        RECT 27.340 28.060 27.520 28.070 ;
        RECT 29.420 28.060 29.760 28.200 ;
        RECT 35.050 28.060 35.230 28.070 ;
        RECT 37.130 28.060 37.470 28.200 ;
        RECT 42.760 28.060 42.940 28.070 ;
        RECT 44.840 28.060 45.180 28.200 ;
        RECT 50.470 28.060 50.650 28.070 ;
        RECT 52.550 28.060 52.890 28.200 ;
        RECT 58.180 28.060 58.360 28.070 ;
        RECT 60.260 28.060 60.600 28.200 ;
        RECT 65.890 28.060 66.070 28.070 ;
        RECT 67.970 28.060 68.310 28.200 ;
        RECT 73.600 28.060 73.780 28.070 ;
        RECT 75.680 28.060 76.020 28.200 ;
        RECT 81.310 28.060 81.490 28.070 ;
        RECT 83.390 28.060 83.730 28.200 ;
        RECT 89.020 28.060 89.200 28.070 ;
        RECT 91.100 28.060 91.440 28.200 ;
        RECT 96.730 28.060 96.910 28.070 ;
        RECT 98.810 28.060 99.150 28.200 ;
        RECT 104.440 28.060 104.620 28.070 ;
        RECT 106.520 28.060 106.860 28.200 ;
        RECT 112.150 28.060 112.330 28.070 ;
        RECT 114.230 28.060 114.570 28.200 ;
        RECT 119.860 28.060 120.040 28.070 ;
        RECT 121.940 28.060 122.280 28.200 ;
        RECT 4.210 27.680 4.570 28.060 ;
        RECT 6.290 27.450 6.430 28.060 ;
        RECT 11.920 27.680 12.280 28.060 ;
        RECT 14.000 27.450 14.140 28.060 ;
        RECT 19.630 27.680 19.990 28.060 ;
        RECT 21.710 27.450 21.850 28.060 ;
        RECT 27.340 27.680 27.700 28.060 ;
        RECT 29.420 27.450 29.560 28.060 ;
        RECT 35.050 27.680 35.410 28.060 ;
        RECT 37.130 27.450 37.270 28.060 ;
        RECT 42.760 27.680 43.120 28.060 ;
        RECT 44.840 27.450 44.980 28.060 ;
        RECT 50.470 27.680 50.830 28.060 ;
        RECT 52.550 27.450 52.690 28.060 ;
        RECT 58.180 27.680 58.540 28.060 ;
        RECT 60.260 27.450 60.400 28.060 ;
        RECT 65.890 27.680 66.250 28.060 ;
        RECT 67.970 27.450 68.110 28.060 ;
        RECT 73.600 27.680 73.960 28.060 ;
        RECT 75.680 27.450 75.820 28.060 ;
        RECT 81.310 27.680 81.670 28.060 ;
        RECT 83.390 27.450 83.530 28.060 ;
        RECT 89.020 27.680 89.380 28.060 ;
        RECT 91.100 27.450 91.240 28.060 ;
        RECT 96.730 27.680 97.090 28.060 ;
        RECT 98.810 27.450 98.950 28.060 ;
        RECT 104.440 27.680 104.800 28.060 ;
        RECT 106.520 27.450 106.660 28.060 ;
        RECT 112.150 27.680 112.510 28.060 ;
        RECT 114.230 27.450 114.370 28.060 ;
        RECT 119.860 27.680 120.220 28.060 ;
        RECT 121.940 27.450 122.080 28.060 ;
        RECT 6.100 27.130 6.430 27.450 ;
        RECT 13.810 27.130 14.140 27.450 ;
        RECT 21.520 27.130 21.850 27.450 ;
        RECT 29.230 27.130 29.560 27.450 ;
        RECT 36.940 27.130 37.270 27.450 ;
        RECT 44.650 27.130 44.980 27.450 ;
        RECT 52.360 27.130 52.690 27.450 ;
        RECT 60.070 27.130 60.400 27.450 ;
        RECT 67.780 27.130 68.110 27.450 ;
        RECT 75.490 27.130 75.820 27.450 ;
        RECT 83.200 27.130 83.530 27.450 ;
        RECT 90.910 27.130 91.240 27.450 ;
        RECT 98.620 27.130 98.950 27.450 ;
        RECT 106.330 27.130 106.660 27.450 ;
        RECT 114.040 27.130 114.370 27.450 ;
        RECT 121.750 27.130 122.080 27.450 ;
        RECT 0.960 6.010 1.290 6.330 ;
        RECT 8.670 6.010 9.000 6.330 ;
        RECT 16.380 6.010 16.710 6.330 ;
        RECT 24.090 6.010 24.420 6.330 ;
        RECT 31.800 6.010 32.130 6.330 ;
        RECT 39.510 6.010 39.840 6.330 ;
        RECT 47.220 6.010 47.550 6.330 ;
        RECT 54.930 6.010 55.260 6.330 ;
        RECT 62.640 6.010 62.970 6.330 ;
        RECT 70.350 6.010 70.680 6.330 ;
        RECT 78.060 6.010 78.390 6.330 ;
        RECT 85.770 6.010 86.100 6.330 ;
        RECT 93.480 6.010 93.810 6.330 ;
        RECT 101.190 6.010 101.520 6.330 ;
        RECT 108.900 6.010 109.230 6.330 ;
        RECT 116.610 6.010 116.940 6.330 ;
        RECT 0.960 5.400 1.100 6.010 ;
        RECT 2.820 5.400 3.180 5.780 ;
        RECT 8.670 5.400 8.810 6.010 ;
        RECT 10.530 5.400 10.890 5.780 ;
        RECT 16.380 5.400 16.520 6.010 ;
        RECT 18.240 5.400 18.600 5.780 ;
        RECT 24.090 5.400 24.230 6.010 ;
        RECT 25.950 5.400 26.310 5.780 ;
        RECT 31.800 5.400 31.940 6.010 ;
        RECT 33.660 5.400 34.020 5.780 ;
        RECT 39.510 5.400 39.650 6.010 ;
        RECT 41.370 5.400 41.730 5.780 ;
        RECT 47.220 5.400 47.360 6.010 ;
        RECT 49.080 5.400 49.440 5.780 ;
        RECT 54.930 5.400 55.070 6.010 ;
        RECT 56.790 5.400 57.150 5.780 ;
        RECT 62.640 5.400 62.780 6.010 ;
        RECT 64.500 5.400 64.860 5.780 ;
        RECT 70.350 5.400 70.490 6.010 ;
        RECT 72.210 5.400 72.570 5.780 ;
        RECT 78.060 5.400 78.200 6.010 ;
        RECT 79.920 5.400 80.280 5.780 ;
        RECT 85.770 5.400 85.910 6.010 ;
        RECT 87.630 5.400 87.990 5.780 ;
        RECT 93.480 5.400 93.620 6.010 ;
        RECT 95.340 5.400 95.700 5.780 ;
        RECT 101.190 5.400 101.330 6.010 ;
        RECT 103.050 5.400 103.410 5.780 ;
        RECT 108.900 5.400 109.040 6.010 ;
        RECT 110.760 5.400 111.120 5.780 ;
        RECT 116.610 5.400 116.750 6.010 ;
        RECT 118.470 5.400 118.830 5.780 ;
        RECT 0.760 5.260 1.100 5.400 ;
        RECT 3.000 5.390 3.180 5.400 ;
        RECT 8.470 5.260 8.810 5.400 ;
        RECT 10.710 5.390 10.890 5.400 ;
        RECT 16.180 5.260 16.520 5.400 ;
        RECT 18.420 5.390 18.600 5.400 ;
        RECT 23.890 5.260 24.230 5.400 ;
        RECT 26.130 5.390 26.310 5.400 ;
        RECT 31.600 5.260 31.940 5.400 ;
        RECT 33.840 5.390 34.020 5.400 ;
        RECT 39.310 5.260 39.650 5.400 ;
        RECT 41.550 5.390 41.730 5.400 ;
        RECT 47.020 5.260 47.360 5.400 ;
        RECT 49.260 5.390 49.440 5.400 ;
        RECT 54.730 5.260 55.070 5.400 ;
        RECT 56.970 5.390 57.150 5.400 ;
        RECT 62.440 5.260 62.780 5.400 ;
        RECT 64.680 5.390 64.860 5.400 ;
        RECT 70.150 5.260 70.490 5.400 ;
        RECT 72.390 5.390 72.570 5.400 ;
        RECT 77.860 5.260 78.200 5.400 ;
        RECT 80.100 5.390 80.280 5.400 ;
        RECT 85.570 5.260 85.910 5.400 ;
        RECT 87.810 5.390 87.990 5.400 ;
        RECT 93.280 5.260 93.620 5.400 ;
        RECT 95.520 5.390 95.700 5.400 ;
        RECT 100.990 5.260 101.330 5.400 ;
        RECT 103.230 5.390 103.410 5.400 ;
        RECT 108.700 5.260 109.040 5.400 ;
        RECT 110.940 5.390 111.120 5.400 ;
        RECT 116.410 5.260 116.750 5.400 ;
        RECT 118.650 5.390 118.830 5.400 ;
        RECT 0.760 2.340 0.900 5.260 ;
        RECT 8.470 2.340 8.610 5.260 ;
        RECT 16.180 2.340 16.320 5.260 ;
        RECT 23.890 2.340 24.030 5.260 ;
        RECT 31.600 2.340 31.740 5.260 ;
        RECT 39.310 2.340 39.450 5.260 ;
        RECT 47.020 2.340 47.160 5.260 ;
        RECT 54.730 2.340 54.870 5.260 ;
        RECT 62.440 2.340 62.580 5.260 ;
        RECT 70.150 2.340 70.290 5.260 ;
        RECT 77.860 2.340 78.000 5.260 ;
        RECT 85.570 2.340 85.710 5.260 ;
        RECT 93.280 2.340 93.420 5.260 ;
        RECT 100.990 2.340 101.130 5.260 ;
        RECT 108.700 2.340 108.840 5.260 ;
        RECT 116.410 2.340 116.550 5.260 ;
        RECT 0.760 1.930 1.080 2.340 ;
        RECT 8.470 1.930 8.790 2.340 ;
        RECT 16.180 1.930 16.500 2.340 ;
        RECT 23.890 1.930 24.210 2.340 ;
        RECT 31.600 1.930 31.920 2.340 ;
        RECT 39.310 1.930 39.630 2.340 ;
        RECT 47.020 1.930 47.340 2.340 ;
        RECT 54.730 1.930 55.050 2.340 ;
        RECT 62.440 1.930 62.760 2.340 ;
        RECT 70.150 1.930 70.470 2.340 ;
        RECT 77.860 1.930 78.180 2.340 ;
        RECT 85.570 1.930 85.890 2.340 ;
        RECT 93.280 1.930 93.600 2.340 ;
        RECT 100.990 1.930 101.310 2.340 ;
        RECT 108.700 1.930 109.020 2.340 ;
        RECT 116.410 1.930 116.730 2.340 ;
    END
  END VSS
  PIN OUT
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 125.425 16.370 125.695 17.275 ;
        RECT 125.515 15.570 125.695 16.370 ;
        RECT 125.435 15.065 125.695 15.570 ;
    END
  END OUT
  PIN C9
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 60.520 29.995 60.850 30.235 ;
      LAYER mcon ;
        RECT 60.630 30.040 60.810 30.220 ;
      LAYER met1 ;
        RECT 60.570 29.990 61.150 30.270 ;
        RECT 60.780 29.910 61.150 29.990 ;
      LAYER via ;
        RECT 60.800 29.950 61.060 30.210 ;
      LAYER met2 ;
        RECT 61.010 30.270 61.150 33.340 ;
        RECT 60.780 29.910 61.150 30.270 ;
    END
  END C9
  PIN C10
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 52.810 29.995 53.140 30.235 ;
      LAYER mcon ;
        RECT 52.910 30.040 53.120 30.210 ;
      LAYER met1 ;
        RECT 53.250 30.260 53.590 30.270 ;
        RECT 52.830 30.010 53.590 30.260 ;
        RECT 53.250 29.950 53.590 30.010 ;
      LAYER via ;
        RECT 53.290 29.980 53.560 30.240 ;
      LAYER met2 ;
        RECT 53.370 30.270 53.590 33.350 ;
        RECT 53.250 29.950 53.590 30.270 ;
    END
  END C10
  PIN C11
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 45.100 29.995 45.430 30.235 ;
      LAYER mcon ;
        RECT 45.200 30.040 45.410 30.210 ;
      LAYER met1 ;
        RECT 45.540 30.260 45.880 30.270 ;
        RECT 45.120 30.010 45.880 30.260 ;
        RECT 45.540 29.950 45.880 30.010 ;
      LAYER via ;
        RECT 45.580 29.980 45.850 30.240 ;
      LAYER met2 ;
        RECT 45.660 30.270 45.880 33.350 ;
        RECT 45.540 29.950 45.880 30.270 ;
    END
  END C11
  PIN C12
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 37.390 29.995 37.720 30.235 ;
      LAYER mcon ;
        RECT 37.490 30.040 37.700 30.210 ;
      LAYER met1 ;
        RECT 37.830 30.260 38.170 30.270 ;
        RECT 37.410 30.010 38.170 30.260 ;
        RECT 37.830 29.950 38.170 30.010 ;
      LAYER via ;
        RECT 37.870 29.980 38.140 30.240 ;
      LAYER met2 ;
        RECT 37.950 30.270 38.170 33.350 ;
        RECT 37.830 29.950 38.170 30.270 ;
    END
  END C12
  PIN C13
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 29.680 29.995 30.010 30.235 ;
      LAYER mcon ;
        RECT 29.780 30.040 29.990 30.210 ;
      LAYER met1 ;
        RECT 30.120 30.260 30.460 30.270 ;
        RECT 29.700 30.010 30.460 30.260 ;
        RECT 30.120 29.950 30.460 30.010 ;
      LAYER via ;
        RECT 30.160 29.980 30.430 30.240 ;
      LAYER met2 ;
        RECT 30.240 30.270 30.460 33.350 ;
        RECT 30.120 29.950 30.460 30.270 ;
    END
  END C13
  PIN C14
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 21.970 29.995 22.300 30.235 ;
      LAYER mcon ;
        RECT 22.070 30.040 22.280 30.210 ;
      LAYER met1 ;
        RECT 22.410 30.260 22.750 30.270 ;
        RECT 21.990 30.010 22.750 30.260 ;
        RECT 22.410 29.950 22.750 30.010 ;
      LAYER via ;
        RECT 22.450 29.980 22.720 30.240 ;
      LAYER met2 ;
        RECT 22.530 30.270 22.750 33.350 ;
        RECT 22.410 29.950 22.750 30.270 ;
    END
  END C14
  PIN C15
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 14.260 29.995 14.590 30.235 ;
      LAYER mcon ;
        RECT 14.360 30.040 14.570 30.210 ;
      LAYER met1 ;
        RECT 14.700 30.260 15.040 30.270 ;
        RECT 14.280 30.010 15.040 30.260 ;
        RECT 14.700 29.950 15.040 30.010 ;
      LAYER via ;
        RECT 14.740 29.980 15.010 30.240 ;
      LAYER met2 ;
        RECT 14.820 30.270 15.040 33.350 ;
        RECT 14.700 29.950 15.040 30.270 ;
    END
  END C15
  PIN C16
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 6.550 29.995 6.880 30.235 ;
      LAYER mcon ;
        RECT 6.650 30.040 6.860 30.210 ;
      LAYER met1 ;
        RECT 6.990 30.260 7.330 30.270 ;
        RECT 6.570 30.010 7.330 30.260 ;
        RECT 6.990 29.950 7.330 30.010 ;
      LAYER via ;
        RECT 7.030 29.980 7.300 30.240 ;
      LAYER met2 ;
        RECT 7.110 30.270 7.330 33.350 ;
        RECT 6.990 29.950 7.330 30.270 ;
    END
  END C16
  PIN C17
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.510 3.225 0.840 3.465 ;
      LAYER mcon ;
        RECT 0.530 3.250 0.740 3.420 ;
      LAYER met1 ;
        RECT 0.060 3.450 0.400 3.510 ;
        RECT 0.060 3.200 0.820 3.450 ;
        RECT 0.060 3.190 0.400 3.200 ;
      LAYER via ;
        RECT 0.090 3.220 0.360 3.480 ;
      LAYER met2 ;
        RECT 0.060 3.190 0.400 3.510 ;
        RECT 0.060 0.110 0.280 3.190 ;
    END
  END C17
  PIN C18
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 8.220 3.225 8.550 3.465 ;
      LAYER mcon ;
        RECT 8.240 3.250 8.450 3.420 ;
      LAYER met1 ;
        RECT 7.770 3.450 8.110 3.510 ;
        RECT 7.770 3.200 8.530 3.450 ;
        RECT 7.770 3.190 8.110 3.200 ;
      LAYER via ;
        RECT 7.800 3.220 8.070 3.480 ;
      LAYER met2 ;
        RECT 7.770 3.190 8.110 3.510 ;
        RECT 7.770 0.110 7.990 3.190 ;
    END
  END C18
  PIN C19
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 15.930 3.225 16.260 3.465 ;
      LAYER mcon ;
        RECT 15.950 3.250 16.160 3.420 ;
      LAYER met1 ;
        RECT 15.480 3.450 15.820 3.510 ;
        RECT 15.480 3.200 16.240 3.450 ;
        RECT 15.480 3.190 15.820 3.200 ;
      LAYER via ;
        RECT 15.510 3.220 15.780 3.480 ;
      LAYER met2 ;
        RECT 15.480 3.190 15.820 3.510 ;
        RECT 15.480 0.110 15.700 3.190 ;
    END
  END C19
  PIN C20
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 23.640 3.225 23.970 3.465 ;
      LAYER mcon ;
        RECT 23.660 3.250 23.870 3.420 ;
      LAYER met1 ;
        RECT 23.190 3.450 23.530 3.510 ;
        RECT 23.190 3.200 23.950 3.450 ;
        RECT 23.190 3.190 23.530 3.200 ;
      LAYER via ;
        RECT 23.220 3.220 23.490 3.480 ;
      LAYER met2 ;
        RECT 23.190 3.190 23.530 3.510 ;
        RECT 23.190 0.110 23.410 3.190 ;
    END
  END C20
  PIN C21
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 31.350 3.225 31.680 3.465 ;
      LAYER mcon ;
        RECT 31.370 3.250 31.580 3.420 ;
      LAYER met1 ;
        RECT 30.900 3.450 31.240 3.510 ;
        RECT 30.900 3.200 31.660 3.450 ;
        RECT 30.900 3.190 31.240 3.200 ;
      LAYER via ;
        RECT 30.930 3.220 31.200 3.480 ;
      LAYER met2 ;
        RECT 30.900 3.190 31.240 3.510 ;
        RECT 30.900 0.110 31.120 3.190 ;
    END
  END C21
  PIN C22
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 39.060 3.225 39.390 3.465 ;
      LAYER mcon ;
        RECT 39.080 3.250 39.290 3.420 ;
      LAYER met1 ;
        RECT 38.610 3.450 38.950 3.510 ;
        RECT 38.610 3.200 39.370 3.450 ;
        RECT 38.610 3.190 38.950 3.200 ;
      LAYER via ;
        RECT 38.640 3.220 38.910 3.480 ;
      LAYER met2 ;
        RECT 38.610 3.190 38.950 3.510 ;
        RECT 38.610 0.110 38.830 3.190 ;
    END
  END C22
  PIN C23
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 46.770 3.225 47.100 3.465 ;
      LAYER mcon ;
        RECT 46.790 3.250 47.000 3.420 ;
      LAYER met1 ;
        RECT 46.320 3.450 46.660 3.510 ;
        RECT 46.320 3.200 47.080 3.450 ;
        RECT 46.320 3.190 46.660 3.200 ;
      LAYER via ;
        RECT 46.350 3.220 46.620 3.480 ;
      LAYER met2 ;
        RECT 46.320 3.190 46.660 3.510 ;
        RECT 46.320 0.110 46.540 3.190 ;
    END
  END C23
  PIN C24
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 54.480 3.225 54.810 3.465 ;
      LAYER mcon ;
        RECT 54.520 3.240 54.700 3.420 ;
      LAYER met1 ;
        RECT 54.180 3.470 54.550 3.550 ;
        RECT 54.180 3.190 54.760 3.470 ;
      LAYER via ;
        RECT 54.270 3.250 54.530 3.510 ;
      LAYER met2 ;
        RECT 54.180 3.190 54.550 3.550 ;
        RECT 54.180 0.120 54.320 3.190 ;
    END
  END C24
  PIN C25
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 62.190 3.225 62.520 3.465 ;
      LAYER mcon ;
        RECT 62.230 3.240 62.410 3.420 ;
      LAYER met1 ;
        RECT 61.890 3.470 62.260 3.550 ;
        RECT 61.890 3.190 62.470 3.470 ;
      LAYER via ;
        RECT 61.980 3.250 62.240 3.510 ;
      LAYER met2 ;
        RECT 61.890 3.190 62.260 3.550 ;
        RECT 61.890 0.120 62.030 3.190 ;
    END
  END C25
  PIN C26
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 69.900 3.225 70.230 3.465 ;
      LAYER mcon ;
        RECT 69.920 3.250 70.130 3.420 ;
      LAYER met1 ;
        RECT 69.450 3.450 69.790 3.510 ;
        RECT 69.450 3.200 70.210 3.450 ;
        RECT 69.450 3.190 69.790 3.200 ;
      LAYER via ;
        RECT 69.480 3.220 69.750 3.480 ;
      LAYER met2 ;
        RECT 69.450 3.190 69.790 3.510 ;
        RECT 69.450 0.110 69.670 3.190 ;
    END
  END C26
  PIN C27
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 77.610 3.225 77.940 3.465 ;
      LAYER mcon ;
        RECT 77.630 3.250 77.840 3.420 ;
      LAYER met1 ;
        RECT 77.160 3.450 77.500 3.510 ;
        RECT 77.160 3.200 77.920 3.450 ;
        RECT 77.160 3.190 77.500 3.200 ;
      LAYER via ;
        RECT 77.190 3.220 77.460 3.480 ;
      LAYER met2 ;
        RECT 77.160 3.190 77.500 3.510 ;
        RECT 77.160 0.110 77.380 3.190 ;
    END
  END C27
  PIN C28
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 85.320 3.225 85.650 3.465 ;
      LAYER mcon ;
        RECT 85.340 3.250 85.550 3.420 ;
      LAYER met1 ;
        RECT 84.870 3.450 85.210 3.510 ;
        RECT 84.870 3.200 85.630 3.450 ;
        RECT 84.870 3.190 85.210 3.200 ;
      LAYER via ;
        RECT 84.900 3.220 85.170 3.480 ;
      LAYER met2 ;
        RECT 84.870 3.190 85.210 3.510 ;
        RECT 84.870 0.110 85.090 3.190 ;
    END
  END C28
  PIN C29
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 93.030 3.225 93.360 3.465 ;
      LAYER mcon ;
        RECT 93.050 3.250 93.260 3.420 ;
      LAYER met1 ;
        RECT 92.580 3.450 92.920 3.510 ;
        RECT 92.580 3.200 93.340 3.450 ;
        RECT 92.580 3.190 92.920 3.200 ;
      LAYER via ;
        RECT 92.610 3.220 92.880 3.480 ;
      LAYER met2 ;
        RECT 92.580 3.190 92.920 3.510 ;
        RECT 92.580 0.110 92.800 3.190 ;
    END
  END C29
  PIN C30
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 100.740 3.225 101.070 3.465 ;
      LAYER mcon ;
        RECT 100.760 3.250 100.970 3.420 ;
      LAYER met1 ;
        RECT 100.290 3.450 100.630 3.510 ;
        RECT 100.290 3.200 101.050 3.450 ;
        RECT 100.290 3.190 100.630 3.200 ;
      LAYER via ;
        RECT 100.320 3.220 100.590 3.480 ;
      LAYER met2 ;
        RECT 100.290 3.190 100.630 3.510 ;
        RECT 100.290 0.110 100.510 3.190 ;
    END
  END C30
  PIN C31
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 108.450 3.225 108.780 3.465 ;
      LAYER mcon ;
        RECT 108.470 3.250 108.680 3.420 ;
      LAYER met1 ;
        RECT 108.000 3.450 108.340 3.510 ;
        RECT 108.000 3.200 108.760 3.450 ;
        RECT 108.000 3.190 108.340 3.200 ;
      LAYER via ;
        RECT 108.030 3.220 108.300 3.480 ;
      LAYER met2 ;
        RECT 108.000 3.190 108.340 3.510 ;
        RECT 108.000 0.110 108.220 3.190 ;
    END
  END C31
  PIN C32
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 116.160 3.225 116.490 3.465 ;
      LAYER mcon ;
        RECT 116.180 3.250 116.390 3.420 ;
      LAYER met1 ;
        RECT 115.710 3.450 116.050 3.510 ;
        RECT 115.710 3.200 116.470 3.450 ;
        RECT 115.710 3.190 116.050 3.200 ;
      LAYER via ;
        RECT 115.740 3.220 116.010 3.480 ;
      LAYER met2 ;
        RECT 115.710 3.190 116.050 3.510 ;
        RECT 115.710 0.110 115.930 3.190 ;
    END
  END C32
  PIN C1
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 122.200 29.995 122.530 30.235 ;
      LAYER mcon ;
        RECT 122.300 30.040 122.510 30.210 ;
      LAYER met1 ;
        RECT 122.640 30.260 122.980 30.270 ;
        RECT 122.220 30.010 122.980 30.260 ;
        RECT 122.640 29.950 122.980 30.010 ;
      LAYER via ;
        RECT 122.680 29.980 122.950 30.240 ;
      LAYER met2 ;
        RECT 122.760 30.270 122.980 33.350 ;
        RECT 122.640 29.950 122.980 30.270 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 114.490 29.995 114.820 30.235 ;
      LAYER mcon ;
        RECT 114.590 30.040 114.800 30.210 ;
      LAYER met1 ;
        RECT 114.930 30.260 115.270 30.270 ;
        RECT 114.510 30.010 115.270 30.260 ;
        RECT 114.930 29.950 115.270 30.010 ;
      LAYER via ;
        RECT 114.970 29.980 115.240 30.240 ;
      LAYER met2 ;
        RECT 115.050 30.270 115.270 33.350 ;
        RECT 114.930 29.950 115.270 30.270 ;
    END
  END C2
  PIN C3
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 106.780 29.995 107.110 30.235 ;
      LAYER mcon ;
        RECT 106.880 30.040 107.090 30.210 ;
      LAYER met1 ;
        RECT 107.220 30.260 107.560 30.270 ;
        RECT 106.800 30.010 107.560 30.260 ;
        RECT 107.220 29.950 107.560 30.010 ;
      LAYER via ;
        RECT 107.260 29.980 107.530 30.240 ;
      LAYER met2 ;
        RECT 107.340 30.270 107.560 33.350 ;
        RECT 107.220 29.950 107.560 30.270 ;
    END
  END C3
  PIN C4
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 99.070 29.995 99.400 30.235 ;
      LAYER mcon ;
        RECT 99.170 30.040 99.380 30.210 ;
      LAYER met1 ;
        RECT 99.510 30.260 99.850 30.270 ;
        RECT 99.090 30.010 99.850 30.260 ;
        RECT 99.510 29.950 99.850 30.010 ;
      LAYER via ;
        RECT 99.550 29.980 99.820 30.240 ;
      LAYER met2 ;
        RECT 99.630 30.270 99.850 33.350 ;
        RECT 99.510 29.950 99.850 30.270 ;
    END
  END C4
  PIN C5
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 91.360 29.995 91.690 30.235 ;
      LAYER mcon ;
        RECT 91.460 30.040 91.670 30.210 ;
      LAYER met1 ;
        RECT 91.800 30.260 92.140 30.270 ;
        RECT 91.380 30.010 92.140 30.260 ;
        RECT 91.800 29.950 92.140 30.010 ;
      LAYER via ;
        RECT 91.840 29.980 92.110 30.240 ;
      LAYER met2 ;
        RECT 91.920 30.270 92.140 33.350 ;
        RECT 91.800 29.950 92.140 30.270 ;
    END
  END C5
  PIN C6
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 83.650 29.995 83.980 30.235 ;
      LAYER mcon ;
        RECT 83.750 30.040 83.960 30.210 ;
      LAYER met1 ;
        RECT 84.090 30.260 84.430 30.270 ;
        RECT 83.670 30.010 84.430 30.260 ;
        RECT 84.090 29.950 84.430 30.010 ;
      LAYER via ;
        RECT 84.130 29.980 84.400 30.240 ;
      LAYER met2 ;
        RECT 84.210 30.270 84.430 33.350 ;
        RECT 84.090 29.950 84.430 30.270 ;
    END
  END C6
  PIN C7
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 75.940 29.995 76.270 30.235 ;
      LAYER mcon ;
        RECT 76.040 30.040 76.250 30.210 ;
      LAYER met1 ;
        RECT 76.380 30.260 76.720 30.270 ;
        RECT 75.960 30.010 76.720 30.260 ;
        RECT 76.380 29.950 76.720 30.010 ;
      LAYER via ;
        RECT 76.420 29.980 76.690 30.240 ;
      LAYER met2 ;
        RECT 76.500 30.270 76.720 33.350 ;
        RECT 76.380 29.950 76.720 30.270 ;
    END
  END C7
  PIN C8
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 68.230 29.995 68.560 30.235 ;
      LAYER mcon ;
        RECT 68.340 30.040 68.520 30.220 ;
      LAYER met1 ;
        RECT 68.280 29.990 68.860 30.270 ;
        RECT 68.490 29.910 68.860 29.990 ;
      LAYER via ;
        RECT 68.510 29.950 68.770 30.210 ;
      LAYER met2 ;
        RECT 68.720 30.270 68.860 33.340 ;
        RECT 68.490 29.910 68.860 30.270 ;
    END
  END C8
  PIN RESET
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 55.770 16.455 56.100 16.695 ;
    END
  END RESET
  OBS
      LAYER pwell ;
        RECT 0.935 31.215 1.105 31.385 ;
        RECT 6.885 31.225 7.055 31.395 ;
        RECT 0.935 31.195 1.040 31.215 ;
        RECT 6.885 31.205 6.990 31.225 ;
        RECT 0.110 30.285 1.040 31.195 ;
        RECT 6.060 30.295 6.990 31.205 ;
        RECT 8.645 31.215 8.815 31.385 ;
        RECT 14.595 31.225 14.765 31.395 ;
        RECT 8.645 31.195 8.750 31.215 ;
        RECT 14.595 31.205 14.700 31.225 ;
        RECT 7.820 30.285 8.750 31.195 ;
        RECT 13.770 30.295 14.700 31.205 ;
        RECT 16.355 31.215 16.525 31.385 ;
        RECT 22.305 31.225 22.475 31.395 ;
        RECT 16.355 31.195 16.460 31.215 ;
        RECT 22.305 31.205 22.410 31.225 ;
        RECT 15.530 30.285 16.460 31.195 ;
        RECT 21.480 30.295 22.410 31.205 ;
        RECT 24.065 31.215 24.235 31.385 ;
        RECT 30.015 31.225 30.185 31.395 ;
        RECT 24.065 31.195 24.170 31.215 ;
        RECT 30.015 31.205 30.120 31.225 ;
        RECT 23.240 30.285 24.170 31.195 ;
        RECT 29.190 30.295 30.120 31.205 ;
        RECT 31.775 31.215 31.945 31.385 ;
        RECT 37.725 31.225 37.895 31.395 ;
        RECT 31.775 31.195 31.880 31.215 ;
        RECT 37.725 31.205 37.830 31.225 ;
        RECT 30.950 30.285 31.880 31.195 ;
        RECT 36.900 30.295 37.830 31.205 ;
        RECT 39.485 31.215 39.655 31.385 ;
        RECT 45.435 31.225 45.605 31.395 ;
        RECT 39.485 31.195 39.590 31.215 ;
        RECT 45.435 31.205 45.540 31.225 ;
        RECT 38.660 30.285 39.590 31.195 ;
        RECT 44.610 30.295 45.540 31.205 ;
        RECT 47.195 31.215 47.365 31.385 ;
        RECT 53.145 31.225 53.315 31.395 ;
        RECT 47.195 31.195 47.300 31.215 ;
        RECT 53.145 31.205 53.250 31.225 ;
        RECT 46.370 30.285 47.300 31.195 ;
        RECT 52.320 30.295 53.250 31.205 ;
        RECT 54.905 31.215 55.075 31.385 ;
        RECT 60.855 31.225 61.025 31.395 ;
        RECT 54.905 31.195 55.010 31.215 ;
        RECT 60.855 31.205 60.960 31.225 ;
        RECT 54.080 30.285 55.010 31.195 ;
        RECT 60.030 30.295 60.960 31.205 ;
        RECT 62.615 31.215 62.785 31.385 ;
        RECT 68.565 31.225 68.735 31.395 ;
        RECT 62.615 31.195 62.720 31.215 ;
        RECT 68.565 31.205 68.670 31.225 ;
        RECT 61.790 30.285 62.720 31.195 ;
        RECT 67.740 30.295 68.670 31.205 ;
        RECT 70.325 31.215 70.495 31.385 ;
        RECT 76.275 31.225 76.445 31.395 ;
        RECT 70.325 31.195 70.430 31.215 ;
        RECT 76.275 31.205 76.380 31.225 ;
        RECT 69.500 30.285 70.430 31.195 ;
        RECT 75.450 30.295 76.380 31.205 ;
        RECT 78.035 31.215 78.205 31.385 ;
        RECT 83.985 31.225 84.155 31.395 ;
        RECT 78.035 31.195 78.140 31.215 ;
        RECT 83.985 31.205 84.090 31.225 ;
        RECT 77.210 30.285 78.140 31.195 ;
        RECT 83.160 30.295 84.090 31.205 ;
        RECT 85.745 31.215 85.915 31.385 ;
        RECT 91.695 31.225 91.865 31.395 ;
        RECT 85.745 31.195 85.850 31.215 ;
        RECT 91.695 31.205 91.800 31.225 ;
        RECT 84.920 30.285 85.850 31.195 ;
        RECT 90.870 30.295 91.800 31.205 ;
        RECT 93.455 31.215 93.625 31.385 ;
        RECT 99.405 31.225 99.575 31.395 ;
        RECT 93.455 31.195 93.560 31.215 ;
        RECT 99.405 31.205 99.510 31.225 ;
        RECT 92.630 30.285 93.560 31.195 ;
        RECT 98.580 30.295 99.510 31.205 ;
        RECT 101.165 31.215 101.335 31.385 ;
        RECT 107.115 31.225 107.285 31.395 ;
        RECT 101.165 31.195 101.270 31.215 ;
        RECT 107.115 31.205 107.220 31.225 ;
        RECT 100.340 30.285 101.270 31.195 ;
        RECT 106.290 30.295 107.220 31.205 ;
        RECT 108.875 31.215 109.045 31.385 ;
        RECT 114.825 31.225 114.995 31.395 ;
        RECT 108.875 31.195 108.980 31.215 ;
        RECT 114.825 31.205 114.930 31.225 ;
        RECT 108.050 30.285 108.980 31.195 ;
        RECT 114.000 30.295 114.930 31.205 ;
        RECT 116.585 31.215 116.755 31.385 ;
        RECT 122.535 31.225 122.705 31.395 ;
        RECT 116.585 31.195 116.690 31.215 ;
        RECT 122.535 31.205 122.640 31.225 ;
        RECT 115.760 30.285 116.690 31.195 ;
        RECT 121.710 30.295 122.640 31.205 ;
        RECT 1.950 25.965 2.120 26.155 ;
        RECT 6.020 25.965 6.190 26.155 ;
        RECT 9.660 25.965 9.830 26.155 ;
        RECT 13.730 25.965 13.900 26.155 ;
        RECT 17.370 25.965 17.540 26.155 ;
        RECT 21.440 25.965 21.610 26.155 ;
        RECT 25.080 25.965 25.250 26.155 ;
        RECT 29.150 25.965 29.320 26.155 ;
        RECT 32.790 25.965 32.960 26.155 ;
        RECT 36.860 25.965 37.030 26.155 ;
        RECT 40.500 25.965 40.670 26.155 ;
        RECT 44.570 25.965 44.740 26.155 ;
        RECT 48.210 25.965 48.380 26.155 ;
        RECT 52.280 25.965 52.450 26.155 ;
        RECT 55.920 25.965 56.090 26.155 ;
        RECT 59.990 25.965 60.160 26.155 ;
        RECT 63.630 25.965 63.800 26.155 ;
        RECT 67.700 25.965 67.870 26.155 ;
        RECT 71.340 25.965 71.510 26.155 ;
        RECT 75.410 25.965 75.580 26.155 ;
        RECT 79.050 25.965 79.220 26.155 ;
        RECT 83.120 25.965 83.290 26.155 ;
        RECT 86.760 25.965 86.930 26.155 ;
        RECT 90.830 25.965 91.000 26.155 ;
        RECT 94.470 25.965 94.640 26.155 ;
        RECT 98.540 25.965 98.710 26.155 ;
        RECT 102.180 25.965 102.350 26.155 ;
        RECT 106.250 25.965 106.420 26.155 ;
        RECT 109.890 25.965 110.060 26.155 ;
        RECT 113.960 25.965 114.130 26.155 ;
        RECT 117.600 25.965 117.770 26.155 ;
        RECT 121.670 25.965 121.840 26.155 ;
        RECT 0.915 25.055 2.265 25.965 ;
        RECT 4.985 25.055 6.335 25.965 ;
        RECT 8.625 25.055 9.975 25.965 ;
        RECT 12.695 25.055 14.045 25.965 ;
        RECT 16.335 25.055 17.685 25.965 ;
        RECT 20.405 25.055 21.755 25.965 ;
        RECT 24.045 25.055 25.395 25.965 ;
        RECT 28.115 25.055 29.465 25.965 ;
        RECT 31.755 25.055 33.105 25.965 ;
        RECT 35.825 25.055 37.175 25.965 ;
        RECT 39.465 25.055 40.815 25.965 ;
        RECT 43.535 25.055 44.885 25.965 ;
        RECT 47.175 25.055 48.525 25.965 ;
        RECT 51.245 25.055 52.595 25.965 ;
        RECT 54.885 25.055 56.235 25.965 ;
        RECT 58.955 25.055 60.305 25.965 ;
        RECT 62.595 25.055 63.945 25.965 ;
        RECT 66.665 25.055 68.015 25.965 ;
        RECT 70.305 25.055 71.655 25.965 ;
        RECT 74.375 25.055 75.725 25.965 ;
        RECT 78.015 25.055 79.365 25.965 ;
        RECT 82.085 25.055 83.435 25.965 ;
        RECT 85.725 25.055 87.075 25.965 ;
        RECT 89.795 25.055 91.145 25.965 ;
        RECT 93.435 25.055 94.785 25.965 ;
        RECT 97.505 25.055 98.855 25.965 ;
        RECT 101.145 25.055 102.495 25.965 ;
        RECT 105.215 25.055 106.565 25.965 ;
        RECT 108.855 25.055 110.205 25.965 ;
        RECT 112.925 25.055 114.275 25.965 ;
        RECT 116.565 25.055 117.915 25.965 ;
        RECT 120.635 25.055 121.985 25.965 ;
        RECT 84.005 21.845 84.175 22.035 ;
        RECT 55.555 21.095 55.725 21.265 ;
        RECT 55.580 21.075 55.725 21.095 ;
        RECT 55.580 20.165 59.450 21.075 ;
        RECT 83.930 20.935 91.160 21.845 ;
        RECT 55.660 15.485 56.590 16.395 ;
        RECT 55.660 15.465 55.765 15.485 ;
        RECT 57.165 15.475 59.355 16.385 ;
        RECT 55.595 15.295 55.765 15.465 ;
        RECT 57.255 15.285 57.425 15.475 ;
        RECT 55.535 14.885 55.705 15.055 ;
        RECT 124.405 14.915 125.775 15.695 ;
        RECT 55.560 14.865 55.705 14.885 ;
        RECT 55.560 13.955 59.430 14.865 ;
        RECT 124.555 14.725 124.725 14.915 ;
        RECT 22.400 11.055 29.630 11.965 ;
        RECT 22.475 10.865 22.645 11.055 ;
        RECT 84.060 11.025 91.290 11.935 ;
        RECT 84.135 10.835 84.305 11.025 ;
        RECT 1.055 7.495 2.405 8.405 ;
        RECT 5.125 7.495 6.475 8.405 ;
        RECT 8.765 7.495 10.115 8.405 ;
        RECT 12.835 7.495 14.185 8.405 ;
        RECT 16.475 7.495 17.825 8.405 ;
        RECT 20.545 7.495 21.895 8.405 ;
        RECT 24.185 7.495 25.535 8.405 ;
        RECT 28.255 7.495 29.605 8.405 ;
        RECT 31.895 7.495 33.245 8.405 ;
        RECT 35.965 7.495 37.315 8.405 ;
        RECT 39.605 7.495 40.955 8.405 ;
        RECT 43.675 7.495 45.025 8.405 ;
        RECT 47.315 7.495 48.665 8.405 ;
        RECT 51.385 7.495 52.735 8.405 ;
        RECT 55.025 7.495 56.375 8.405 ;
        RECT 59.095 7.495 60.445 8.405 ;
        RECT 62.735 7.495 64.085 8.405 ;
        RECT 66.805 7.495 68.155 8.405 ;
        RECT 70.445 7.495 71.795 8.405 ;
        RECT 74.515 7.495 75.865 8.405 ;
        RECT 78.155 7.495 79.505 8.405 ;
        RECT 82.225 7.495 83.575 8.405 ;
        RECT 85.865 7.495 87.215 8.405 ;
        RECT 89.935 7.495 91.285 8.405 ;
        RECT 93.575 7.495 94.925 8.405 ;
        RECT 97.645 7.495 98.995 8.405 ;
        RECT 101.285 7.495 102.635 8.405 ;
        RECT 105.355 7.495 106.705 8.405 ;
        RECT 108.995 7.495 110.345 8.405 ;
        RECT 113.065 7.495 114.415 8.405 ;
        RECT 116.705 7.495 118.055 8.405 ;
        RECT 120.775 7.495 122.125 8.405 ;
        RECT 1.200 7.305 1.370 7.495 ;
        RECT 5.270 7.305 5.440 7.495 ;
        RECT 8.910 7.305 9.080 7.495 ;
        RECT 12.980 7.305 13.150 7.495 ;
        RECT 16.620 7.305 16.790 7.495 ;
        RECT 20.690 7.305 20.860 7.495 ;
        RECT 24.330 7.305 24.500 7.495 ;
        RECT 28.400 7.305 28.570 7.495 ;
        RECT 32.040 7.305 32.210 7.495 ;
        RECT 36.110 7.305 36.280 7.495 ;
        RECT 39.750 7.305 39.920 7.495 ;
        RECT 43.820 7.305 43.990 7.495 ;
        RECT 47.460 7.305 47.630 7.495 ;
        RECT 51.530 7.305 51.700 7.495 ;
        RECT 55.170 7.305 55.340 7.495 ;
        RECT 59.240 7.305 59.410 7.495 ;
        RECT 62.880 7.305 63.050 7.495 ;
        RECT 66.950 7.305 67.120 7.495 ;
        RECT 70.590 7.305 70.760 7.495 ;
        RECT 74.660 7.305 74.830 7.495 ;
        RECT 78.300 7.305 78.470 7.495 ;
        RECT 82.370 7.305 82.540 7.495 ;
        RECT 86.010 7.305 86.180 7.495 ;
        RECT 90.080 7.305 90.250 7.495 ;
        RECT 93.720 7.305 93.890 7.495 ;
        RECT 97.790 7.305 97.960 7.495 ;
        RECT 101.430 7.305 101.600 7.495 ;
        RECT 105.500 7.305 105.670 7.495 ;
        RECT 109.140 7.305 109.310 7.495 ;
        RECT 113.210 7.305 113.380 7.495 ;
        RECT 116.850 7.305 117.020 7.495 ;
        RECT 120.920 7.305 121.090 7.495 ;
        RECT 0.400 2.255 1.330 3.165 ;
        RECT 6.350 2.265 7.280 3.175 ;
        RECT 0.400 2.235 0.505 2.255 ;
        RECT 6.350 2.245 6.455 2.265 ;
        RECT 0.335 2.065 0.505 2.235 ;
        RECT 6.285 2.075 6.455 2.245 ;
        RECT 8.110 2.255 9.040 3.165 ;
        RECT 14.060 2.265 14.990 3.175 ;
        RECT 8.110 2.235 8.215 2.255 ;
        RECT 14.060 2.245 14.165 2.265 ;
        RECT 8.045 2.065 8.215 2.235 ;
        RECT 13.995 2.075 14.165 2.245 ;
        RECT 15.820 2.255 16.750 3.165 ;
        RECT 21.770 2.265 22.700 3.175 ;
        RECT 15.820 2.235 15.925 2.255 ;
        RECT 21.770 2.245 21.875 2.265 ;
        RECT 15.755 2.065 15.925 2.235 ;
        RECT 21.705 2.075 21.875 2.245 ;
        RECT 23.530 2.255 24.460 3.165 ;
        RECT 29.480 2.265 30.410 3.175 ;
        RECT 23.530 2.235 23.635 2.255 ;
        RECT 29.480 2.245 29.585 2.265 ;
        RECT 23.465 2.065 23.635 2.235 ;
        RECT 29.415 2.075 29.585 2.245 ;
        RECT 31.240 2.255 32.170 3.165 ;
        RECT 37.190 2.265 38.120 3.175 ;
        RECT 31.240 2.235 31.345 2.255 ;
        RECT 37.190 2.245 37.295 2.265 ;
        RECT 31.175 2.065 31.345 2.235 ;
        RECT 37.125 2.075 37.295 2.245 ;
        RECT 38.950 2.255 39.880 3.165 ;
        RECT 44.900 2.265 45.830 3.175 ;
        RECT 38.950 2.235 39.055 2.255 ;
        RECT 44.900 2.245 45.005 2.265 ;
        RECT 38.885 2.065 39.055 2.235 ;
        RECT 44.835 2.075 45.005 2.245 ;
        RECT 46.660 2.255 47.590 3.165 ;
        RECT 52.610 2.265 53.540 3.175 ;
        RECT 46.660 2.235 46.765 2.255 ;
        RECT 52.610 2.245 52.715 2.265 ;
        RECT 46.595 2.065 46.765 2.235 ;
        RECT 52.545 2.075 52.715 2.245 ;
        RECT 54.370 2.255 55.300 3.165 ;
        RECT 60.320 2.265 61.250 3.175 ;
        RECT 54.370 2.235 54.475 2.255 ;
        RECT 60.320 2.245 60.425 2.265 ;
        RECT 54.305 2.065 54.475 2.235 ;
        RECT 60.255 2.075 60.425 2.245 ;
        RECT 62.080 2.255 63.010 3.165 ;
        RECT 68.030 2.265 68.960 3.175 ;
        RECT 62.080 2.235 62.185 2.255 ;
        RECT 68.030 2.245 68.135 2.265 ;
        RECT 62.015 2.065 62.185 2.235 ;
        RECT 67.965 2.075 68.135 2.245 ;
        RECT 69.790 2.255 70.720 3.165 ;
        RECT 75.740 2.265 76.670 3.175 ;
        RECT 69.790 2.235 69.895 2.255 ;
        RECT 75.740 2.245 75.845 2.265 ;
        RECT 69.725 2.065 69.895 2.235 ;
        RECT 75.675 2.075 75.845 2.245 ;
        RECT 77.500 2.255 78.430 3.165 ;
        RECT 83.450 2.265 84.380 3.175 ;
        RECT 77.500 2.235 77.605 2.255 ;
        RECT 83.450 2.245 83.555 2.265 ;
        RECT 77.435 2.065 77.605 2.235 ;
        RECT 83.385 2.075 83.555 2.245 ;
        RECT 85.210 2.255 86.140 3.165 ;
        RECT 91.160 2.265 92.090 3.175 ;
        RECT 85.210 2.235 85.315 2.255 ;
        RECT 91.160 2.245 91.265 2.265 ;
        RECT 85.145 2.065 85.315 2.235 ;
        RECT 91.095 2.075 91.265 2.245 ;
        RECT 92.920 2.255 93.850 3.165 ;
        RECT 98.870 2.265 99.800 3.175 ;
        RECT 92.920 2.235 93.025 2.255 ;
        RECT 98.870 2.245 98.975 2.265 ;
        RECT 92.855 2.065 93.025 2.235 ;
        RECT 98.805 2.075 98.975 2.245 ;
        RECT 100.630 2.255 101.560 3.165 ;
        RECT 106.580 2.265 107.510 3.175 ;
        RECT 100.630 2.235 100.735 2.255 ;
        RECT 106.580 2.245 106.685 2.265 ;
        RECT 100.565 2.065 100.735 2.235 ;
        RECT 106.515 2.075 106.685 2.245 ;
        RECT 108.340 2.255 109.270 3.165 ;
        RECT 114.290 2.265 115.220 3.175 ;
        RECT 108.340 2.235 108.445 2.255 ;
        RECT 114.290 2.245 114.395 2.265 ;
        RECT 108.275 2.065 108.445 2.235 ;
        RECT 114.225 2.075 114.395 2.245 ;
        RECT 116.050 2.255 116.980 3.165 ;
        RECT 122.000 2.265 122.930 3.175 ;
        RECT 116.050 2.235 116.155 2.255 ;
        RECT 122.000 2.245 122.105 2.265 ;
        RECT 115.985 2.065 116.155 2.235 ;
        RECT 121.935 2.075 122.105 2.245 ;
      LAYER li1 ;
        RECT 3.840 32.530 4.170 32.700 ;
        RECT 11.550 32.530 11.880 32.700 ;
        RECT 19.260 32.530 19.590 32.700 ;
        RECT 26.970 32.530 27.300 32.700 ;
        RECT 34.680 32.530 35.010 32.700 ;
        RECT 42.390 32.530 42.720 32.700 ;
        RECT 50.100 32.530 50.430 32.700 ;
        RECT 57.810 32.530 58.140 32.700 ;
        RECT 65.520 32.530 65.850 32.700 ;
        RECT 73.230 32.530 73.560 32.700 ;
        RECT 80.940 32.530 81.270 32.700 ;
        RECT 88.650 32.530 88.980 32.700 ;
        RECT 96.360 32.530 96.690 32.700 ;
        RECT 104.070 32.530 104.400 32.700 ;
        RECT 111.780 32.530 112.110 32.700 ;
        RECT 119.490 32.530 119.820 32.700 ;
        RECT 3.200 31.670 3.370 32.360 ;
        RECT 3.680 31.670 3.850 32.360 ;
        RECT 4.160 31.670 4.330 32.360 ;
        RECT 10.910 31.670 11.080 32.360 ;
        RECT 11.390 31.670 11.560 32.360 ;
        RECT 11.870 31.670 12.040 32.360 ;
        RECT 18.620 31.670 18.790 32.360 ;
        RECT 19.100 31.670 19.270 32.360 ;
        RECT 19.580 31.670 19.750 32.360 ;
        RECT 26.330 31.670 26.500 32.360 ;
        RECT 26.810 31.670 26.980 32.360 ;
        RECT 27.290 31.670 27.460 32.360 ;
        RECT 34.040 31.670 34.210 32.360 ;
        RECT 34.520 31.670 34.690 32.360 ;
        RECT 35.000 31.670 35.170 32.360 ;
        RECT 41.750 31.670 41.920 32.360 ;
        RECT 42.230 31.670 42.400 32.360 ;
        RECT 42.710 31.670 42.880 32.360 ;
        RECT 49.460 31.670 49.630 32.360 ;
        RECT 49.940 31.670 50.110 32.360 ;
        RECT 50.420 31.670 50.590 32.360 ;
        RECT 57.170 31.670 57.340 32.360 ;
        RECT 57.650 31.670 57.820 32.360 ;
        RECT 58.130 31.670 58.300 32.360 ;
        RECT 64.880 31.670 65.050 32.360 ;
        RECT 65.360 31.670 65.530 32.360 ;
        RECT 65.840 31.670 66.010 32.360 ;
        RECT 72.590 31.670 72.760 32.360 ;
        RECT 73.070 31.670 73.240 32.360 ;
        RECT 73.550 31.670 73.720 32.360 ;
        RECT 80.300 31.670 80.470 32.360 ;
        RECT 80.780 31.670 80.950 32.360 ;
        RECT 81.260 31.670 81.430 32.360 ;
        RECT 88.010 31.670 88.180 32.360 ;
        RECT 88.490 31.670 88.660 32.360 ;
        RECT 88.970 31.670 89.140 32.360 ;
        RECT 95.720 31.670 95.890 32.360 ;
        RECT 96.200 31.670 96.370 32.360 ;
        RECT 96.680 31.670 96.850 32.360 ;
        RECT 103.430 31.670 103.600 32.360 ;
        RECT 103.910 31.670 104.080 32.360 ;
        RECT 104.390 31.670 104.560 32.360 ;
        RECT 111.140 31.670 111.310 32.360 ;
        RECT 111.620 31.670 111.790 32.360 ;
        RECT 112.100 31.670 112.270 32.360 ;
        RECT 118.850 31.670 119.020 32.360 ;
        RECT 119.330 31.670 119.500 32.360 ;
        RECT 119.810 31.670 119.980 32.360 ;
        RECT 0.200 30.415 0.530 31.045 ;
        RECT 2.050 30.700 2.290 31.370 ;
        RECT 3.360 31.330 3.690 31.500 ;
        RECT 3.920 31.090 4.250 31.095 ;
        RECT 3.920 30.930 4.980 31.090 ;
        RECT 6.150 30.930 6.480 31.055 ;
        RECT 3.920 30.910 6.480 30.930 ;
        RECT 4.800 30.750 6.480 30.910 ;
        RECT 3.280 30.700 3.450 30.710 ;
        RECT 2.050 30.530 3.450 30.700 ;
        RECT 0.200 29.815 0.430 30.415 ;
        RECT 1.790 30.290 2.120 30.295 ;
        RECT 0.600 30.190 0.930 30.225 ;
        RECT 1.190 30.190 2.120 30.290 ;
        RECT 0.600 30.120 2.120 30.190 ;
        RECT 0.600 30.020 1.380 30.120 ;
        RECT 1.790 30.110 2.120 30.120 ;
        RECT 0.600 29.985 0.930 30.020 ;
        RECT 0.200 28.835 0.530 29.815 ;
        RECT 1.650 29.070 1.820 29.910 ;
        RECT 3.280 29.670 3.450 30.530 ;
        RECT 3.760 29.670 3.930 30.710 ;
        RECT 4.240 29.670 4.410 30.710 ;
        RECT 6.150 30.425 6.480 30.750 ;
        RECT 5.020 30.125 5.350 30.295 ;
        RECT 3.440 29.285 3.770 29.455 ;
        RECT 1.450 28.870 1.830 29.070 ;
        RECT 5.320 28.870 5.490 29.910 ;
        RECT 6.150 29.825 6.380 30.425 ;
        RECT 7.910 30.415 8.240 31.045 ;
        RECT 9.760 30.700 10.000 31.370 ;
        RECT 11.070 31.330 11.400 31.500 ;
        RECT 11.630 31.090 11.960 31.095 ;
        RECT 11.630 30.930 12.690 31.090 ;
        RECT 13.860 30.930 14.190 31.055 ;
        RECT 11.630 30.910 14.190 30.930 ;
        RECT 12.510 30.750 14.190 30.910 ;
        RECT 10.990 30.700 11.160 30.710 ;
        RECT 9.760 30.530 11.160 30.700 ;
        RECT 1.450 27.080 1.620 28.870 ;
        RECT 6.150 28.845 6.480 29.825 ;
        RECT 7.910 29.815 8.140 30.415 ;
        RECT 9.500 30.290 9.830 30.295 ;
        RECT 8.310 30.190 8.640 30.225 ;
        RECT 8.900 30.190 9.830 30.290 ;
        RECT 8.310 30.120 9.830 30.190 ;
        RECT 8.310 30.020 9.090 30.120 ;
        RECT 9.500 30.110 9.830 30.120 ;
        RECT 8.310 29.985 8.640 30.020 ;
        RECT 7.910 28.835 8.240 29.815 ;
        RECT 9.360 29.070 9.530 29.910 ;
        RECT 10.990 29.670 11.160 30.530 ;
        RECT 11.470 29.670 11.640 30.710 ;
        RECT 11.950 29.670 12.120 30.710 ;
        RECT 13.860 30.425 14.190 30.750 ;
        RECT 12.730 30.125 13.060 30.295 ;
        RECT 11.150 29.285 11.480 29.455 ;
        RECT 9.160 28.870 9.540 29.070 ;
        RECT 13.030 28.870 13.200 29.910 ;
        RECT 13.860 29.825 14.090 30.425 ;
        RECT 15.620 30.415 15.950 31.045 ;
        RECT 17.470 30.700 17.710 31.370 ;
        RECT 18.780 31.330 19.110 31.500 ;
        RECT 19.340 31.090 19.670 31.095 ;
        RECT 19.340 30.930 20.400 31.090 ;
        RECT 21.570 30.930 21.900 31.055 ;
        RECT 19.340 30.910 21.900 30.930 ;
        RECT 20.220 30.750 21.900 30.910 ;
        RECT 18.700 30.700 18.870 30.710 ;
        RECT 17.470 30.530 18.870 30.700 ;
        RECT 1.790 28.485 2.120 28.655 ;
        RECT 5.020 28.485 5.350 28.655 ;
        RECT 3.830 27.250 4.160 27.420 ;
        RECT 9.160 27.080 9.330 28.870 ;
        RECT 13.860 28.845 14.190 29.825 ;
        RECT 15.620 29.815 15.850 30.415 ;
        RECT 17.210 30.290 17.540 30.295 ;
        RECT 16.020 30.190 16.350 30.225 ;
        RECT 16.610 30.190 17.540 30.290 ;
        RECT 16.020 30.120 17.540 30.190 ;
        RECT 16.020 30.020 16.800 30.120 ;
        RECT 17.210 30.110 17.540 30.120 ;
        RECT 16.020 29.985 16.350 30.020 ;
        RECT 15.620 28.835 15.950 29.815 ;
        RECT 17.070 29.070 17.240 29.910 ;
        RECT 18.700 29.670 18.870 30.530 ;
        RECT 19.180 29.670 19.350 30.710 ;
        RECT 19.660 29.670 19.830 30.710 ;
        RECT 21.570 30.425 21.900 30.750 ;
        RECT 20.440 30.125 20.770 30.295 ;
        RECT 18.860 29.285 19.190 29.455 ;
        RECT 16.870 28.870 17.250 29.070 ;
        RECT 20.740 28.870 20.910 29.910 ;
        RECT 21.570 29.825 21.800 30.425 ;
        RECT 23.330 30.415 23.660 31.045 ;
        RECT 25.180 30.700 25.420 31.370 ;
        RECT 26.490 31.330 26.820 31.500 ;
        RECT 27.050 31.090 27.380 31.095 ;
        RECT 27.050 30.930 28.110 31.090 ;
        RECT 29.280 30.930 29.610 31.055 ;
        RECT 27.050 30.910 29.610 30.930 ;
        RECT 27.930 30.750 29.610 30.910 ;
        RECT 26.410 30.700 26.580 30.710 ;
        RECT 25.180 30.530 26.580 30.700 ;
        RECT 9.500 28.485 9.830 28.655 ;
        RECT 12.730 28.485 13.060 28.655 ;
        RECT 11.540 27.250 11.870 27.420 ;
        RECT 16.870 27.080 17.040 28.870 ;
        RECT 21.570 28.845 21.900 29.825 ;
        RECT 23.330 29.815 23.560 30.415 ;
        RECT 24.920 30.290 25.250 30.295 ;
        RECT 23.730 30.190 24.060 30.225 ;
        RECT 24.320 30.190 25.250 30.290 ;
        RECT 23.730 30.120 25.250 30.190 ;
        RECT 23.730 30.020 24.510 30.120 ;
        RECT 24.920 30.110 25.250 30.120 ;
        RECT 23.730 29.985 24.060 30.020 ;
        RECT 23.330 28.835 23.660 29.815 ;
        RECT 24.780 29.070 24.950 29.910 ;
        RECT 26.410 29.670 26.580 30.530 ;
        RECT 26.890 29.670 27.060 30.710 ;
        RECT 27.370 29.670 27.540 30.710 ;
        RECT 29.280 30.425 29.610 30.750 ;
        RECT 28.150 30.125 28.480 30.295 ;
        RECT 26.570 29.285 26.900 29.455 ;
        RECT 24.580 28.870 24.960 29.070 ;
        RECT 28.450 28.870 28.620 29.910 ;
        RECT 29.280 29.825 29.510 30.425 ;
        RECT 31.040 30.415 31.370 31.045 ;
        RECT 32.890 30.700 33.130 31.370 ;
        RECT 34.200 31.330 34.530 31.500 ;
        RECT 34.760 31.090 35.090 31.095 ;
        RECT 34.760 30.930 35.820 31.090 ;
        RECT 36.990 30.930 37.320 31.055 ;
        RECT 34.760 30.910 37.320 30.930 ;
        RECT 35.640 30.750 37.320 30.910 ;
        RECT 34.120 30.700 34.290 30.710 ;
        RECT 32.890 30.530 34.290 30.700 ;
        RECT 17.210 28.485 17.540 28.655 ;
        RECT 20.440 28.485 20.770 28.655 ;
        RECT 19.250 27.250 19.580 27.420 ;
        RECT 24.580 27.080 24.750 28.870 ;
        RECT 29.280 28.845 29.610 29.825 ;
        RECT 31.040 29.815 31.270 30.415 ;
        RECT 32.630 30.290 32.960 30.295 ;
        RECT 31.440 30.190 31.770 30.225 ;
        RECT 32.030 30.190 32.960 30.290 ;
        RECT 31.440 30.120 32.960 30.190 ;
        RECT 31.440 30.020 32.220 30.120 ;
        RECT 32.630 30.110 32.960 30.120 ;
        RECT 31.440 29.985 31.770 30.020 ;
        RECT 31.040 28.835 31.370 29.815 ;
        RECT 32.490 29.070 32.660 29.910 ;
        RECT 34.120 29.670 34.290 30.530 ;
        RECT 34.600 29.670 34.770 30.710 ;
        RECT 35.080 29.670 35.250 30.710 ;
        RECT 36.990 30.425 37.320 30.750 ;
        RECT 35.860 30.125 36.190 30.295 ;
        RECT 34.280 29.285 34.610 29.455 ;
        RECT 32.290 28.870 32.670 29.070 ;
        RECT 36.160 28.870 36.330 29.910 ;
        RECT 36.990 29.825 37.220 30.425 ;
        RECT 38.750 30.415 39.080 31.045 ;
        RECT 40.600 30.700 40.840 31.370 ;
        RECT 41.910 31.330 42.240 31.500 ;
        RECT 42.470 31.090 42.800 31.095 ;
        RECT 42.470 30.930 43.530 31.090 ;
        RECT 44.700 30.930 45.030 31.055 ;
        RECT 42.470 30.910 45.030 30.930 ;
        RECT 43.350 30.750 45.030 30.910 ;
        RECT 41.830 30.700 42.000 30.710 ;
        RECT 40.600 30.530 42.000 30.700 ;
        RECT 24.920 28.485 25.250 28.655 ;
        RECT 28.150 28.485 28.480 28.655 ;
        RECT 26.960 27.250 27.290 27.420 ;
        RECT 32.290 27.080 32.460 28.870 ;
        RECT 36.990 28.845 37.320 29.825 ;
        RECT 38.750 29.815 38.980 30.415 ;
        RECT 40.340 30.290 40.670 30.295 ;
        RECT 39.150 30.190 39.480 30.225 ;
        RECT 39.740 30.190 40.670 30.290 ;
        RECT 39.150 30.120 40.670 30.190 ;
        RECT 39.150 30.020 39.930 30.120 ;
        RECT 40.340 30.110 40.670 30.120 ;
        RECT 39.150 29.985 39.480 30.020 ;
        RECT 38.750 28.835 39.080 29.815 ;
        RECT 40.200 29.070 40.370 29.910 ;
        RECT 41.830 29.670 42.000 30.530 ;
        RECT 42.310 29.670 42.480 30.710 ;
        RECT 42.790 29.670 42.960 30.710 ;
        RECT 44.700 30.425 45.030 30.750 ;
        RECT 43.570 30.125 43.900 30.295 ;
        RECT 41.990 29.285 42.320 29.455 ;
        RECT 40.000 28.870 40.380 29.070 ;
        RECT 43.870 28.870 44.040 29.910 ;
        RECT 44.700 29.825 44.930 30.425 ;
        RECT 46.460 30.415 46.790 31.045 ;
        RECT 48.310 30.700 48.550 31.370 ;
        RECT 49.620 31.330 49.950 31.500 ;
        RECT 50.180 31.090 50.510 31.095 ;
        RECT 50.180 30.930 51.240 31.090 ;
        RECT 52.410 30.930 52.740 31.055 ;
        RECT 50.180 30.910 52.740 30.930 ;
        RECT 51.060 30.750 52.740 30.910 ;
        RECT 49.540 30.700 49.710 30.710 ;
        RECT 48.310 30.530 49.710 30.700 ;
        RECT 32.630 28.485 32.960 28.655 ;
        RECT 35.860 28.485 36.190 28.655 ;
        RECT 34.670 27.250 35.000 27.420 ;
        RECT 40.000 27.080 40.170 28.870 ;
        RECT 44.700 28.845 45.030 29.825 ;
        RECT 46.460 29.815 46.690 30.415 ;
        RECT 48.050 30.290 48.380 30.295 ;
        RECT 46.860 30.190 47.190 30.225 ;
        RECT 47.450 30.190 48.380 30.290 ;
        RECT 46.860 30.120 48.380 30.190 ;
        RECT 46.860 30.020 47.640 30.120 ;
        RECT 48.050 30.110 48.380 30.120 ;
        RECT 46.860 29.985 47.190 30.020 ;
        RECT 46.460 28.835 46.790 29.815 ;
        RECT 47.910 29.070 48.080 29.910 ;
        RECT 49.540 29.670 49.710 30.530 ;
        RECT 50.020 29.670 50.190 30.710 ;
        RECT 50.500 29.670 50.670 30.710 ;
        RECT 52.410 30.425 52.740 30.750 ;
        RECT 51.280 30.125 51.610 30.295 ;
        RECT 49.700 29.285 50.030 29.455 ;
        RECT 47.710 28.870 48.090 29.070 ;
        RECT 51.580 28.870 51.750 29.910 ;
        RECT 52.410 29.825 52.640 30.425 ;
        RECT 54.170 30.415 54.500 31.045 ;
        RECT 56.020 30.700 56.260 31.370 ;
        RECT 57.330 31.330 57.660 31.500 ;
        RECT 57.890 31.090 58.220 31.095 ;
        RECT 57.890 30.930 58.950 31.090 ;
        RECT 60.120 30.930 60.450 31.055 ;
        RECT 57.890 30.910 60.450 30.930 ;
        RECT 58.770 30.750 60.450 30.910 ;
        RECT 57.250 30.700 57.420 30.710 ;
        RECT 56.020 30.530 57.420 30.700 ;
        RECT 40.340 28.485 40.670 28.655 ;
        RECT 43.570 28.485 43.900 28.655 ;
        RECT 42.380 27.250 42.710 27.420 ;
        RECT 47.710 27.080 47.880 28.870 ;
        RECT 52.410 28.845 52.740 29.825 ;
        RECT 54.170 29.815 54.400 30.415 ;
        RECT 55.760 30.290 56.090 30.295 ;
        RECT 54.570 30.190 54.900 30.225 ;
        RECT 55.160 30.190 56.090 30.290 ;
        RECT 54.570 30.120 56.090 30.190 ;
        RECT 54.570 30.020 55.350 30.120 ;
        RECT 55.760 30.110 56.090 30.120 ;
        RECT 54.570 29.985 54.900 30.020 ;
        RECT 54.170 28.835 54.500 29.815 ;
        RECT 55.620 29.070 55.790 29.910 ;
        RECT 57.250 29.670 57.420 30.530 ;
        RECT 57.730 29.670 57.900 30.710 ;
        RECT 58.210 29.670 58.380 30.710 ;
        RECT 60.120 30.425 60.450 30.750 ;
        RECT 58.990 30.125 59.320 30.295 ;
        RECT 57.410 29.285 57.740 29.455 ;
        RECT 55.420 28.870 55.800 29.070 ;
        RECT 59.290 28.870 59.460 29.910 ;
        RECT 60.120 29.825 60.350 30.425 ;
        RECT 61.880 30.415 62.210 31.045 ;
        RECT 63.730 30.700 63.970 31.370 ;
        RECT 65.040 31.330 65.370 31.500 ;
        RECT 65.600 31.090 65.930 31.095 ;
        RECT 65.600 30.930 66.660 31.090 ;
        RECT 67.830 30.930 68.160 31.055 ;
        RECT 65.600 30.910 68.160 30.930 ;
        RECT 66.480 30.750 68.160 30.910 ;
        RECT 64.960 30.700 65.130 30.710 ;
        RECT 63.730 30.530 65.130 30.700 ;
        RECT 48.050 28.485 48.380 28.655 ;
        RECT 51.280 28.485 51.610 28.655 ;
        RECT 50.090 27.250 50.420 27.420 ;
        RECT 55.420 27.080 55.590 28.870 ;
        RECT 60.120 28.845 60.450 29.825 ;
        RECT 61.880 29.815 62.110 30.415 ;
        RECT 63.470 30.290 63.800 30.295 ;
        RECT 62.280 30.190 62.610 30.225 ;
        RECT 62.870 30.190 63.800 30.290 ;
        RECT 62.280 30.120 63.800 30.190 ;
        RECT 62.280 30.020 63.060 30.120 ;
        RECT 63.470 30.110 63.800 30.120 ;
        RECT 62.280 29.985 62.610 30.020 ;
        RECT 61.880 28.835 62.210 29.815 ;
        RECT 63.330 29.070 63.500 29.910 ;
        RECT 64.960 29.670 65.130 30.530 ;
        RECT 65.440 29.670 65.610 30.710 ;
        RECT 65.920 29.670 66.090 30.710 ;
        RECT 67.830 30.425 68.160 30.750 ;
        RECT 66.700 30.125 67.030 30.295 ;
        RECT 65.120 29.285 65.450 29.455 ;
        RECT 63.130 28.870 63.510 29.070 ;
        RECT 67.000 28.870 67.170 29.910 ;
        RECT 67.830 29.825 68.060 30.425 ;
        RECT 69.590 30.415 69.920 31.045 ;
        RECT 71.440 30.700 71.680 31.370 ;
        RECT 72.750 31.330 73.080 31.500 ;
        RECT 73.310 31.090 73.640 31.095 ;
        RECT 73.310 30.930 74.370 31.090 ;
        RECT 75.540 30.930 75.870 31.055 ;
        RECT 73.310 30.910 75.870 30.930 ;
        RECT 74.190 30.750 75.870 30.910 ;
        RECT 72.670 30.700 72.840 30.710 ;
        RECT 71.440 30.530 72.840 30.700 ;
        RECT 55.760 28.485 56.090 28.655 ;
        RECT 58.990 28.485 59.320 28.655 ;
        RECT 57.800 27.250 58.130 27.420 ;
        RECT 63.130 27.080 63.300 28.870 ;
        RECT 67.830 28.845 68.160 29.825 ;
        RECT 69.590 29.815 69.820 30.415 ;
        RECT 71.180 30.290 71.510 30.295 ;
        RECT 69.990 30.190 70.320 30.225 ;
        RECT 70.580 30.190 71.510 30.290 ;
        RECT 69.990 30.120 71.510 30.190 ;
        RECT 69.990 30.020 70.770 30.120 ;
        RECT 71.180 30.110 71.510 30.120 ;
        RECT 69.990 29.985 70.320 30.020 ;
        RECT 69.590 28.835 69.920 29.815 ;
        RECT 71.040 29.070 71.210 29.910 ;
        RECT 72.670 29.670 72.840 30.530 ;
        RECT 73.150 29.670 73.320 30.710 ;
        RECT 73.630 29.670 73.800 30.710 ;
        RECT 75.540 30.425 75.870 30.750 ;
        RECT 74.410 30.125 74.740 30.295 ;
        RECT 72.830 29.285 73.160 29.455 ;
        RECT 70.840 28.870 71.220 29.070 ;
        RECT 74.710 28.870 74.880 29.910 ;
        RECT 75.540 29.825 75.770 30.425 ;
        RECT 77.300 30.415 77.630 31.045 ;
        RECT 79.150 30.700 79.390 31.370 ;
        RECT 80.460 31.330 80.790 31.500 ;
        RECT 81.020 31.090 81.350 31.095 ;
        RECT 81.020 30.930 82.080 31.090 ;
        RECT 83.250 30.930 83.580 31.055 ;
        RECT 81.020 30.910 83.580 30.930 ;
        RECT 81.900 30.750 83.580 30.910 ;
        RECT 80.380 30.700 80.550 30.710 ;
        RECT 79.150 30.530 80.550 30.700 ;
        RECT 63.470 28.485 63.800 28.655 ;
        RECT 66.700 28.485 67.030 28.655 ;
        RECT 65.510 27.250 65.840 27.420 ;
        RECT 70.840 27.080 71.010 28.870 ;
        RECT 75.540 28.845 75.870 29.825 ;
        RECT 77.300 29.815 77.530 30.415 ;
        RECT 78.890 30.290 79.220 30.295 ;
        RECT 77.700 30.190 78.030 30.225 ;
        RECT 78.290 30.190 79.220 30.290 ;
        RECT 77.700 30.120 79.220 30.190 ;
        RECT 77.700 30.020 78.480 30.120 ;
        RECT 78.890 30.110 79.220 30.120 ;
        RECT 77.700 29.985 78.030 30.020 ;
        RECT 77.300 28.835 77.630 29.815 ;
        RECT 78.750 29.070 78.920 29.910 ;
        RECT 80.380 29.670 80.550 30.530 ;
        RECT 80.860 29.670 81.030 30.710 ;
        RECT 81.340 29.670 81.510 30.710 ;
        RECT 83.250 30.425 83.580 30.750 ;
        RECT 82.120 30.125 82.450 30.295 ;
        RECT 80.540 29.285 80.870 29.455 ;
        RECT 78.550 28.870 78.930 29.070 ;
        RECT 82.420 28.870 82.590 29.910 ;
        RECT 83.250 29.825 83.480 30.425 ;
        RECT 85.010 30.415 85.340 31.045 ;
        RECT 86.860 30.700 87.100 31.370 ;
        RECT 88.170 31.330 88.500 31.500 ;
        RECT 88.730 31.090 89.060 31.095 ;
        RECT 88.730 30.930 89.790 31.090 ;
        RECT 90.960 30.930 91.290 31.055 ;
        RECT 88.730 30.910 91.290 30.930 ;
        RECT 89.610 30.750 91.290 30.910 ;
        RECT 88.090 30.700 88.260 30.710 ;
        RECT 86.860 30.530 88.260 30.700 ;
        RECT 71.180 28.485 71.510 28.655 ;
        RECT 74.410 28.485 74.740 28.655 ;
        RECT 73.220 27.250 73.550 27.420 ;
        RECT 78.550 27.080 78.720 28.870 ;
        RECT 83.250 28.845 83.580 29.825 ;
        RECT 85.010 29.815 85.240 30.415 ;
        RECT 86.600 30.290 86.930 30.295 ;
        RECT 85.410 30.190 85.740 30.225 ;
        RECT 86.000 30.190 86.930 30.290 ;
        RECT 85.410 30.120 86.930 30.190 ;
        RECT 85.410 30.020 86.190 30.120 ;
        RECT 86.600 30.110 86.930 30.120 ;
        RECT 85.410 29.985 85.740 30.020 ;
        RECT 85.010 28.835 85.340 29.815 ;
        RECT 86.460 29.070 86.630 29.910 ;
        RECT 88.090 29.670 88.260 30.530 ;
        RECT 88.570 29.670 88.740 30.710 ;
        RECT 89.050 29.670 89.220 30.710 ;
        RECT 90.960 30.425 91.290 30.750 ;
        RECT 89.830 30.125 90.160 30.295 ;
        RECT 88.250 29.285 88.580 29.455 ;
        RECT 86.260 28.870 86.640 29.070 ;
        RECT 90.130 28.870 90.300 29.910 ;
        RECT 90.960 29.825 91.190 30.425 ;
        RECT 92.720 30.415 93.050 31.045 ;
        RECT 94.570 30.700 94.810 31.370 ;
        RECT 95.880 31.330 96.210 31.500 ;
        RECT 96.440 31.090 96.770 31.095 ;
        RECT 96.440 30.930 97.500 31.090 ;
        RECT 98.670 30.930 99.000 31.055 ;
        RECT 96.440 30.910 99.000 30.930 ;
        RECT 97.320 30.750 99.000 30.910 ;
        RECT 95.800 30.700 95.970 30.710 ;
        RECT 94.570 30.530 95.970 30.700 ;
        RECT 78.890 28.485 79.220 28.655 ;
        RECT 82.120 28.485 82.450 28.655 ;
        RECT 80.930 27.250 81.260 27.420 ;
        RECT 86.260 27.080 86.430 28.870 ;
        RECT 90.960 28.845 91.290 29.825 ;
        RECT 92.720 29.815 92.950 30.415 ;
        RECT 94.310 30.290 94.640 30.295 ;
        RECT 93.120 30.190 93.450 30.225 ;
        RECT 93.710 30.190 94.640 30.290 ;
        RECT 93.120 30.120 94.640 30.190 ;
        RECT 93.120 30.020 93.900 30.120 ;
        RECT 94.310 30.110 94.640 30.120 ;
        RECT 93.120 29.985 93.450 30.020 ;
        RECT 92.720 28.835 93.050 29.815 ;
        RECT 94.170 29.070 94.340 29.910 ;
        RECT 95.800 29.670 95.970 30.530 ;
        RECT 96.280 29.670 96.450 30.710 ;
        RECT 96.760 29.670 96.930 30.710 ;
        RECT 98.670 30.425 99.000 30.750 ;
        RECT 97.540 30.125 97.870 30.295 ;
        RECT 95.960 29.285 96.290 29.455 ;
        RECT 93.970 28.870 94.350 29.070 ;
        RECT 97.840 28.870 98.010 29.910 ;
        RECT 98.670 29.825 98.900 30.425 ;
        RECT 100.430 30.415 100.760 31.045 ;
        RECT 102.280 30.700 102.520 31.370 ;
        RECT 103.590 31.330 103.920 31.500 ;
        RECT 104.150 31.090 104.480 31.095 ;
        RECT 104.150 30.930 105.210 31.090 ;
        RECT 106.380 30.930 106.710 31.055 ;
        RECT 104.150 30.910 106.710 30.930 ;
        RECT 105.030 30.750 106.710 30.910 ;
        RECT 103.510 30.700 103.680 30.710 ;
        RECT 102.280 30.530 103.680 30.700 ;
        RECT 86.600 28.485 86.930 28.655 ;
        RECT 89.830 28.485 90.160 28.655 ;
        RECT 88.640 27.250 88.970 27.420 ;
        RECT 93.970 27.080 94.140 28.870 ;
        RECT 98.670 28.845 99.000 29.825 ;
        RECT 100.430 29.815 100.660 30.415 ;
        RECT 102.020 30.290 102.350 30.295 ;
        RECT 100.830 30.190 101.160 30.225 ;
        RECT 101.420 30.190 102.350 30.290 ;
        RECT 100.830 30.120 102.350 30.190 ;
        RECT 100.830 30.020 101.610 30.120 ;
        RECT 102.020 30.110 102.350 30.120 ;
        RECT 100.830 29.985 101.160 30.020 ;
        RECT 100.430 28.835 100.760 29.815 ;
        RECT 101.880 29.070 102.050 29.910 ;
        RECT 103.510 29.670 103.680 30.530 ;
        RECT 103.990 29.670 104.160 30.710 ;
        RECT 104.470 29.670 104.640 30.710 ;
        RECT 106.380 30.425 106.710 30.750 ;
        RECT 105.250 30.125 105.580 30.295 ;
        RECT 103.670 29.285 104.000 29.455 ;
        RECT 101.680 28.870 102.060 29.070 ;
        RECT 105.550 28.870 105.720 29.910 ;
        RECT 106.380 29.825 106.610 30.425 ;
        RECT 108.140 30.415 108.470 31.045 ;
        RECT 109.990 30.700 110.230 31.370 ;
        RECT 111.300 31.330 111.630 31.500 ;
        RECT 111.860 31.090 112.190 31.095 ;
        RECT 111.860 30.930 112.920 31.090 ;
        RECT 114.090 30.930 114.420 31.055 ;
        RECT 111.860 30.910 114.420 30.930 ;
        RECT 112.740 30.750 114.420 30.910 ;
        RECT 111.220 30.700 111.390 30.710 ;
        RECT 109.990 30.530 111.390 30.700 ;
        RECT 94.310 28.485 94.640 28.655 ;
        RECT 97.540 28.485 97.870 28.655 ;
        RECT 96.350 27.250 96.680 27.420 ;
        RECT 101.680 27.080 101.850 28.870 ;
        RECT 106.380 28.845 106.710 29.825 ;
        RECT 108.140 29.815 108.370 30.415 ;
        RECT 109.730 30.290 110.060 30.295 ;
        RECT 108.540 30.190 108.870 30.225 ;
        RECT 109.130 30.190 110.060 30.290 ;
        RECT 108.540 30.120 110.060 30.190 ;
        RECT 108.540 30.020 109.320 30.120 ;
        RECT 109.730 30.110 110.060 30.120 ;
        RECT 108.540 29.985 108.870 30.020 ;
        RECT 108.140 28.835 108.470 29.815 ;
        RECT 109.590 29.070 109.760 29.910 ;
        RECT 111.220 29.670 111.390 30.530 ;
        RECT 111.700 29.670 111.870 30.710 ;
        RECT 112.180 29.670 112.350 30.710 ;
        RECT 114.090 30.425 114.420 30.750 ;
        RECT 112.960 30.125 113.290 30.295 ;
        RECT 111.380 29.285 111.710 29.455 ;
        RECT 109.390 28.870 109.770 29.070 ;
        RECT 113.260 28.870 113.430 29.910 ;
        RECT 114.090 29.825 114.320 30.425 ;
        RECT 115.850 30.415 116.180 31.045 ;
        RECT 117.700 30.700 117.940 31.370 ;
        RECT 119.010 31.330 119.340 31.500 ;
        RECT 119.570 31.090 119.900 31.095 ;
        RECT 119.570 30.930 120.630 31.090 ;
        RECT 121.800 30.930 122.130 31.055 ;
        RECT 119.570 30.910 122.130 30.930 ;
        RECT 120.450 30.750 122.130 30.910 ;
        RECT 118.930 30.700 119.100 30.710 ;
        RECT 117.700 30.530 119.100 30.700 ;
        RECT 102.020 28.485 102.350 28.655 ;
        RECT 105.250 28.485 105.580 28.655 ;
        RECT 104.060 27.250 104.390 27.420 ;
        RECT 109.390 27.080 109.560 28.870 ;
        RECT 114.090 28.845 114.420 29.825 ;
        RECT 115.850 29.815 116.080 30.415 ;
        RECT 117.440 30.290 117.770 30.295 ;
        RECT 116.250 30.190 116.580 30.225 ;
        RECT 116.840 30.190 117.770 30.290 ;
        RECT 116.250 30.120 117.770 30.190 ;
        RECT 116.250 30.020 117.030 30.120 ;
        RECT 117.440 30.110 117.770 30.120 ;
        RECT 116.250 29.985 116.580 30.020 ;
        RECT 115.850 28.835 116.180 29.815 ;
        RECT 117.300 29.070 117.470 29.910 ;
        RECT 118.930 29.670 119.100 30.530 ;
        RECT 119.410 29.670 119.580 30.710 ;
        RECT 119.890 29.670 120.060 30.710 ;
        RECT 121.800 30.425 122.130 30.750 ;
        RECT 120.670 30.125 121.000 30.295 ;
        RECT 119.090 29.285 119.420 29.455 ;
        RECT 117.100 28.870 117.480 29.070 ;
        RECT 120.970 28.870 121.140 29.910 ;
        RECT 121.800 29.825 122.030 30.425 ;
        RECT 109.730 28.485 110.060 28.655 ;
        RECT 112.960 28.485 113.290 28.655 ;
        RECT 111.770 27.250 112.100 27.420 ;
        RECT 117.100 27.080 117.270 28.870 ;
        RECT 121.800 28.845 122.130 29.825 ;
        RECT 117.440 28.485 117.770 28.655 ;
        RECT 120.670 28.485 121.000 28.655 ;
        RECT 119.480 27.250 119.810 27.420 ;
        RECT 1.450 26.880 3.360 27.080 ;
        RECT 3.190 26.390 3.360 26.880 ;
        RECT 3.670 26.390 3.840 27.080 ;
        RECT 4.150 26.390 4.320 27.080 ;
        RECT 9.160 26.880 11.070 27.080 ;
        RECT 10.900 26.390 11.070 26.880 ;
        RECT 11.380 26.390 11.550 27.080 ;
        RECT 11.860 26.390 12.030 27.080 ;
        RECT 16.870 26.880 18.780 27.080 ;
        RECT 18.610 26.390 18.780 26.880 ;
        RECT 19.090 26.390 19.260 27.080 ;
        RECT 19.570 26.390 19.740 27.080 ;
        RECT 24.580 26.880 26.490 27.080 ;
        RECT 26.320 26.390 26.490 26.880 ;
        RECT 26.800 26.390 26.970 27.080 ;
        RECT 27.280 26.390 27.450 27.080 ;
        RECT 32.290 26.880 34.200 27.080 ;
        RECT 34.030 26.390 34.200 26.880 ;
        RECT 34.510 26.390 34.680 27.080 ;
        RECT 34.990 26.390 35.160 27.080 ;
        RECT 40.000 26.880 41.910 27.080 ;
        RECT 41.740 26.390 41.910 26.880 ;
        RECT 42.220 26.390 42.390 27.080 ;
        RECT 42.700 26.390 42.870 27.080 ;
        RECT 47.710 26.880 49.620 27.080 ;
        RECT 49.450 26.390 49.620 26.880 ;
        RECT 49.930 26.390 50.100 27.080 ;
        RECT 50.410 26.390 50.580 27.080 ;
        RECT 55.420 26.880 57.330 27.080 ;
        RECT 57.160 26.390 57.330 26.880 ;
        RECT 57.640 26.390 57.810 27.080 ;
        RECT 58.120 26.390 58.290 27.080 ;
        RECT 63.130 26.880 65.040 27.080 ;
        RECT 64.870 26.390 65.040 26.880 ;
        RECT 65.350 26.390 65.520 27.080 ;
        RECT 65.830 26.390 66.000 27.080 ;
        RECT 70.840 26.880 72.750 27.080 ;
        RECT 72.580 26.390 72.750 26.880 ;
        RECT 73.060 26.390 73.230 27.080 ;
        RECT 73.540 26.390 73.710 27.080 ;
        RECT 78.550 26.880 80.460 27.080 ;
        RECT 80.290 26.390 80.460 26.880 ;
        RECT 80.770 26.390 80.940 27.080 ;
        RECT 81.250 26.390 81.420 27.080 ;
        RECT 86.260 26.880 88.170 27.080 ;
        RECT 88.000 26.390 88.170 26.880 ;
        RECT 88.480 26.390 88.650 27.080 ;
        RECT 88.960 26.390 89.130 27.080 ;
        RECT 93.970 26.880 95.880 27.080 ;
        RECT 95.710 26.390 95.880 26.880 ;
        RECT 96.190 26.390 96.360 27.080 ;
        RECT 96.670 26.390 96.840 27.080 ;
        RECT 101.680 26.880 103.590 27.080 ;
        RECT 103.420 26.390 103.590 26.880 ;
        RECT 103.900 26.390 104.070 27.080 ;
        RECT 104.380 26.390 104.550 27.080 ;
        RECT 109.390 26.880 111.300 27.080 ;
        RECT 111.130 26.390 111.300 26.880 ;
        RECT 111.610 26.390 111.780 27.080 ;
        RECT 112.090 26.390 112.260 27.080 ;
        RECT 117.100 26.880 119.010 27.080 ;
        RECT 118.840 26.390 119.010 26.880 ;
        RECT 119.320 26.390 119.490 27.080 ;
        RECT 119.800 26.390 119.970 27.080 ;
        RECT 3.350 26.050 3.680 26.220 ;
        RECT 11.060 26.050 11.390 26.220 ;
        RECT 18.770 26.050 19.100 26.220 ;
        RECT 26.480 26.050 26.810 26.220 ;
        RECT 34.190 26.050 34.520 26.220 ;
        RECT 41.900 26.050 42.230 26.220 ;
        RECT 49.610 26.050 49.940 26.220 ;
        RECT 57.320 26.050 57.650 26.220 ;
        RECT 65.030 26.050 65.360 26.220 ;
        RECT 72.740 26.050 73.070 26.220 ;
        RECT 80.450 26.050 80.780 26.220 ;
        RECT 88.160 26.050 88.490 26.220 ;
        RECT 95.870 26.050 96.200 26.220 ;
        RECT 103.580 26.050 103.910 26.220 ;
        RECT 111.290 26.050 111.620 26.220 ;
        RECT 119.000 26.050 119.330 26.220 ;
        RECT 1.425 25.175 1.755 25.815 ;
        RECT 3.910 25.645 4.240 25.815 ;
        RECT 0.975 24.745 1.325 24.995 ;
        RECT 1.495 24.575 1.665 25.175 ;
        RECT 1.835 24.990 2.185 24.995 ;
        RECT 3.270 24.990 3.440 25.430 ;
        RECT 1.835 24.820 3.440 24.990 ;
        RECT 1.835 24.745 2.185 24.820 ;
        RECT 1.495 24.405 2.175 24.575 ;
        RECT 1.845 23.620 2.175 24.405 ;
        RECT 3.270 24.390 3.440 24.820 ;
        RECT 3.750 24.390 3.920 25.430 ;
        RECT 4.230 24.390 4.400 25.430 ;
        RECT 5.495 25.175 5.825 25.815 ;
        RECT 9.135 25.175 9.465 25.815 ;
        RECT 11.620 25.645 11.950 25.815 ;
        RECT 5.045 24.745 5.395 24.995 ;
        RECT 5.565 24.575 5.735 25.175 ;
        RECT 5.905 24.745 6.255 24.995 ;
        RECT 8.685 24.745 9.035 24.995 ;
        RECT 9.205 24.575 9.375 25.175 ;
        RECT 9.545 24.990 9.895 24.995 ;
        RECT 10.980 24.990 11.150 25.430 ;
        RECT 9.545 24.820 11.150 24.990 ;
        RECT 9.545 24.745 9.895 24.820 ;
        RECT 5.565 24.405 6.245 24.575 ;
        RECT 9.205 24.405 9.885 24.575 ;
        RECT 3.430 24.005 3.760 24.175 ;
        RECT 5.915 23.620 6.245 24.405 ;
        RECT 9.555 23.620 9.885 24.405 ;
        RECT 10.980 24.390 11.150 24.820 ;
        RECT 11.460 24.390 11.630 25.430 ;
        RECT 11.940 24.390 12.110 25.430 ;
        RECT 13.205 25.175 13.535 25.815 ;
        RECT 16.845 25.175 17.175 25.815 ;
        RECT 19.330 25.645 19.660 25.815 ;
        RECT 12.755 24.745 13.105 24.995 ;
        RECT 13.275 24.575 13.445 25.175 ;
        RECT 13.615 24.745 13.965 24.995 ;
        RECT 16.395 24.745 16.745 24.995 ;
        RECT 16.915 24.575 17.085 25.175 ;
        RECT 17.255 24.990 17.605 24.995 ;
        RECT 18.690 24.990 18.860 25.430 ;
        RECT 17.255 24.820 18.860 24.990 ;
        RECT 17.255 24.745 17.605 24.820 ;
        RECT 13.275 24.405 13.955 24.575 ;
        RECT 16.915 24.405 17.595 24.575 ;
        RECT 11.140 24.005 11.470 24.175 ;
        RECT 13.625 23.620 13.955 24.405 ;
        RECT 17.265 23.620 17.595 24.405 ;
        RECT 18.690 24.390 18.860 24.820 ;
        RECT 19.170 24.390 19.340 25.430 ;
        RECT 19.650 24.390 19.820 25.430 ;
        RECT 20.915 25.175 21.245 25.815 ;
        RECT 24.555 25.175 24.885 25.815 ;
        RECT 27.040 25.645 27.370 25.815 ;
        RECT 20.465 24.745 20.815 24.995 ;
        RECT 20.985 24.575 21.155 25.175 ;
        RECT 21.325 24.745 21.675 24.995 ;
        RECT 24.105 24.745 24.455 24.995 ;
        RECT 24.625 24.575 24.795 25.175 ;
        RECT 24.965 24.990 25.315 24.995 ;
        RECT 26.400 24.990 26.570 25.430 ;
        RECT 24.965 24.820 26.570 24.990 ;
        RECT 24.965 24.745 25.315 24.820 ;
        RECT 20.985 24.405 21.665 24.575 ;
        RECT 24.625 24.405 25.305 24.575 ;
        RECT 18.850 24.005 19.180 24.175 ;
        RECT 21.335 23.620 21.665 24.405 ;
        RECT 24.975 23.620 25.305 24.405 ;
        RECT 26.400 24.390 26.570 24.820 ;
        RECT 26.880 24.390 27.050 25.430 ;
        RECT 27.360 24.390 27.530 25.430 ;
        RECT 28.625 25.175 28.955 25.815 ;
        RECT 32.265 25.175 32.595 25.815 ;
        RECT 34.750 25.645 35.080 25.815 ;
        RECT 28.175 24.745 28.525 24.995 ;
        RECT 28.695 24.575 28.865 25.175 ;
        RECT 29.035 24.745 29.385 24.995 ;
        RECT 31.815 24.745 32.165 24.995 ;
        RECT 32.335 24.575 32.505 25.175 ;
        RECT 32.675 24.990 33.025 24.995 ;
        RECT 34.110 24.990 34.280 25.430 ;
        RECT 32.675 24.820 34.280 24.990 ;
        RECT 32.675 24.745 33.025 24.820 ;
        RECT 28.695 24.405 29.375 24.575 ;
        RECT 32.335 24.405 33.015 24.575 ;
        RECT 26.560 24.005 26.890 24.175 ;
        RECT 29.045 23.620 29.375 24.405 ;
        RECT 32.685 23.620 33.015 24.405 ;
        RECT 34.110 24.390 34.280 24.820 ;
        RECT 34.590 24.390 34.760 25.430 ;
        RECT 35.070 24.390 35.240 25.430 ;
        RECT 36.335 25.175 36.665 25.815 ;
        RECT 39.975 25.175 40.305 25.815 ;
        RECT 42.460 25.645 42.790 25.815 ;
        RECT 35.885 24.745 36.235 24.995 ;
        RECT 36.405 24.575 36.575 25.175 ;
        RECT 36.745 24.745 37.095 24.995 ;
        RECT 39.525 24.745 39.875 24.995 ;
        RECT 40.045 24.575 40.215 25.175 ;
        RECT 40.385 24.990 40.735 24.995 ;
        RECT 41.820 24.990 41.990 25.430 ;
        RECT 40.385 24.820 41.990 24.990 ;
        RECT 40.385 24.745 40.735 24.820 ;
        RECT 36.405 24.405 37.085 24.575 ;
        RECT 40.045 24.405 40.725 24.575 ;
        RECT 34.270 24.005 34.600 24.175 ;
        RECT 36.755 23.620 37.085 24.405 ;
        RECT 40.395 23.620 40.725 24.405 ;
        RECT 41.820 24.390 41.990 24.820 ;
        RECT 42.300 24.390 42.470 25.430 ;
        RECT 42.780 24.390 42.950 25.430 ;
        RECT 44.045 25.175 44.375 25.815 ;
        RECT 47.685 25.175 48.015 25.815 ;
        RECT 50.170 25.645 50.500 25.815 ;
        RECT 43.595 24.745 43.945 24.995 ;
        RECT 44.115 24.575 44.285 25.175 ;
        RECT 44.455 24.745 44.805 24.995 ;
        RECT 47.235 24.745 47.585 24.995 ;
        RECT 47.755 24.575 47.925 25.175 ;
        RECT 48.095 24.990 48.445 24.995 ;
        RECT 49.530 24.990 49.700 25.430 ;
        RECT 48.095 24.820 49.700 24.990 ;
        RECT 48.095 24.745 48.445 24.820 ;
        RECT 44.115 24.405 44.795 24.575 ;
        RECT 47.755 24.405 48.435 24.575 ;
        RECT 41.980 24.005 42.310 24.175 ;
        RECT 44.465 23.620 44.795 24.405 ;
        RECT 48.105 23.620 48.435 24.405 ;
        RECT 49.530 24.390 49.700 24.820 ;
        RECT 50.010 24.390 50.180 25.430 ;
        RECT 50.490 24.390 50.660 25.430 ;
        RECT 51.755 25.175 52.085 25.815 ;
        RECT 55.395 25.175 55.725 25.815 ;
        RECT 57.880 25.645 58.210 25.815 ;
        RECT 51.305 24.745 51.655 24.995 ;
        RECT 51.825 24.575 51.995 25.175 ;
        RECT 52.165 24.745 52.515 24.995 ;
        RECT 54.945 24.745 55.295 24.995 ;
        RECT 55.465 24.575 55.635 25.175 ;
        RECT 55.805 24.990 56.155 24.995 ;
        RECT 57.240 24.990 57.410 25.430 ;
        RECT 55.805 24.820 57.410 24.990 ;
        RECT 55.805 24.745 56.155 24.820 ;
        RECT 51.825 24.405 52.505 24.575 ;
        RECT 55.465 24.405 56.145 24.575 ;
        RECT 49.690 24.005 50.020 24.175 ;
        RECT 52.175 23.620 52.505 24.405 ;
        RECT 55.815 23.620 56.145 24.405 ;
        RECT 57.240 24.390 57.410 24.820 ;
        RECT 57.720 24.390 57.890 25.430 ;
        RECT 58.200 24.390 58.370 25.430 ;
        RECT 59.465 25.175 59.795 25.815 ;
        RECT 63.105 25.175 63.435 25.815 ;
        RECT 65.590 25.645 65.920 25.815 ;
        RECT 59.015 24.745 59.365 24.995 ;
        RECT 59.535 24.575 59.705 25.175 ;
        RECT 59.875 24.745 60.225 24.995 ;
        RECT 62.655 24.745 63.005 24.995 ;
        RECT 63.175 24.575 63.345 25.175 ;
        RECT 63.515 24.990 63.865 24.995 ;
        RECT 64.950 24.990 65.120 25.430 ;
        RECT 63.515 24.820 65.120 24.990 ;
        RECT 63.515 24.745 63.865 24.820 ;
        RECT 59.535 24.405 60.215 24.575 ;
        RECT 63.175 24.405 63.855 24.575 ;
        RECT 57.400 24.005 57.730 24.175 ;
        RECT 59.885 23.620 60.215 24.405 ;
        RECT 63.525 23.620 63.855 24.405 ;
        RECT 64.950 24.390 65.120 24.820 ;
        RECT 65.430 24.390 65.600 25.430 ;
        RECT 65.910 24.390 66.080 25.430 ;
        RECT 67.175 25.175 67.505 25.815 ;
        RECT 70.815 25.175 71.145 25.815 ;
        RECT 73.300 25.645 73.630 25.815 ;
        RECT 66.725 24.745 67.075 24.995 ;
        RECT 67.245 24.575 67.415 25.175 ;
        RECT 67.585 24.745 67.935 24.995 ;
        RECT 70.365 24.745 70.715 24.995 ;
        RECT 70.885 24.575 71.055 25.175 ;
        RECT 71.225 24.990 71.575 24.995 ;
        RECT 72.660 24.990 72.830 25.430 ;
        RECT 71.225 24.820 72.830 24.990 ;
        RECT 71.225 24.745 71.575 24.820 ;
        RECT 67.245 24.405 67.925 24.575 ;
        RECT 70.885 24.405 71.565 24.575 ;
        RECT 65.110 24.005 65.440 24.175 ;
        RECT 67.595 23.620 67.925 24.405 ;
        RECT 71.235 23.620 71.565 24.405 ;
        RECT 72.660 24.390 72.830 24.820 ;
        RECT 73.140 24.390 73.310 25.430 ;
        RECT 73.620 24.390 73.790 25.430 ;
        RECT 74.885 25.175 75.215 25.815 ;
        RECT 78.525 25.175 78.855 25.815 ;
        RECT 81.010 25.645 81.340 25.815 ;
        RECT 74.435 24.745 74.785 24.995 ;
        RECT 74.955 24.575 75.125 25.175 ;
        RECT 75.295 24.745 75.645 24.995 ;
        RECT 78.075 24.745 78.425 24.995 ;
        RECT 78.595 24.575 78.765 25.175 ;
        RECT 78.935 24.990 79.285 24.995 ;
        RECT 80.370 24.990 80.540 25.430 ;
        RECT 78.935 24.820 80.540 24.990 ;
        RECT 78.935 24.745 79.285 24.820 ;
        RECT 74.955 24.405 75.635 24.575 ;
        RECT 78.595 24.405 79.275 24.575 ;
        RECT 72.820 24.005 73.150 24.175 ;
        RECT 75.305 23.620 75.635 24.405 ;
        RECT 78.945 23.620 79.275 24.405 ;
        RECT 80.370 24.390 80.540 24.820 ;
        RECT 80.850 24.390 81.020 25.430 ;
        RECT 81.330 24.390 81.500 25.430 ;
        RECT 82.595 25.175 82.925 25.815 ;
        RECT 86.235 25.175 86.565 25.815 ;
        RECT 88.720 25.645 89.050 25.815 ;
        RECT 82.145 24.745 82.495 24.995 ;
        RECT 82.665 24.575 82.835 25.175 ;
        RECT 83.005 24.745 83.355 24.995 ;
        RECT 85.785 24.745 86.135 24.995 ;
        RECT 86.305 24.575 86.475 25.175 ;
        RECT 86.645 24.990 86.995 24.995 ;
        RECT 88.080 24.990 88.250 25.430 ;
        RECT 86.645 24.820 88.250 24.990 ;
        RECT 86.645 24.745 86.995 24.820 ;
        RECT 82.665 24.405 83.345 24.575 ;
        RECT 86.305 24.405 86.985 24.575 ;
        RECT 80.530 24.005 80.860 24.175 ;
        RECT 83.015 23.620 83.345 24.405 ;
        RECT 86.655 23.620 86.985 24.405 ;
        RECT 88.080 24.390 88.250 24.820 ;
        RECT 88.560 24.390 88.730 25.430 ;
        RECT 89.040 24.390 89.210 25.430 ;
        RECT 90.305 25.175 90.635 25.815 ;
        RECT 93.945 25.175 94.275 25.815 ;
        RECT 96.430 25.645 96.760 25.815 ;
        RECT 89.855 24.745 90.205 24.995 ;
        RECT 90.375 24.575 90.545 25.175 ;
        RECT 90.715 24.745 91.065 24.995 ;
        RECT 93.495 24.745 93.845 24.995 ;
        RECT 94.015 24.575 94.185 25.175 ;
        RECT 94.355 24.990 94.705 24.995 ;
        RECT 95.790 24.990 95.960 25.430 ;
        RECT 94.355 24.820 95.960 24.990 ;
        RECT 94.355 24.745 94.705 24.820 ;
        RECT 90.375 24.405 91.055 24.575 ;
        RECT 94.015 24.405 94.695 24.575 ;
        RECT 88.240 24.005 88.570 24.175 ;
        RECT 90.725 23.620 91.055 24.405 ;
        RECT 94.365 23.620 94.695 24.405 ;
        RECT 95.790 24.390 95.960 24.820 ;
        RECT 96.270 24.390 96.440 25.430 ;
        RECT 96.750 24.390 96.920 25.430 ;
        RECT 98.015 25.175 98.345 25.815 ;
        RECT 101.655 25.175 101.985 25.815 ;
        RECT 104.140 25.645 104.470 25.815 ;
        RECT 97.565 24.745 97.915 24.995 ;
        RECT 98.085 24.575 98.255 25.175 ;
        RECT 98.425 24.745 98.775 24.995 ;
        RECT 101.205 24.745 101.555 24.995 ;
        RECT 101.725 24.575 101.895 25.175 ;
        RECT 102.065 24.990 102.415 24.995 ;
        RECT 103.500 24.990 103.670 25.430 ;
        RECT 102.065 24.820 103.670 24.990 ;
        RECT 102.065 24.745 102.415 24.820 ;
        RECT 98.085 24.405 98.765 24.575 ;
        RECT 101.725 24.405 102.405 24.575 ;
        RECT 95.950 24.005 96.280 24.175 ;
        RECT 98.435 23.620 98.765 24.405 ;
        RECT 102.075 23.620 102.405 24.405 ;
        RECT 103.500 24.390 103.670 24.820 ;
        RECT 103.980 24.390 104.150 25.430 ;
        RECT 104.460 24.390 104.630 25.430 ;
        RECT 105.725 25.175 106.055 25.815 ;
        RECT 109.365 25.175 109.695 25.815 ;
        RECT 111.850 25.645 112.180 25.815 ;
        RECT 105.275 24.745 105.625 24.995 ;
        RECT 105.795 24.575 105.965 25.175 ;
        RECT 106.135 24.745 106.485 24.995 ;
        RECT 108.915 24.745 109.265 24.995 ;
        RECT 109.435 24.575 109.605 25.175 ;
        RECT 109.775 24.990 110.125 24.995 ;
        RECT 111.210 24.990 111.380 25.430 ;
        RECT 109.775 24.820 111.380 24.990 ;
        RECT 109.775 24.745 110.125 24.820 ;
        RECT 105.795 24.405 106.475 24.575 ;
        RECT 109.435 24.405 110.115 24.575 ;
        RECT 103.660 24.005 103.990 24.175 ;
        RECT 106.145 23.620 106.475 24.405 ;
        RECT 109.785 23.620 110.115 24.405 ;
        RECT 111.210 24.390 111.380 24.820 ;
        RECT 111.690 24.390 111.860 25.430 ;
        RECT 112.170 24.390 112.340 25.430 ;
        RECT 113.435 25.175 113.765 25.815 ;
        RECT 117.075 25.175 117.405 25.815 ;
        RECT 119.560 25.645 119.890 25.815 ;
        RECT 112.985 24.745 113.335 24.995 ;
        RECT 113.505 24.575 113.675 25.175 ;
        RECT 113.845 24.745 114.195 24.995 ;
        RECT 116.625 24.745 116.975 24.995 ;
        RECT 117.145 24.575 117.315 25.175 ;
        RECT 117.485 24.990 117.835 24.995 ;
        RECT 118.920 24.990 119.090 25.430 ;
        RECT 117.485 24.820 119.090 24.990 ;
        RECT 117.485 24.745 117.835 24.820 ;
        RECT 113.505 24.405 114.185 24.575 ;
        RECT 117.145 24.405 117.825 24.575 ;
        RECT 111.370 24.005 111.700 24.175 ;
        RECT 113.855 23.620 114.185 24.405 ;
        RECT 117.495 23.620 117.825 24.405 ;
        RECT 118.920 24.390 119.090 24.820 ;
        RECT 119.400 24.390 119.570 25.430 ;
        RECT 119.880 24.390 120.050 25.430 ;
        RECT 121.145 25.175 121.475 25.815 ;
        RECT 120.695 24.745 121.045 24.995 ;
        RECT 121.215 24.575 121.385 25.175 ;
        RECT 121.555 24.745 121.905 24.995 ;
        RECT 121.215 24.405 121.895 24.575 ;
        RECT 119.080 24.005 119.410 24.175 ;
        RECT 121.565 23.620 121.895 24.405 ;
        RECT 22.780 21.205 23.110 21.665 ;
        RECT 23.620 21.205 23.950 21.665 ;
        RECT 24.460 21.205 24.790 21.665 ;
        RECT 25.300 21.205 25.630 21.665 ;
        RECT 26.140 21.205 26.470 21.665 ;
        RECT 26.980 21.205 27.310 21.665 ;
        RECT 27.820 21.205 28.150 21.665 ;
        RECT 28.660 21.205 28.990 21.665 ;
        RECT 22.780 21.015 28.990 21.205 ;
        RECT 84.440 21.235 84.770 21.695 ;
        RECT 85.280 21.235 85.610 21.695 ;
        RECT 86.120 21.235 86.450 21.695 ;
        RECT 86.960 21.235 87.290 21.695 ;
        RECT 87.800 21.235 88.130 21.695 ;
        RECT 88.640 21.235 88.970 21.695 ;
        RECT 89.480 21.235 89.810 21.695 ;
        RECT 90.320 21.235 90.650 21.695 ;
        RECT 84.440 21.045 90.650 21.235 ;
        RECT 21.490 20.850 21.835 20.910 ;
        RECT 21.490 20.845 22.700 20.850 ;
        RECT 21.490 20.610 27.725 20.845 ;
        RECT 21.490 18.535 21.835 20.610 ;
        RECT 22.285 20.605 27.725 20.610 ;
        RECT 28.660 20.425 28.990 21.015 ;
        RECT 56.090 20.465 56.420 20.925 ;
        RECT 56.930 20.465 57.260 20.925 ;
        RECT 57.770 20.465 58.100 20.925 ;
        RECT 58.610 20.465 58.940 20.925 ;
        RECT 83.160 20.875 83.950 20.880 ;
        RECT 83.160 20.870 89.385 20.875 ;
        RECT 83.140 20.640 89.385 20.870 ;
        RECT 22.780 20.255 28.990 20.425 ;
        RECT 22.780 19.455 23.110 20.255 ;
        RECT 23.620 19.455 23.950 20.255 ;
        RECT 24.460 19.455 24.790 20.255 ;
        RECT 25.300 19.455 25.630 20.255 ;
        RECT 26.140 19.455 26.470 20.255 ;
        RECT 26.980 19.455 27.310 20.255 ;
        RECT 27.820 19.455 28.150 20.255 ;
        RECT 28.660 19.455 28.990 20.255 ;
        RECT 55.495 20.280 59.465 20.465 ;
        RECT 83.140 20.280 83.460 20.640 ;
        RECT 83.945 20.635 89.385 20.640 ;
        RECT 90.320 20.455 90.650 21.045 ;
        RECT 55.495 20.275 83.460 20.280 ;
        RECT 55.495 20.245 55.840 20.275 ;
        RECT 29.920 19.900 55.840 20.245 ;
        RECT 29.920 18.535 30.265 19.900 ;
        RECT 55.495 19.685 55.840 19.900 ;
        RECT 56.090 19.855 58.945 20.105 ;
        RECT 59.145 19.960 83.460 20.275 ;
        RECT 84.440 20.285 90.650 20.455 ;
        RECT 59.145 19.685 59.465 19.960 ;
        RECT 55.495 19.515 59.465 19.685 ;
        RECT 56.090 18.715 56.420 19.515 ;
        RECT 56.930 18.715 57.260 19.515 ;
        RECT 57.770 18.715 58.100 19.515 ;
        RECT 58.610 18.715 58.940 19.515 ;
        RECT 84.440 19.485 84.770 20.285 ;
        RECT 85.280 19.485 85.610 20.285 ;
        RECT 86.120 19.485 86.450 20.285 ;
        RECT 86.960 19.485 87.290 20.285 ;
        RECT 87.800 19.485 88.130 20.285 ;
        RECT 88.640 19.485 88.970 20.285 ;
        RECT 89.480 19.485 89.810 20.285 ;
        RECT 90.320 19.485 90.650 20.285 ;
        RECT 21.490 18.190 30.265 18.535 ;
        RECT 56.170 16.865 56.500 17.845 ;
        RECT 57.675 17.035 58.005 17.835 ;
        RECT 58.515 17.055 58.845 17.835 ;
        RECT 58.515 17.035 59.280 17.055 ;
        RECT 57.675 16.865 59.280 17.035 ;
        RECT 56.270 16.670 56.500 16.865 ;
        RECT 57.215 16.670 58.845 16.695 ;
        RECT 56.270 16.460 58.845 16.670 ;
        RECT 56.270 16.265 56.500 16.460 ;
        RECT 57.215 16.445 58.845 16.460 ;
        RECT 59.015 16.275 59.280 16.865 ;
        RECT 124.565 16.515 124.745 17.275 ;
        RECT 124.565 16.345 125.240 16.515 ;
        RECT 21.640 15.645 21.985 15.670 ;
        RECT 30.540 15.645 30.885 15.660 ;
        RECT 21.630 15.300 30.885 15.645 ;
        RECT 56.170 15.635 56.500 16.265 ;
        RECT 57.675 16.095 59.280 16.275 ;
        RECT 125.070 16.200 125.240 16.345 ;
        RECT 57.675 15.625 58.005 16.095 ;
        RECT 58.515 15.625 58.845 16.095 ;
        RECT 124.505 15.795 124.845 16.165 ;
        RECT 125.070 15.870 125.345 16.200 ;
        RECT 125.070 15.615 125.240 15.870 ;
        RECT 21.640 12.260 21.985 15.300 ;
        RECT 30.540 14.045 30.885 15.300 ;
        RECT 124.575 15.445 125.240 15.615 ;
        RECT 124.575 15.065 124.745 15.445 ;
        RECT 56.070 14.255 56.400 14.715 ;
        RECT 56.910 14.255 57.240 14.715 ;
        RECT 57.750 14.255 58.080 14.715 ;
        RECT 58.590 14.255 58.920 14.715 ;
        RECT 55.475 14.065 59.445 14.255 ;
        RECT 55.475 14.045 55.820 14.065 ;
        RECT 30.540 13.700 55.820 14.045 ;
        RECT 59.125 13.990 59.445 14.065 ;
        RECT 55.475 13.475 55.820 13.700 ;
        RECT 56.070 13.645 58.925 13.895 ;
        RECT 59.125 13.670 83.480 13.990 ;
        RECT 59.125 13.475 59.445 13.670 ;
        RECT 22.910 12.615 23.240 13.415 ;
        RECT 23.750 12.615 24.080 13.415 ;
        RECT 24.590 12.615 24.920 13.415 ;
        RECT 25.430 12.615 25.760 13.415 ;
        RECT 26.270 12.615 26.600 13.415 ;
        RECT 27.110 12.615 27.440 13.415 ;
        RECT 27.950 12.615 28.280 13.415 ;
        RECT 28.790 12.615 29.120 13.415 ;
        RECT 55.475 13.305 59.445 13.475 ;
        RECT 22.910 12.445 29.120 12.615 ;
        RECT 56.070 12.505 56.400 13.305 ;
        RECT 56.910 12.505 57.240 13.305 ;
        RECT 57.750 12.505 58.080 13.305 ;
        RECT 58.590 12.505 58.920 13.305 ;
        RECT 22.415 12.260 27.855 12.265 ;
        RECT 21.640 12.030 27.855 12.260 ;
        RECT 22.415 12.025 27.855 12.030 ;
        RECT 28.790 11.855 29.120 12.445 ;
        RECT 83.160 12.230 83.480 13.670 ;
        RECT 84.570 12.585 84.900 13.385 ;
        RECT 85.410 12.585 85.740 13.385 ;
        RECT 86.250 12.585 86.580 13.385 ;
        RECT 87.090 12.585 87.420 13.385 ;
        RECT 87.930 12.585 88.260 13.385 ;
        RECT 88.770 12.585 89.100 13.385 ;
        RECT 89.610 12.585 89.940 13.385 ;
        RECT 90.450 12.585 90.780 13.385 ;
        RECT 84.570 12.415 90.780 12.585 ;
        RECT 84.075 12.230 89.515 12.235 ;
        RECT 83.160 12.020 89.515 12.230 ;
        RECT 83.170 12.000 89.515 12.020 ;
        RECT 84.075 11.995 89.515 12.000 ;
        RECT 22.910 11.665 29.120 11.855 ;
        RECT 90.450 11.825 90.780 12.415 ;
        RECT 22.910 11.205 23.240 11.665 ;
        RECT 23.750 11.205 24.080 11.665 ;
        RECT 24.590 11.205 24.920 11.665 ;
        RECT 25.430 11.205 25.760 11.665 ;
        RECT 26.270 11.205 26.600 11.665 ;
        RECT 27.110 11.205 27.440 11.665 ;
        RECT 27.950 11.205 28.280 11.665 ;
        RECT 28.790 11.205 29.120 11.665 ;
        RECT 84.570 11.635 90.780 11.825 ;
        RECT 84.570 11.175 84.900 11.635 ;
        RECT 85.410 11.175 85.740 11.635 ;
        RECT 86.250 11.175 86.580 11.635 ;
        RECT 87.090 11.175 87.420 11.635 ;
        RECT 87.930 11.175 88.260 11.635 ;
        RECT 88.770 11.175 89.100 11.635 ;
        RECT 89.610 11.175 89.940 11.635 ;
        RECT 90.450 11.175 90.780 11.635 ;
        RECT 1.145 9.055 1.475 9.840 ;
        RECT 3.630 9.285 3.960 9.455 ;
        RECT 1.145 8.885 1.825 9.055 ;
        RECT 1.135 8.465 1.485 8.715 ;
        RECT 1.655 8.285 1.825 8.885 ;
        RECT 1.995 8.465 2.345 8.715 ;
        RECT 1.565 7.645 1.895 8.285 ;
        RECT 2.990 8.030 3.160 9.070 ;
        RECT 3.470 8.030 3.640 9.070 ;
        RECT 3.950 8.640 4.120 9.070 ;
        RECT 5.215 9.055 5.545 9.840 ;
        RECT 8.855 9.055 9.185 9.840 ;
        RECT 11.340 9.285 11.670 9.455 ;
        RECT 5.215 8.885 5.895 9.055 ;
        RECT 8.855 8.885 9.535 9.055 ;
        RECT 5.205 8.640 5.555 8.715 ;
        RECT 3.950 8.470 5.555 8.640 ;
        RECT 3.950 8.030 4.120 8.470 ;
        RECT 5.205 8.465 5.555 8.470 ;
        RECT 5.725 8.285 5.895 8.885 ;
        RECT 6.065 8.465 6.415 8.715 ;
        RECT 8.845 8.465 9.195 8.715 ;
        RECT 9.365 8.285 9.535 8.885 ;
        RECT 9.705 8.465 10.055 8.715 ;
        RECT 3.150 7.645 3.480 7.815 ;
        RECT 5.635 7.645 5.965 8.285 ;
        RECT 9.275 7.645 9.605 8.285 ;
        RECT 10.700 8.030 10.870 9.070 ;
        RECT 11.180 8.030 11.350 9.070 ;
        RECT 11.660 8.640 11.830 9.070 ;
        RECT 12.925 9.055 13.255 9.840 ;
        RECT 16.565 9.055 16.895 9.840 ;
        RECT 19.050 9.285 19.380 9.455 ;
        RECT 12.925 8.885 13.605 9.055 ;
        RECT 16.565 8.885 17.245 9.055 ;
        RECT 12.915 8.640 13.265 8.715 ;
        RECT 11.660 8.470 13.265 8.640 ;
        RECT 11.660 8.030 11.830 8.470 ;
        RECT 12.915 8.465 13.265 8.470 ;
        RECT 13.435 8.285 13.605 8.885 ;
        RECT 13.775 8.465 14.125 8.715 ;
        RECT 16.555 8.465 16.905 8.715 ;
        RECT 17.075 8.285 17.245 8.885 ;
        RECT 17.415 8.465 17.765 8.715 ;
        RECT 10.860 7.645 11.190 7.815 ;
        RECT 13.345 7.645 13.675 8.285 ;
        RECT 16.985 7.645 17.315 8.285 ;
        RECT 18.410 8.030 18.580 9.070 ;
        RECT 18.890 8.030 19.060 9.070 ;
        RECT 19.370 8.640 19.540 9.070 ;
        RECT 20.635 9.055 20.965 9.840 ;
        RECT 24.275 9.055 24.605 9.840 ;
        RECT 26.760 9.285 27.090 9.455 ;
        RECT 20.635 8.885 21.315 9.055 ;
        RECT 24.275 8.885 24.955 9.055 ;
        RECT 20.625 8.640 20.975 8.715 ;
        RECT 19.370 8.470 20.975 8.640 ;
        RECT 19.370 8.030 19.540 8.470 ;
        RECT 20.625 8.465 20.975 8.470 ;
        RECT 21.145 8.285 21.315 8.885 ;
        RECT 21.485 8.465 21.835 8.715 ;
        RECT 24.265 8.465 24.615 8.715 ;
        RECT 24.785 8.285 24.955 8.885 ;
        RECT 25.125 8.465 25.475 8.715 ;
        RECT 18.570 7.645 18.900 7.815 ;
        RECT 21.055 7.645 21.385 8.285 ;
        RECT 24.695 7.645 25.025 8.285 ;
        RECT 26.120 8.030 26.290 9.070 ;
        RECT 26.600 8.030 26.770 9.070 ;
        RECT 27.080 8.640 27.250 9.070 ;
        RECT 28.345 9.055 28.675 9.840 ;
        RECT 31.985 9.055 32.315 9.840 ;
        RECT 34.470 9.285 34.800 9.455 ;
        RECT 28.345 8.885 29.025 9.055 ;
        RECT 31.985 8.885 32.665 9.055 ;
        RECT 28.335 8.640 28.685 8.715 ;
        RECT 27.080 8.470 28.685 8.640 ;
        RECT 27.080 8.030 27.250 8.470 ;
        RECT 28.335 8.465 28.685 8.470 ;
        RECT 28.855 8.285 29.025 8.885 ;
        RECT 29.195 8.465 29.545 8.715 ;
        RECT 31.975 8.465 32.325 8.715 ;
        RECT 32.495 8.285 32.665 8.885 ;
        RECT 32.835 8.465 33.185 8.715 ;
        RECT 26.280 7.645 26.610 7.815 ;
        RECT 28.765 7.645 29.095 8.285 ;
        RECT 32.405 7.645 32.735 8.285 ;
        RECT 33.830 8.030 34.000 9.070 ;
        RECT 34.310 8.030 34.480 9.070 ;
        RECT 34.790 8.640 34.960 9.070 ;
        RECT 36.055 9.055 36.385 9.840 ;
        RECT 39.695 9.055 40.025 9.840 ;
        RECT 42.180 9.285 42.510 9.455 ;
        RECT 36.055 8.885 36.735 9.055 ;
        RECT 39.695 8.885 40.375 9.055 ;
        RECT 36.045 8.640 36.395 8.715 ;
        RECT 34.790 8.470 36.395 8.640 ;
        RECT 34.790 8.030 34.960 8.470 ;
        RECT 36.045 8.465 36.395 8.470 ;
        RECT 36.565 8.285 36.735 8.885 ;
        RECT 36.905 8.465 37.255 8.715 ;
        RECT 39.685 8.465 40.035 8.715 ;
        RECT 40.205 8.285 40.375 8.885 ;
        RECT 40.545 8.465 40.895 8.715 ;
        RECT 33.990 7.645 34.320 7.815 ;
        RECT 36.475 7.645 36.805 8.285 ;
        RECT 40.115 7.645 40.445 8.285 ;
        RECT 41.540 8.030 41.710 9.070 ;
        RECT 42.020 8.030 42.190 9.070 ;
        RECT 42.500 8.640 42.670 9.070 ;
        RECT 43.765 9.055 44.095 9.840 ;
        RECT 47.405 9.055 47.735 9.840 ;
        RECT 49.890 9.285 50.220 9.455 ;
        RECT 43.765 8.885 44.445 9.055 ;
        RECT 47.405 8.885 48.085 9.055 ;
        RECT 43.755 8.640 44.105 8.715 ;
        RECT 42.500 8.470 44.105 8.640 ;
        RECT 42.500 8.030 42.670 8.470 ;
        RECT 43.755 8.465 44.105 8.470 ;
        RECT 44.275 8.285 44.445 8.885 ;
        RECT 44.615 8.465 44.965 8.715 ;
        RECT 47.395 8.465 47.745 8.715 ;
        RECT 47.915 8.285 48.085 8.885 ;
        RECT 48.255 8.465 48.605 8.715 ;
        RECT 41.700 7.645 42.030 7.815 ;
        RECT 44.185 7.645 44.515 8.285 ;
        RECT 47.825 7.645 48.155 8.285 ;
        RECT 49.250 8.030 49.420 9.070 ;
        RECT 49.730 8.030 49.900 9.070 ;
        RECT 50.210 8.640 50.380 9.070 ;
        RECT 51.475 9.055 51.805 9.840 ;
        RECT 55.115 9.055 55.445 9.840 ;
        RECT 57.600 9.285 57.930 9.455 ;
        RECT 51.475 8.885 52.155 9.055 ;
        RECT 55.115 8.885 55.795 9.055 ;
        RECT 51.465 8.640 51.815 8.715 ;
        RECT 50.210 8.470 51.815 8.640 ;
        RECT 50.210 8.030 50.380 8.470 ;
        RECT 51.465 8.465 51.815 8.470 ;
        RECT 51.985 8.285 52.155 8.885 ;
        RECT 52.325 8.465 52.675 8.715 ;
        RECT 55.105 8.465 55.455 8.715 ;
        RECT 55.625 8.285 55.795 8.885 ;
        RECT 55.965 8.465 56.315 8.715 ;
        RECT 49.410 7.645 49.740 7.815 ;
        RECT 51.895 7.645 52.225 8.285 ;
        RECT 55.535 7.645 55.865 8.285 ;
        RECT 56.960 8.030 57.130 9.070 ;
        RECT 57.440 8.030 57.610 9.070 ;
        RECT 57.920 8.640 58.090 9.070 ;
        RECT 59.185 9.055 59.515 9.840 ;
        RECT 62.825 9.055 63.155 9.840 ;
        RECT 65.310 9.285 65.640 9.455 ;
        RECT 59.185 8.885 59.865 9.055 ;
        RECT 62.825 8.885 63.505 9.055 ;
        RECT 59.175 8.640 59.525 8.715 ;
        RECT 57.920 8.470 59.525 8.640 ;
        RECT 57.920 8.030 58.090 8.470 ;
        RECT 59.175 8.465 59.525 8.470 ;
        RECT 59.695 8.285 59.865 8.885 ;
        RECT 60.035 8.465 60.385 8.715 ;
        RECT 62.815 8.465 63.165 8.715 ;
        RECT 63.335 8.285 63.505 8.885 ;
        RECT 63.675 8.465 64.025 8.715 ;
        RECT 57.120 7.645 57.450 7.815 ;
        RECT 59.605 7.645 59.935 8.285 ;
        RECT 63.245 7.645 63.575 8.285 ;
        RECT 64.670 8.030 64.840 9.070 ;
        RECT 65.150 8.030 65.320 9.070 ;
        RECT 65.630 8.640 65.800 9.070 ;
        RECT 66.895 9.055 67.225 9.840 ;
        RECT 70.535 9.055 70.865 9.840 ;
        RECT 73.020 9.285 73.350 9.455 ;
        RECT 66.895 8.885 67.575 9.055 ;
        RECT 70.535 8.885 71.215 9.055 ;
        RECT 66.885 8.640 67.235 8.715 ;
        RECT 65.630 8.470 67.235 8.640 ;
        RECT 65.630 8.030 65.800 8.470 ;
        RECT 66.885 8.465 67.235 8.470 ;
        RECT 67.405 8.285 67.575 8.885 ;
        RECT 67.745 8.465 68.095 8.715 ;
        RECT 70.525 8.465 70.875 8.715 ;
        RECT 71.045 8.285 71.215 8.885 ;
        RECT 71.385 8.465 71.735 8.715 ;
        RECT 64.830 7.645 65.160 7.815 ;
        RECT 67.315 7.645 67.645 8.285 ;
        RECT 70.955 7.645 71.285 8.285 ;
        RECT 72.380 8.030 72.550 9.070 ;
        RECT 72.860 8.030 73.030 9.070 ;
        RECT 73.340 8.640 73.510 9.070 ;
        RECT 74.605 9.055 74.935 9.840 ;
        RECT 78.245 9.055 78.575 9.840 ;
        RECT 80.730 9.285 81.060 9.455 ;
        RECT 74.605 8.885 75.285 9.055 ;
        RECT 78.245 8.885 78.925 9.055 ;
        RECT 74.595 8.640 74.945 8.715 ;
        RECT 73.340 8.470 74.945 8.640 ;
        RECT 73.340 8.030 73.510 8.470 ;
        RECT 74.595 8.465 74.945 8.470 ;
        RECT 75.115 8.285 75.285 8.885 ;
        RECT 75.455 8.465 75.805 8.715 ;
        RECT 78.235 8.465 78.585 8.715 ;
        RECT 78.755 8.285 78.925 8.885 ;
        RECT 79.095 8.465 79.445 8.715 ;
        RECT 72.540 7.645 72.870 7.815 ;
        RECT 75.025 7.645 75.355 8.285 ;
        RECT 78.665 7.645 78.995 8.285 ;
        RECT 80.090 8.030 80.260 9.070 ;
        RECT 80.570 8.030 80.740 9.070 ;
        RECT 81.050 8.640 81.220 9.070 ;
        RECT 82.315 9.055 82.645 9.840 ;
        RECT 85.955 9.055 86.285 9.840 ;
        RECT 88.440 9.285 88.770 9.455 ;
        RECT 82.315 8.885 82.995 9.055 ;
        RECT 85.955 8.885 86.635 9.055 ;
        RECT 82.305 8.640 82.655 8.715 ;
        RECT 81.050 8.470 82.655 8.640 ;
        RECT 81.050 8.030 81.220 8.470 ;
        RECT 82.305 8.465 82.655 8.470 ;
        RECT 82.825 8.285 82.995 8.885 ;
        RECT 83.165 8.465 83.515 8.715 ;
        RECT 85.945 8.465 86.295 8.715 ;
        RECT 86.465 8.285 86.635 8.885 ;
        RECT 86.805 8.465 87.155 8.715 ;
        RECT 80.250 7.645 80.580 7.815 ;
        RECT 82.735 7.645 83.065 8.285 ;
        RECT 86.375 7.645 86.705 8.285 ;
        RECT 87.800 8.030 87.970 9.070 ;
        RECT 88.280 8.030 88.450 9.070 ;
        RECT 88.760 8.640 88.930 9.070 ;
        RECT 90.025 9.055 90.355 9.840 ;
        RECT 93.665 9.055 93.995 9.840 ;
        RECT 96.150 9.285 96.480 9.455 ;
        RECT 90.025 8.885 90.705 9.055 ;
        RECT 93.665 8.885 94.345 9.055 ;
        RECT 90.015 8.640 90.365 8.715 ;
        RECT 88.760 8.470 90.365 8.640 ;
        RECT 88.760 8.030 88.930 8.470 ;
        RECT 90.015 8.465 90.365 8.470 ;
        RECT 90.535 8.285 90.705 8.885 ;
        RECT 90.875 8.465 91.225 8.715 ;
        RECT 93.655 8.465 94.005 8.715 ;
        RECT 94.175 8.285 94.345 8.885 ;
        RECT 94.515 8.465 94.865 8.715 ;
        RECT 87.960 7.645 88.290 7.815 ;
        RECT 90.445 7.645 90.775 8.285 ;
        RECT 94.085 7.645 94.415 8.285 ;
        RECT 95.510 8.030 95.680 9.070 ;
        RECT 95.990 8.030 96.160 9.070 ;
        RECT 96.470 8.640 96.640 9.070 ;
        RECT 97.735 9.055 98.065 9.840 ;
        RECT 101.375 9.055 101.705 9.840 ;
        RECT 103.860 9.285 104.190 9.455 ;
        RECT 97.735 8.885 98.415 9.055 ;
        RECT 101.375 8.885 102.055 9.055 ;
        RECT 97.725 8.640 98.075 8.715 ;
        RECT 96.470 8.470 98.075 8.640 ;
        RECT 96.470 8.030 96.640 8.470 ;
        RECT 97.725 8.465 98.075 8.470 ;
        RECT 98.245 8.285 98.415 8.885 ;
        RECT 98.585 8.465 98.935 8.715 ;
        RECT 101.365 8.465 101.715 8.715 ;
        RECT 101.885 8.285 102.055 8.885 ;
        RECT 102.225 8.465 102.575 8.715 ;
        RECT 95.670 7.645 96.000 7.815 ;
        RECT 98.155 7.645 98.485 8.285 ;
        RECT 101.795 7.645 102.125 8.285 ;
        RECT 103.220 8.030 103.390 9.070 ;
        RECT 103.700 8.030 103.870 9.070 ;
        RECT 104.180 8.640 104.350 9.070 ;
        RECT 105.445 9.055 105.775 9.840 ;
        RECT 109.085 9.055 109.415 9.840 ;
        RECT 111.570 9.285 111.900 9.455 ;
        RECT 105.445 8.885 106.125 9.055 ;
        RECT 109.085 8.885 109.765 9.055 ;
        RECT 105.435 8.640 105.785 8.715 ;
        RECT 104.180 8.470 105.785 8.640 ;
        RECT 104.180 8.030 104.350 8.470 ;
        RECT 105.435 8.465 105.785 8.470 ;
        RECT 105.955 8.285 106.125 8.885 ;
        RECT 106.295 8.465 106.645 8.715 ;
        RECT 109.075 8.465 109.425 8.715 ;
        RECT 109.595 8.285 109.765 8.885 ;
        RECT 109.935 8.465 110.285 8.715 ;
        RECT 103.380 7.645 103.710 7.815 ;
        RECT 105.865 7.645 106.195 8.285 ;
        RECT 109.505 7.645 109.835 8.285 ;
        RECT 110.930 8.030 111.100 9.070 ;
        RECT 111.410 8.030 111.580 9.070 ;
        RECT 111.890 8.640 112.060 9.070 ;
        RECT 113.155 9.055 113.485 9.840 ;
        RECT 116.795 9.055 117.125 9.840 ;
        RECT 119.280 9.285 119.610 9.455 ;
        RECT 113.155 8.885 113.835 9.055 ;
        RECT 116.795 8.885 117.475 9.055 ;
        RECT 113.145 8.640 113.495 8.715 ;
        RECT 111.890 8.470 113.495 8.640 ;
        RECT 111.890 8.030 112.060 8.470 ;
        RECT 113.145 8.465 113.495 8.470 ;
        RECT 113.665 8.285 113.835 8.885 ;
        RECT 114.005 8.465 114.355 8.715 ;
        RECT 116.785 8.465 117.135 8.715 ;
        RECT 117.305 8.285 117.475 8.885 ;
        RECT 117.645 8.465 117.995 8.715 ;
        RECT 111.090 7.645 111.420 7.815 ;
        RECT 113.575 7.645 113.905 8.285 ;
        RECT 117.215 7.645 117.545 8.285 ;
        RECT 118.640 8.030 118.810 9.070 ;
        RECT 119.120 8.030 119.290 9.070 ;
        RECT 119.600 8.640 119.770 9.070 ;
        RECT 120.865 9.055 121.195 9.840 ;
        RECT 120.865 8.885 121.545 9.055 ;
        RECT 120.855 8.640 121.205 8.715 ;
        RECT 119.600 8.470 121.205 8.640 ;
        RECT 119.600 8.030 119.770 8.470 ;
        RECT 120.855 8.465 121.205 8.470 ;
        RECT 121.375 8.285 121.545 8.885 ;
        RECT 121.715 8.465 122.065 8.715 ;
        RECT 118.800 7.645 119.130 7.815 ;
        RECT 121.285 7.645 121.615 8.285 ;
        RECT 3.710 7.240 4.040 7.410 ;
        RECT 11.420 7.240 11.750 7.410 ;
        RECT 19.130 7.240 19.460 7.410 ;
        RECT 26.840 7.240 27.170 7.410 ;
        RECT 34.550 7.240 34.880 7.410 ;
        RECT 42.260 7.240 42.590 7.410 ;
        RECT 49.970 7.240 50.300 7.410 ;
        RECT 57.680 7.240 58.010 7.410 ;
        RECT 65.390 7.240 65.720 7.410 ;
        RECT 73.100 7.240 73.430 7.410 ;
        RECT 80.810 7.240 81.140 7.410 ;
        RECT 88.520 7.240 88.850 7.410 ;
        RECT 96.230 7.240 96.560 7.410 ;
        RECT 103.940 7.240 104.270 7.410 ;
        RECT 111.650 7.240 111.980 7.410 ;
        RECT 119.360 7.240 119.690 7.410 ;
        RECT 3.070 6.380 3.240 7.070 ;
        RECT 3.550 6.380 3.720 7.070 ;
        RECT 4.030 6.580 4.200 7.070 ;
        RECT 4.030 6.380 5.940 6.580 ;
        RECT 10.780 6.380 10.950 7.070 ;
        RECT 11.260 6.380 11.430 7.070 ;
        RECT 11.740 6.580 11.910 7.070 ;
        RECT 11.740 6.380 13.650 6.580 ;
        RECT 18.490 6.380 18.660 7.070 ;
        RECT 18.970 6.380 19.140 7.070 ;
        RECT 19.450 6.580 19.620 7.070 ;
        RECT 19.450 6.380 21.360 6.580 ;
        RECT 26.200 6.380 26.370 7.070 ;
        RECT 26.680 6.380 26.850 7.070 ;
        RECT 27.160 6.580 27.330 7.070 ;
        RECT 27.160 6.380 29.070 6.580 ;
        RECT 33.910 6.380 34.080 7.070 ;
        RECT 34.390 6.380 34.560 7.070 ;
        RECT 34.870 6.580 35.040 7.070 ;
        RECT 34.870 6.380 36.780 6.580 ;
        RECT 41.620 6.380 41.790 7.070 ;
        RECT 42.100 6.380 42.270 7.070 ;
        RECT 42.580 6.580 42.750 7.070 ;
        RECT 42.580 6.380 44.490 6.580 ;
        RECT 49.330 6.380 49.500 7.070 ;
        RECT 49.810 6.380 49.980 7.070 ;
        RECT 50.290 6.580 50.460 7.070 ;
        RECT 50.290 6.380 52.200 6.580 ;
        RECT 57.040 6.380 57.210 7.070 ;
        RECT 57.520 6.380 57.690 7.070 ;
        RECT 58.000 6.580 58.170 7.070 ;
        RECT 58.000 6.380 59.910 6.580 ;
        RECT 64.750 6.380 64.920 7.070 ;
        RECT 65.230 6.380 65.400 7.070 ;
        RECT 65.710 6.580 65.880 7.070 ;
        RECT 65.710 6.380 67.620 6.580 ;
        RECT 72.460 6.380 72.630 7.070 ;
        RECT 72.940 6.380 73.110 7.070 ;
        RECT 73.420 6.580 73.590 7.070 ;
        RECT 73.420 6.380 75.330 6.580 ;
        RECT 80.170 6.380 80.340 7.070 ;
        RECT 80.650 6.380 80.820 7.070 ;
        RECT 81.130 6.580 81.300 7.070 ;
        RECT 81.130 6.380 83.040 6.580 ;
        RECT 87.880 6.380 88.050 7.070 ;
        RECT 88.360 6.380 88.530 7.070 ;
        RECT 88.840 6.580 89.010 7.070 ;
        RECT 88.840 6.380 90.750 6.580 ;
        RECT 95.590 6.380 95.760 7.070 ;
        RECT 96.070 6.380 96.240 7.070 ;
        RECT 96.550 6.580 96.720 7.070 ;
        RECT 96.550 6.380 98.460 6.580 ;
        RECT 103.300 6.380 103.470 7.070 ;
        RECT 103.780 6.380 103.950 7.070 ;
        RECT 104.260 6.580 104.430 7.070 ;
        RECT 104.260 6.380 106.170 6.580 ;
        RECT 111.010 6.380 111.180 7.070 ;
        RECT 111.490 6.380 111.660 7.070 ;
        RECT 111.970 6.580 112.140 7.070 ;
        RECT 111.970 6.380 113.880 6.580 ;
        RECT 118.720 6.380 118.890 7.070 ;
        RECT 119.200 6.380 119.370 7.070 ;
        RECT 119.680 6.580 119.850 7.070 ;
        RECT 119.680 6.380 121.590 6.580 ;
        RECT 3.230 6.040 3.560 6.210 ;
        RECT 2.040 4.805 2.370 4.975 ;
        RECT 5.270 4.805 5.600 4.975 ;
        RECT 0.910 3.635 1.240 4.615 ;
        RECT 5.770 4.590 5.940 6.380 ;
        RECT 10.940 6.040 11.270 6.210 ;
        RECT 9.750 4.805 10.080 4.975 ;
        RECT 12.980 4.805 13.310 4.975 ;
        RECT 1.010 3.035 1.240 3.635 ;
        RECT 1.900 3.550 2.070 4.590 ;
        RECT 5.560 4.390 5.940 4.590 ;
        RECT 3.620 4.005 3.950 4.175 ;
        RECT 2.040 3.165 2.370 3.335 ;
        RECT 0.910 2.710 1.240 3.035 ;
        RECT 2.980 2.750 3.150 3.790 ;
        RECT 3.460 2.750 3.630 3.790 ;
        RECT 3.940 2.930 4.110 3.790 ;
        RECT 5.570 3.550 5.740 4.390 ;
        RECT 6.860 3.645 7.190 4.625 ;
        RECT 6.460 3.440 6.790 3.475 ;
        RECT 5.270 3.340 5.600 3.350 ;
        RECT 6.010 3.340 6.790 3.440 ;
        RECT 5.270 3.270 6.790 3.340 ;
        RECT 5.270 3.170 6.200 3.270 ;
        RECT 6.460 3.235 6.790 3.270 ;
        RECT 5.270 3.165 5.600 3.170 ;
        RECT 6.960 3.045 7.190 3.645 ;
        RECT 8.620 3.635 8.950 4.615 ;
        RECT 13.480 4.590 13.650 6.380 ;
        RECT 18.650 6.040 18.980 6.210 ;
        RECT 17.460 4.805 17.790 4.975 ;
        RECT 20.690 4.805 21.020 4.975 ;
        RECT 3.940 2.760 5.340 2.930 ;
        RECT 3.940 2.750 4.110 2.760 ;
        RECT 0.910 2.550 2.590 2.710 ;
        RECT 0.910 2.530 3.470 2.550 ;
        RECT 0.910 2.405 1.240 2.530 ;
        RECT 2.410 2.370 3.470 2.530 ;
        RECT 3.140 2.365 3.470 2.370 ;
        RECT 3.700 1.960 4.030 2.130 ;
        RECT 5.100 2.090 5.340 2.760 ;
        RECT 6.860 2.415 7.190 3.045 ;
        RECT 8.720 3.035 8.950 3.635 ;
        RECT 9.610 3.550 9.780 4.590 ;
        RECT 13.270 4.390 13.650 4.590 ;
        RECT 11.330 4.005 11.660 4.175 ;
        RECT 9.750 3.165 10.080 3.335 ;
        RECT 8.620 2.710 8.950 3.035 ;
        RECT 10.690 2.750 10.860 3.790 ;
        RECT 11.170 2.750 11.340 3.790 ;
        RECT 11.650 2.930 11.820 3.790 ;
        RECT 13.280 3.550 13.450 4.390 ;
        RECT 14.570 3.645 14.900 4.625 ;
        RECT 14.170 3.440 14.500 3.475 ;
        RECT 12.980 3.340 13.310 3.350 ;
        RECT 13.720 3.340 14.500 3.440 ;
        RECT 12.980 3.270 14.500 3.340 ;
        RECT 12.980 3.170 13.910 3.270 ;
        RECT 14.170 3.235 14.500 3.270 ;
        RECT 12.980 3.165 13.310 3.170 ;
        RECT 14.670 3.045 14.900 3.645 ;
        RECT 16.330 3.635 16.660 4.615 ;
        RECT 21.190 4.590 21.360 6.380 ;
        RECT 26.360 6.040 26.690 6.210 ;
        RECT 25.170 4.805 25.500 4.975 ;
        RECT 28.400 4.805 28.730 4.975 ;
        RECT 11.650 2.760 13.050 2.930 ;
        RECT 11.650 2.750 11.820 2.760 ;
        RECT 8.620 2.550 10.300 2.710 ;
        RECT 8.620 2.530 11.180 2.550 ;
        RECT 8.620 2.405 8.950 2.530 ;
        RECT 10.120 2.370 11.180 2.530 ;
        RECT 10.850 2.365 11.180 2.370 ;
        RECT 11.410 1.960 11.740 2.130 ;
        RECT 12.810 2.090 13.050 2.760 ;
        RECT 14.570 2.415 14.900 3.045 ;
        RECT 16.430 3.035 16.660 3.635 ;
        RECT 17.320 3.550 17.490 4.590 ;
        RECT 20.980 4.390 21.360 4.590 ;
        RECT 19.040 4.005 19.370 4.175 ;
        RECT 17.460 3.165 17.790 3.335 ;
        RECT 16.330 2.710 16.660 3.035 ;
        RECT 18.400 2.750 18.570 3.790 ;
        RECT 18.880 2.750 19.050 3.790 ;
        RECT 19.360 2.930 19.530 3.790 ;
        RECT 20.990 3.550 21.160 4.390 ;
        RECT 22.280 3.645 22.610 4.625 ;
        RECT 21.880 3.440 22.210 3.475 ;
        RECT 20.690 3.340 21.020 3.350 ;
        RECT 21.430 3.340 22.210 3.440 ;
        RECT 20.690 3.270 22.210 3.340 ;
        RECT 20.690 3.170 21.620 3.270 ;
        RECT 21.880 3.235 22.210 3.270 ;
        RECT 20.690 3.165 21.020 3.170 ;
        RECT 22.380 3.045 22.610 3.645 ;
        RECT 24.040 3.635 24.370 4.615 ;
        RECT 28.900 4.590 29.070 6.380 ;
        RECT 34.070 6.040 34.400 6.210 ;
        RECT 32.880 4.805 33.210 4.975 ;
        RECT 36.110 4.805 36.440 4.975 ;
        RECT 19.360 2.760 20.760 2.930 ;
        RECT 19.360 2.750 19.530 2.760 ;
        RECT 16.330 2.550 18.010 2.710 ;
        RECT 16.330 2.530 18.890 2.550 ;
        RECT 16.330 2.405 16.660 2.530 ;
        RECT 17.830 2.370 18.890 2.530 ;
        RECT 18.560 2.365 18.890 2.370 ;
        RECT 19.120 1.960 19.450 2.130 ;
        RECT 20.520 2.090 20.760 2.760 ;
        RECT 22.280 2.415 22.610 3.045 ;
        RECT 24.140 3.035 24.370 3.635 ;
        RECT 25.030 3.550 25.200 4.590 ;
        RECT 28.690 4.390 29.070 4.590 ;
        RECT 26.750 4.005 27.080 4.175 ;
        RECT 25.170 3.165 25.500 3.335 ;
        RECT 24.040 2.710 24.370 3.035 ;
        RECT 26.110 2.750 26.280 3.790 ;
        RECT 26.590 2.750 26.760 3.790 ;
        RECT 27.070 2.930 27.240 3.790 ;
        RECT 28.700 3.550 28.870 4.390 ;
        RECT 29.990 3.645 30.320 4.625 ;
        RECT 29.590 3.440 29.920 3.475 ;
        RECT 28.400 3.340 28.730 3.350 ;
        RECT 29.140 3.340 29.920 3.440 ;
        RECT 28.400 3.270 29.920 3.340 ;
        RECT 28.400 3.170 29.330 3.270 ;
        RECT 29.590 3.235 29.920 3.270 ;
        RECT 28.400 3.165 28.730 3.170 ;
        RECT 30.090 3.045 30.320 3.645 ;
        RECT 31.750 3.635 32.080 4.615 ;
        RECT 36.610 4.590 36.780 6.380 ;
        RECT 41.780 6.040 42.110 6.210 ;
        RECT 40.590 4.805 40.920 4.975 ;
        RECT 43.820 4.805 44.150 4.975 ;
        RECT 27.070 2.760 28.470 2.930 ;
        RECT 27.070 2.750 27.240 2.760 ;
        RECT 24.040 2.550 25.720 2.710 ;
        RECT 24.040 2.530 26.600 2.550 ;
        RECT 24.040 2.405 24.370 2.530 ;
        RECT 25.540 2.370 26.600 2.530 ;
        RECT 26.270 2.365 26.600 2.370 ;
        RECT 26.830 1.960 27.160 2.130 ;
        RECT 28.230 2.090 28.470 2.760 ;
        RECT 29.990 2.415 30.320 3.045 ;
        RECT 31.850 3.035 32.080 3.635 ;
        RECT 32.740 3.550 32.910 4.590 ;
        RECT 36.400 4.390 36.780 4.590 ;
        RECT 34.460 4.005 34.790 4.175 ;
        RECT 32.880 3.165 33.210 3.335 ;
        RECT 31.750 2.710 32.080 3.035 ;
        RECT 33.820 2.750 33.990 3.790 ;
        RECT 34.300 2.750 34.470 3.790 ;
        RECT 34.780 2.930 34.950 3.790 ;
        RECT 36.410 3.550 36.580 4.390 ;
        RECT 37.700 3.645 38.030 4.625 ;
        RECT 37.300 3.440 37.630 3.475 ;
        RECT 36.110 3.340 36.440 3.350 ;
        RECT 36.850 3.340 37.630 3.440 ;
        RECT 36.110 3.270 37.630 3.340 ;
        RECT 36.110 3.170 37.040 3.270 ;
        RECT 37.300 3.235 37.630 3.270 ;
        RECT 36.110 3.165 36.440 3.170 ;
        RECT 37.800 3.045 38.030 3.645 ;
        RECT 39.460 3.635 39.790 4.615 ;
        RECT 44.320 4.590 44.490 6.380 ;
        RECT 49.490 6.040 49.820 6.210 ;
        RECT 48.300 4.805 48.630 4.975 ;
        RECT 51.530 4.805 51.860 4.975 ;
        RECT 34.780 2.760 36.180 2.930 ;
        RECT 34.780 2.750 34.950 2.760 ;
        RECT 31.750 2.550 33.430 2.710 ;
        RECT 31.750 2.530 34.310 2.550 ;
        RECT 31.750 2.405 32.080 2.530 ;
        RECT 33.250 2.370 34.310 2.530 ;
        RECT 33.980 2.365 34.310 2.370 ;
        RECT 34.540 1.960 34.870 2.130 ;
        RECT 35.940 2.090 36.180 2.760 ;
        RECT 37.700 2.415 38.030 3.045 ;
        RECT 39.560 3.035 39.790 3.635 ;
        RECT 40.450 3.550 40.620 4.590 ;
        RECT 44.110 4.390 44.490 4.590 ;
        RECT 42.170 4.005 42.500 4.175 ;
        RECT 40.590 3.165 40.920 3.335 ;
        RECT 39.460 2.710 39.790 3.035 ;
        RECT 41.530 2.750 41.700 3.790 ;
        RECT 42.010 2.750 42.180 3.790 ;
        RECT 42.490 2.930 42.660 3.790 ;
        RECT 44.120 3.550 44.290 4.390 ;
        RECT 45.410 3.645 45.740 4.625 ;
        RECT 45.010 3.440 45.340 3.475 ;
        RECT 43.820 3.340 44.150 3.350 ;
        RECT 44.560 3.340 45.340 3.440 ;
        RECT 43.820 3.270 45.340 3.340 ;
        RECT 43.820 3.170 44.750 3.270 ;
        RECT 45.010 3.235 45.340 3.270 ;
        RECT 43.820 3.165 44.150 3.170 ;
        RECT 45.510 3.045 45.740 3.645 ;
        RECT 47.170 3.635 47.500 4.615 ;
        RECT 52.030 4.590 52.200 6.380 ;
        RECT 57.200 6.040 57.530 6.210 ;
        RECT 56.010 4.805 56.340 4.975 ;
        RECT 59.240 4.805 59.570 4.975 ;
        RECT 42.490 2.760 43.890 2.930 ;
        RECT 42.490 2.750 42.660 2.760 ;
        RECT 39.460 2.550 41.140 2.710 ;
        RECT 39.460 2.530 42.020 2.550 ;
        RECT 39.460 2.405 39.790 2.530 ;
        RECT 40.960 2.370 42.020 2.530 ;
        RECT 41.690 2.365 42.020 2.370 ;
        RECT 42.250 1.960 42.580 2.130 ;
        RECT 43.650 2.090 43.890 2.760 ;
        RECT 45.410 2.415 45.740 3.045 ;
        RECT 47.270 3.035 47.500 3.635 ;
        RECT 48.160 3.550 48.330 4.590 ;
        RECT 51.820 4.390 52.200 4.590 ;
        RECT 49.880 4.005 50.210 4.175 ;
        RECT 48.300 3.165 48.630 3.335 ;
        RECT 47.170 2.710 47.500 3.035 ;
        RECT 49.240 2.750 49.410 3.790 ;
        RECT 49.720 2.750 49.890 3.790 ;
        RECT 50.200 2.930 50.370 3.790 ;
        RECT 51.830 3.550 52.000 4.390 ;
        RECT 53.120 3.645 53.450 4.625 ;
        RECT 52.720 3.440 53.050 3.475 ;
        RECT 51.530 3.340 51.860 3.350 ;
        RECT 52.270 3.340 53.050 3.440 ;
        RECT 51.530 3.270 53.050 3.340 ;
        RECT 51.530 3.170 52.460 3.270 ;
        RECT 52.720 3.235 53.050 3.270 ;
        RECT 51.530 3.165 51.860 3.170 ;
        RECT 53.220 3.045 53.450 3.645 ;
        RECT 54.880 3.635 55.210 4.615 ;
        RECT 59.740 4.590 59.910 6.380 ;
        RECT 64.910 6.040 65.240 6.210 ;
        RECT 63.720 4.805 64.050 4.975 ;
        RECT 66.950 4.805 67.280 4.975 ;
        RECT 50.200 2.760 51.600 2.930 ;
        RECT 50.200 2.750 50.370 2.760 ;
        RECT 47.170 2.550 48.850 2.710 ;
        RECT 47.170 2.530 49.730 2.550 ;
        RECT 47.170 2.405 47.500 2.530 ;
        RECT 48.670 2.370 49.730 2.530 ;
        RECT 49.400 2.365 49.730 2.370 ;
        RECT 49.960 1.960 50.290 2.130 ;
        RECT 51.360 2.090 51.600 2.760 ;
        RECT 53.120 2.415 53.450 3.045 ;
        RECT 54.980 3.035 55.210 3.635 ;
        RECT 55.870 3.550 56.040 4.590 ;
        RECT 59.530 4.390 59.910 4.590 ;
        RECT 57.590 4.005 57.920 4.175 ;
        RECT 56.010 3.165 56.340 3.335 ;
        RECT 54.880 2.710 55.210 3.035 ;
        RECT 56.950 2.750 57.120 3.790 ;
        RECT 57.430 2.750 57.600 3.790 ;
        RECT 57.910 2.930 58.080 3.790 ;
        RECT 59.540 3.550 59.710 4.390 ;
        RECT 60.830 3.645 61.160 4.625 ;
        RECT 60.430 3.440 60.760 3.475 ;
        RECT 59.240 3.340 59.570 3.350 ;
        RECT 59.980 3.340 60.760 3.440 ;
        RECT 59.240 3.270 60.760 3.340 ;
        RECT 59.240 3.170 60.170 3.270 ;
        RECT 60.430 3.235 60.760 3.270 ;
        RECT 59.240 3.165 59.570 3.170 ;
        RECT 60.930 3.045 61.160 3.645 ;
        RECT 62.590 3.635 62.920 4.615 ;
        RECT 67.450 4.590 67.620 6.380 ;
        RECT 72.620 6.040 72.950 6.210 ;
        RECT 71.430 4.805 71.760 4.975 ;
        RECT 74.660 4.805 74.990 4.975 ;
        RECT 57.910 2.760 59.310 2.930 ;
        RECT 57.910 2.750 58.080 2.760 ;
        RECT 54.880 2.550 56.560 2.710 ;
        RECT 54.880 2.530 57.440 2.550 ;
        RECT 54.880 2.405 55.210 2.530 ;
        RECT 56.380 2.370 57.440 2.530 ;
        RECT 57.110 2.365 57.440 2.370 ;
        RECT 57.670 1.960 58.000 2.130 ;
        RECT 59.070 2.090 59.310 2.760 ;
        RECT 60.830 2.415 61.160 3.045 ;
        RECT 62.690 3.035 62.920 3.635 ;
        RECT 63.580 3.550 63.750 4.590 ;
        RECT 67.240 4.390 67.620 4.590 ;
        RECT 65.300 4.005 65.630 4.175 ;
        RECT 63.720 3.165 64.050 3.335 ;
        RECT 62.590 2.710 62.920 3.035 ;
        RECT 64.660 2.750 64.830 3.790 ;
        RECT 65.140 2.750 65.310 3.790 ;
        RECT 65.620 2.930 65.790 3.790 ;
        RECT 67.250 3.550 67.420 4.390 ;
        RECT 68.540 3.645 68.870 4.625 ;
        RECT 68.140 3.440 68.470 3.475 ;
        RECT 66.950 3.340 67.280 3.350 ;
        RECT 67.690 3.340 68.470 3.440 ;
        RECT 66.950 3.270 68.470 3.340 ;
        RECT 66.950 3.170 67.880 3.270 ;
        RECT 68.140 3.235 68.470 3.270 ;
        RECT 66.950 3.165 67.280 3.170 ;
        RECT 68.640 3.045 68.870 3.645 ;
        RECT 70.300 3.635 70.630 4.615 ;
        RECT 75.160 4.590 75.330 6.380 ;
        RECT 80.330 6.040 80.660 6.210 ;
        RECT 79.140 4.805 79.470 4.975 ;
        RECT 82.370 4.805 82.700 4.975 ;
        RECT 65.620 2.760 67.020 2.930 ;
        RECT 65.620 2.750 65.790 2.760 ;
        RECT 62.590 2.550 64.270 2.710 ;
        RECT 62.590 2.530 65.150 2.550 ;
        RECT 62.590 2.405 62.920 2.530 ;
        RECT 64.090 2.370 65.150 2.530 ;
        RECT 64.820 2.365 65.150 2.370 ;
        RECT 65.380 1.960 65.710 2.130 ;
        RECT 66.780 2.090 67.020 2.760 ;
        RECT 68.540 2.415 68.870 3.045 ;
        RECT 70.400 3.035 70.630 3.635 ;
        RECT 71.290 3.550 71.460 4.590 ;
        RECT 74.950 4.390 75.330 4.590 ;
        RECT 73.010 4.005 73.340 4.175 ;
        RECT 71.430 3.165 71.760 3.335 ;
        RECT 70.300 2.710 70.630 3.035 ;
        RECT 72.370 2.750 72.540 3.790 ;
        RECT 72.850 2.750 73.020 3.790 ;
        RECT 73.330 2.930 73.500 3.790 ;
        RECT 74.960 3.550 75.130 4.390 ;
        RECT 76.250 3.645 76.580 4.625 ;
        RECT 75.850 3.440 76.180 3.475 ;
        RECT 74.660 3.340 74.990 3.350 ;
        RECT 75.400 3.340 76.180 3.440 ;
        RECT 74.660 3.270 76.180 3.340 ;
        RECT 74.660 3.170 75.590 3.270 ;
        RECT 75.850 3.235 76.180 3.270 ;
        RECT 74.660 3.165 74.990 3.170 ;
        RECT 76.350 3.045 76.580 3.645 ;
        RECT 78.010 3.635 78.340 4.615 ;
        RECT 82.870 4.590 83.040 6.380 ;
        RECT 88.040 6.040 88.370 6.210 ;
        RECT 86.850 4.805 87.180 4.975 ;
        RECT 90.080 4.805 90.410 4.975 ;
        RECT 73.330 2.760 74.730 2.930 ;
        RECT 73.330 2.750 73.500 2.760 ;
        RECT 70.300 2.550 71.980 2.710 ;
        RECT 70.300 2.530 72.860 2.550 ;
        RECT 70.300 2.405 70.630 2.530 ;
        RECT 71.800 2.370 72.860 2.530 ;
        RECT 72.530 2.365 72.860 2.370 ;
        RECT 73.090 1.960 73.420 2.130 ;
        RECT 74.490 2.090 74.730 2.760 ;
        RECT 76.250 2.415 76.580 3.045 ;
        RECT 78.110 3.035 78.340 3.635 ;
        RECT 79.000 3.550 79.170 4.590 ;
        RECT 82.660 4.390 83.040 4.590 ;
        RECT 80.720 4.005 81.050 4.175 ;
        RECT 79.140 3.165 79.470 3.335 ;
        RECT 78.010 2.710 78.340 3.035 ;
        RECT 80.080 2.750 80.250 3.790 ;
        RECT 80.560 2.750 80.730 3.790 ;
        RECT 81.040 2.930 81.210 3.790 ;
        RECT 82.670 3.550 82.840 4.390 ;
        RECT 83.960 3.645 84.290 4.625 ;
        RECT 83.560 3.440 83.890 3.475 ;
        RECT 82.370 3.340 82.700 3.350 ;
        RECT 83.110 3.340 83.890 3.440 ;
        RECT 82.370 3.270 83.890 3.340 ;
        RECT 82.370 3.170 83.300 3.270 ;
        RECT 83.560 3.235 83.890 3.270 ;
        RECT 82.370 3.165 82.700 3.170 ;
        RECT 84.060 3.045 84.290 3.645 ;
        RECT 85.720 3.635 86.050 4.615 ;
        RECT 90.580 4.590 90.750 6.380 ;
        RECT 95.750 6.040 96.080 6.210 ;
        RECT 94.560 4.805 94.890 4.975 ;
        RECT 97.790 4.805 98.120 4.975 ;
        RECT 81.040 2.760 82.440 2.930 ;
        RECT 81.040 2.750 81.210 2.760 ;
        RECT 78.010 2.550 79.690 2.710 ;
        RECT 78.010 2.530 80.570 2.550 ;
        RECT 78.010 2.405 78.340 2.530 ;
        RECT 79.510 2.370 80.570 2.530 ;
        RECT 80.240 2.365 80.570 2.370 ;
        RECT 80.800 1.960 81.130 2.130 ;
        RECT 82.200 2.090 82.440 2.760 ;
        RECT 83.960 2.415 84.290 3.045 ;
        RECT 85.820 3.035 86.050 3.635 ;
        RECT 86.710 3.550 86.880 4.590 ;
        RECT 90.370 4.390 90.750 4.590 ;
        RECT 88.430 4.005 88.760 4.175 ;
        RECT 86.850 3.165 87.180 3.335 ;
        RECT 85.720 2.710 86.050 3.035 ;
        RECT 87.790 2.750 87.960 3.790 ;
        RECT 88.270 2.750 88.440 3.790 ;
        RECT 88.750 2.930 88.920 3.790 ;
        RECT 90.380 3.550 90.550 4.390 ;
        RECT 91.670 3.645 92.000 4.625 ;
        RECT 91.270 3.440 91.600 3.475 ;
        RECT 90.080 3.340 90.410 3.350 ;
        RECT 90.820 3.340 91.600 3.440 ;
        RECT 90.080 3.270 91.600 3.340 ;
        RECT 90.080 3.170 91.010 3.270 ;
        RECT 91.270 3.235 91.600 3.270 ;
        RECT 90.080 3.165 90.410 3.170 ;
        RECT 91.770 3.045 92.000 3.645 ;
        RECT 93.430 3.635 93.760 4.615 ;
        RECT 98.290 4.590 98.460 6.380 ;
        RECT 103.460 6.040 103.790 6.210 ;
        RECT 102.270 4.805 102.600 4.975 ;
        RECT 105.500 4.805 105.830 4.975 ;
        RECT 88.750 2.760 90.150 2.930 ;
        RECT 88.750 2.750 88.920 2.760 ;
        RECT 85.720 2.550 87.400 2.710 ;
        RECT 85.720 2.530 88.280 2.550 ;
        RECT 85.720 2.405 86.050 2.530 ;
        RECT 87.220 2.370 88.280 2.530 ;
        RECT 87.950 2.365 88.280 2.370 ;
        RECT 88.510 1.960 88.840 2.130 ;
        RECT 89.910 2.090 90.150 2.760 ;
        RECT 91.670 2.415 92.000 3.045 ;
        RECT 93.530 3.035 93.760 3.635 ;
        RECT 94.420 3.550 94.590 4.590 ;
        RECT 98.080 4.390 98.460 4.590 ;
        RECT 96.140 4.005 96.470 4.175 ;
        RECT 94.560 3.165 94.890 3.335 ;
        RECT 93.430 2.710 93.760 3.035 ;
        RECT 95.500 2.750 95.670 3.790 ;
        RECT 95.980 2.750 96.150 3.790 ;
        RECT 96.460 2.930 96.630 3.790 ;
        RECT 98.090 3.550 98.260 4.390 ;
        RECT 99.380 3.645 99.710 4.625 ;
        RECT 98.980 3.440 99.310 3.475 ;
        RECT 97.790 3.340 98.120 3.350 ;
        RECT 98.530 3.340 99.310 3.440 ;
        RECT 97.790 3.270 99.310 3.340 ;
        RECT 97.790 3.170 98.720 3.270 ;
        RECT 98.980 3.235 99.310 3.270 ;
        RECT 97.790 3.165 98.120 3.170 ;
        RECT 99.480 3.045 99.710 3.645 ;
        RECT 101.140 3.635 101.470 4.615 ;
        RECT 106.000 4.590 106.170 6.380 ;
        RECT 111.170 6.040 111.500 6.210 ;
        RECT 109.980 4.805 110.310 4.975 ;
        RECT 113.210 4.805 113.540 4.975 ;
        RECT 96.460 2.760 97.860 2.930 ;
        RECT 96.460 2.750 96.630 2.760 ;
        RECT 93.430 2.550 95.110 2.710 ;
        RECT 93.430 2.530 95.990 2.550 ;
        RECT 93.430 2.405 93.760 2.530 ;
        RECT 94.930 2.370 95.990 2.530 ;
        RECT 95.660 2.365 95.990 2.370 ;
        RECT 96.220 1.960 96.550 2.130 ;
        RECT 97.620 2.090 97.860 2.760 ;
        RECT 99.380 2.415 99.710 3.045 ;
        RECT 101.240 3.035 101.470 3.635 ;
        RECT 102.130 3.550 102.300 4.590 ;
        RECT 105.790 4.390 106.170 4.590 ;
        RECT 103.850 4.005 104.180 4.175 ;
        RECT 102.270 3.165 102.600 3.335 ;
        RECT 101.140 2.710 101.470 3.035 ;
        RECT 103.210 2.750 103.380 3.790 ;
        RECT 103.690 2.750 103.860 3.790 ;
        RECT 104.170 2.930 104.340 3.790 ;
        RECT 105.800 3.550 105.970 4.390 ;
        RECT 107.090 3.645 107.420 4.625 ;
        RECT 106.690 3.440 107.020 3.475 ;
        RECT 105.500 3.340 105.830 3.350 ;
        RECT 106.240 3.340 107.020 3.440 ;
        RECT 105.500 3.270 107.020 3.340 ;
        RECT 105.500 3.170 106.430 3.270 ;
        RECT 106.690 3.235 107.020 3.270 ;
        RECT 105.500 3.165 105.830 3.170 ;
        RECT 107.190 3.045 107.420 3.645 ;
        RECT 108.850 3.635 109.180 4.615 ;
        RECT 113.710 4.590 113.880 6.380 ;
        RECT 118.880 6.040 119.210 6.210 ;
        RECT 117.690 4.805 118.020 4.975 ;
        RECT 120.920 4.805 121.250 4.975 ;
        RECT 104.170 2.760 105.570 2.930 ;
        RECT 104.170 2.750 104.340 2.760 ;
        RECT 101.140 2.550 102.820 2.710 ;
        RECT 101.140 2.530 103.700 2.550 ;
        RECT 101.140 2.405 101.470 2.530 ;
        RECT 102.640 2.370 103.700 2.530 ;
        RECT 103.370 2.365 103.700 2.370 ;
        RECT 103.930 1.960 104.260 2.130 ;
        RECT 105.330 2.090 105.570 2.760 ;
        RECT 107.090 2.415 107.420 3.045 ;
        RECT 108.950 3.035 109.180 3.635 ;
        RECT 109.840 3.550 110.010 4.590 ;
        RECT 113.500 4.390 113.880 4.590 ;
        RECT 111.560 4.005 111.890 4.175 ;
        RECT 109.980 3.165 110.310 3.335 ;
        RECT 108.850 2.710 109.180 3.035 ;
        RECT 110.920 2.750 111.090 3.790 ;
        RECT 111.400 2.750 111.570 3.790 ;
        RECT 111.880 2.930 112.050 3.790 ;
        RECT 113.510 3.550 113.680 4.390 ;
        RECT 114.800 3.645 115.130 4.625 ;
        RECT 114.400 3.440 114.730 3.475 ;
        RECT 113.210 3.340 113.540 3.350 ;
        RECT 113.950 3.340 114.730 3.440 ;
        RECT 113.210 3.270 114.730 3.340 ;
        RECT 113.210 3.170 114.140 3.270 ;
        RECT 114.400 3.235 114.730 3.270 ;
        RECT 113.210 3.165 113.540 3.170 ;
        RECT 114.900 3.045 115.130 3.645 ;
        RECT 116.560 3.635 116.890 4.615 ;
        RECT 121.420 4.590 121.590 6.380 ;
        RECT 111.880 2.760 113.280 2.930 ;
        RECT 111.880 2.750 112.050 2.760 ;
        RECT 108.850 2.550 110.530 2.710 ;
        RECT 108.850 2.530 111.410 2.550 ;
        RECT 108.850 2.405 109.180 2.530 ;
        RECT 110.350 2.370 111.410 2.530 ;
        RECT 111.080 2.365 111.410 2.370 ;
        RECT 111.640 1.960 111.970 2.130 ;
        RECT 113.040 2.090 113.280 2.760 ;
        RECT 114.800 2.415 115.130 3.045 ;
        RECT 116.660 3.035 116.890 3.635 ;
        RECT 117.550 3.550 117.720 4.590 ;
        RECT 121.210 4.390 121.590 4.590 ;
        RECT 119.270 4.005 119.600 4.175 ;
        RECT 117.690 3.165 118.020 3.335 ;
        RECT 116.560 2.710 116.890 3.035 ;
        RECT 118.630 2.750 118.800 3.790 ;
        RECT 119.110 2.750 119.280 3.790 ;
        RECT 119.590 2.930 119.760 3.790 ;
        RECT 121.220 3.550 121.390 4.390 ;
        RECT 122.510 3.645 122.840 4.625 ;
        RECT 122.110 3.440 122.440 3.475 ;
        RECT 120.920 3.340 121.250 3.350 ;
        RECT 121.660 3.340 122.440 3.440 ;
        RECT 120.920 3.270 122.440 3.340 ;
        RECT 120.920 3.170 121.850 3.270 ;
        RECT 122.110 3.235 122.440 3.270 ;
        RECT 120.920 3.165 121.250 3.170 ;
        RECT 122.610 3.045 122.840 3.645 ;
        RECT 119.590 2.760 120.990 2.930 ;
        RECT 119.590 2.750 119.760 2.760 ;
        RECT 116.560 2.550 118.240 2.710 ;
        RECT 116.560 2.530 119.120 2.550 ;
        RECT 116.560 2.405 116.890 2.530 ;
        RECT 118.060 2.370 119.120 2.530 ;
        RECT 118.790 2.365 119.120 2.370 ;
        RECT 119.350 1.960 119.680 2.130 ;
        RECT 120.750 2.090 120.990 2.760 ;
        RECT 122.510 2.415 122.840 3.045 ;
        RECT 3.060 1.100 3.230 1.790 ;
        RECT 3.540 1.100 3.710 1.790 ;
        RECT 4.020 1.100 4.190 1.790 ;
        RECT 10.770 1.100 10.940 1.790 ;
        RECT 11.250 1.100 11.420 1.790 ;
        RECT 11.730 1.100 11.900 1.790 ;
        RECT 18.480 1.100 18.650 1.790 ;
        RECT 18.960 1.100 19.130 1.790 ;
        RECT 19.440 1.100 19.610 1.790 ;
        RECT 26.190 1.100 26.360 1.790 ;
        RECT 26.670 1.100 26.840 1.790 ;
        RECT 27.150 1.100 27.320 1.790 ;
        RECT 33.900 1.100 34.070 1.790 ;
        RECT 34.380 1.100 34.550 1.790 ;
        RECT 34.860 1.100 35.030 1.790 ;
        RECT 41.610 1.100 41.780 1.790 ;
        RECT 42.090 1.100 42.260 1.790 ;
        RECT 42.570 1.100 42.740 1.790 ;
        RECT 49.320 1.100 49.490 1.790 ;
        RECT 49.800 1.100 49.970 1.790 ;
        RECT 50.280 1.100 50.450 1.790 ;
        RECT 57.030 1.100 57.200 1.790 ;
        RECT 57.510 1.100 57.680 1.790 ;
        RECT 57.990 1.100 58.160 1.790 ;
        RECT 64.740 1.100 64.910 1.790 ;
        RECT 65.220 1.100 65.390 1.790 ;
        RECT 65.700 1.100 65.870 1.790 ;
        RECT 72.450 1.100 72.620 1.790 ;
        RECT 72.930 1.100 73.100 1.790 ;
        RECT 73.410 1.100 73.580 1.790 ;
        RECT 80.160 1.100 80.330 1.790 ;
        RECT 80.640 1.100 80.810 1.790 ;
        RECT 81.120 1.100 81.290 1.790 ;
        RECT 87.870 1.100 88.040 1.790 ;
        RECT 88.350 1.100 88.520 1.790 ;
        RECT 88.830 1.100 89.000 1.790 ;
        RECT 95.580 1.100 95.750 1.790 ;
        RECT 96.060 1.100 96.230 1.790 ;
        RECT 96.540 1.100 96.710 1.790 ;
        RECT 103.290 1.100 103.460 1.790 ;
        RECT 103.770 1.100 103.940 1.790 ;
        RECT 104.250 1.100 104.420 1.790 ;
        RECT 111.000 1.100 111.170 1.790 ;
        RECT 111.480 1.100 111.650 1.790 ;
        RECT 111.960 1.100 112.130 1.790 ;
        RECT 118.710 1.100 118.880 1.790 ;
        RECT 119.190 1.100 119.360 1.790 ;
        RECT 119.670 1.100 119.840 1.790 ;
        RECT 3.220 0.760 3.550 0.930 ;
        RECT 10.930 0.760 11.260 0.930 ;
        RECT 18.640 0.760 18.970 0.930 ;
        RECT 26.350 0.760 26.680 0.930 ;
        RECT 34.060 0.760 34.390 0.930 ;
        RECT 41.770 0.760 42.100 0.930 ;
        RECT 49.480 0.760 49.810 0.930 ;
        RECT 57.190 0.760 57.520 0.930 ;
        RECT 64.900 0.760 65.230 0.930 ;
        RECT 72.610 0.760 72.940 0.930 ;
        RECT 80.320 0.760 80.650 0.930 ;
        RECT 88.030 0.760 88.360 0.930 ;
        RECT 95.740 0.760 96.070 0.930 ;
        RECT 103.450 0.760 103.780 0.930 ;
        RECT 111.160 0.760 111.490 0.930 ;
        RECT 118.870 0.760 119.200 0.930 ;
      LAYER mcon ;
        RECT 3.920 32.530 4.090 32.700 ;
        RECT 11.630 32.530 11.800 32.700 ;
        RECT 19.340 32.530 19.510 32.700 ;
        RECT 27.050 32.530 27.220 32.700 ;
        RECT 34.760 32.530 34.930 32.700 ;
        RECT 42.470 32.530 42.640 32.700 ;
        RECT 50.180 32.530 50.350 32.700 ;
        RECT 57.890 32.530 58.060 32.700 ;
        RECT 65.600 32.530 65.770 32.700 ;
        RECT 73.310 32.530 73.480 32.700 ;
        RECT 81.020 32.530 81.190 32.700 ;
        RECT 88.730 32.530 88.900 32.700 ;
        RECT 96.440 32.530 96.610 32.700 ;
        RECT 104.150 32.530 104.320 32.700 ;
        RECT 111.860 32.530 112.030 32.700 ;
        RECT 119.570 32.530 119.740 32.700 ;
        RECT 3.200 31.750 3.370 32.280 ;
        RECT 3.680 31.750 3.850 32.280 ;
        RECT 4.160 31.750 4.330 32.280 ;
        RECT 10.910 31.750 11.080 32.280 ;
        RECT 11.390 31.750 11.560 32.280 ;
        RECT 11.870 31.750 12.040 32.280 ;
        RECT 18.620 31.750 18.790 32.280 ;
        RECT 19.100 31.750 19.270 32.280 ;
        RECT 19.580 31.750 19.750 32.280 ;
        RECT 26.330 31.750 26.500 32.280 ;
        RECT 26.810 31.750 26.980 32.280 ;
        RECT 27.290 31.750 27.460 32.280 ;
        RECT 34.040 31.750 34.210 32.280 ;
        RECT 34.520 31.750 34.690 32.280 ;
        RECT 35.000 31.750 35.170 32.280 ;
        RECT 41.750 31.750 41.920 32.280 ;
        RECT 42.230 31.750 42.400 32.280 ;
        RECT 42.710 31.750 42.880 32.280 ;
        RECT 49.460 31.750 49.630 32.280 ;
        RECT 49.940 31.750 50.110 32.280 ;
        RECT 50.420 31.750 50.590 32.280 ;
        RECT 57.170 31.750 57.340 32.280 ;
        RECT 57.650 31.750 57.820 32.280 ;
        RECT 58.130 31.750 58.300 32.280 ;
        RECT 64.880 31.750 65.050 32.280 ;
        RECT 65.360 31.750 65.530 32.280 ;
        RECT 65.840 31.750 66.010 32.280 ;
        RECT 72.590 31.750 72.760 32.280 ;
        RECT 73.070 31.750 73.240 32.280 ;
        RECT 73.550 31.750 73.720 32.280 ;
        RECT 80.300 31.750 80.470 32.280 ;
        RECT 80.780 31.750 80.950 32.280 ;
        RECT 81.260 31.750 81.430 32.280 ;
        RECT 88.010 31.750 88.180 32.280 ;
        RECT 88.490 31.750 88.660 32.280 ;
        RECT 88.970 31.750 89.140 32.280 ;
        RECT 95.720 31.750 95.890 32.280 ;
        RECT 96.200 31.750 96.370 32.280 ;
        RECT 96.680 31.750 96.850 32.280 ;
        RECT 103.430 31.750 103.600 32.280 ;
        RECT 103.910 31.750 104.080 32.280 ;
        RECT 104.390 31.750 104.560 32.280 ;
        RECT 111.140 31.750 111.310 32.280 ;
        RECT 111.620 31.750 111.790 32.280 ;
        RECT 112.100 31.750 112.270 32.280 ;
        RECT 118.850 31.750 119.020 32.280 ;
        RECT 119.330 31.750 119.500 32.280 ;
        RECT 119.810 31.750 119.980 32.280 ;
        RECT 3.440 31.330 3.610 31.500 ;
        RECT 2.070 31.140 2.260 31.310 ;
        RECT 0.280 30.560 0.450 30.730 ;
        RECT 11.150 31.330 11.320 31.500 ;
        RECT 9.780 31.140 9.970 31.310 ;
        RECT 4.000 30.925 4.170 31.095 ;
        RECT 1.870 30.125 2.040 30.295 ;
        RECT 1.650 28.950 1.820 29.830 ;
        RECT 3.280 29.750 3.450 30.630 ;
        RECT 3.760 29.750 3.930 30.630 ;
        RECT 4.240 29.750 4.410 30.630 ;
        RECT 7.990 30.560 8.160 30.730 ;
        RECT 5.100 30.125 5.270 30.295 ;
        RECT 3.520 29.285 3.690 29.455 ;
        RECT 5.320 28.950 5.490 29.830 ;
        RECT 18.860 31.330 19.030 31.500 ;
        RECT 17.490 31.140 17.680 31.310 ;
        RECT 11.710 30.925 11.880 31.095 ;
        RECT 9.580 30.125 9.750 30.295 ;
        RECT 9.360 28.950 9.530 29.830 ;
        RECT 10.990 29.750 11.160 30.630 ;
        RECT 11.470 29.750 11.640 30.630 ;
        RECT 11.950 29.750 12.120 30.630 ;
        RECT 15.700 30.560 15.870 30.730 ;
        RECT 12.810 30.125 12.980 30.295 ;
        RECT 11.230 29.285 11.400 29.455 ;
        RECT 13.030 28.950 13.200 29.830 ;
        RECT 26.570 31.330 26.740 31.500 ;
        RECT 25.200 31.140 25.390 31.310 ;
        RECT 19.420 30.925 19.590 31.095 ;
        RECT 1.870 28.485 2.040 28.655 ;
        RECT 5.100 28.485 5.270 28.655 ;
        RECT 3.910 27.250 4.080 27.420 ;
        RECT 17.290 30.125 17.460 30.295 ;
        RECT 17.070 28.950 17.240 29.830 ;
        RECT 18.700 29.750 18.870 30.630 ;
        RECT 19.180 29.750 19.350 30.630 ;
        RECT 19.660 29.750 19.830 30.630 ;
        RECT 23.410 30.560 23.580 30.730 ;
        RECT 20.520 30.125 20.690 30.295 ;
        RECT 18.940 29.285 19.110 29.455 ;
        RECT 20.740 28.950 20.910 29.830 ;
        RECT 34.280 31.330 34.450 31.500 ;
        RECT 32.910 31.140 33.100 31.310 ;
        RECT 27.130 30.925 27.300 31.095 ;
        RECT 9.580 28.485 9.750 28.655 ;
        RECT 12.810 28.485 12.980 28.655 ;
        RECT 11.620 27.250 11.790 27.420 ;
        RECT 25.000 30.125 25.170 30.295 ;
        RECT 24.780 28.950 24.950 29.830 ;
        RECT 26.410 29.750 26.580 30.630 ;
        RECT 26.890 29.750 27.060 30.630 ;
        RECT 27.370 29.750 27.540 30.630 ;
        RECT 31.120 30.560 31.290 30.730 ;
        RECT 28.230 30.125 28.400 30.295 ;
        RECT 26.650 29.285 26.820 29.455 ;
        RECT 28.450 28.950 28.620 29.830 ;
        RECT 41.990 31.330 42.160 31.500 ;
        RECT 40.620 31.140 40.810 31.310 ;
        RECT 34.840 30.925 35.010 31.095 ;
        RECT 17.290 28.485 17.460 28.655 ;
        RECT 20.520 28.485 20.690 28.655 ;
        RECT 19.330 27.250 19.500 27.420 ;
        RECT 32.710 30.125 32.880 30.295 ;
        RECT 32.490 28.950 32.660 29.830 ;
        RECT 34.120 29.750 34.290 30.630 ;
        RECT 34.600 29.750 34.770 30.630 ;
        RECT 35.080 29.750 35.250 30.630 ;
        RECT 38.830 30.560 39.000 30.730 ;
        RECT 35.940 30.125 36.110 30.295 ;
        RECT 34.360 29.285 34.530 29.455 ;
        RECT 36.160 28.950 36.330 29.830 ;
        RECT 49.700 31.330 49.870 31.500 ;
        RECT 48.330 31.140 48.520 31.310 ;
        RECT 42.550 30.925 42.720 31.095 ;
        RECT 25.000 28.485 25.170 28.655 ;
        RECT 28.230 28.485 28.400 28.655 ;
        RECT 27.040 27.250 27.210 27.420 ;
        RECT 40.420 30.125 40.590 30.295 ;
        RECT 40.200 28.950 40.370 29.830 ;
        RECT 41.830 29.750 42.000 30.630 ;
        RECT 42.310 29.750 42.480 30.630 ;
        RECT 42.790 29.750 42.960 30.630 ;
        RECT 46.540 30.560 46.710 30.730 ;
        RECT 43.650 30.125 43.820 30.295 ;
        RECT 42.070 29.285 42.240 29.455 ;
        RECT 43.870 28.950 44.040 29.830 ;
        RECT 57.410 31.330 57.580 31.500 ;
        RECT 56.040 31.140 56.230 31.310 ;
        RECT 50.260 30.925 50.430 31.095 ;
        RECT 32.710 28.485 32.880 28.655 ;
        RECT 35.940 28.485 36.110 28.655 ;
        RECT 34.750 27.250 34.920 27.420 ;
        RECT 48.130 30.125 48.300 30.295 ;
        RECT 47.910 28.950 48.080 29.830 ;
        RECT 49.540 29.750 49.710 30.630 ;
        RECT 50.020 29.750 50.190 30.630 ;
        RECT 50.500 29.750 50.670 30.630 ;
        RECT 54.250 30.560 54.420 30.730 ;
        RECT 51.360 30.125 51.530 30.295 ;
        RECT 49.780 29.285 49.950 29.455 ;
        RECT 51.580 28.950 51.750 29.830 ;
        RECT 65.120 31.330 65.290 31.500 ;
        RECT 63.750 31.140 63.940 31.310 ;
        RECT 57.970 30.925 58.140 31.095 ;
        RECT 40.420 28.485 40.590 28.655 ;
        RECT 43.650 28.485 43.820 28.655 ;
        RECT 42.460 27.250 42.630 27.420 ;
        RECT 55.840 30.125 56.010 30.295 ;
        RECT 55.620 28.950 55.790 29.830 ;
        RECT 57.250 29.750 57.420 30.630 ;
        RECT 57.730 29.750 57.900 30.630 ;
        RECT 58.210 29.750 58.380 30.630 ;
        RECT 61.960 30.560 62.130 30.730 ;
        RECT 59.070 30.125 59.240 30.295 ;
        RECT 57.490 29.285 57.660 29.455 ;
        RECT 59.290 28.950 59.460 29.830 ;
        RECT 72.830 31.330 73.000 31.500 ;
        RECT 71.460 31.140 71.650 31.310 ;
        RECT 65.680 30.925 65.850 31.095 ;
        RECT 48.130 28.485 48.300 28.655 ;
        RECT 51.360 28.485 51.530 28.655 ;
        RECT 50.170 27.250 50.340 27.420 ;
        RECT 63.550 30.125 63.720 30.295 ;
        RECT 63.330 28.950 63.500 29.830 ;
        RECT 64.960 29.750 65.130 30.630 ;
        RECT 65.440 29.750 65.610 30.630 ;
        RECT 65.920 29.750 66.090 30.630 ;
        RECT 69.670 30.560 69.840 30.730 ;
        RECT 66.780 30.125 66.950 30.295 ;
        RECT 65.200 29.285 65.370 29.455 ;
        RECT 67.000 28.950 67.170 29.830 ;
        RECT 80.540 31.330 80.710 31.500 ;
        RECT 79.170 31.140 79.360 31.310 ;
        RECT 73.390 30.925 73.560 31.095 ;
        RECT 55.840 28.485 56.010 28.655 ;
        RECT 59.070 28.485 59.240 28.655 ;
        RECT 57.880 27.250 58.050 27.420 ;
        RECT 71.260 30.125 71.430 30.295 ;
        RECT 71.040 28.950 71.210 29.830 ;
        RECT 72.670 29.750 72.840 30.630 ;
        RECT 73.150 29.750 73.320 30.630 ;
        RECT 73.630 29.750 73.800 30.630 ;
        RECT 77.380 30.560 77.550 30.730 ;
        RECT 74.490 30.125 74.660 30.295 ;
        RECT 72.910 29.285 73.080 29.455 ;
        RECT 74.710 28.950 74.880 29.830 ;
        RECT 88.250 31.330 88.420 31.500 ;
        RECT 86.880 31.140 87.070 31.310 ;
        RECT 81.100 30.925 81.270 31.095 ;
        RECT 63.550 28.485 63.720 28.655 ;
        RECT 66.780 28.485 66.950 28.655 ;
        RECT 65.590 27.250 65.760 27.420 ;
        RECT 78.970 30.125 79.140 30.295 ;
        RECT 78.750 28.950 78.920 29.830 ;
        RECT 80.380 29.750 80.550 30.630 ;
        RECT 80.860 29.750 81.030 30.630 ;
        RECT 81.340 29.750 81.510 30.630 ;
        RECT 85.090 30.560 85.260 30.730 ;
        RECT 82.200 30.125 82.370 30.295 ;
        RECT 80.620 29.285 80.790 29.455 ;
        RECT 82.420 28.950 82.590 29.830 ;
        RECT 95.960 31.330 96.130 31.500 ;
        RECT 94.590 31.140 94.780 31.310 ;
        RECT 88.810 30.925 88.980 31.095 ;
        RECT 71.260 28.485 71.430 28.655 ;
        RECT 74.490 28.485 74.660 28.655 ;
        RECT 73.300 27.250 73.470 27.420 ;
        RECT 86.680 30.125 86.850 30.295 ;
        RECT 86.460 28.950 86.630 29.830 ;
        RECT 88.090 29.750 88.260 30.630 ;
        RECT 88.570 29.750 88.740 30.630 ;
        RECT 89.050 29.750 89.220 30.630 ;
        RECT 92.800 30.560 92.970 30.730 ;
        RECT 89.910 30.125 90.080 30.295 ;
        RECT 88.330 29.285 88.500 29.455 ;
        RECT 90.130 28.950 90.300 29.830 ;
        RECT 103.670 31.330 103.840 31.500 ;
        RECT 102.300 31.140 102.490 31.310 ;
        RECT 96.520 30.925 96.690 31.095 ;
        RECT 78.970 28.485 79.140 28.655 ;
        RECT 82.200 28.485 82.370 28.655 ;
        RECT 81.010 27.250 81.180 27.420 ;
        RECT 94.390 30.125 94.560 30.295 ;
        RECT 94.170 28.950 94.340 29.830 ;
        RECT 95.800 29.750 95.970 30.630 ;
        RECT 96.280 29.750 96.450 30.630 ;
        RECT 96.760 29.750 96.930 30.630 ;
        RECT 100.510 30.560 100.680 30.730 ;
        RECT 97.620 30.125 97.790 30.295 ;
        RECT 96.040 29.285 96.210 29.455 ;
        RECT 97.840 28.950 98.010 29.830 ;
        RECT 111.380 31.330 111.550 31.500 ;
        RECT 110.010 31.140 110.200 31.310 ;
        RECT 104.230 30.925 104.400 31.095 ;
        RECT 86.680 28.485 86.850 28.655 ;
        RECT 89.910 28.485 90.080 28.655 ;
        RECT 88.720 27.250 88.890 27.420 ;
        RECT 102.100 30.125 102.270 30.295 ;
        RECT 101.880 28.950 102.050 29.830 ;
        RECT 103.510 29.750 103.680 30.630 ;
        RECT 103.990 29.750 104.160 30.630 ;
        RECT 104.470 29.750 104.640 30.630 ;
        RECT 108.220 30.560 108.390 30.730 ;
        RECT 105.330 30.125 105.500 30.295 ;
        RECT 103.750 29.285 103.920 29.455 ;
        RECT 105.550 28.950 105.720 29.830 ;
        RECT 119.090 31.330 119.260 31.500 ;
        RECT 117.720 31.140 117.910 31.310 ;
        RECT 111.940 30.925 112.110 31.095 ;
        RECT 94.390 28.485 94.560 28.655 ;
        RECT 97.620 28.485 97.790 28.655 ;
        RECT 96.430 27.250 96.600 27.420 ;
        RECT 109.810 30.125 109.980 30.295 ;
        RECT 109.590 28.950 109.760 29.830 ;
        RECT 111.220 29.750 111.390 30.630 ;
        RECT 111.700 29.750 111.870 30.630 ;
        RECT 112.180 29.750 112.350 30.630 ;
        RECT 115.930 30.560 116.100 30.730 ;
        RECT 113.040 30.125 113.210 30.295 ;
        RECT 111.460 29.285 111.630 29.455 ;
        RECT 113.260 28.950 113.430 29.830 ;
        RECT 119.650 30.925 119.820 31.095 ;
        RECT 102.100 28.485 102.270 28.655 ;
        RECT 105.330 28.485 105.500 28.655 ;
        RECT 104.140 27.250 104.310 27.420 ;
        RECT 117.520 30.125 117.690 30.295 ;
        RECT 117.300 28.950 117.470 29.830 ;
        RECT 118.930 29.750 119.100 30.630 ;
        RECT 119.410 29.750 119.580 30.630 ;
        RECT 119.890 29.750 120.060 30.630 ;
        RECT 120.750 30.125 120.920 30.295 ;
        RECT 119.170 29.285 119.340 29.455 ;
        RECT 120.970 28.950 121.140 29.830 ;
        RECT 109.810 28.485 109.980 28.655 ;
        RECT 113.040 28.485 113.210 28.655 ;
        RECT 111.850 27.250 112.020 27.420 ;
        RECT 117.520 28.485 117.690 28.655 ;
        RECT 120.750 28.485 120.920 28.655 ;
        RECT 119.560 27.250 119.730 27.420 ;
        RECT 3.190 26.470 3.360 27.000 ;
        RECT 3.670 26.470 3.840 27.000 ;
        RECT 4.150 26.470 4.320 27.000 ;
        RECT 10.900 26.470 11.070 27.000 ;
        RECT 11.380 26.470 11.550 27.000 ;
        RECT 11.860 26.470 12.030 27.000 ;
        RECT 18.610 26.470 18.780 27.000 ;
        RECT 19.090 26.470 19.260 27.000 ;
        RECT 19.570 26.470 19.740 27.000 ;
        RECT 26.320 26.470 26.490 27.000 ;
        RECT 26.800 26.470 26.970 27.000 ;
        RECT 27.280 26.470 27.450 27.000 ;
        RECT 34.030 26.470 34.200 27.000 ;
        RECT 34.510 26.470 34.680 27.000 ;
        RECT 34.990 26.470 35.160 27.000 ;
        RECT 41.740 26.470 41.910 27.000 ;
        RECT 42.220 26.470 42.390 27.000 ;
        RECT 42.700 26.470 42.870 27.000 ;
        RECT 49.450 26.470 49.620 27.000 ;
        RECT 49.930 26.470 50.100 27.000 ;
        RECT 50.410 26.470 50.580 27.000 ;
        RECT 57.160 26.470 57.330 27.000 ;
        RECT 57.640 26.470 57.810 27.000 ;
        RECT 58.120 26.470 58.290 27.000 ;
        RECT 64.870 26.470 65.040 27.000 ;
        RECT 65.350 26.470 65.520 27.000 ;
        RECT 65.830 26.470 66.000 27.000 ;
        RECT 72.580 26.470 72.750 27.000 ;
        RECT 73.060 26.470 73.230 27.000 ;
        RECT 73.540 26.470 73.710 27.000 ;
        RECT 80.290 26.470 80.460 27.000 ;
        RECT 80.770 26.470 80.940 27.000 ;
        RECT 81.250 26.470 81.420 27.000 ;
        RECT 88.000 26.470 88.170 27.000 ;
        RECT 88.480 26.470 88.650 27.000 ;
        RECT 88.960 26.470 89.130 27.000 ;
        RECT 95.710 26.470 95.880 27.000 ;
        RECT 96.190 26.470 96.360 27.000 ;
        RECT 96.670 26.470 96.840 27.000 ;
        RECT 103.420 26.470 103.590 27.000 ;
        RECT 103.900 26.470 104.070 27.000 ;
        RECT 104.380 26.470 104.550 27.000 ;
        RECT 111.130 26.470 111.300 27.000 ;
        RECT 111.610 26.470 111.780 27.000 ;
        RECT 112.090 26.470 112.260 27.000 ;
        RECT 118.840 26.470 119.010 27.000 ;
        RECT 119.320 26.470 119.490 27.000 ;
        RECT 119.800 26.470 119.970 27.000 ;
        RECT 3.430 26.050 3.600 26.220 ;
        RECT 11.140 26.050 11.310 26.220 ;
        RECT 18.850 26.050 19.020 26.220 ;
        RECT 26.560 26.050 26.730 26.220 ;
        RECT 34.270 26.050 34.440 26.220 ;
        RECT 41.980 26.050 42.150 26.220 ;
        RECT 49.690 26.050 49.860 26.220 ;
        RECT 57.400 26.050 57.570 26.220 ;
        RECT 65.110 26.050 65.280 26.220 ;
        RECT 72.820 26.050 72.990 26.220 ;
        RECT 80.530 26.050 80.700 26.220 ;
        RECT 88.240 26.050 88.410 26.220 ;
        RECT 95.950 26.050 96.120 26.220 ;
        RECT 103.660 26.050 103.830 26.220 ;
        RECT 111.370 26.050 111.540 26.220 ;
        RECT 119.080 26.050 119.250 26.220 ;
        RECT 3.990 25.645 4.160 25.815 ;
        RECT 1.490 25.400 1.670 25.580 ;
        RECT 1.060 24.790 1.240 24.960 ;
        RECT 3.270 24.470 3.440 25.350 ;
        RECT 3.750 24.470 3.920 25.350 ;
        RECT 4.230 24.470 4.400 25.350 ;
        RECT 5.580 25.370 5.760 25.560 ;
        RECT 11.700 25.645 11.870 25.815 ;
        RECT 9.200 25.400 9.380 25.580 ;
        RECT 5.120 24.800 5.310 24.970 ;
        RECT 5.990 24.780 6.170 24.950 ;
        RECT 8.770 24.790 8.950 24.960 ;
        RECT 3.510 24.005 3.680 24.175 ;
        RECT 10.980 24.470 11.150 25.350 ;
        RECT 11.460 24.470 11.630 25.350 ;
        RECT 11.940 24.470 12.110 25.350 ;
        RECT 13.290 25.370 13.470 25.560 ;
        RECT 19.410 25.645 19.580 25.815 ;
        RECT 16.910 25.400 17.090 25.580 ;
        RECT 12.830 24.800 13.020 24.970 ;
        RECT 13.700 24.780 13.880 24.950 ;
        RECT 16.480 24.790 16.660 24.960 ;
        RECT 11.220 24.005 11.390 24.175 ;
        RECT 18.690 24.470 18.860 25.350 ;
        RECT 19.170 24.470 19.340 25.350 ;
        RECT 19.650 24.470 19.820 25.350 ;
        RECT 21.000 25.370 21.180 25.560 ;
        RECT 27.120 25.645 27.290 25.815 ;
        RECT 24.620 25.400 24.800 25.580 ;
        RECT 20.540 24.800 20.730 24.970 ;
        RECT 21.410 24.780 21.590 24.950 ;
        RECT 24.190 24.790 24.370 24.960 ;
        RECT 18.930 24.005 19.100 24.175 ;
        RECT 26.400 24.470 26.570 25.350 ;
        RECT 26.880 24.470 27.050 25.350 ;
        RECT 27.360 24.470 27.530 25.350 ;
        RECT 28.710 25.370 28.890 25.560 ;
        RECT 34.830 25.645 35.000 25.815 ;
        RECT 32.330 25.400 32.510 25.580 ;
        RECT 28.250 24.800 28.440 24.970 ;
        RECT 29.120 24.780 29.300 24.950 ;
        RECT 31.900 24.790 32.080 24.960 ;
        RECT 26.640 24.005 26.810 24.175 ;
        RECT 34.110 24.470 34.280 25.350 ;
        RECT 34.590 24.470 34.760 25.350 ;
        RECT 35.070 24.470 35.240 25.350 ;
        RECT 36.420 25.370 36.600 25.560 ;
        RECT 42.540 25.645 42.710 25.815 ;
        RECT 40.040 25.400 40.220 25.580 ;
        RECT 35.960 24.800 36.150 24.970 ;
        RECT 36.830 24.780 37.010 24.950 ;
        RECT 39.610 24.790 39.790 24.960 ;
        RECT 34.350 24.005 34.520 24.175 ;
        RECT 41.820 24.470 41.990 25.350 ;
        RECT 42.300 24.470 42.470 25.350 ;
        RECT 42.780 24.470 42.950 25.350 ;
        RECT 44.130 25.370 44.310 25.560 ;
        RECT 50.250 25.645 50.420 25.815 ;
        RECT 47.750 25.400 47.930 25.580 ;
        RECT 43.670 24.800 43.860 24.970 ;
        RECT 44.540 24.780 44.720 24.950 ;
        RECT 47.320 24.790 47.500 24.960 ;
        RECT 42.060 24.005 42.230 24.175 ;
        RECT 49.530 24.470 49.700 25.350 ;
        RECT 50.010 24.470 50.180 25.350 ;
        RECT 50.490 24.470 50.660 25.350 ;
        RECT 51.840 25.370 52.020 25.560 ;
        RECT 57.960 25.645 58.130 25.815 ;
        RECT 55.460 25.400 55.640 25.580 ;
        RECT 51.380 24.800 51.570 24.970 ;
        RECT 52.250 24.780 52.430 24.950 ;
        RECT 55.030 24.790 55.210 24.960 ;
        RECT 49.770 24.005 49.940 24.175 ;
        RECT 57.240 24.470 57.410 25.350 ;
        RECT 57.720 24.470 57.890 25.350 ;
        RECT 58.200 24.470 58.370 25.350 ;
        RECT 59.550 25.370 59.730 25.560 ;
        RECT 65.670 25.645 65.840 25.815 ;
        RECT 63.170 25.400 63.350 25.580 ;
        RECT 59.090 24.800 59.280 24.970 ;
        RECT 59.960 24.780 60.140 24.950 ;
        RECT 62.740 24.790 62.920 24.960 ;
        RECT 57.480 24.005 57.650 24.175 ;
        RECT 64.950 24.470 65.120 25.350 ;
        RECT 65.430 24.470 65.600 25.350 ;
        RECT 65.910 24.470 66.080 25.350 ;
        RECT 67.260 25.370 67.440 25.560 ;
        RECT 73.380 25.645 73.550 25.815 ;
        RECT 70.880 25.400 71.060 25.580 ;
        RECT 66.800 24.800 66.990 24.970 ;
        RECT 67.670 24.780 67.850 24.950 ;
        RECT 70.450 24.790 70.630 24.960 ;
        RECT 65.190 24.005 65.360 24.175 ;
        RECT 72.660 24.470 72.830 25.350 ;
        RECT 73.140 24.470 73.310 25.350 ;
        RECT 73.620 24.470 73.790 25.350 ;
        RECT 74.970 25.370 75.150 25.560 ;
        RECT 81.090 25.645 81.260 25.815 ;
        RECT 78.590 25.400 78.770 25.580 ;
        RECT 74.510 24.800 74.700 24.970 ;
        RECT 75.380 24.780 75.560 24.950 ;
        RECT 78.160 24.790 78.340 24.960 ;
        RECT 72.900 24.005 73.070 24.175 ;
        RECT 80.370 24.470 80.540 25.350 ;
        RECT 80.850 24.470 81.020 25.350 ;
        RECT 81.330 24.470 81.500 25.350 ;
        RECT 82.680 25.370 82.860 25.560 ;
        RECT 88.800 25.645 88.970 25.815 ;
        RECT 86.300 25.400 86.480 25.580 ;
        RECT 82.220 24.800 82.410 24.970 ;
        RECT 83.090 24.780 83.270 24.950 ;
        RECT 85.870 24.790 86.050 24.960 ;
        RECT 80.610 24.005 80.780 24.175 ;
        RECT 88.080 24.470 88.250 25.350 ;
        RECT 88.560 24.470 88.730 25.350 ;
        RECT 89.040 24.470 89.210 25.350 ;
        RECT 90.390 25.370 90.570 25.560 ;
        RECT 96.510 25.645 96.680 25.815 ;
        RECT 94.010 25.400 94.190 25.580 ;
        RECT 89.930 24.800 90.120 24.970 ;
        RECT 90.800 24.780 90.980 24.950 ;
        RECT 93.580 24.790 93.760 24.960 ;
        RECT 88.320 24.005 88.490 24.175 ;
        RECT 95.790 24.470 95.960 25.350 ;
        RECT 96.270 24.470 96.440 25.350 ;
        RECT 96.750 24.470 96.920 25.350 ;
        RECT 98.100 25.370 98.280 25.560 ;
        RECT 104.220 25.645 104.390 25.815 ;
        RECT 101.720 25.400 101.900 25.580 ;
        RECT 97.640 24.800 97.830 24.970 ;
        RECT 98.510 24.780 98.690 24.950 ;
        RECT 101.290 24.790 101.470 24.960 ;
        RECT 96.030 24.005 96.200 24.175 ;
        RECT 103.500 24.470 103.670 25.350 ;
        RECT 103.980 24.470 104.150 25.350 ;
        RECT 104.460 24.470 104.630 25.350 ;
        RECT 105.810 25.370 105.990 25.560 ;
        RECT 111.930 25.645 112.100 25.815 ;
        RECT 109.430 25.400 109.610 25.580 ;
        RECT 105.350 24.800 105.540 24.970 ;
        RECT 106.220 24.780 106.400 24.950 ;
        RECT 109.000 24.790 109.180 24.960 ;
        RECT 103.740 24.005 103.910 24.175 ;
        RECT 111.210 24.470 111.380 25.350 ;
        RECT 111.690 24.470 111.860 25.350 ;
        RECT 112.170 24.470 112.340 25.350 ;
        RECT 113.520 25.370 113.700 25.560 ;
        RECT 119.640 25.645 119.810 25.815 ;
        RECT 117.140 25.400 117.320 25.580 ;
        RECT 113.060 24.800 113.250 24.970 ;
        RECT 113.930 24.780 114.110 24.950 ;
        RECT 116.710 24.790 116.890 24.960 ;
        RECT 111.450 24.005 111.620 24.175 ;
        RECT 118.920 24.470 119.090 25.350 ;
        RECT 119.400 24.470 119.570 25.350 ;
        RECT 119.880 24.470 120.050 25.350 ;
        RECT 121.230 25.370 121.410 25.560 ;
        RECT 120.770 24.800 120.960 24.970 ;
        RECT 121.640 24.780 121.820 24.950 ;
        RECT 119.160 24.005 119.330 24.175 ;
        RECT 28.720 20.610 28.950 20.840 ;
        RECT 90.380 20.620 90.600 20.820 ;
        RECT 58.570 19.890 58.740 20.060 ;
        RECT 59.060 16.490 59.240 16.680 ;
        RECT 58.570 15.860 58.760 16.040 ;
        RECT 124.580 15.880 124.800 16.070 ;
        RECT 58.500 13.680 58.670 13.860 ;
        RECT 28.840 11.940 29.070 12.230 ;
        RECT 90.490 11.990 90.750 12.220 ;
        RECT 3.710 9.285 3.880 9.455 ;
        RECT 1.220 8.510 1.400 8.680 ;
        RECT 2.080 8.490 2.270 8.660 ;
        RECT 1.630 7.900 1.810 8.090 ;
        RECT 2.990 8.110 3.160 8.990 ;
        RECT 3.470 8.110 3.640 8.990 ;
        RECT 3.950 8.110 4.120 8.990 ;
        RECT 11.420 9.285 11.590 9.455 ;
        RECT 6.150 8.500 6.330 8.670 ;
        RECT 8.930 8.510 9.110 8.680 ;
        RECT 9.790 8.490 9.980 8.660 ;
        RECT 5.720 7.880 5.900 8.060 ;
        RECT 3.230 7.645 3.400 7.815 ;
        RECT 9.340 7.900 9.520 8.090 ;
        RECT 10.700 8.110 10.870 8.990 ;
        RECT 11.180 8.110 11.350 8.990 ;
        RECT 11.660 8.110 11.830 8.990 ;
        RECT 19.130 9.285 19.300 9.455 ;
        RECT 13.860 8.500 14.040 8.670 ;
        RECT 16.640 8.510 16.820 8.680 ;
        RECT 17.500 8.490 17.690 8.660 ;
        RECT 13.430 7.880 13.610 8.060 ;
        RECT 10.940 7.645 11.110 7.815 ;
        RECT 17.050 7.900 17.230 8.090 ;
        RECT 18.410 8.110 18.580 8.990 ;
        RECT 18.890 8.110 19.060 8.990 ;
        RECT 19.370 8.110 19.540 8.990 ;
        RECT 26.840 9.285 27.010 9.455 ;
        RECT 21.570 8.500 21.750 8.670 ;
        RECT 24.350 8.510 24.530 8.680 ;
        RECT 25.210 8.490 25.400 8.660 ;
        RECT 21.140 7.880 21.320 8.060 ;
        RECT 18.650 7.645 18.820 7.815 ;
        RECT 24.760 7.900 24.940 8.090 ;
        RECT 26.120 8.110 26.290 8.990 ;
        RECT 26.600 8.110 26.770 8.990 ;
        RECT 27.080 8.110 27.250 8.990 ;
        RECT 34.550 9.285 34.720 9.455 ;
        RECT 29.280 8.500 29.460 8.670 ;
        RECT 32.060 8.510 32.240 8.680 ;
        RECT 32.920 8.490 33.110 8.660 ;
        RECT 28.850 7.880 29.030 8.060 ;
        RECT 26.360 7.645 26.530 7.815 ;
        RECT 32.470 7.900 32.650 8.090 ;
        RECT 33.830 8.110 34.000 8.990 ;
        RECT 34.310 8.110 34.480 8.990 ;
        RECT 34.790 8.110 34.960 8.990 ;
        RECT 42.260 9.285 42.430 9.455 ;
        RECT 36.990 8.500 37.170 8.670 ;
        RECT 39.770 8.510 39.950 8.680 ;
        RECT 40.630 8.490 40.820 8.660 ;
        RECT 36.560 7.880 36.740 8.060 ;
        RECT 34.070 7.645 34.240 7.815 ;
        RECT 40.180 7.900 40.360 8.090 ;
        RECT 41.540 8.110 41.710 8.990 ;
        RECT 42.020 8.110 42.190 8.990 ;
        RECT 42.500 8.110 42.670 8.990 ;
        RECT 49.970 9.285 50.140 9.455 ;
        RECT 44.700 8.500 44.880 8.670 ;
        RECT 47.480 8.510 47.660 8.680 ;
        RECT 48.340 8.490 48.530 8.660 ;
        RECT 44.270 7.880 44.450 8.060 ;
        RECT 41.780 7.645 41.950 7.815 ;
        RECT 47.890 7.900 48.070 8.090 ;
        RECT 49.250 8.110 49.420 8.990 ;
        RECT 49.730 8.110 49.900 8.990 ;
        RECT 50.210 8.110 50.380 8.990 ;
        RECT 57.680 9.285 57.850 9.455 ;
        RECT 52.410 8.500 52.590 8.670 ;
        RECT 55.190 8.510 55.370 8.680 ;
        RECT 56.050 8.490 56.240 8.660 ;
        RECT 51.980 7.880 52.160 8.060 ;
        RECT 49.490 7.645 49.660 7.815 ;
        RECT 55.600 7.900 55.780 8.090 ;
        RECT 56.960 8.110 57.130 8.990 ;
        RECT 57.440 8.110 57.610 8.990 ;
        RECT 57.920 8.110 58.090 8.990 ;
        RECT 65.390 9.285 65.560 9.455 ;
        RECT 60.120 8.500 60.300 8.670 ;
        RECT 62.900 8.510 63.080 8.680 ;
        RECT 63.760 8.490 63.950 8.660 ;
        RECT 59.690 7.880 59.870 8.060 ;
        RECT 57.200 7.645 57.370 7.815 ;
        RECT 63.310 7.900 63.490 8.090 ;
        RECT 64.670 8.110 64.840 8.990 ;
        RECT 65.150 8.110 65.320 8.990 ;
        RECT 65.630 8.110 65.800 8.990 ;
        RECT 73.100 9.285 73.270 9.455 ;
        RECT 67.830 8.500 68.010 8.670 ;
        RECT 70.610 8.510 70.790 8.680 ;
        RECT 71.470 8.490 71.660 8.660 ;
        RECT 67.400 7.880 67.580 8.060 ;
        RECT 64.910 7.645 65.080 7.815 ;
        RECT 71.020 7.900 71.200 8.090 ;
        RECT 72.380 8.110 72.550 8.990 ;
        RECT 72.860 8.110 73.030 8.990 ;
        RECT 73.340 8.110 73.510 8.990 ;
        RECT 80.810 9.285 80.980 9.455 ;
        RECT 75.540 8.500 75.720 8.670 ;
        RECT 78.320 8.510 78.500 8.680 ;
        RECT 79.180 8.490 79.370 8.660 ;
        RECT 75.110 7.880 75.290 8.060 ;
        RECT 72.620 7.645 72.790 7.815 ;
        RECT 78.730 7.900 78.910 8.090 ;
        RECT 80.090 8.110 80.260 8.990 ;
        RECT 80.570 8.110 80.740 8.990 ;
        RECT 81.050 8.110 81.220 8.990 ;
        RECT 88.520 9.285 88.690 9.455 ;
        RECT 83.250 8.500 83.430 8.670 ;
        RECT 86.030 8.510 86.210 8.680 ;
        RECT 86.890 8.490 87.080 8.660 ;
        RECT 82.820 7.880 83.000 8.060 ;
        RECT 80.330 7.645 80.500 7.815 ;
        RECT 86.440 7.900 86.620 8.090 ;
        RECT 87.800 8.110 87.970 8.990 ;
        RECT 88.280 8.110 88.450 8.990 ;
        RECT 88.760 8.110 88.930 8.990 ;
        RECT 96.230 9.285 96.400 9.455 ;
        RECT 90.960 8.500 91.140 8.670 ;
        RECT 93.740 8.510 93.920 8.680 ;
        RECT 94.600 8.490 94.790 8.660 ;
        RECT 90.530 7.880 90.710 8.060 ;
        RECT 88.040 7.645 88.210 7.815 ;
        RECT 94.150 7.900 94.330 8.090 ;
        RECT 95.510 8.110 95.680 8.990 ;
        RECT 95.990 8.110 96.160 8.990 ;
        RECT 96.470 8.110 96.640 8.990 ;
        RECT 103.940 9.285 104.110 9.455 ;
        RECT 98.670 8.500 98.850 8.670 ;
        RECT 101.450 8.510 101.630 8.680 ;
        RECT 102.310 8.490 102.500 8.660 ;
        RECT 98.240 7.880 98.420 8.060 ;
        RECT 95.750 7.645 95.920 7.815 ;
        RECT 101.860 7.900 102.040 8.090 ;
        RECT 103.220 8.110 103.390 8.990 ;
        RECT 103.700 8.110 103.870 8.990 ;
        RECT 104.180 8.110 104.350 8.990 ;
        RECT 111.650 9.285 111.820 9.455 ;
        RECT 106.380 8.500 106.560 8.670 ;
        RECT 109.160 8.510 109.340 8.680 ;
        RECT 110.020 8.490 110.210 8.660 ;
        RECT 105.950 7.880 106.130 8.060 ;
        RECT 103.460 7.645 103.630 7.815 ;
        RECT 109.570 7.900 109.750 8.090 ;
        RECT 110.930 8.110 111.100 8.990 ;
        RECT 111.410 8.110 111.580 8.990 ;
        RECT 111.890 8.110 112.060 8.990 ;
        RECT 119.360 9.285 119.530 9.455 ;
        RECT 114.090 8.500 114.270 8.670 ;
        RECT 116.870 8.510 117.050 8.680 ;
        RECT 117.730 8.490 117.920 8.660 ;
        RECT 113.660 7.880 113.840 8.060 ;
        RECT 111.170 7.645 111.340 7.815 ;
        RECT 117.280 7.900 117.460 8.090 ;
        RECT 118.640 8.110 118.810 8.990 ;
        RECT 119.120 8.110 119.290 8.990 ;
        RECT 119.600 8.110 119.770 8.990 ;
        RECT 121.800 8.500 121.980 8.670 ;
        RECT 121.370 7.880 121.550 8.060 ;
        RECT 118.880 7.645 119.050 7.815 ;
        RECT 3.790 7.240 3.960 7.410 ;
        RECT 11.500 7.240 11.670 7.410 ;
        RECT 19.210 7.240 19.380 7.410 ;
        RECT 26.920 7.240 27.090 7.410 ;
        RECT 34.630 7.240 34.800 7.410 ;
        RECT 42.340 7.240 42.510 7.410 ;
        RECT 50.050 7.240 50.220 7.410 ;
        RECT 57.760 7.240 57.930 7.410 ;
        RECT 65.470 7.240 65.640 7.410 ;
        RECT 73.180 7.240 73.350 7.410 ;
        RECT 80.890 7.240 81.060 7.410 ;
        RECT 88.600 7.240 88.770 7.410 ;
        RECT 96.310 7.240 96.480 7.410 ;
        RECT 104.020 7.240 104.190 7.410 ;
        RECT 111.730 7.240 111.900 7.410 ;
        RECT 119.440 7.240 119.610 7.410 ;
        RECT 3.070 6.460 3.240 6.990 ;
        RECT 3.550 6.460 3.720 6.990 ;
        RECT 4.030 6.460 4.200 6.990 ;
        RECT 10.780 6.460 10.950 6.990 ;
        RECT 11.260 6.460 11.430 6.990 ;
        RECT 11.740 6.460 11.910 6.990 ;
        RECT 18.490 6.460 18.660 6.990 ;
        RECT 18.970 6.460 19.140 6.990 ;
        RECT 19.450 6.460 19.620 6.990 ;
        RECT 26.200 6.460 26.370 6.990 ;
        RECT 26.680 6.460 26.850 6.990 ;
        RECT 27.160 6.460 27.330 6.990 ;
        RECT 33.910 6.460 34.080 6.990 ;
        RECT 34.390 6.460 34.560 6.990 ;
        RECT 34.870 6.460 35.040 6.990 ;
        RECT 41.620 6.460 41.790 6.990 ;
        RECT 42.100 6.460 42.270 6.990 ;
        RECT 42.580 6.460 42.750 6.990 ;
        RECT 49.330 6.460 49.500 6.990 ;
        RECT 49.810 6.460 49.980 6.990 ;
        RECT 50.290 6.460 50.460 6.990 ;
        RECT 57.040 6.460 57.210 6.990 ;
        RECT 57.520 6.460 57.690 6.990 ;
        RECT 58.000 6.460 58.170 6.990 ;
        RECT 64.750 6.460 64.920 6.990 ;
        RECT 65.230 6.460 65.400 6.990 ;
        RECT 65.710 6.460 65.880 6.990 ;
        RECT 72.460 6.460 72.630 6.990 ;
        RECT 72.940 6.460 73.110 6.990 ;
        RECT 73.420 6.460 73.590 6.990 ;
        RECT 80.170 6.460 80.340 6.990 ;
        RECT 80.650 6.460 80.820 6.990 ;
        RECT 81.130 6.460 81.300 6.990 ;
        RECT 87.880 6.460 88.050 6.990 ;
        RECT 88.360 6.460 88.530 6.990 ;
        RECT 88.840 6.460 89.010 6.990 ;
        RECT 95.590 6.460 95.760 6.990 ;
        RECT 96.070 6.460 96.240 6.990 ;
        RECT 96.550 6.460 96.720 6.990 ;
        RECT 103.300 6.460 103.470 6.990 ;
        RECT 103.780 6.460 103.950 6.990 ;
        RECT 104.260 6.460 104.430 6.990 ;
        RECT 111.010 6.460 111.180 6.990 ;
        RECT 111.490 6.460 111.660 6.990 ;
        RECT 111.970 6.460 112.140 6.990 ;
        RECT 118.720 6.460 118.890 6.990 ;
        RECT 119.200 6.460 119.370 6.990 ;
        RECT 119.680 6.460 119.850 6.990 ;
        RECT 3.310 6.040 3.480 6.210 ;
        RECT 2.120 4.805 2.290 4.975 ;
        RECT 5.350 4.805 5.520 4.975 ;
        RECT 11.020 6.040 11.190 6.210 ;
        RECT 9.830 4.805 10.000 4.975 ;
        RECT 13.060 4.805 13.230 4.975 ;
        RECT 1.900 3.630 2.070 4.510 ;
        RECT 3.700 4.005 3.870 4.175 ;
        RECT 2.120 3.165 2.290 3.335 ;
        RECT 2.980 2.830 3.150 3.710 ;
        RECT 3.460 2.830 3.630 3.710 ;
        RECT 3.940 2.830 4.110 3.710 ;
        RECT 5.570 3.630 5.740 4.510 ;
        RECT 5.350 3.165 5.520 3.335 ;
        RECT 18.730 6.040 18.900 6.210 ;
        RECT 17.540 4.805 17.710 4.975 ;
        RECT 20.770 4.805 20.940 4.975 ;
        RECT 3.220 2.365 3.390 2.535 ;
        RECT 9.610 3.630 9.780 4.510 ;
        RECT 11.410 4.005 11.580 4.175 ;
        RECT 9.830 3.165 10.000 3.335 ;
        RECT 6.940 2.730 7.110 2.900 ;
        RECT 10.690 2.830 10.860 3.710 ;
        RECT 11.170 2.830 11.340 3.710 ;
        RECT 11.650 2.830 11.820 3.710 ;
        RECT 13.280 3.630 13.450 4.510 ;
        RECT 13.060 3.165 13.230 3.335 ;
        RECT 26.440 6.040 26.610 6.210 ;
        RECT 25.250 4.805 25.420 4.975 ;
        RECT 28.480 4.805 28.650 4.975 ;
        RECT 10.930 2.365 11.100 2.535 ;
        RECT 5.130 2.150 5.320 2.320 ;
        RECT 3.780 1.960 3.950 2.130 ;
        RECT 17.320 3.630 17.490 4.510 ;
        RECT 19.120 4.005 19.290 4.175 ;
        RECT 17.540 3.165 17.710 3.335 ;
        RECT 14.650 2.730 14.820 2.900 ;
        RECT 18.400 2.830 18.570 3.710 ;
        RECT 18.880 2.830 19.050 3.710 ;
        RECT 19.360 2.830 19.530 3.710 ;
        RECT 20.990 3.630 21.160 4.510 ;
        RECT 20.770 3.165 20.940 3.335 ;
        RECT 34.150 6.040 34.320 6.210 ;
        RECT 32.960 4.805 33.130 4.975 ;
        RECT 36.190 4.805 36.360 4.975 ;
        RECT 18.640 2.365 18.810 2.535 ;
        RECT 12.840 2.150 13.030 2.320 ;
        RECT 11.490 1.960 11.660 2.130 ;
        RECT 25.030 3.630 25.200 4.510 ;
        RECT 26.830 4.005 27.000 4.175 ;
        RECT 25.250 3.165 25.420 3.335 ;
        RECT 22.360 2.730 22.530 2.900 ;
        RECT 26.110 2.830 26.280 3.710 ;
        RECT 26.590 2.830 26.760 3.710 ;
        RECT 27.070 2.830 27.240 3.710 ;
        RECT 28.700 3.630 28.870 4.510 ;
        RECT 28.480 3.165 28.650 3.335 ;
        RECT 41.860 6.040 42.030 6.210 ;
        RECT 40.670 4.805 40.840 4.975 ;
        RECT 43.900 4.805 44.070 4.975 ;
        RECT 26.350 2.365 26.520 2.535 ;
        RECT 20.550 2.150 20.740 2.320 ;
        RECT 19.200 1.960 19.370 2.130 ;
        RECT 32.740 3.630 32.910 4.510 ;
        RECT 34.540 4.005 34.710 4.175 ;
        RECT 32.960 3.165 33.130 3.335 ;
        RECT 30.070 2.730 30.240 2.900 ;
        RECT 33.820 2.830 33.990 3.710 ;
        RECT 34.300 2.830 34.470 3.710 ;
        RECT 34.780 2.830 34.950 3.710 ;
        RECT 36.410 3.630 36.580 4.510 ;
        RECT 36.190 3.165 36.360 3.335 ;
        RECT 49.570 6.040 49.740 6.210 ;
        RECT 48.380 4.805 48.550 4.975 ;
        RECT 51.610 4.805 51.780 4.975 ;
        RECT 34.060 2.365 34.230 2.535 ;
        RECT 28.260 2.150 28.450 2.320 ;
        RECT 26.910 1.960 27.080 2.130 ;
        RECT 40.450 3.630 40.620 4.510 ;
        RECT 42.250 4.005 42.420 4.175 ;
        RECT 40.670 3.165 40.840 3.335 ;
        RECT 37.780 2.730 37.950 2.900 ;
        RECT 41.530 2.830 41.700 3.710 ;
        RECT 42.010 2.830 42.180 3.710 ;
        RECT 42.490 2.830 42.660 3.710 ;
        RECT 44.120 3.630 44.290 4.510 ;
        RECT 43.900 3.165 44.070 3.335 ;
        RECT 57.280 6.040 57.450 6.210 ;
        RECT 56.090 4.805 56.260 4.975 ;
        RECT 59.320 4.805 59.490 4.975 ;
        RECT 41.770 2.365 41.940 2.535 ;
        RECT 35.970 2.150 36.160 2.320 ;
        RECT 34.620 1.960 34.790 2.130 ;
        RECT 48.160 3.630 48.330 4.510 ;
        RECT 49.960 4.005 50.130 4.175 ;
        RECT 48.380 3.165 48.550 3.335 ;
        RECT 45.490 2.730 45.660 2.900 ;
        RECT 49.240 2.830 49.410 3.710 ;
        RECT 49.720 2.830 49.890 3.710 ;
        RECT 50.200 2.830 50.370 3.710 ;
        RECT 51.830 3.630 52.000 4.510 ;
        RECT 51.610 3.165 51.780 3.335 ;
        RECT 64.990 6.040 65.160 6.210 ;
        RECT 63.800 4.805 63.970 4.975 ;
        RECT 67.030 4.805 67.200 4.975 ;
        RECT 49.480 2.365 49.650 2.535 ;
        RECT 43.680 2.150 43.870 2.320 ;
        RECT 42.330 1.960 42.500 2.130 ;
        RECT 55.870 3.630 56.040 4.510 ;
        RECT 57.670 4.005 57.840 4.175 ;
        RECT 56.090 3.165 56.260 3.335 ;
        RECT 53.200 2.730 53.370 2.900 ;
        RECT 56.950 2.830 57.120 3.710 ;
        RECT 57.430 2.830 57.600 3.710 ;
        RECT 57.910 2.830 58.080 3.710 ;
        RECT 59.540 3.630 59.710 4.510 ;
        RECT 59.320 3.165 59.490 3.335 ;
        RECT 72.700 6.040 72.870 6.210 ;
        RECT 71.510 4.805 71.680 4.975 ;
        RECT 74.740 4.805 74.910 4.975 ;
        RECT 57.190 2.365 57.360 2.535 ;
        RECT 51.390 2.150 51.580 2.320 ;
        RECT 50.040 1.960 50.210 2.130 ;
        RECT 63.580 3.630 63.750 4.510 ;
        RECT 65.380 4.005 65.550 4.175 ;
        RECT 63.800 3.165 63.970 3.335 ;
        RECT 60.910 2.730 61.080 2.900 ;
        RECT 64.660 2.830 64.830 3.710 ;
        RECT 65.140 2.830 65.310 3.710 ;
        RECT 65.620 2.830 65.790 3.710 ;
        RECT 67.250 3.630 67.420 4.510 ;
        RECT 67.030 3.165 67.200 3.335 ;
        RECT 80.410 6.040 80.580 6.210 ;
        RECT 79.220 4.805 79.390 4.975 ;
        RECT 82.450 4.805 82.620 4.975 ;
        RECT 64.900 2.365 65.070 2.535 ;
        RECT 59.100 2.150 59.290 2.320 ;
        RECT 57.750 1.960 57.920 2.130 ;
        RECT 71.290 3.630 71.460 4.510 ;
        RECT 73.090 4.005 73.260 4.175 ;
        RECT 71.510 3.165 71.680 3.335 ;
        RECT 68.620 2.730 68.790 2.900 ;
        RECT 72.370 2.830 72.540 3.710 ;
        RECT 72.850 2.830 73.020 3.710 ;
        RECT 73.330 2.830 73.500 3.710 ;
        RECT 74.960 3.630 75.130 4.510 ;
        RECT 74.740 3.165 74.910 3.335 ;
        RECT 88.120 6.040 88.290 6.210 ;
        RECT 86.930 4.805 87.100 4.975 ;
        RECT 90.160 4.805 90.330 4.975 ;
        RECT 72.610 2.365 72.780 2.535 ;
        RECT 66.810 2.150 67.000 2.320 ;
        RECT 65.460 1.960 65.630 2.130 ;
        RECT 79.000 3.630 79.170 4.510 ;
        RECT 80.800 4.005 80.970 4.175 ;
        RECT 79.220 3.165 79.390 3.335 ;
        RECT 76.330 2.730 76.500 2.900 ;
        RECT 80.080 2.830 80.250 3.710 ;
        RECT 80.560 2.830 80.730 3.710 ;
        RECT 81.040 2.830 81.210 3.710 ;
        RECT 82.670 3.630 82.840 4.510 ;
        RECT 82.450 3.165 82.620 3.335 ;
        RECT 95.830 6.040 96.000 6.210 ;
        RECT 94.640 4.805 94.810 4.975 ;
        RECT 97.870 4.805 98.040 4.975 ;
        RECT 80.320 2.365 80.490 2.535 ;
        RECT 74.520 2.150 74.710 2.320 ;
        RECT 73.170 1.960 73.340 2.130 ;
        RECT 86.710 3.630 86.880 4.510 ;
        RECT 88.510 4.005 88.680 4.175 ;
        RECT 86.930 3.165 87.100 3.335 ;
        RECT 84.040 2.730 84.210 2.900 ;
        RECT 87.790 2.830 87.960 3.710 ;
        RECT 88.270 2.830 88.440 3.710 ;
        RECT 88.750 2.830 88.920 3.710 ;
        RECT 90.380 3.630 90.550 4.510 ;
        RECT 90.160 3.165 90.330 3.335 ;
        RECT 103.540 6.040 103.710 6.210 ;
        RECT 102.350 4.805 102.520 4.975 ;
        RECT 105.580 4.805 105.750 4.975 ;
        RECT 88.030 2.365 88.200 2.535 ;
        RECT 82.230 2.150 82.420 2.320 ;
        RECT 80.880 1.960 81.050 2.130 ;
        RECT 94.420 3.630 94.590 4.510 ;
        RECT 96.220 4.005 96.390 4.175 ;
        RECT 94.640 3.165 94.810 3.335 ;
        RECT 91.750 2.730 91.920 2.900 ;
        RECT 95.500 2.830 95.670 3.710 ;
        RECT 95.980 2.830 96.150 3.710 ;
        RECT 96.460 2.830 96.630 3.710 ;
        RECT 98.090 3.630 98.260 4.510 ;
        RECT 97.870 3.165 98.040 3.335 ;
        RECT 111.250 6.040 111.420 6.210 ;
        RECT 110.060 4.805 110.230 4.975 ;
        RECT 113.290 4.805 113.460 4.975 ;
        RECT 95.740 2.365 95.910 2.535 ;
        RECT 89.940 2.150 90.130 2.320 ;
        RECT 88.590 1.960 88.760 2.130 ;
        RECT 102.130 3.630 102.300 4.510 ;
        RECT 103.930 4.005 104.100 4.175 ;
        RECT 102.350 3.165 102.520 3.335 ;
        RECT 99.460 2.730 99.630 2.900 ;
        RECT 103.210 2.830 103.380 3.710 ;
        RECT 103.690 2.830 103.860 3.710 ;
        RECT 104.170 2.830 104.340 3.710 ;
        RECT 105.800 3.630 105.970 4.510 ;
        RECT 105.580 3.165 105.750 3.335 ;
        RECT 118.960 6.040 119.130 6.210 ;
        RECT 117.770 4.805 117.940 4.975 ;
        RECT 121.000 4.805 121.170 4.975 ;
        RECT 103.450 2.365 103.620 2.535 ;
        RECT 97.650 2.150 97.840 2.320 ;
        RECT 96.300 1.960 96.470 2.130 ;
        RECT 109.840 3.630 110.010 4.510 ;
        RECT 111.640 4.005 111.810 4.175 ;
        RECT 110.060 3.165 110.230 3.335 ;
        RECT 107.170 2.730 107.340 2.900 ;
        RECT 110.920 2.830 111.090 3.710 ;
        RECT 111.400 2.830 111.570 3.710 ;
        RECT 111.880 2.830 112.050 3.710 ;
        RECT 113.510 3.630 113.680 4.510 ;
        RECT 113.290 3.165 113.460 3.335 ;
        RECT 111.160 2.365 111.330 2.535 ;
        RECT 105.360 2.150 105.550 2.320 ;
        RECT 104.010 1.960 104.180 2.130 ;
        RECT 117.550 3.630 117.720 4.510 ;
        RECT 119.350 4.005 119.520 4.175 ;
        RECT 117.770 3.165 117.940 3.335 ;
        RECT 114.880 2.730 115.050 2.900 ;
        RECT 118.630 2.830 118.800 3.710 ;
        RECT 119.110 2.830 119.280 3.710 ;
        RECT 119.590 2.830 119.760 3.710 ;
        RECT 121.220 3.630 121.390 4.510 ;
        RECT 121.000 3.165 121.170 3.335 ;
        RECT 118.870 2.365 119.040 2.535 ;
        RECT 113.070 2.150 113.260 2.320 ;
        RECT 111.720 1.960 111.890 2.130 ;
        RECT 122.590 2.730 122.760 2.900 ;
        RECT 120.780 2.150 120.970 2.320 ;
        RECT 119.430 1.960 119.600 2.130 ;
        RECT 3.060 1.180 3.230 1.710 ;
        RECT 3.540 1.180 3.710 1.710 ;
        RECT 4.020 1.180 4.190 1.710 ;
        RECT 10.770 1.180 10.940 1.710 ;
        RECT 11.250 1.180 11.420 1.710 ;
        RECT 11.730 1.180 11.900 1.710 ;
        RECT 18.480 1.180 18.650 1.710 ;
        RECT 18.960 1.180 19.130 1.710 ;
        RECT 19.440 1.180 19.610 1.710 ;
        RECT 26.190 1.180 26.360 1.710 ;
        RECT 26.670 1.180 26.840 1.710 ;
        RECT 27.150 1.180 27.320 1.710 ;
        RECT 33.900 1.180 34.070 1.710 ;
        RECT 34.380 1.180 34.550 1.710 ;
        RECT 34.860 1.180 35.030 1.710 ;
        RECT 41.610 1.180 41.780 1.710 ;
        RECT 42.090 1.180 42.260 1.710 ;
        RECT 42.570 1.180 42.740 1.710 ;
        RECT 49.320 1.180 49.490 1.710 ;
        RECT 49.800 1.180 49.970 1.710 ;
        RECT 50.280 1.180 50.450 1.710 ;
        RECT 57.030 1.180 57.200 1.710 ;
        RECT 57.510 1.180 57.680 1.710 ;
        RECT 57.990 1.180 58.160 1.710 ;
        RECT 64.740 1.180 64.910 1.710 ;
        RECT 65.220 1.180 65.390 1.710 ;
        RECT 65.700 1.180 65.870 1.710 ;
        RECT 72.450 1.180 72.620 1.710 ;
        RECT 72.930 1.180 73.100 1.710 ;
        RECT 73.410 1.180 73.580 1.710 ;
        RECT 80.160 1.180 80.330 1.710 ;
        RECT 80.640 1.180 80.810 1.710 ;
        RECT 81.120 1.180 81.290 1.710 ;
        RECT 87.870 1.180 88.040 1.710 ;
        RECT 88.350 1.180 88.520 1.710 ;
        RECT 88.830 1.180 89.000 1.710 ;
        RECT 95.580 1.180 95.750 1.710 ;
        RECT 96.060 1.180 96.230 1.710 ;
        RECT 96.540 1.180 96.710 1.710 ;
        RECT 103.290 1.180 103.460 1.710 ;
        RECT 103.770 1.180 103.940 1.710 ;
        RECT 104.250 1.180 104.420 1.710 ;
        RECT 111.000 1.180 111.170 1.710 ;
        RECT 111.480 1.180 111.650 1.710 ;
        RECT 111.960 1.180 112.130 1.710 ;
        RECT 118.710 1.180 118.880 1.710 ;
        RECT 119.190 1.180 119.360 1.710 ;
        RECT 119.670 1.180 119.840 1.710 ;
        RECT 3.300 0.760 3.470 0.930 ;
        RECT 11.010 0.760 11.180 0.930 ;
        RECT 18.720 0.760 18.890 0.930 ;
        RECT 26.430 0.760 26.600 0.930 ;
        RECT 34.140 0.760 34.310 0.930 ;
        RECT 41.850 0.760 42.020 0.930 ;
        RECT 49.560 0.760 49.730 0.930 ;
        RECT 57.270 0.760 57.440 0.930 ;
        RECT 64.980 0.760 65.150 0.930 ;
        RECT 72.690 0.760 72.860 0.930 ;
        RECT 80.400 0.760 80.570 0.930 ;
        RECT 88.110 0.760 88.280 0.930 ;
        RECT 95.820 0.760 95.990 0.930 ;
        RECT 103.530 0.760 103.700 0.930 ;
        RECT 111.240 0.760 111.410 0.930 ;
        RECT 118.950 0.760 119.120 0.930 ;
      LAYER met1 ;
        RECT 2.560 32.480 4.160 32.790 ;
        RECT 10.270 32.480 11.870 32.790 ;
        RECT 17.980 32.480 19.580 32.790 ;
        RECT 25.690 32.480 27.290 32.790 ;
        RECT 33.400 32.480 35.000 32.790 ;
        RECT 41.110 32.480 42.710 32.790 ;
        RECT 48.820 32.480 50.420 32.790 ;
        RECT 56.530 32.480 58.130 32.790 ;
        RECT 64.240 32.480 65.840 32.790 ;
        RECT 71.950 32.480 73.550 32.790 ;
        RECT 79.660 32.480 81.260 32.790 ;
        RECT 87.370 32.480 88.970 32.790 ;
        RECT 95.080 32.480 96.680 32.790 ;
        RECT 102.790 32.480 104.390 32.790 ;
        RECT 110.500 32.480 112.100 32.790 ;
        RECT 118.210 32.480 119.810 32.790 ;
        RECT 1.950 31.050 2.330 31.370 ;
        RECT 2.560 30.830 2.860 32.480 ;
        RECT 3.170 32.280 3.400 32.340 ;
        RECT 0.220 30.660 2.860 30.830 ;
        RECT 0.220 30.490 0.510 30.660 ;
        RECT 1.790 30.060 2.120 30.340 ;
        RECT 1.620 28.890 1.850 29.890 ;
        RECT 2.560 29.500 2.860 30.660 ;
        RECT 3.000 31.690 3.400 32.280 ;
        RECT 3.600 32.020 3.930 32.340 ;
        RECT 3.650 31.690 3.880 32.020 ;
        RECT 4.130 31.690 4.640 32.340 ;
        RECT 3.000 30.690 3.230 31.690 ;
        RECT 3.380 31.240 3.670 31.550 ;
        RECT 4.390 31.290 4.640 31.690 ;
        RECT 3.940 30.850 4.230 31.180 ;
        RECT 4.390 30.960 4.740 31.290 ;
        RECT 9.660 31.050 10.040 31.370 ;
        RECT 4.390 30.690 4.640 30.960 ;
        RECT 10.270 30.830 10.570 32.480 ;
        RECT 10.880 32.280 11.110 32.340 ;
        RECT 3.000 29.690 3.480 30.690 ;
        RECT 3.730 29.990 3.960 30.690 ;
        RECT 3.680 29.650 4.010 29.990 ;
        RECT 4.210 29.710 4.640 30.690 ;
        RECT 7.930 30.660 10.570 30.830 ;
        RECT 7.930 30.490 8.220 30.660 ;
        RECT 5.020 30.070 5.350 30.360 ;
        RECT 9.500 30.060 9.830 30.340 ;
        RECT 4.210 29.690 4.440 29.710 ;
        RECT 2.560 29.340 3.750 29.500 ;
        RECT 2.550 29.200 3.750 29.340 ;
        RECT 1.790 28.430 2.120 28.710 ;
        RECT 2.550 28.470 2.720 29.200 ;
        RECT 3.460 29.190 3.750 29.200 ;
        RECT 5.290 29.020 5.520 29.890 ;
        RECT 5.290 28.880 5.650 29.020 ;
        RECT 9.330 28.890 9.560 29.890 ;
        RECT 10.270 29.500 10.570 30.660 ;
        RECT 10.710 31.690 11.110 32.280 ;
        RECT 11.310 32.020 11.640 32.340 ;
        RECT 11.360 31.690 11.590 32.020 ;
        RECT 11.840 31.690 12.350 32.340 ;
        RECT 10.710 30.690 10.940 31.690 ;
        RECT 11.090 31.240 11.380 31.550 ;
        RECT 12.100 31.290 12.350 31.690 ;
        RECT 11.650 30.850 11.940 31.180 ;
        RECT 12.100 30.960 12.450 31.290 ;
        RECT 17.370 31.050 17.750 31.370 ;
        RECT 12.100 30.690 12.350 30.960 ;
        RECT 17.980 30.830 18.280 32.480 ;
        RECT 18.590 32.280 18.820 32.340 ;
        RECT 10.710 29.690 11.190 30.690 ;
        RECT 11.440 29.990 11.670 30.690 ;
        RECT 11.390 29.650 11.720 29.990 ;
        RECT 11.920 29.710 12.350 30.690 ;
        RECT 15.640 30.660 18.280 30.830 ;
        RECT 15.640 30.490 15.930 30.660 ;
        RECT 12.730 30.070 13.060 30.360 ;
        RECT 17.210 30.060 17.540 30.340 ;
        RECT 11.920 29.690 12.150 29.710 ;
        RECT 10.270 29.340 11.460 29.500 ;
        RECT 10.260 29.200 11.460 29.340 ;
        RECT 5.020 28.470 5.350 28.700 ;
        RECT 2.550 28.330 5.350 28.470 ;
        RECT 2.550 27.510 2.720 28.330 ;
        RECT 2.550 27.200 4.150 27.510 ;
        RECT 1.420 25.300 1.740 25.620 ;
        RECT 0.980 24.720 1.300 25.040 ;
        RECT 2.550 24.220 2.850 27.200 ;
        RECT 5.510 27.130 5.650 28.880 ;
        RECT 9.500 28.430 9.830 28.710 ;
        RECT 10.260 28.470 10.430 29.200 ;
        RECT 11.170 29.190 11.460 29.200 ;
        RECT 13.000 29.020 13.230 29.890 ;
        RECT 13.000 28.880 13.360 29.020 ;
        RECT 17.040 28.890 17.270 29.890 ;
        RECT 17.980 29.500 18.280 30.660 ;
        RECT 18.420 31.690 18.820 32.280 ;
        RECT 19.020 32.020 19.350 32.340 ;
        RECT 19.070 31.690 19.300 32.020 ;
        RECT 19.550 31.690 20.060 32.340 ;
        RECT 18.420 30.690 18.650 31.690 ;
        RECT 18.800 31.240 19.090 31.550 ;
        RECT 19.810 31.290 20.060 31.690 ;
        RECT 19.360 30.850 19.650 31.180 ;
        RECT 19.810 30.960 20.160 31.290 ;
        RECT 25.080 31.050 25.460 31.370 ;
        RECT 19.810 30.690 20.060 30.960 ;
        RECT 25.690 30.830 25.990 32.480 ;
        RECT 26.300 32.280 26.530 32.340 ;
        RECT 18.420 29.690 18.900 30.690 ;
        RECT 19.150 29.990 19.380 30.690 ;
        RECT 19.100 29.650 19.430 29.990 ;
        RECT 19.630 29.710 20.060 30.690 ;
        RECT 23.350 30.660 25.990 30.830 ;
        RECT 23.350 30.490 23.640 30.660 ;
        RECT 20.440 30.070 20.770 30.360 ;
        RECT 24.920 30.060 25.250 30.340 ;
        RECT 19.630 29.690 19.860 29.710 ;
        RECT 17.980 29.340 19.170 29.500 ;
        RECT 17.970 29.200 19.170 29.340 ;
        RECT 12.730 28.470 13.060 28.700 ;
        RECT 4.380 27.060 5.650 27.130 ;
        RECT 3.160 27.000 3.390 27.060 ;
        RECT 2.990 26.410 3.390 27.000 ;
        RECT 3.590 26.740 3.920 27.060 ;
        RECT 4.120 26.990 5.650 27.060 ;
        RECT 10.260 28.330 13.060 28.470 ;
        RECT 10.260 27.510 10.430 28.330 ;
        RECT 10.260 27.200 11.860 27.510 ;
        RECT 3.640 26.410 3.870 26.740 ;
        RECT 4.120 26.410 4.630 26.990 ;
        RECT 5.230 26.660 6.400 26.800 ;
        RECT 5.230 26.460 5.550 26.660 ;
        RECT 6.110 26.460 6.430 26.660 ;
        RECT 2.990 25.410 3.220 26.410 ;
        RECT 3.370 25.960 3.660 26.270 ;
        RECT 3.930 25.570 4.220 25.900 ;
        RECT 4.380 25.410 4.630 26.410 ;
        RECT 2.990 24.410 3.470 25.410 ;
        RECT 3.720 24.710 3.950 25.410 ;
        RECT 3.670 24.370 4.000 24.710 ;
        RECT 4.200 24.550 4.630 25.410 ;
        RECT 5.490 25.290 5.830 25.630 ;
        RECT 9.130 25.300 9.450 25.620 ;
        RECT 5.040 24.730 5.380 25.050 ;
        RECT 5.910 24.740 6.240 25.010 ;
        RECT 6.100 24.550 6.240 24.740 ;
        RECT 8.690 24.720 9.010 25.040 ;
        RECT 4.200 24.410 6.240 24.550 ;
        RECT 4.410 24.390 6.240 24.410 ;
        RECT 10.260 24.220 10.560 27.200 ;
        RECT 13.220 27.130 13.360 28.880 ;
        RECT 17.210 28.430 17.540 28.710 ;
        RECT 17.970 28.470 18.140 29.200 ;
        RECT 18.880 29.190 19.170 29.200 ;
        RECT 20.710 29.020 20.940 29.890 ;
        RECT 20.710 28.880 21.070 29.020 ;
        RECT 24.750 28.890 24.980 29.890 ;
        RECT 25.690 29.500 25.990 30.660 ;
        RECT 26.130 31.690 26.530 32.280 ;
        RECT 26.730 32.020 27.060 32.340 ;
        RECT 26.780 31.690 27.010 32.020 ;
        RECT 27.260 31.690 27.770 32.340 ;
        RECT 26.130 30.690 26.360 31.690 ;
        RECT 26.510 31.240 26.800 31.550 ;
        RECT 27.520 31.290 27.770 31.690 ;
        RECT 27.070 30.850 27.360 31.180 ;
        RECT 27.520 30.960 27.870 31.290 ;
        RECT 32.790 31.050 33.170 31.370 ;
        RECT 27.520 30.690 27.770 30.960 ;
        RECT 33.400 30.830 33.700 32.480 ;
        RECT 34.010 32.280 34.240 32.340 ;
        RECT 26.130 29.690 26.610 30.690 ;
        RECT 26.860 29.990 27.090 30.690 ;
        RECT 26.810 29.650 27.140 29.990 ;
        RECT 27.340 29.710 27.770 30.690 ;
        RECT 31.060 30.660 33.700 30.830 ;
        RECT 31.060 30.490 31.350 30.660 ;
        RECT 28.150 30.070 28.480 30.360 ;
        RECT 32.630 30.060 32.960 30.340 ;
        RECT 27.340 29.690 27.570 29.710 ;
        RECT 25.690 29.340 26.880 29.500 ;
        RECT 25.680 29.200 26.880 29.340 ;
        RECT 20.440 28.470 20.770 28.700 ;
        RECT 12.090 27.060 13.360 27.130 ;
        RECT 10.870 27.000 11.100 27.060 ;
        RECT 10.700 26.410 11.100 27.000 ;
        RECT 11.300 26.740 11.630 27.060 ;
        RECT 11.830 26.990 13.360 27.060 ;
        RECT 17.970 28.330 20.770 28.470 ;
        RECT 17.970 27.510 18.140 28.330 ;
        RECT 17.970 27.200 19.570 27.510 ;
        RECT 11.350 26.410 11.580 26.740 ;
        RECT 11.830 26.410 12.340 26.990 ;
        RECT 12.940 26.660 14.110 26.800 ;
        RECT 12.940 26.460 13.260 26.660 ;
        RECT 13.820 26.460 14.140 26.660 ;
        RECT 10.700 25.410 10.930 26.410 ;
        RECT 11.080 25.960 11.370 26.270 ;
        RECT 11.640 25.570 11.930 25.900 ;
        RECT 12.090 25.410 12.340 26.410 ;
        RECT 10.700 24.410 11.180 25.410 ;
        RECT 11.430 24.710 11.660 25.410 ;
        RECT 11.380 24.370 11.710 24.710 ;
        RECT 11.910 24.550 12.340 25.410 ;
        RECT 13.200 25.290 13.540 25.630 ;
        RECT 16.840 25.300 17.160 25.620 ;
        RECT 12.750 24.730 13.090 25.050 ;
        RECT 13.620 24.740 13.950 25.010 ;
        RECT 13.810 24.550 13.950 24.740 ;
        RECT 16.400 24.720 16.720 25.040 ;
        RECT 11.910 24.410 13.950 24.550 ;
        RECT 12.120 24.390 13.950 24.410 ;
        RECT 17.970 24.220 18.270 27.200 ;
        RECT 20.930 27.130 21.070 28.880 ;
        RECT 24.920 28.430 25.250 28.710 ;
        RECT 25.680 28.470 25.850 29.200 ;
        RECT 26.590 29.190 26.880 29.200 ;
        RECT 28.420 29.020 28.650 29.890 ;
        RECT 28.420 28.880 28.780 29.020 ;
        RECT 32.460 28.890 32.690 29.890 ;
        RECT 33.400 29.500 33.700 30.660 ;
        RECT 33.840 31.690 34.240 32.280 ;
        RECT 34.440 32.020 34.770 32.340 ;
        RECT 34.490 31.690 34.720 32.020 ;
        RECT 34.970 31.690 35.480 32.340 ;
        RECT 33.840 30.690 34.070 31.690 ;
        RECT 34.220 31.240 34.510 31.550 ;
        RECT 35.230 31.290 35.480 31.690 ;
        RECT 34.780 30.850 35.070 31.180 ;
        RECT 35.230 30.960 35.580 31.290 ;
        RECT 40.500 31.050 40.880 31.370 ;
        RECT 35.230 30.690 35.480 30.960 ;
        RECT 41.110 30.830 41.410 32.480 ;
        RECT 41.720 32.280 41.950 32.340 ;
        RECT 33.840 29.690 34.320 30.690 ;
        RECT 34.570 29.990 34.800 30.690 ;
        RECT 34.520 29.650 34.850 29.990 ;
        RECT 35.050 29.710 35.480 30.690 ;
        RECT 38.770 30.660 41.410 30.830 ;
        RECT 38.770 30.490 39.060 30.660 ;
        RECT 35.860 30.070 36.190 30.360 ;
        RECT 40.340 30.060 40.670 30.340 ;
        RECT 35.050 29.690 35.280 29.710 ;
        RECT 33.400 29.340 34.590 29.500 ;
        RECT 33.390 29.200 34.590 29.340 ;
        RECT 28.150 28.470 28.480 28.700 ;
        RECT 19.800 27.060 21.070 27.130 ;
        RECT 18.580 27.000 18.810 27.060 ;
        RECT 18.410 26.410 18.810 27.000 ;
        RECT 19.010 26.740 19.340 27.060 ;
        RECT 19.540 26.990 21.070 27.060 ;
        RECT 25.680 28.330 28.480 28.470 ;
        RECT 25.680 27.510 25.850 28.330 ;
        RECT 25.680 27.200 27.280 27.510 ;
        RECT 19.060 26.410 19.290 26.740 ;
        RECT 19.540 26.410 20.050 26.990 ;
        RECT 20.650 26.660 21.820 26.800 ;
        RECT 20.650 26.460 20.970 26.660 ;
        RECT 21.530 26.460 21.850 26.660 ;
        RECT 18.410 25.410 18.640 26.410 ;
        RECT 18.790 25.960 19.080 26.270 ;
        RECT 19.350 25.570 19.640 25.900 ;
        RECT 19.800 25.410 20.050 26.410 ;
        RECT 18.410 24.410 18.890 25.410 ;
        RECT 19.140 24.710 19.370 25.410 ;
        RECT 19.090 24.370 19.420 24.710 ;
        RECT 19.620 24.550 20.050 25.410 ;
        RECT 20.910 25.290 21.250 25.630 ;
        RECT 24.550 25.300 24.870 25.620 ;
        RECT 20.460 24.730 20.800 25.050 ;
        RECT 21.330 24.740 21.660 25.010 ;
        RECT 21.520 24.550 21.660 24.740 ;
        RECT 24.110 24.720 24.430 25.040 ;
        RECT 19.620 24.410 21.660 24.550 ;
        RECT 19.830 24.390 21.660 24.410 ;
        RECT 25.680 24.220 25.980 27.200 ;
        RECT 28.640 27.130 28.780 28.880 ;
        RECT 32.630 28.430 32.960 28.710 ;
        RECT 33.390 28.470 33.560 29.200 ;
        RECT 34.300 29.190 34.590 29.200 ;
        RECT 36.130 29.020 36.360 29.890 ;
        RECT 36.130 28.880 36.490 29.020 ;
        RECT 40.170 28.890 40.400 29.890 ;
        RECT 41.110 29.500 41.410 30.660 ;
        RECT 41.550 31.690 41.950 32.280 ;
        RECT 42.150 32.020 42.480 32.340 ;
        RECT 42.200 31.690 42.430 32.020 ;
        RECT 42.680 31.690 43.190 32.340 ;
        RECT 41.550 30.690 41.780 31.690 ;
        RECT 41.930 31.240 42.220 31.550 ;
        RECT 42.940 31.290 43.190 31.690 ;
        RECT 42.490 30.850 42.780 31.180 ;
        RECT 42.940 30.960 43.290 31.290 ;
        RECT 48.210 31.050 48.590 31.370 ;
        RECT 42.940 30.690 43.190 30.960 ;
        RECT 48.820 30.830 49.120 32.480 ;
        RECT 49.430 32.280 49.660 32.340 ;
        RECT 41.550 29.690 42.030 30.690 ;
        RECT 42.280 29.990 42.510 30.690 ;
        RECT 42.230 29.650 42.560 29.990 ;
        RECT 42.760 29.710 43.190 30.690 ;
        RECT 46.480 30.660 49.120 30.830 ;
        RECT 46.480 30.490 46.770 30.660 ;
        RECT 43.570 30.070 43.900 30.360 ;
        RECT 48.050 30.060 48.380 30.340 ;
        RECT 42.760 29.690 42.990 29.710 ;
        RECT 41.110 29.340 42.300 29.500 ;
        RECT 41.100 29.200 42.300 29.340 ;
        RECT 35.860 28.470 36.190 28.700 ;
        RECT 27.510 27.060 28.780 27.130 ;
        RECT 26.290 27.000 26.520 27.060 ;
        RECT 26.120 26.410 26.520 27.000 ;
        RECT 26.720 26.740 27.050 27.060 ;
        RECT 27.250 26.990 28.780 27.060 ;
        RECT 33.390 28.330 36.190 28.470 ;
        RECT 33.390 27.510 33.560 28.330 ;
        RECT 33.390 27.200 34.990 27.510 ;
        RECT 26.770 26.410 27.000 26.740 ;
        RECT 27.250 26.410 27.760 26.990 ;
        RECT 28.360 26.660 29.530 26.800 ;
        RECT 28.360 26.460 28.680 26.660 ;
        RECT 29.240 26.460 29.560 26.660 ;
        RECT 26.120 25.410 26.350 26.410 ;
        RECT 26.500 25.960 26.790 26.270 ;
        RECT 27.060 25.570 27.350 25.900 ;
        RECT 27.510 25.410 27.760 26.410 ;
        RECT 26.120 24.410 26.600 25.410 ;
        RECT 26.850 24.710 27.080 25.410 ;
        RECT 26.800 24.370 27.130 24.710 ;
        RECT 27.330 24.550 27.760 25.410 ;
        RECT 28.620 25.290 28.960 25.630 ;
        RECT 32.260 25.300 32.580 25.620 ;
        RECT 28.170 24.730 28.510 25.050 ;
        RECT 29.040 24.740 29.370 25.010 ;
        RECT 29.230 24.550 29.370 24.740 ;
        RECT 31.820 24.720 32.140 25.040 ;
        RECT 27.330 24.410 29.370 24.550 ;
        RECT 27.540 24.390 29.370 24.410 ;
        RECT 33.390 24.220 33.690 27.200 ;
        RECT 36.350 27.130 36.490 28.880 ;
        RECT 40.340 28.430 40.670 28.710 ;
        RECT 41.100 28.470 41.270 29.200 ;
        RECT 42.010 29.190 42.300 29.200 ;
        RECT 43.840 29.020 44.070 29.890 ;
        RECT 43.840 28.880 44.200 29.020 ;
        RECT 47.880 28.890 48.110 29.890 ;
        RECT 48.820 29.500 49.120 30.660 ;
        RECT 49.260 31.690 49.660 32.280 ;
        RECT 49.860 32.020 50.190 32.340 ;
        RECT 49.910 31.690 50.140 32.020 ;
        RECT 50.390 31.690 50.900 32.340 ;
        RECT 49.260 30.690 49.490 31.690 ;
        RECT 49.640 31.240 49.930 31.550 ;
        RECT 50.650 31.290 50.900 31.690 ;
        RECT 50.200 30.850 50.490 31.180 ;
        RECT 50.650 30.960 51.000 31.290 ;
        RECT 55.920 31.050 56.300 31.370 ;
        RECT 50.650 30.690 50.900 30.960 ;
        RECT 56.530 30.830 56.830 32.480 ;
        RECT 57.140 32.280 57.370 32.340 ;
        RECT 49.260 29.690 49.740 30.690 ;
        RECT 49.990 29.990 50.220 30.690 ;
        RECT 49.940 29.650 50.270 29.990 ;
        RECT 50.470 29.710 50.900 30.690 ;
        RECT 54.190 30.660 56.830 30.830 ;
        RECT 54.190 30.490 54.480 30.660 ;
        RECT 51.280 30.070 51.610 30.360 ;
        RECT 55.760 30.060 56.090 30.340 ;
        RECT 50.470 29.690 50.700 29.710 ;
        RECT 48.820 29.340 50.010 29.500 ;
        RECT 48.810 29.200 50.010 29.340 ;
        RECT 43.570 28.470 43.900 28.700 ;
        RECT 35.220 27.060 36.490 27.130 ;
        RECT 34.000 27.000 34.230 27.060 ;
        RECT 33.830 26.410 34.230 27.000 ;
        RECT 34.430 26.740 34.760 27.060 ;
        RECT 34.960 26.990 36.490 27.060 ;
        RECT 41.100 28.330 43.900 28.470 ;
        RECT 41.100 27.510 41.270 28.330 ;
        RECT 41.100 27.200 42.700 27.510 ;
        RECT 34.480 26.410 34.710 26.740 ;
        RECT 34.960 26.410 35.470 26.990 ;
        RECT 36.070 26.660 37.240 26.800 ;
        RECT 36.070 26.460 36.390 26.660 ;
        RECT 36.950 26.460 37.270 26.660 ;
        RECT 33.830 25.410 34.060 26.410 ;
        RECT 34.210 25.960 34.500 26.270 ;
        RECT 34.770 25.570 35.060 25.900 ;
        RECT 35.220 25.410 35.470 26.410 ;
        RECT 33.830 24.410 34.310 25.410 ;
        RECT 34.560 24.710 34.790 25.410 ;
        RECT 34.510 24.370 34.840 24.710 ;
        RECT 35.040 24.550 35.470 25.410 ;
        RECT 36.330 25.290 36.670 25.630 ;
        RECT 39.970 25.300 40.290 25.620 ;
        RECT 35.880 24.730 36.220 25.050 ;
        RECT 36.750 24.740 37.080 25.010 ;
        RECT 36.940 24.550 37.080 24.740 ;
        RECT 39.530 24.720 39.850 25.040 ;
        RECT 35.040 24.410 37.080 24.550 ;
        RECT 35.250 24.390 37.080 24.410 ;
        RECT 41.100 24.220 41.400 27.200 ;
        RECT 44.060 27.130 44.200 28.880 ;
        RECT 48.050 28.430 48.380 28.710 ;
        RECT 48.810 28.470 48.980 29.200 ;
        RECT 49.720 29.190 50.010 29.200 ;
        RECT 51.550 29.020 51.780 29.890 ;
        RECT 51.550 28.880 51.910 29.020 ;
        RECT 55.590 28.890 55.820 29.890 ;
        RECT 56.530 29.500 56.830 30.660 ;
        RECT 56.970 31.690 57.370 32.280 ;
        RECT 57.570 32.020 57.900 32.340 ;
        RECT 57.620 31.690 57.850 32.020 ;
        RECT 58.100 31.690 58.610 32.340 ;
        RECT 56.970 30.690 57.200 31.690 ;
        RECT 57.350 31.240 57.640 31.550 ;
        RECT 58.360 31.290 58.610 31.690 ;
        RECT 57.910 30.850 58.200 31.180 ;
        RECT 58.360 30.960 58.710 31.290 ;
        RECT 63.630 31.050 64.010 31.370 ;
        RECT 58.360 30.690 58.610 30.960 ;
        RECT 64.240 30.830 64.540 32.480 ;
        RECT 64.850 32.280 65.080 32.340 ;
        RECT 56.970 29.690 57.450 30.690 ;
        RECT 57.700 29.990 57.930 30.690 ;
        RECT 57.650 29.650 57.980 29.990 ;
        RECT 58.180 29.710 58.610 30.690 ;
        RECT 61.900 30.660 64.540 30.830 ;
        RECT 61.900 30.490 62.190 30.660 ;
        RECT 58.990 30.070 59.320 30.360 ;
        RECT 63.470 30.060 63.800 30.340 ;
        RECT 58.180 29.690 58.410 29.710 ;
        RECT 56.530 29.340 57.720 29.500 ;
        RECT 56.520 29.200 57.720 29.340 ;
        RECT 51.280 28.470 51.610 28.700 ;
        RECT 42.930 27.060 44.200 27.130 ;
        RECT 41.710 27.000 41.940 27.060 ;
        RECT 41.540 26.410 41.940 27.000 ;
        RECT 42.140 26.740 42.470 27.060 ;
        RECT 42.670 26.990 44.200 27.060 ;
        RECT 48.810 28.330 51.610 28.470 ;
        RECT 48.810 27.510 48.980 28.330 ;
        RECT 48.810 27.200 50.410 27.510 ;
        RECT 42.190 26.410 42.420 26.740 ;
        RECT 42.670 26.410 43.180 26.990 ;
        RECT 43.780 26.660 44.950 26.800 ;
        RECT 43.780 26.460 44.100 26.660 ;
        RECT 44.660 26.460 44.980 26.660 ;
        RECT 41.540 25.410 41.770 26.410 ;
        RECT 41.920 25.960 42.210 26.270 ;
        RECT 42.480 25.570 42.770 25.900 ;
        RECT 42.930 25.410 43.180 26.410 ;
        RECT 41.540 24.410 42.020 25.410 ;
        RECT 42.270 24.710 42.500 25.410 ;
        RECT 42.220 24.370 42.550 24.710 ;
        RECT 42.750 24.550 43.180 25.410 ;
        RECT 44.040 25.290 44.380 25.630 ;
        RECT 47.680 25.300 48.000 25.620 ;
        RECT 43.590 24.730 43.930 25.050 ;
        RECT 44.460 24.740 44.790 25.010 ;
        RECT 44.650 24.550 44.790 24.740 ;
        RECT 47.240 24.720 47.560 25.040 ;
        RECT 42.750 24.410 44.790 24.550 ;
        RECT 42.960 24.390 44.790 24.410 ;
        RECT 48.810 24.220 49.110 27.200 ;
        RECT 51.770 27.130 51.910 28.880 ;
        RECT 55.760 28.430 56.090 28.710 ;
        RECT 56.520 28.470 56.690 29.200 ;
        RECT 57.430 29.190 57.720 29.200 ;
        RECT 59.260 29.020 59.490 29.890 ;
        RECT 59.260 28.880 59.620 29.020 ;
        RECT 63.300 28.890 63.530 29.890 ;
        RECT 64.240 29.500 64.540 30.660 ;
        RECT 64.680 31.690 65.080 32.280 ;
        RECT 65.280 32.020 65.610 32.340 ;
        RECT 65.330 31.690 65.560 32.020 ;
        RECT 65.810 31.690 66.320 32.340 ;
        RECT 64.680 30.690 64.910 31.690 ;
        RECT 65.060 31.240 65.350 31.550 ;
        RECT 66.070 31.290 66.320 31.690 ;
        RECT 65.620 30.850 65.910 31.180 ;
        RECT 66.070 30.960 66.420 31.290 ;
        RECT 71.340 31.050 71.720 31.370 ;
        RECT 66.070 30.690 66.320 30.960 ;
        RECT 71.950 30.830 72.250 32.480 ;
        RECT 72.560 32.280 72.790 32.340 ;
        RECT 64.680 29.690 65.160 30.690 ;
        RECT 65.410 29.990 65.640 30.690 ;
        RECT 65.360 29.650 65.690 29.990 ;
        RECT 65.890 29.710 66.320 30.690 ;
        RECT 69.610 30.660 72.250 30.830 ;
        RECT 69.610 30.490 69.900 30.660 ;
        RECT 66.700 30.070 67.030 30.360 ;
        RECT 71.180 30.060 71.510 30.340 ;
        RECT 65.890 29.690 66.120 29.710 ;
        RECT 64.240 29.340 65.430 29.500 ;
        RECT 64.230 29.200 65.430 29.340 ;
        RECT 58.990 28.470 59.320 28.700 ;
        RECT 50.640 27.060 51.910 27.130 ;
        RECT 49.420 27.000 49.650 27.060 ;
        RECT 49.250 26.410 49.650 27.000 ;
        RECT 49.850 26.740 50.180 27.060 ;
        RECT 50.380 26.990 51.910 27.060 ;
        RECT 56.520 28.330 59.320 28.470 ;
        RECT 56.520 27.510 56.690 28.330 ;
        RECT 56.520 27.200 58.120 27.510 ;
        RECT 49.900 26.410 50.130 26.740 ;
        RECT 50.380 26.410 50.890 26.990 ;
        RECT 51.490 26.660 52.660 26.800 ;
        RECT 51.490 26.460 51.810 26.660 ;
        RECT 52.370 26.460 52.690 26.660 ;
        RECT 49.250 25.410 49.480 26.410 ;
        RECT 49.630 25.960 49.920 26.270 ;
        RECT 50.190 25.570 50.480 25.900 ;
        RECT 50.640 25.410 50.890 26.410 ;
        RECT 49.250 24.410 49.730 25.410 ;
        RECT 49.980 24.710 50.210 25.410 ;
        RECT 49.930 24.370 50.260 24.710 ;
        RECT 50.460 24.550 50.890 25.410 ;
        RECT 51.750 25.290 52.090 25.630 ;
        RECT 55.390 25.300 55.710 25.620 ;
        RECT 51.300 24.730 51.640 25.050 ;
        RECT 52.170 24.740 52.500 25.010 ;
        RECT 52.360 24.550 52.500 24.740 ;
        RECT 54.950 24.720 55.270 25.040 ;
        RECT 50.460 24.410 52.500 24.550 ;
        RECT 50.670 24.390 52.500 24.410 ;
        RECT 56.520 24.220 56.820 27.200 ;
        RECT 59.480 27.130 59.620 28.880 ;
        RECT 63.470 28.430 63.800 28.710 ;
        RECT 64.230 28.470 64.400 29.200 ;
        RECT 65.140 29.190 65.430 29.200 ;
        RECT 66.970 29.020 67.200 29.890 ;
        RECT 66.970 28.880 67.330 29.020 ;
        RECT 71.010 28.890 71.240 29.890 ;
        RECT 71.950 29.500 72.250 30.660 ;
        RECT 72.390 31.690 72.790 32.280 ;
        RECT 72.990 32.020 73.320 32.340 ;
        RECT 73.040 31.690 73.270 32.020 ;
        RECT 73.520 31.690 74.030 32.340 ;
        RECT 72.390 30.690 72.620 31.690 ;
        RECT 72.770 31.240 73.060 31.550 ;
        RECT 73.780 31.290 74.030 31.690 ;
        RECT 73.330 30.850 73.620 31.180 ;
        RECT 73.780 30.960 74.130 31.290 ;
        RECT 79.050 31.050 79.430 31.370 ;
        RECT 73.780 30.690 74.030 30.960 ;
        RECT 79.660 30.830 79.960 32.480 ;
        RECT 80.270 32.280 80.500 32.340 ;
        RECT 72.390 29.690 72.870 30.690 ;
        RECT 73.120 29.990 73.350 30.690 ;
        RECT 73.070 29.650 73.400 29.990 ;
        RECT 73.600 29.710 74.030 30.690 ;
        RECT 77.320 30.660 79.960 30.830 ;
        RECT 77.320 30.490 77.610 30.660 ;
        RECT 74.410 30.070 74.740 30.360 ;
        RECT 78.890 30.060 79.220 30.340 ;
        RECT 73.600 29.690 73.830 29.710 ;
        RECT 71.950 29.340 73.140 29.500 ;
        RECT 71.940 29.200 73.140 29.340 ;
        RECT 66.700 28.470 67.030 28.700 ;
        RECT 58.350 27.060 59.620 27.130 ;
        RECT 57.130 27.000 57.360 27.060 ;
        RECT 56.960 26.410 57.360 27.000 ;
        RECT 57.560 26.740 57.890 27.060 ;
        RECT 58.090 26.990 59.620 27.060 ;
        RECT 64.230 28.330 67.030 28.470 ;
        RECT 64.230 27.510 64.400 28.330 ;
        RECT 64.230 27.200 65.830 27.510 ;
        RECT 57.610 26.410 57.840 26.740 ;
        RECT 58.090 26.410 58.600 26.990 ;
        RECT 59.200 26.660 60.370 26.800 ;
        RECT 59.200 26.460 59.520 26.660 ;
        RECT 60.080 26.460 60.400 26.660 ;
        RECT 56.960 25.410 57.190 26.410 ;
        RECT 57.340 25.960 57.630 26.270 ;
        RECT 57.900 25.570 58.190 25.900 ;
        RECT 58.350 25.410 58.600 26.410 ;
        RECT 56.960 24.410 57.440 25.410 ;
        RECT 57.690 24.710 57.920 25.410 ;
        RECT 57.640 24.370 57.970 24.710 ;
        RECT 58.170 24.550 58.600 25.410 ;
        RECT 59.460 25.290 59.800 25.630 ;
        RECT 63.100 25.300 63.420 25.620 ;
        RECT 59.010 24.730 59.350 25.050 ;
        RECT 59.880 24.740 60.210 25.010 ;
        RECT 60.070 24.550 60.210 24.740 ;
        RECT 62.660 24.720 62.980 25.040 ;
        RECT 58.170 24.410 60.210 24.550 ;
        RECT 58.380 24.390 60.210 24.410 ;
        RECT 64.230 24.220 64.530 27.200 ;
        RECT 67.190 27.130 67.330 28.880 ;
        RECT 71.180 28.430 71.510 28.710 ;
        RECT 71.940 28.470 72.110 29.200 ;
        RECT 72.850 29.190 73.140 29.200 ;
        RECT 74.680 29.020 74.910 29.890 ;
        RECT 74.680 28.880 75.040 29.020 ;
        RECT 78.720 28.890 78.950 29.890 ;
        RECT 79.660 29.500 79.960 30.660 ;
        RECT 80.100 31.690 80.500 32.280 ;
        RECT 80.700 32.020 81.030 32.340 ;
        RECT 80.750 31.690 80.980 32.020 ;
        RECT 81.230 31.690 81.740 32.340 ;
        RECT 80.100 30.690 80.330 31.690 ;
        RECT 80.480 31.240 80.770 31.550 ;
        RECT 81.490 31.290 81.740 31.690 ;
        RECT 81.040 30.850 81.330 31.180 ;
        RECT 81.490 30.960 81.840 31.290 ;
        RECT 86.760 31.050 87.140 31.370 ;
        RECT 81.490 30.690 81.740 30.960 ;
        RECT 87.370 30.830 87.670 32.480 ;
        RECT 87.980 32.280 88.210 32.340 ;
        RECT 80.100 29.690 80.580 30.690 ;
        RECT 80.830 29.990 81.060 30.690 ;
        RECT 80.780 29.650 81.110 29.990 ;
        RECT 81.310 29.710 81.740 30.690 ;
        RECT 85.030 30.660 87.670 30.830 ;
        RECT 85.030 30.490 85.320 30.660 ;
        RECT 82.120 30.070 82.450 30.360 ;
        RECT 86.600 30.060 86.930 30.340 ;
        RECT 81.310 29.690 81.540 29.710 ;
        RECT 79.660 29.340 80.850 29.500 ;
        RECT 79.650 29.200 80.850 29.340 ;
        RECT 74.410 28.470 74.740 28.700 ;
        RECT 66.060 27.060 67.330 27.130 ;
        RECT 64.840 27.000 65.070 27.060 ;
        RECT 64.670 26.410 65.070 27.000 ;
        RECT 65.270 26.740 65.600 27.060 ;
        RECT 65.800 26.990 67.330 27.060 ;
        RECT 71.940 28.330 74.740 28.470 ;
        RECT 71.940 27.510 72.110 28.330 ;
        RECT 71.940 27.200 73.540 27.510 ;
        RECT 65.320 26.410 65.550 26.740 ;
        RECT 65.800 26.410 66.310 26.990 ;
        RECT 66.910 26.660 68.080 26.800 ;
        RECT 66.910 26.460 67.230 26.660 ;
        RECT 67.790 26.460 68.110 26.660 ;
        RECT 64.670 25.410 64.900 26.410 ;
        RECT 65.050 25.960 65.340 26.270 ;
        RECT 65.610 25.570 65.900 25.900 ;
        RECT 66.060 25.410 66.310 26.410 ;
        RECT 64.670 24.410 65.150 25.410 ;
        RECT 65.400 24.710 65.630 25.410 ;
        RECT 65.350 24.370 65.680 24.710 ;
        RECT 65.880 24.550 66.310 25.410 ;
        RECT 67.170 25.290 67.510 25.630 ;
        RECT 70.810 25.300 71.130 25.620 ;
        RECT 66.720 24.730 67.060 25.050 ;
        RECT 67.590 24.740 67.920 25.010 ;
        RECT 67.780 24.550 67.920 24.740 ;
        RECT 70.370 24.720 70.690 25.040 ;
        RECT 65.880 24.410 67.920 24.550 ;
        RECT 66.090 24.390 67.920 24.410 ;
        RECT 71.940 24.220 72.240 27.200 ;
        RECT 74.900 27.130 75.040 28.880 ;
        RECT 78.890 28.430 79.220 28.710 ;
        RECT 79.650 28.470 79.820 29.200 ;
        RECT 80.560 29.190 80.850 29.200 ;
        RECT 82.390 29.020 82.620 29.890 ;
        RECT 82.390 28.880 82.750 29.020 ;
        RECT 86.430 28.890 86.660 29.890 ;
        RECT 87.370 29.500 87.670 30.660 ;
        RECT 87.810 31.690 88.210 32.280 ;
        RECT 88.410 32.020 88.740 32.340 ;
        RECT 88.460 31.690 88.690 32.020 ;
        RECT 88.940 31.690 89.450 32.340 ;
        RECT 87.810 30.690 88.040 31.690 ;
        RECT 88.190 31.240 88.480 31.550 ;
        RECT 89.200 31.290 89.450 31.690 ;
        RECT 88.750 30.850 89.040 31.180 ;
        RECT 89.200 30.960 89.550 31.290 ;
        RECT 94.470 31.050 94.850 31.370 ;
        RECT 89.200 30.690 89.450 30.960 ;
        RECT 95.080 30.830 95.380 32.480 ;
        RECT 95.690 32.280 95.920 32.340 ;
        RECT 87.810 29.690 88.290 30.690 ;
        RECT 88.540 29.990 88.770 30.690 ;
        RECT 88.490 29.650 88.820 29.990 ;
        RECT 89.020 29.710 89.450 30.690 ;
        RECT 92.740 30.660 95.380 30.830 ;
        RECT 92.740 30.490 93.030 30.660 ;
        RECT 89.830 30.070 90.160 30.360 ;
        RECT 94.310 30.060 94.640 30.340 ;
        RECT 89.020 29.690 89.250 29.710 ;
        RECT 87.370 29.340 88.560 29.500 ;
        RECT 87.360 29.200 88.560 29.340 ;
        RECT 82.120 28.470 82.450 28.700 ;
        RECT 73.770 27.060 75.040 27.130 ;
        RECT 72.550 27.000 72.780 27.060 ;
        RECT 72.380 26.410 72.780 27.000 ;
        RECT 72.980 26.740 73.310 27.060 ;
        RECT 73.510 26.990 75.040 27.060 ;
        RECT 79.650 28.330 82.450 28.470 ;
        RECT 79.650 27.510 79.820 28.330 ;
        RECT 79.650 27.200 81.250 27.510 ;
        RECT 73.030 26.410 73.260 26.740 ;
        RECT 73.510 26.410 74.020 26.990 ;
        RECT 74.620 26.660 75.790 26.800 ;
        RECT 74.620 26.460 74.940 26.660 ;
        RECT 75.500 26.460 75.820 26.660 ;
        RECT 72.380 25.410 72.610 26.410 ;
        RECT 72.760 25.960 73.050 26.270 ;
        RECT 73.320 25.570 73.610 25.900 ;
        RECT 73.770 25.410 74.020 26.410 ;
        RECT 72.380 24.410 72.860 25.410 ;
        RECT 73.110 24.710 73.340 25.410 ;
        RECT 73.060 24.370 73.390 24.710 ;
        RECT 73.590 24.550 74.020 25.410 ;
        RECT 74.880 25.290 75.220 25.630 ;
        RECT 78.520 25.300 78.840 25.620 ;
        RECT 74.430 24.730 74.770 25.050 ;
        RECT 75.300 24.740 75.630 25.010 ;
        RECT 75.490 24.550 75.630 24.740 ;
        RECT 78.080 24.720 78.400 25.040 ;
        RECT 73.590 24.410 75.630 24.550 ;
        RECT 73.800 24.390 75.630 24.410 ;
        RECT 79.650 24.220 79.950 27.200 ;
        RECT 82.610 27.130 82.750 28.880 ;
        RECT 86.600 28.430 86.930 28.710 ;
        RECT 87.360 28.470 87.530 29.200 ;
        RECT 88.270 29.190 88.560 29.200 ;
        RECT 90.100 29.020 90.330 29.890 ;
        RECT 90.100 28.880 90.460 29.020 ;
        RECT 94.140 28.890 94.370 29.890 ;
        RECT 95.080 29.500 95.380 30.660 ;
        RECT 95.520 31.690 95.920 32.280 ;
        RECT 96.120 32.020 96.450 32.340 ;
        RECT 96.170 31.690 96.400 32.020 ;
        RECT 96.650 31.690 97.160 32.340 ;
        RECT 95.520 30.690 95.750 31.690 ;
        RECT 95.900 31.240 96.190 31.550 ;
        RECT 96.910 31.290 97.160 31.690 ;
        RECT 96.460 30.850 96.750 31.180 ;
        RECT 96.910 30.960 97.260 31.290 ;
        RECT 102.180 31.050 102.560 31.370 ;
        RECT 96.910 30.690 97.160 30.960 ;
        RECT 102.790 30.830 103.090 32.480 ;
        RECT 103.400 32.280 103.630 32.340 ;
        RECT 95.520 29.690 96.000 30.690 ;
        RECT 96.250 29.990 96.480 30.690 ;
        RECT 96.200 29.650 96.530 29.990 ;
        RECT 96.730 29.710 97.160 30.690 ;
        RECT 100.450 30.660 103.090 30.830 ;
        RECT 100.450 30.490 100.740 30.660 ;
        RECT 97.540 30.070 97.870 30.360 ;
        RECT 102.020 30.060 102.350 30.340 ;
        RECT 96.730 29.690 96.960 29.710 ;
        RECT 95.080 29.340 96.270 29.500 ;
        RECT 95.070 29.200 96.270 29.340 ;
        RECT 89.830 28.470 90.160 28.700 ;
        RECT 81.480 27.060 82.750 27.130 ;
        RECT 80.260 27.000 80.490 27.060 ;
        RECT 80.090 26.410 80.490 27.000 ;
        RECT 80.690 26.740 81.020 27.060 ;
        RECT 81.220 26.990 82.750 27.060 ;
        RECT 87.360 28.330 90.160 28.470 ;
        RECT 87.360 27.510 87.530 28.330 ;
        RECT 87.360 27.200 88.960 27.510 ;
        RECT 80.740 26.410 80.970 26.740 ;
        RECT 81.220 26.410 81.730 26.990 ;
        RECT 82.330 26.660 83.500 26.800 ;
        RECT 82.330 26.460 82.650 26.660 ;
        RECT 83.210 26.460 83.530 26.660 ;
        RECT 80.090 25.410 80.320 26.410 ;
        RECT 80.470 25.960 80.760 26.270 ;
        RECT 81.030 25.570 81.320 25.900 ;
        RECT 81.480 25.410 81.730 26.410 ;
        RECT 80.090 24.410 80.570 25.410 ;
        RECT 80.820 24.710 81.050 25.410 ;
        RECT 80.770 24.370 81.100 24.710 ;
        RECT 81.300 24.550 81.730 25.410 ;
        RECT 82.590 25.290 82.930 25.630 ;
        RECT 86.230 25.300 86.550 25.620 ;
        RECT 82.140 24.730 82.480 25.050 ;
        RECT 83.010 24.740 83.340 25.010 ;
        RECT 83.200 24.550 83.340 24.740 ;
        RECT 85.790 24.720 86.110 25.040 ;
        RECT 81.300 24.410 83.340 24.550 ;
        RECT 81.510 24.390 83.340 24.410 ;
        RECT 87.360 24.220 87.660 27.200 ;
        RECT 90.320 27.130 90.460 28.880 ;
        RECT 94.310 28.430 94.640 28.710 ;
        RECT 95.070 28.470 95.240 29.200 ;
        RECT 95.980 29.190 96.270 29.200 ;
        RECT 97.810 29.020 98.040 29.890 ;
        RECT 97.810 28.880 98.170 29.020 ;
        RECT 101.850 28.890 102.080 29.890 ;
        RECT 102.790 29.500 103.090 30.660 ;
        RECT 103.230 31.690 103.630 32.280 ;
        RECT 103.830 32.020 104.160 32.340 ;
        RECT 103.880 31.690 104.110 32.020 ;
        RECT 104.360 31.690 104.870 32.340 ;
        RECT 103.230 30.690 103.460 31.690 ;
        RECT 103.610 31.240 103.900 31.550 ;
        RECT 104.620 31.290 104.870 31.690 ;
        RECT 104.170 30.850 104.460 31.180 ;
        RECT 104.620 30.960 104.970 31.290 ;
        RECT 109.890 31.050 110.270 31.370 ;
        RECT 104.620 30.690 104.870 30.960 ;
        RECT 110.500 30.830 110.800 32.480 ;
        RECT 111.110 32.280 111.340 32.340 ;
        RECT 103.230 29.690 103.710 30.690 ;
        RECT 103.960 29.990 104.190 30.690 ;
        RECT 103.910 29.650 104.240 29.990 ;
        RECT 104.440 29.710 104.870 30.690 ;
        RECT 108.160 30.660 110.800 30.830 ;
        RECT 108.160 30.490 108.450 30.660 ;
        RECT 105.250 30.070 105.580 30.360 ;
        RECT 109.730 30.060 110.060 30.340 ;
        RECT 104.440 29.690 104.670 29.710 ;
        RECT 102.790 29.340 103.980 29.500 ;
        RECT 102.780 29.200 103.980 29.340 ;
        RECT 97.540 28.470 97.870 28.700 ;
        RECT 89.190 27.060 90.460 27.130 ;
        RECT 87.970 27.000 88.200 27.060 ;
        RECT 87.800 26.410 88.200 27.000 ;
        RECT 88.400 26.740 88.730 27.060 ;
        RECT 88.930 26.990 90.460 27.060 ;
        RECT 95.070 28.330 97.870 28.470 ;
        RECT 95.070 27.510 95.240 28.330 ;
        RECT 95.070 27.200 96.670 27.510 ;
        RECT 88.450 26.410 88.680 26.740 ;
        RECT 88.930 26.410 89.440 26.990 ;
        RECT 90.040 26.660 91.210 26.800 ;
        RECT 90.040 26.460 90.360 26.660 ;
        RECT 90.920 26.460 91.240 26.660 ;
        RECT 87.800 25.410 88.030 26.410 ;
        RECT 88.180 25.960 88.470 26.270 ;
        RECT 88.740 25.570 89.030 25.900 ;
        RECT 89.190 25.410 89.440 26.410 ;
        RECT 87.800 24.410 88.280 25.410 ;
        RECT 88.530 24.710 88.760 25.410 ;
        RECT 88.480 24.370 88.810 24.710 ;
        RECT 89.010 24.550 89.440 25.410 ;
        RECT 90.300 25.290 90.640 25.630 ;
        RECT 93.940 25.300 94.260 25.620 ;
        RECT 89.850 24.730 90.190 25.050 ;
        RECT 90.720 24.740 91.050 25.010 ;
        RECT 90.910 24.550 91.050 24.740 ;
        RECT 93.500 24.720 93.820 25.040 ;
        RECT 89.010 24.410 91.050 24.550 ;
        RECT 89.220 24.390 91.050 24.410 ;
        RECT 95.070 24.220 95.370 27.200 ;
        RECT 98.030 27.130 98.170 28.880 ;
        RECT 102.020 28.430 102.350 28.710 ;
        RECT 102.780 28.470 102.950 29.200 ;
        RECT 103.690 29.190 103.980 29.200 ;
        RECT 105.520 29.020 105.750 29.890 ;
        RECT 105.520 28.880 105.880 29.020 ;
        RECT 109.560 28.890 109.790 29.890 ;
        RECT 110.500 29.500 110.800 30.660 ;
        RECT 110.940 31.690 111.340 32.280 ;
        RECT 111.540 32.020 111.870 32.340 ;
        RECT 111.590 31.690 111.820 32.020 ;
        RECT 112.070 31.690 112.580 32.340 ;
        RECT 110.940 30.690 111.170 31.690 ;
        RECT 111.320 31.240 111.610 31.550 ;
        RECT 112.330 31.290 112.580 31.690 ;
        RECT 111.880 30.850 112.170 31.180 ;
        RECT 112.330 30.960 112.680 31.290 ;
        RECT 117.600 31.050 117.980 31.370 ;
        RECT 112.330 30.690 112.580 30.960 ;
        RECT 118.210 30.830 118.510 32.480 ;
        RECT 118.820 32.280 119.050 32.340 ;
        RECT 110.940 29.690 111.420 30.690 ;
        RECT 111.670 29.990 111.900 30.690 ;
        RECT 111.620 29.650 111.950 29.990 ;
        RECT 112.150 29.710 112.580 30.690 ;
        RECT 115.870 30.660 118.510 30.830 ;
        RECT 115.870 30.490 116.160 30.660 ;
        RECT 112.960 30.070 113.290 30.360 ;
        RECT 117.440 30.060 117.770 30.340 ;
        RECT 112.150 29.690 112.380 29.710 ;
        RECT 110.500 29.340 111.690 29.500 ;
        RECT 110.490 29.200 111.690 29.340 ;
        RECT 105.250 28.470 105.580 28.700 ;
        RECT 96.900 27.060 98.170 27.130 ;
        RECT 95.680 27.000 95.910 27.060 ;
        RECT 95.510 26.410 95.910 27.000 ;
        RECT 96.110 26.740 96.440 27.060 ;
        RECT 96.640 26.990 98.170 27.060 ;
        RECT 102.780 28.330 105.580 28.470 ;
        RECT 102.780 27.510 102.950 28.330 ;
        RECT 102.780 27.200 104.380 27.510 ;
        RECT 96.160 26.410 96.390 26.740 ;
        RECT 96.640 26.410 97.150 26.990 ;
        RECT 97.750 26.660 98.920 26.800 ;
        RECT 97.750 26.460 98.070 26.660 ;
        RECT 98.630 26.460 98.950 26.660 ;
        RECT 95.510 25.410 95.740 26.410 ;
        RECT 95.890 25.960 96.180 26.270 ;
        RECT 96.450 25.570 96.740 25.900 ;
        RECT 96.900 25.410 97.150 26.410 ;
        RECT 95.510 24.410 95.990 25.410 ;
        RECT 96.240 24.710 96.470 25.410 ;
        RECT 96.190 24.370 96.520 24.710 ;
        RECT 96.720 24.550 97.150 25.410 ;
        RECT 98.010 25.290 98.350 25.630 ;
        RECT 101.650 25.300 101.970 25.620 ;
        RECT 97.560 24.730 97.900 25.050 ;
        RECT 98.430 24.740 98.760 25.010 ;
        RECT 98.620 24.550 98.760 24.740 ;
        RECT 101.210 24.720 101.530 25.040 ;
        RECT 96.720 24.410 98.760 24.550 ;
        RECT 96.930 24.390 98.760 24.410 ;
        RECT 102.780 24.220 103.080 27.200 ;
        RECT 105.740 27.130 105.880 28.880 ;
        RECT 109.730 28.430 110.060 28.710 ;
        RECT 110.490 28.470 110.660 29.200 ;
        RECT 111.400 29.190 111.690 29.200 ;
        RECT 113.230 29.020 113.460 29.890 ;
        RECT 113.230 28.880 113.590 29.020 ;
        RECT 117.270 28.890 117.500 29.890 ;
        RECT 118.210 29.500 118.510 30.660 ;
        RECT 118.650 31.690 119.050 32.280 ;
        RECT 119.250 32.020 119.580 32.340 ;
        RECT 119.300 31.690 119.530 32.020 ;
        RECT 119.780 31.690 120.290 32.340 ;
        RECT 118.650 30.690 118.880 31.690 ;
        RECT 119.030 31.240 119.320 31.550 ;
        RECT 120.040 31.290 120.290 31.690 ;
        RECT 119.590 30.850 119.880 31.180 ;
        RECT 120.040 30.960 120.390 31.290 ;
        RECT 120.040 30.690 120.290 30.960 ;
        RECT 118.650 29.690 119.130 30.690 ;
        RECT 119.380 29.990 119.610 30.690 ;
        RECT 119.330 29.650 119.660 29.990 ;
        RECT 119.860 29.710 120.290 30.690 ;
        RECT 120.670 30.070 121.000 30.360 ;
        RECT 119.860 29.690 120.090 29.710 ;
        RECT 118.210 29.340 119.400 29.500 ;
        RECT 118.200 29.200 119.400 29.340 ;
        RECT 112.960 28.470 113.290 28.700 ;
        RECT 104.610 27.060 105.880 27.130 ;
        RECT 103.390 27.000 103.620 27.060 ;
        RECT 103.220 26.410 103.620 27.000 ;
        RECT 103.820 26.740 104.150 27.060 ;
        RECT 104.350 26.990 105.880 27.060 ;
        RECT 110.490 28.330 113.290 28.470 ;
        RECT 110.490 27.510 110.660 28.330 ;
        RECT 110.490 27.200 112.090 27.510 ;
        RECT 103.870 26.410 104.100 26.740 ;
        RECT 104.350 26.410 104.860 26.990 ;
        RECT 105.460 26.660 106.630 26.800 ;
        RECT 105.460 26.460 105.780 26.660 ;
        RECT 106.340 26.460 106.660 26.660 ;
        RECT 103.220 25.410 103.450 26.410 ;
        RECT 103.600 25.960 103.890 26.270 ;
        RECT 104.160 25.570 104.450 25.900 ;
        RECT 104.610 25.410 104.860 26.410 ;
        RECT 103.220 24.410 103.700 25.410 ;
        RECT 103.950 24.710 104.180 25.410 ;
        RECT 103.900 24.370 104.230 24.710 ;
        RECT 104.430 24.550 104.860 25.410 ;
        RECT 105.720 25.290 106.060 25.630 ;
        RECT 109.360 25.300 109.680 25.620 ;
        RECT 105.270 24.730 105.610 25.050 ;
        RECT 106.140 24.740 106.470 25.010 ;
        RECT 106.330 24.550 106.470 24.740 ;
        RECT 108.920 24.720 109.240 25.040 ;
        RECT 104.430 24.410 106.470 24.550 ;
        RECT 104.640 24.390 106.470 24.410 ;
        RECT 110.490 24.220 110.790 27.200 ;
        RECT 113.450 27.130 113.590 28.880 ;
        RECT 117.440 28.430 117.770 28.710 ;
        RECT 118.200 28.470 118.370 29.200 ;
        RECT 119.110 29.190 119.400 29.200 ;
        RECT 120.940 29.020 121.170 29.890 ;
        RECT 120.940 28.880 121.300 29.020 ;
        RECT 120.670 28.470 121.000 28.700 ;
        RECT 112.320 27.060 113.590 27.130 ;
        RECT 111.100 27.000 111.330 27.060 ;
        RECT 110.930 26.410 111.330 27.000 ;
        RECT 111.530 26.740 111.860 27.060 ;
        RECT 112.060 26.990 113.590 27.060 ;
        RECT 118.200 28.330 121.000 28.470 ;
        RECT 118.200 27.510 118.370 28.330 ;
        RECT 118.200 27.200 119.800 27.510 ;
        RECT 111.580 26.410 111.810 26.740 ;
        RECT 112.060 26.410 112.570 26.990 ;
        RECT 113.170 26.660 114.340 26.800 ;
        RECT 113.170 26.460 113.490 26.660 ;
        RECT 114.050 26.460 114.370 26.660 ;
        RECT 110.930 25.410 111.160 26.410 ;
        RECT 111.310 25.960 111.600 26.270 ;
        RECT 111.870 25.570 112.160 25.900 ;
        RECT 112.320 25.410 112.570 26.410 ;
        RECT 110.930 24.410 111.410 25.410 ;
        RECT 111.660 24.710 111.890 25.410 ;
        RECT 111.610 24.370 111.940 24.710 ;
        RECT 112.140 24.550 112.570 25.410 ;
        RECT 113.430 25.290 113.770 25.630 ;
        RECT 117.070 25.300 117.390 25.620 ;
        RECT 112.980 24.730 113.320 25.050 ;
        RECT 113.850 24.740 114.180 25.010 ;
        RECT 114.040 24.550 114.180 24.740 ;
        RECT 116.630 24.720 116.950 25.040 ;
        RECT 112.140 24.410 114.180 24.550 ;
        RECT 112.350 24.390 114.180 24.410 ;
        RECT 118.200 24.220 118.500 27.200 ;
        RECT 121.160 27.130 121.300 28.880 ;
        RECT 120.030 27.060 121.300 27.130 ;
        RECT 118.810 27.000 119.040 27.060 ;
        RECT 118.640 26.410 119.040 27.000 ;
        RECT 119.240 26.740 119.570 27.060 ;
        RECT 119.770 26.990 121.300 27.060 ;
        RECT 119.290 26.410 119.520 26.740 ;
        RECT 119.770 26.410 120.280 26.990 ;
        RECT 120.880 26.660 122.050 26.800 ;
        RECT 120.880 26.460 121.200 26.660 ;
        RECT 121.760 26.460 122.080 26.660 ;
        RECT 118.640 25.410 118.870 26.410 ;
        RECT 119.020 25.960 119.310 26.270 ;
        RECT 119.580 25.570 119.870 25.900 ;
        RECT 120.030 25.410 120.280 26.410 ;
        RECT 118.640 24.410 119.120 25.410 ;
        RECT 119.370 24.710 119.600 25.410 ;
        RECT 119.320 24.370 119.650 24.710 ;
        RECT 119.850 24.550 120.280 25.410 ;
        RECT 121.140 25.290 121.480 25.630 ;
        RECT 120.690 24.730 121.030 25.050 ;
        RECT 121.560 24.740 121.890 25.010 ;
        RECT 121.750 24.550 121.890 24.740 ;
        RECT 119.850 24.410 121.890 24.550 ;
        RECT 120.060 24.390 121.890 24.410 ;
        RECT 2.550 23.920 3.740 24.220 ;
        RECT 10.260 23.920 11.450 24.220 ;
        RECT 17.970 23.920 19.160 24.220 ;
        RECT 25.680 23.920 26.870 24.220 ;
        RECT 33.390 23.920 34.580 24.220 ;
        RECT 41.100 23.920 42.290 24.220 ;
        RECT 48.810 23.920 50.000 24.220 ;
        RECT 56.520 23.920 57.710 24.220 ;
        RECT 64.230 23.920 65.420 24.220 ;
        RECT 71.940 23.920 73.130 24.220 ;
        RECT 79.650 23.920 80.840 24.220 ;
        RECT 87.360 23.920 88.550 24.220 ;
        RECT 95.070 23.920 96.260 24.220 ;
        RECT 102.780 23.920 103.970 24.220 ;
        RECT 110.490 23.920 111.680 24.220 ;
        RECT 118.200 23.920 119.390 24.220 ;
        RECT 3.450 23.910 3.740 23.920 ;
        RECT 11.160 23.910 11.450 23.920 ;
        RECT 18.870 23.910 19.160 23.920 ;
        RECT 26.580 23.910 26.870 23.920 ;
        RECT 34.290 23.910 34.580 23.920 ;
        RECT 42.000 23.910 42.290 23.920 ;
        RECT 49.710 23.910 50.000 23.920 ;
        RECT 57.420 23.910 57.710 23.920 ;
        RECT 65.130 23.910 65.420 23.920 ;
        RECT 72.840 23.910 73.130 23.920 ;
        RECT 80.550 23.910 80.840 23.920 ;
        RECT 88.260 23.910 88.550 23.920 ;
        RECT 95.970 23.910 96.260 23.920 ;
        RECT 103.680 23.910 103.970 23.920 ;
        RECT 111.390 23.910 111.680 23.920 ;
        RECT 119.100 23.910 119.390 23.920 ;
        RECT 28.660 20.540 29.010 20.930 ;
        RECT 90.310 20.560 90.660 20.890 ;
        RECT 58.500 20.110 58.820 20.160 ;
        RECT 58.490 19.850 58.820 20.110 ;
        RECT 58.500 19.840 58.820 19.850 ;
        RECT 58.980 16.420 59.320 16.750 ;
        RECT 58.510 15.800 58.840 16.120 ;
        RECT 124.510 15.830 124.860 16.150 ;
        RECT 124.510 15.810 124.850 15.830 ;
        RECT 58.400 13.900 58.740 13.940 ;
        RECT 58.400 13.640 58.760 13.900 ;
        RECT 58.400 13.610 58.740 13.640 ;
        RECT 28.780 11.890 29.150 12.290 ;
        RECT 90.430 11.910 90.810 12.280 ;
        RECT 28.790 11.880 29.140 11.890 ;
        RECT 3.650 9.540 3.940 9.550 ;
        RECT 11.360 9.540 11.650 9.550 ;
        RECT 19.070 9.540 19.360 9.550 ;
        RECT 26.780 9.540 27.070 9.550 ;
        RECT 34.490 9.540 34.780 9.550 ;
        RECT 42.200 9.540 42.490 9.550 ;
        RECT 49.910 9.540 50.200 9.550 ;
        RECT 57.620 9.540 57.910 9.550 ;
        RECT 65.330 9.540 65.620 9.550 ;
        RECT 73.040 9.540 73.330 9.550 ;
        RECT 80.750 9.540 81.040 9.550 ;
        RECT 88.460 9.540 88.750 9.550 ;
        RECT 96.170 9.540 96.460 9.550 ;
        RECT 103.880 9.540 104.170 9.550 ;
        RECT 111.590 9.540 111.880 9.550 ;
        RECT 119.300 9.540 119.590 9.550 ;
        RECT 3.650 9.240 4.840 9.540 ;
        RECT 11.360 9.240 12.550 9.540 ;
        RECT 19.070 9.240 20.260 9.540 ;
        RECT 26.780 9.240 27.970 9.540 ;
        RECT 34.490 9.240 35.680 9.540 ;
        RECT 42.200 9.240 43.390 9.540 ;
        RECT 49.910 9.240 51.100 9.540 ;
        RECT 57.620 9.240 58.810 9.540 ;
        RECT 65.330 9.240 66.520 9.540 ;
        RECT 73.040 9.240 74.230 9.540 ;
        RECT 80.750 9.240 81.940 9.540 ;
        RECT 88.460 9.240 89.650 9.540 ;
        RECT 96.170 9.240 97.360 9.540 ;
        RECT 103.880 9.240 105.070 9.540 ;
        RECT 111.590 9.240 112.780 9.540 ;
        RECT 119.300 9.240 120.490 9.540 ;
        RECT 1.150 9.050 2.980 9.070 ;
        RECT 1.150 8.910 3.190 9.050 ;
        RECT 1.150 8.720 1.290 8.910 ;
        RECT 1.150 8.450 1.480 8.720 ;
        RECT 2.010 8.410 2.350 8.730 ;
        RECT 1.560 7.830 1.900 8.170 ;
        RECT 2.760 8.050 3.190 8.910 ;
        RECT 3.390 8.750 3.720 9.090 ;
        RECT 3.440 8.050 3.670 8.750 ;
        RECT 3.920 8.050 4.400 9.050 ;
        RECT 2.760 7.050 3.010 8.050 ;
        RECT 3.170 7.560 3.460 7.890 ;
        RECT 3.730 7.190 4.020 7.500 ;
        RECT 4.170 7.050 4.400 8.050 ;
        RECT 0.960 6.800 1.280 7.000 ;
        RECT 1.840 6.800 2.160 7.000 ;
        RECT 0.990 6.660 2.160 6.800 ;
        RECT 2.760 6.470 3.270 7.050 ;
        RECT 3.520 6.720 3.750 7.050 ;
        RECT 1.740 6.400 3.270 6.470 ;
        RECT 3.470 6.400 3.800 6.720 ;
        RECT 4.000 6.460 4.400 7.050 ;
        RECT 4.000 6.400 4.230 6.460 ;
        RECT 1.740 6.330 3.010 6.400 ;
        RECT 1.740 4.580 1.880 6.330 ;
        RECT 4.540 6.260 4.840 9.240 ;
        RECT 8.860 9.050 10.690 9.070 ;
        RECT 8.860 8.910 10.900 9.050 ;
        RECT 6.090 8.420 6.410 8.740 ;
        RECT 8.860 8.720 9.000 8.910 ;
        RECT 8.860 8.450 9.190 8.720 ;
        RECT 9.720 8.410 10.060 8.730 ;
        RECT 5.650 7.840 5.970 8.160 ;
        RECT 9.270 7.830 9.610 8.170 ;
        RECT 10.470 8.050 10.900 8.910 ;
        RECT 11.100 8.750 11.430 9.090 ;
        RECT 11.150 8.050 11.380 8.750 ;
        RECT 11.630 8.050 12.110 9.050 ;
        RECT 10.470 7.050 10.720 8.050 ;
        RECT 10.880 7.560 11.170 7.890 ;
        RECT 11.440 7.190 11.730 7.500 ;
        RECT 11.880 7.050 12.110 8.050 ;
        RECT 8.670 6.800 8.990 7.000 ;
        RECT 9.550 6.800 9.870 7.000 ;
        RECT 8.700 6.660 9.870 6.800 ;
        RECT 10.470 6.470 10.980 7.050 ;
        RECT 11.230 6.720 11.460 7.050 ;
        RECT 3.240 5.950 4.840 6.260 ;
        RECT 4.670 5.130 4.840 5.950 ;
        RECT 2.040 4.990 4.840 5.130 ;
        RECT 9.450 6.400 10.980 6.470 ;
        RECT 11.180 6.400 11.510 6.720 ;
        RECT 11.710 6.460 12.110 7.050 ;
        RECT 11.710 6.400 11.940 6.460 ;
        RECT 9.450 6.330 10.720 6.400 ;
        RECT 2.040 4.760 2.370 4.990 ;
        RECT 1.740 4.440 2.100 4.580 ;
        RECT 1.870 3.570 2.100 4.440 ;
        RECT 3.640 4.260 3.930 4.270 ;
        RECT 4.670 4.260 4.840 4.990 ;
        RECT 5.270 4.750 5.600 5.030 ;
        RECT 9.450 4.580 9.590 6.330 ;
        RECT 12.250 6.260 12.550 9.240 ;
        RECT 16.570 9.050 18.400 9.070 ;
        RECT 16.570 8.910 18.610 9.050 ;
        RECT 13.800 8.420 14.120 8.740 ;
        RECT 16.570 8.720 16.710 8.910 ;
        RECT 16.570 8.450 16.900 8.720 ;
        RECT 17.430 8.410 17.770 8.730 ;
        RECT 13.360 7.840 13.680 8.160 ;
        RECT 16.980 7.830 17.320 8.170 ;
        RECT 18.180 8.050 18.610 8.910 ;
        RECT 18.810 8.750 19.140 9.090 ;
        RECT 18.860 8.050 19.090 8.750 ;
        RECT 19.340 8.050 19.820 9.050 ;
        RECT 18.180 7.050 18.430 8.050 ;
        RECT 18.590 7.560 18.880 7.890 ;
        RECT 19.150 7.190 19.440 7.500 ;
        RECT 19.590 7.050 19.820 8.050 ;
        RECT 16.380 6.800 16.700 7.000 ;
        RECT 17.260 6.800 17.580 7.000 ;
        RECT 16.410 6.660 17.580 6.800 ;
        RECT 18.180 6.470 18.690 7.050 ;
        RECT 18.940 6.720 19.170 7.050 ;
        RECT 10.950 5.950 12.550 6.260 ;
        RECT 12.380 5.130 12.550 5.950 ;
        RECT 9.750 4.990 12.550 5.130 ;
        RECT 17.160 6.400 18.690 6.470 ;
        RECT 18.890 6.400 19.220 6.720 ;
        RECT 19.420 6.460 19.820 7.050 ;
        RECT 19.420 6.400 19.650 6.460 ;
        RECT 17.160 6.330 18.430 6.400 ;
        RECT 9.750 4.760 10.080 4.990 ;
        RECT 3.640 4.120 4.840 4.260 ;
        RECT 3.640 3.960 4.830 4.120 ;
        RECT 2.950 3.750 3.180 3.770 ;
        RECT 2.040 3.100 2.370 3.390 ;
        RECT 2.750 2.770 3.180 3.750 ;
        RECT 3.380 3.470 3.710 3.810 ;
        RECT 3.430 2.770 3.660 3.470 ;
        RECT 3.910 2.770 4.390 3.770 ;
        RECT 2.750 2.500 3.000 2.770 ;
        RECT 2.650 2.170 3.000 2.500 ;
        RECT 3.160 2.280 3.450 2.610 ;
        RECT 2.750 1.770 3.000 2.170 ;
        RECT 3.720 1.910 4.010 2.220 ;
        RECT 4.160 1.770 4.390 2.770 ;
        RECT 2.750 1.120 3.260 1.770 ;
        RECT 3.510 1.440 3.740 1.770 ;
        RECT 3.460 1.120 3.790 1.440 ;
        RECT 3.990 1.180 4.390 1.770 ;
        RECT 4.530 2.800 4.830 3.960 ;
        RECT 5.540 3.570 5.770 4.570 ;
        RECT 9.450 4.440 9.810 4.580 ;
        RECT 9.580 3.570 9.810 4.440 ;
        RECT 11.350 4.260 11.640 4.270 ;
        RECT 12.380 4.260 12.550 4.990 ;
        RECT 12.980 4.750 13.310 5.030 ;
        RECT 17.160 4.580 17.300 6.330 ;
        RECT 19.960 6.260 20.260 9.240 ;
        RECT 24.280 9.050 26.110 9.070 ;
        RECT 24.280 8.910 26.320 9.050 ;
        RECT 21.510 8.420 21.830 8.740 ;
        RECT 24.280 8.720 24.420 8.910 ;
        RECT 24.280 8.450 24.610 8.720 ;
        RECT 25.140 8.410 25.480 8.730 ;
        RECT 21.070 7.840 21.390 8.160 ;
        RECT 24.690 7.830 25.030 8.170 ;
        RECT 25.890 8.050 26.320 8.910 ;
        RECT 26.520 8.750 26.850 9.090 ;
        RECT 26.570 8.050 26.800 8.750 ;
        RECT 27.050 8.050 27.530 9.050 ;
        RECT 25.890 7.050 26.140 8.050 ;
        RECT 26.300 7.560 26.590 7.890 ;
        RECT 26.860 7.190 27.150 7.500 ;
        RECT 27.300 7.050 27.530 8.050 ;
        RECT 24.090 6.800 24.410 7.000 ;
        RECT 24.970 6.800 25.290 7.000 ;
        RECT 24.120 6.660 25.290 6.800 ;
        RECT 25.890 6.470 26.400 7.050 ;
        RECT 26.650 6.720 26.880 7.050 ;
        RECT 18.660 5.950 20.260 6.260 ;
        RECT 20.090 5.130 20.260 5.950 ;
        RECT 17.460 4.990 20.260 5.130 ;
        RECT 24.870 6.400 26.400 6.470 ;
        RECT 26.600 6.400 26.930 6.720 ;
        RECT 27.130 6.460 27.530 7.050 ;
        RECT 27.130 6.400 27.360 6.460 ;
        RECT 24.870 6.330 26.140 6.400 ;
        RECT 17.460 4.760 17.790 4.990 ;
        RECT 11.350 4.120 12.550 4.260 ;
        RECT 11.350 3.960 12.540 4.120 ;
        RECT 10.660 3.750 10.890 3.770 ;
        RECT 5.270 3.120 5.600 3.400 ;
        RECT 9.750 3.100 10.080 3.390 ;
        RECT 6.880 2.800 7.170 2.970 ;
        RECT 4.530 2.630 7.170 2.800 ;
        RECT 10.460 2.770 10.890 3.750 ;
        RECT 11.090 3.470 11.420 3.810 ;
        RECT 11.140 2.770 11.370 3.470 ;
        RECT 11.620 2.770 12.100 3.770 ;
        RECT 3.990 1.120 4.220 1.180 ;
        RECT 4.530 0.980 4.830 2.630 ;
        RECT 10.460 2.500 10.710 2.770 ;
        RECT 5.060 2.090 5.440 2.410 ;
        RECT 10.360 2.170 10.710 2.500 ;
        RECT 10.870 2.280 11.160 2.610 ;
        RECT 10.460 1.770 10.710 2.170 ;
        RECT 11.430 1.910 11.720 2.220 ;
        RECT 11.870 1.770 12.100 2.770 ;
        RECT 10.460 1.120 10.970 1.770 ;
        RECT 11.220 1.440 11.450 1.770 ;
        RECT 11.170 1.120 11.500 1.440 ;
        RECT 11.700 1.180 12.100 1.770 ;
        RECT 12.240 2.800 12.540 3.960 ;
        RECT 13.250 3.570 13.480 4.570 ;
        RECT 17.160 4.440 17.520 4.580 ;
        RECT 17.290 3.570 17.520 4.440 ;
        RECT 19.060 4.260 19.350 4.270 ;
        RECT 20.090 4.260 20.260 4.990 ;
        RECT 20.690 4.750 21.020 5.030 ;
        RECT 24.870 4.580 25.010 6.330 ;
        RECT 27.670 6.260 27.970 9.240 ;
        RECT 31.990 9.050 33.820 9.070 ;
        RECT 31.990 8.910 34.030 9.050 ;
        RECT 29.220 8.420 29.540 8.740 ;
        RECT 31.990 8.720 32.130 8.910 ;
        RECT 31.990 8.450 32.320 8.720 ;
        RECT 32.850 8.410 33.190 8.730 ;
        RECT 28.780 7.840 29.100 8.160 ;
        RECT 32.400 7.830 32.740 8.170 ;
        RECT 33.600 8.050 34.030 8.910 ;
        RECT 34.230 8.750 34.560 9.090 ;
        RECT 34.280 8.050 34.510 8.750 ;
        RECT 34.760 8.050 35.240 9.050 ;
        RECT 33.600 7.050 33.850 8.050 ;
        RECT 34.010 7.560 34.300 7.890 ;
        RECT 34.570 7.190 34.860 7.500 ;
        RECT 35.010 7.050 35.240 8.050 ;
        RECT 31.800 6.800 32.120 7.000 ;
        RECT 32.680 6.800 33.000 7.000 ;
        RECT 31.830 6.660 33.000 6.800 ;
        RECT 33.600 6.470 34.110 7.050 ;
        RECT 34.360 6.720 34.590 7.050 ;
        RECT 26.370 5.950 27.970 6.260 ;
        RECT 27.800 5.130 27.970 5.950 ;
        RECT 25.170 4.990 27.970 5.130 ;
        RECT 32.580 6.400 34.110 6.470 ;
        RECT 34.310 6.400 34.640 6.720 ;
        RECT 34.840 6.460 35.240 7.050 ;
        RECT 34.840 6.400 35.070 6.460 ;
        RECT 32.580 6.330 33.850 6.400 ;
        RECT 25.170 4.760 25.500 4.990 ;
        RECT 19.060 4.120 20.260 4.260 ;
        RECT 19.060 3.960 20.250 4.120 ;
        RECT 18.370 3.750 18.600 3.770 ;
        RECT 12.980 3.120 13.310 3.400 ;
        RECT 17.460 3.100 17.790 3.390 ;
        RECT 14.590 2.800 14.880 2.970 ;
        RECT 12.240 2.630 14.880 2.800 ;
        RECT 18.170 2.770 18.600 3.750 ;
        RECT 18.800 3.470 19.130 3.810 ;
        RECT 18.850 2.770 19.080 3.470 ;
        RECT 19.330 2.770 19.810 3.770 ;
        RECT 11.700 1.120 11.930 1.180 ;
        RECT 12.240 0.980 12.540 2.630 ;
        RECT 18.170 2.500 18.420 2.770 ;
        RECT 12.770 2.090 13.150 2.410 ;
        RECT 18.070 2.170 18.420 2.500 ;
        RECT 18.580 2.280 18.870 2.610 ;
        RECT 18.170 1.770 18.420 2.170 ;
        RECT 19.140 1.910 19.430 2.220 ;
        RECT 19.580 1.770 19.810 2.770 ;
        RECT 18.170 1.120 18.680 1.770 ;
        RECT 18.930 1.440 19.160 1.770 ;
        RECT 18.880 1.120 19.210 1.440 ;
        RECT 19.410 1.180 19.810 1.770 ;
        RECT 19.950 2.800 20.250 3.960 ;
        RECT 20.960 3.570 21.190 4.570 ;
        RECT 24.870 4.440 25.230 4.580 ;
        RECT 25.000 3.570 25.230 4.440 ;
        RECT 26.770 4.260 27.060 4.270 ;
        RECT 27.800 4.260 27.970 4.990 ;
        RECT 28.400 4.750 28.730 5.030 ;
        RECT 32.580 4.580 32.720 6.330 ;
        RECT 35.380 6.260 35.680 9.240 ;
        RECT 39.700 9.050 41.530 9.070 ;
        RECT 39.700 8.910 41.740 9.050 ;
        RECT 36.930 8.420 37.250 8.740 ;
        RECT 39.700 8.720 39.840 8.910 ;
        RECT 39.700 8.450 40.030 8.720 ;
        RECT 40.560 8.410 40.900 8.730 ;
        RECT 36.490 7.840 36.810 8.160 ;
        RECT 40.110 7.830 40.450 8.170 ;
        RECT 41.310 8.050 41.740 8.910 ;
        RECT 41.940 8.750 42.270 9.090 ;
        RECT 41.990 8.050 42.220 8.750 ;
        RECT 42.470 8.050 42.950 9.050 ;
        RECT 41.310 7.050 41.560 8.050 ;
        RECT 41.720 7.560 42.010 7.890 ;
        RECT 42.280 7.190 42.570 7.500 ;
        RECT 42.720 7.050 42.950 8.050 ;
        RECT 39.510 6.800 39.830 7.000 ;
        RECT 40.390 6.800 40.710 7.000 ;
        RECT 39.540 6.660 40.710 6.800 ;
        RECT 41.310 6.470 41.820 7.050 ;
        RECT 42.070 6.720 42.300 7.050 ;
        RECT 34.080 5.950 35.680 6.260 ;
        RECT 35.510 5.130 35.680 5.950 ;
        RECT 32.880 4.990 35.680 5.130 ;
        RECT 40.290 6.400 41.820 6.470 ;
        RECT 42.020 6.400 42.350 6.720 ;
        RECT 42.550 6.460 42.950 7.050 ;
        RECT 42.550 6.400 42.780 6.460 ;
        RECT 40.290 6.330 41.560 6.400 ;
        RECT 32.880 4.760 33.210 4.990 ;
        RECT 26.770 4.120 27.970 4.260 ;
        RECT 26.770 3.960 27.960 4.120 ;
        RECT 26.080 3.750 26.310 3.770 ;
        RECT 20.690 3.120 21.020 3.400 ;
        RECT 25.170 3.100 25.500 3.390 ;
        RECT 22.300 2.800 22.590 2.970 ;
        RECT 19.950 2.630 22.590 2.800 ;
        RECT 25.880 2.770 26.310 3.750 ;
        RECT 26.510 3.470 26.840 3.810 ;
        RECT 26.560 2.770 26.790 3.470 ;
        RECT 27.040 2.770 27.520 3.770 ;
        RECT 19.410 1.120 19.640 1.180 ;
        RECT 19.950 0.980 20.250 2.630 ;
        RECT 25.880 2.500 26.130 2.770 ;
        RECT 20.480 2.090 20.860 2.410 ;
        RECT 25.780 2.170 26.130 2.500 ;
        RECT 26.290 2.280 26.580 2.610 ;
        RECT 25.880 1.770 26.130 2.170 ;
        RECT 26.850 1.910 27.140 2.220 ;
        RECT 27.290 1.770 27.520 2.770 ;
        RECT 25.880 1.120 26.390 1.770 ;
        RECT 26.640 1.440 26.870 1.770 ;
        RECT 26.590 1.120 26.920 1.440 ;
        RECT 27.120 1.180 27.520 1.770 ;
        RECT 27.660 2.800 27.960 3.960 ;
        RECT 28.670 3.570 28.900 4.570 ;
        RECT 32.580 4.440 32.940 4.580 ;
        RECT 32.710 3.570 32.940 4.440 ;
        RECT 34.480 4.260 34.770 4.270 ;
        RECT 35.510 4.260 35.680 4.990 ;
        RECT 36.110 4.750 36.440 5.030 ;
        RECT 40.290 4.580 40.430 6.330 ;
        RECT 43.090 6.260 43.390 9.240 ;
        RECT 47.410 9.050 49.240 9.070 ;
        RECT 47.410 8.910 49.450 9.050 ;
        RECT 44.640 8.420 44.960 8.740 ;
        RECT 47.410 8.720 47.550 8.910 ;
        RECT 47.410 8.450 47.740 8.720 ;
        RECT 48.270 8.410 48.610 8.730 ;
        RECT 44.200 7.840 44.520 8.160 ;
        RECT 47.820 7.830 48.160 8.170 ;
        RECT 49.020 8.050 49.450 8.910 ;
        RECT 49.650 8.750 49.980 9.090 ;
        RECT 49.700 8.050 49.930 8.750 ;
        RECT 50.180 8.050 50.660 9.050 ;
        RECT 49.020 7.050 49.270 8.050 ;
        RECT 49.430 7.560 49.720 7.890 ;
        RECT 49.990 7.190 50.280 7.500 ;
        RECT 50.430 7.050 50.660 8.050 ;
        RECT 47.220 6.800 47.540 7.000 ;
        RECT 48.100 6.800 48.420 7.000 ;
        RECT 47.250 6.660 48.420 6.800 ;
        RECT 49.020 6.470 49.530 7.050 ;
        RECT 49.780 6.720 50.010 7.050 ;
        RECT 41.790 5.950 43.390 6.260 ;
        RECT 43.220 5.130 43.390 5.950 ;
        RECT 40.590 4.990 43.390 5.130 ;
        RECT 48.000 6.400 49.530 6.470 ;
        RECT 49.730 6.400 50.060 6.720 ;
        RECT 50.260 6.460 50.660 7.050 ;
        RECT 50.260 6.400 50.490 6.460 ;
        RECT 48.000 6.330 49.270 6.400 ;
        RECT 40.590 4.760 40.920 4.990 ;
        RECT 34.480 4.120 35.680 4.260 ;
        RECT 34.480 3.960 35.670 4.120 ;
        RECT 33.790 3.750 34.020 3.770 ;
        RECT 28.400 3.120 28.730 3.400 ;
        RECT 32.880 3.100 33.210 3.390 ;
        RECT 30.010 2.800 30.300 2.970 ;
        RECT 27.660 2.630 30.300 2.800 ;
        RECT 33.590 2.770 34.020 3.750 ;
        RECT 34.220 3.470 34.550 3.810 ;
        RECT 34.270 2.770 34.500 3.470 ;
        RECT 34.750 2.770 35.230 3.770 ;
        RECT 27.120 1.120 27.350 1.180 ;
        RECT 27.660 0.980 27.960 2.630 ;
        RECT 33.590 2.500 33.840 2.770 ;
        RECT 28.190 2.090 28.570 2.410 ;
        RECT 33.490 2.170 33.840 2.500 ;
        RECT 34.000 2.280 34.290 2.610 ;
        RECT 33.590 1.770 33.840 2.170 ;
        RECT 34.560 1.910 34.850 2.220 ;
        RECT 35.000 1.770 35.230 2.770 ;
        RECT 33.590 1.120 34.100 1.770 ;
        RECT 34.350 1.440 34.580 1.770 ;
        RECT 34.300 1.120 34.630 1.440 ;
        RECT 34.830 1.180 35.230 1.770 ;
        RECT 35.370 2.800 35.670 3.960 ;
        RECT 36.380 3.570 36.610 4.570 ;
        RECT 40.290 4.440 40.650 4.580 ;
        RECT 40.420 3.570 40.650 4.440 ;
        RECT 42.190 4.260 42.480 4.270 ;
        RECT 43.220 4.260 43.390 4.990 ;
        RECT 43.820 4.750 44.150 5.030 ;
        RECT 48.000 4.580 48.140 6.330 ;
        RECT 50.800 6.260 51.100 9.240 ;
        RECT 55.120 9.050 56.950 9.070 ;
        RECT 55.120 8.910 57.160 9.050 ;
        RECT 52.350 8.420 52.670 8.740 ;
        RECT 55.120 8.720 55.260 8.910 ;
        RECT 55.120 8.450 55.450 8.720 ;
        RECT 55.980 8.410 56.320 8.730 ;
        RECT 51.910 7.840 52.230 8.160 ;
        RECT 55.530 7.830 55.870 8.170 ;
        RECT 56.730 8.050 57.160 8.910 ;
        RECT 57.360 8.750 57.690 9.090 ;
        RECT 57.410 8.050 57.640 8.750 ;
        RECT 57.890 8.050 58.370 9.050 ;
        RECT 56.730 7.050 56.980 8.050 ;
        RECT 57.140 7.560 57.430 7.890 ;
        RECT 57.700 7.190 57.990 7.500 ;
        RECT 58.140 7.050 58.370 8.050 ;
        RECT 54.930 6.800 55.250 7.000 ;
        RECT 55.810 6.800 56.130 7.000 ;
        RECT 54.960 6.660 56.130 6.800 ;
        RECT 56.730 6.470 57.240 7.050 ;
        RECT 57.490 6.720 57.720 7.050 ;
        RECT 49.500 5.950 51.100 6.260 ;
        RECT 50.930 5.130 51.100 5.950 ;
        RECT 48.300 4.990 51.100 5.130 ;
        RECT 55.710 6.400 57.240 6.470 ;
        RECT 57.440 6.400 57.770 6.720 ;
        RECT 57.970 6.460 58.370 7.050 ;
        RECT 57.970 6.400 58.200 6.460 ;
        RECT 55.710 6.330 56.980 6.400 ;
        RECT 48.300 4.760 48.630 4.990 ;
        RECT 42.190 4.120 43.390 4.260 ;
        RECT 42.190 3.960 43.380 4.120 ;
        RECT 41.500 3.750 41.730 3.770 ;
        RECT 36.110 3.120 36.440 3.400 ;
        RECT 40.590 3.100 40.920 3.390 ;
        RECT 37.720 2.800 38.010 2.970 ;
        RECT 35.370 2.630 38.010 2.800 ;
        RECT 41.300 2.770 41.730 3.750 ;
        RECT 41.930 3.470 42.260 3.810 ;
        RECT 41.980 2.770 42.210 3.470 ;
        RECT 42.460 2.770 42.940 3.770 ;
        RECT 34.830 1.120 35.060 1.180 ;
        RECT 35.370 0.980 35.670 2.630 ;
        RECT 41.300 2.500 41.550 2.770 ;
        RECT 35.900 2.090 36.280 2.410 ;
        RECT 41.200 2.170 41.550 2.500 ;
        RECT 41.710 2.280 42.000 2.610 ;
        RECT 41.300 1.770 41.550 2.170 ;
        RECT 42.270 1.910 42.560 2.220 ;
        RECT 42.710 1.770 42.940 2.770 ;
        RECT 41.300 1.120 41.810 1.770 ;
        RECT 42.060 1.440 42.290 1.770 ;
        RECT 42.010 1.120 42.340 1.440 ;
        RECT 42.540 1.180 42.940 1.770 ;
        RECT 43.080 2.800 43.380 3.960 ;
        RECT 44.090 3.570 44.320 4.570 ;
        RECT 48.000 4.440 48.360 4.580 ;
        RECT 48.130 3.570 48.360 4.440 ;
        RECT 49.900 4.260 50.190 4.270 ;
        RECT 50.930 4.260 51.100 4.990 ;
        RECT 51.530 4.750 51.860 5.030 ;
        RECT 55.710 4.580 55.850 6.330 ;
        RECT 58.510 6.260 58.810 9.240 ;
        RECT 62.830 9.050 64.660 9.070 ;
        RECT 62.830 8.910 64.870 9.050 ;
        RECT 60.060 8.420 60.380 8.740 ;
        RECT 62.830 8.720 62.970 8.910 ;
        RECT 62.830 8.450 63.160 8.720 ;
        RECT 63.690 8.410 64.030 8.730 ;
        RECT 59.620 7.840 59.940 8.160 ;
        RECT 63.240 7.830 63.580 8.170 ;
        RECT 64.440 8.050 64.870 8.910 ;
        RECT 65.070 8.750 65.400 9.090 ;
        RECT 65.120 8.050 65.350 8.750 ;
        RECT 65.600 8.050 66.080 9.050 ;
        RECT 64.440 7.050 64.690 8.050 ;
        RECT 64.850 7.560 65.140 7.890 ;
        RECT 65.410 7.190 65.700 7.500 ;
        RECT 65.850 7.050 66.080 8.050 ;
        RECT 62.640 6.800 62.960 7.000 ;
        RECT 63.520 6.800 63.840 7.000 ;
        RECT 62.670 6.660 63.840 6.800 ;
        RECT 64.440 6.470 64.950 7.050 ;
        RECT 65.200 6.720 65.430 7.050 ;
        RECT 57.210 5.950 58.810 6.260 ;
        RECT 58.640 5.130 58.810 5.950 ;
        RECT 56.010 4.990 58.810 5.130 ;
        RECT 63.420 6.400 64.950 6.470 ;
        RECT 65.150 6.400 65.480 6.720 ;
        RECT 65.680 6.460 66.080 7.050 ;
        RECT 65.680 6.400 65.910 6.460 ;
        RECT 63.420 6.330 64.690 6.400 ;
        RECT 56.010 4.760 56.340 4.990 ;
        RECT 49.900 4.120 51.100 4.260 ;
        RECT 49.900 3.960 51.090 4.120 ;
        RECT 49.210 3.750 49.440 3.770 ;
        RECT 43.820 3.120 44.150 3.400 ;
        RECT 48.300 3.100 48.630 3.390 ;
        RECT 45.430 2.800 45.720 2.970 ;
        RECT 43.080 2.630 45.720 2.800 ;
        RECT 49.010 2.770 49.440 3.750 ;
        RECT 49.640 3.470 49.970 3.810 ;
        RECT 49.690 2.770 49.920 3.470 ;
        RECT 50.170 2.770 50.650 3.770 ;
        RECT 42.540 1.120 42.770 1.180 ;
        RECT 43.080 0.980 43.380 2.630 ;
        RECT 49.010 2.500 49.260 2.770 ;
        RECT 43.610 2.090 43.990 2.410 ;
        RECT 48.910 2.170 49.260 2.500 ;
        RECT 49.420 2.280 49.710 2.610 ;
        RECT 49.010 1.770 49.260 2.170 ;
        RECT 49.980 1.910 50.270 2.220 ;
        RECT 50.420 1.770 50.650 2.770 ;
        RECT 49.010 1.120 49.520 1.770 ;
        RECT 49.770 1.440 50.000 1.770 ;
        RECT 49.720 1.120 50.050 1.440 ;
        RECT 50.250 1.180 50.650 1.770 ;
        RECT 50.790 2.800 51.090 3.960 ;
        RECT 51.800 3.570 52.030 4.570 ;
        RECT 55.710 4.440 56.070 4.580 ;
        RECT 55.840 3.570 56.070 4.440 ;
        RECT 57.610 4.260 57.900 4.270 ;
        RECT 58.640 4.260 58.810 4.990 ;
        RECT 59.240 4.750 59.570 5.030 ;
        RECT 63.420 4.580 63.560 6.330 ;
        RECT 66.220 6.260 66.520 9.240 ;
        RECT 70.540 9.050 72.370 9.070 ;
        RECT 70.540 8.910 72.580 9.050 ;
        RECT 67.770 8.420 68.090 8.740 ;
        RECT 70.540 8.720 70.680 8.910 ;
        RECT 70.540 8.450 70.870 8.720 ;
        RECT 71.400 8.410 71.740 8.730 ;
        RECT 67.330 7.840 67.650 8.160 ;
        RECT 70.950 7.830 71.290 8.170 ;
        RECT 72.150 8.050 72.580 8.910 ;
        RECT 72.780 8.750 73.110 9.090 ;
        RECT 72.830 8.050 73.060 8.750 ;
        RECT 73.310 8.050 73.790 9.050 ;
        RECT 72.150 7.050 72.400 8.050 ;
        RECT 72.560 7.560 72.850 7.890 ;
        RECT 73.120 7.190 73.410 7.500 ;
        RECT 73.560 7.050 73.790 8.050 ;
        RECT 70.350 6.800 70.670 7.000 ;
        RECT 71.230 6.800 71.550 7.000 ;
        RECT 70.380 6.660 71.550 6.800 ;
        RECT 72.150 6.470 72.660 7.050 ;
        RECT 72.910 6.720 73.140 7.050 ;
        RECT 64.920 5.950 66.520 6.260 ;
        RECT 66.350 5.130 66.520 5.950 ;
        RECT 63.720 4.990 66.520 5.130 ;
        RECT 71.130 6.400 72.660 6.470 ;
        RECT 72.860 6.400 73.190 6.720 ;
        RECT 73.390 6.460 73.790 7.050 ;
        RECT 73.390 6.400 73.620 6.460 ;
        RECT 71.130 6.330 72.400 6.400 ;
        RECT 63.720 4.760 64.050 4.990 ;
        RECT 57.610 4.120 58.810 4.260 ;
        RECT 57.610 3.960 58.800 4.120 ;
        RECT 56.920 3.750 57.150 3.770 ;
        RECT 51.530 3.120 51.860 3.400 ;
        RECT 56.010 3.100 56.340 3.390 ;
        RECT 53.140 2.800 53.430 2.970 ;
        RECT 50.790 2.630 53.430 2.800 ;
        RECT 56.720 2.770 57.150 3.750 ;
        RECT 57.350 3.470 57.680 3.810 ;
        RECT 57.400 2.770 57.630 3.470 ;
        RECT 57.880 2.770 58.360 3.770 ;
        RECT 50.250 1.120 50.480 1.180 ;
        RECT 50.790 0.980 51.090 2.630 ;
        RECT 56.720 2.500 56.970 2.770 ;
        RECT 51.320 2.090 51.700 2.410 ;
        RECT 56.620 2.170 56.970 2.500 ;
        RECT 57.130 2.280 57.420 2.610 ;
        RECT 56.720 1.770 56.970 2.170 ;
        RECT 57.690 1.910 57.980 2.220 ;
        RECT 58.130 1.770 58.360 2.770 ;
        RECT 56.720 1.120 57.230 1.770 ;
        RECT 57.480 1.440 57.710 1.770 ;
        RECT 57.430 1.120 57.760 1.440 ;
        RECT 57.960 1.180 58.360 1.770 ;
        RECT 58.500 2.800 58.800 3.960 ;
        RECT 59.510 3.570 59.740 4.570 ;
        RECT 63.420 4.440 63.780 4.580 ;
        RECT 63.550 3.570 63.780 4.440 ;
        RECT 65.320 4.260 65.610 4.270 ;
        RECT 66.350 4.260 66.520 4.990 ;
        RECT 66.950 4.750 67.280 5.030 ;
        RECT 71.130 4.580 71.270 6.330 ;
        RECT 73.930 6.260 74.230 9.240 ;
        RECT 78.250 9.050 80.080 9.070 ;
        RECT 78.250 8.910 80.290 9.050 ;
        RECT 75.480 8.420 75.800 8.740 ;
        RECT 78.250 8.720 78.390 8.910 ;
        RECT 78.250 8.450 78.580 8.720 ;
        RECT 79.110 8.410 79.450 8.730 ;
        RECT 75.040 7.840 75.360 8.160 ;
        RECT 78.660 7.830 79.000 8.170 ;
        RECT 79.860 8.050 80.290 8.910 ;
        RECT 80.490 8.750 80.820 9.090 ;
        RECT 80.540 8.050 80.770 8.750 ;
        RECT 81.020 8.050 81.500 9.050 ;
        RECT 79.860 7.050 80.110 8.050 ;
        RECT 80.270 7.560 80.560 7.890 ;
        RECT 80.830 7.190 81.120 7.500 ;
        RECT 81.270 7.050 81.500 8.050 ;
        RECT 78.060 6.800 78.380 7.000 ;
        RECT 78.940 6.800 79.260 7.000 ;
        RECT 78.090 6.660 79.260 6.800 ;
        RECT 79.860 6.470 80.370 7.050 ;
        RECT 80.620 6.720 80.850 7.050 ;
        RECT 72.630 5.950 74.230 6.260 ;
        RECT 74.060 5.130 74.230 5.950 ;
        RECT 71.430 4.990 74.230 5.130 ;
        RECT 78.840 6.400 80.370 6.470 ;
        RECT 80.570 6.400 80.900 6.720 ;
        RECT 81.100 6.460 81.500 7.050 ;
        RECT 81.100 6.400 81.330 6.460 ;
        RECT 78.840 6.330 80.110 6.400 ;
        RECT 71.430 4.760 71.760 4.990 ;
        RECT 65.320 4.120 66.520 4.260 ;
        RECT 65.320 3.960 66.510 4.120 ;
        RECT 64.630 3.750 64.860 3.770 ;
        RECT 59.240 3.120 59.570 3.400 ;
        RECT 63.720 3.100 64.050 3.390 ;
        RECT 60.850 2.800 61.140 2.970 ;
        RECT 58.500 2.630 61.140 2.800 ;
        RECT 64.430 2.770 64.860 3.750 ;
        RECT 65.060 3.470 65.390 3.810 ;
        RECT 65.110 2.770 65.340 3.470 ;
        RECT 65.590 2.770 66.070 3.770 ;
        RECT 57.960 1.120 58.190 1.180 ;
        RECT 58.500 0.980 58.800 2.630 ;
        RECT 64.430 2.500 64.680 2.770 ;
        RECT 59.030 2.090 59.410 2.410 ;
        RECT 64.330 2.170 64.680 2.500 ;
        RECT 64.840 2.280 65.130 2.610 ;
        RECT 64.430 1.770 64.680 2.170 ;
        RECT 65.400 1.910 65.690 2.220 ;
        RECT 65.840 1.770 66.070 2.770 ;
        RECT 64.430 1.120 64.940 1.770 ;
        RECT 65.190 1.440 65.420 1.770 ;
        RECT 65.140 1.120 65.470 1.440 ;
        RECT 65.670 1.180 66.070 1.770 ;
        RECT 66.210 2.800 66.510 3.960 ;
        RECT 67.220 3.570 67.450 4.570 ;
        RECT 71.130 4.440 71.490 4.580 ;
        RECT 71.260 3.570 71.490 4.440 ;
        RECT 73.030 4.260 73.320 4.270 ;
        RECT 74.060 4.260 74.230 4.990 ;
        RECT 74.660 4.750 74.990 5.030 ;
        RECT 78.840 4.580 78.980 6.330 ;
        RECT 81.640 6.260 81.940 9.240 ;
        RECT 85.960 9.050 87.790 9.070 ;
        RECT 85.960 8.910 88.000 9.050 ;
        RECT 83.190 8.420 83.510 8.740 ;
        RECT 85.960 8.720 86.100 8.910 ;
        RECT 85.960 8.450 86.290 8.720 ;
        RECT 86.820 8.410 87.160 8.730 ;
        RECT 82.750 7.840 83.070 8.160 ;
        RECT 86.370 7.830 86.710 8.170 ;
        RECT 87.570 8.050 88.000 8.910 ;
        RECT 88.200 8.750 88.530 9.090 ;
        RECT 88.250 8.050 88.480 8.750 ;
        RECT 88.730 8.050 89.210 9.050 ;
        RECT 87.570 7.050 87.820 8.050 ;
        RECT 87.980 7.560 88.270 7.890 ;
        RECT 88.540 7.190 88.830 7.500 ;
        RECT 88.980 7.050 89.210 8.050 ;
        RECT 85.770 6.800 86.090 7.000 ;
        RECT 86.650 6.800 86.970 7.000 ;
        RECT 85.800 6.660 86.970 6.800 ;
        RECT 87.570 6.470 88.080 7.050 ;
        RECT 88.330 6.720 88.560 7.050 ;
        RECT 80.340 5.950 81.940 6.260 ;
        RECT 81.770 5.130 81.940 5.950 ;
        RECT 79.140 4.990 81.940 5.130 ;
        RECT 86.550 6.400 88.080 6.470 ;
        RECT 88.280 6.400 88.610 6.720 ;
        RECT 88.810 6.460 89.210 7.050 ;
        RECT 88.810 6.400 89.040 6.460 ;
        RECT 86.550 6.330 87.820 6.400 ;
        RECT 79.140 4.760 79.470 4.990 ;
        RECT 73.030 4.120 74.230 4.260 ;
        RECT 73.030 3.960 74.220 4.120 ;
        RECT 72.340 3.750 72.570 3.770 ;
        RECT 66.950 3.120 67.280 3.400 ;
        RECT 71.430 3.100 71.760 3.390 ;
        RECT 68.560 2.800 68.850 2.970 ;
        RECT 66.210 2.630 68.850 2.800 ;
        RECT 72.140 2.770 72.570 3.750 ;
        RECT 72.770 3.470 73.100 3.810 ;
        RECT 72.820 2.770 73.050 3.470 ;
        RECT 73.300 2.770 73.780 3.770 ;
        RECT 65.670 1.120 65.900 1.180 ;
        RECT 66.210 0.980 66.510 2.630 ;
        RECT 72.140 2.500 72.390 2.770 ;
        RECT 66.740 2.090 67.120 2.410 ;
        RECT 72.040 2.170 72.390 2.500 ;
        RECT 72.550 2.280 72.840 2.610 ;
        RECT 72.140 1.770 72.390 2.170 ;
        RECT 73.110 1.910 73.400 2.220 ;
        RECT 73.550 1.770 73.780 2.770 ;
        RECT 72.140 1.120 72.650 1.770 ;
        RECT 72.900 1.440 73.130 1.770 ;
        RECT 72.850 1.120 73.180 1.440 ;
        RECT 73.380 1.180 73.780 1.770 ;
        RECT 73.920 2.800 74.220 3.960 ;
        RECT 74.930 3.570 75.160 4.570 ;
        RECT 78.840 4.440 79.200 4.580 ;
        RECT 78.970 3.570 79.200 4.440 ;
        RECT 80.740 4.260 81.030 4.270 ;
        RECT 81.770 4.260 81.940 4.990 ;
        RECT 82.370 4.750 82.700 5.030 ;
        RECT 86.550 4.580 86.690 6.330 ;
        RECT 89.350 6.260 89.650 9.240 ;
        RECT 93.670 9.050 95.500 9.070 ;
        RECT 93.670 8.910 95.710 9.050 ;
        RECT 90.900 8.420 91.220 8.740 ;
        RECT 93.670 8.720 93.810 8.910 ;
        RECT 93.670 8.450 94.000 8.720 ;
        RECT 94.530 8.410 94.870 8.730 ;
        RECT 90.460 7.840 90.780 8.160 ;
        RECT 94.080 7.830 94.420 8.170 ;
        RECT 95.280 8.050 95.710 8.910 ;
        RECT 95.910 8.750 96.240 9.090 ;
        RECT 95.960 8.050 96.190 8.750 ;
        RECT 96.440 8.050 96.920 9.050 ;
        RECT 95.280 7.050 95.530 8.050 ;
        RECT 95.690 7.560 95.980 7.890 ;
        RECT 96.250 7.190 96.540 7.500 ;
        RECT 96.690 7.050 96.920 8.050 ;
        RECT 93.480 6.800 93.800 7.000 ;
        RECT 94.360 6.800 94.680 7.000 ;
        RECT 93.510 6.660 94.680 6.800 ;
        RECT 95.280 6.470 95.790 7.050 ;
        RECT 96.040 6.720 96.270 7.050 ;
        RECT 88.050 5.950 89.650 6.260 ;
        RECT 89.480 5.130 89.650 5.950 ;
        RECT 86.850 4.990 89.650 5.130 ;
        RECT 94.260 6.400 95.790 6.470 ;
        RECT 95.990 6.400 96.320 6.720 ;
        RECT 96.520 6.460 96.920 7.050 ;
        RECT 96.520 6.400 96.750 6.460 ;
        RECT 94.260 6.330 95.530 6.400 ;
        RECT 86.850 4.760 87.180 4.990 ;
        RECT 80.740 4.120 81.940 4.260 ;
        RECT 80.740 3.960 81.930 4.120 ;
        RECT 80.050 3.750 80.280 3.770 ;
        RECT 74.660 3.120 74.990 3.400 ;
        RECT 79.140 3.100 79.470 3.390 ;
        RECT 76.270 2.800 76.560 2.970 ;
        RECT 73.920 2.630 76.560 2.800 ;
        RECT 79.850 2.770 80.280 3.750 ;
        RECT 80.480 3.470 80.810 3.810 ;
        RECT 80.530 2.770 80.760 3.470 ;
        RECT 81.010 2.770 81.490 3.770 ;
        RECT 73.380 1.120 73.610 1.180 ;
        RECT 73.920 0.980 74.220 2.630 ;
        RECT 79.850 2.500 80.100 2.770 ;
        RECT 74.450 2.090 74.830 2.410 ;
        RECT 79.750 2.170 80.100 2.500 ;
        RECT 80.260 2.280 80.550 2.610 ;
        RECT 79.850 1.770 80.100 2.170 ;
        RECT 80.820 1.910 81.110 2.220 ;
        RECT 81.260 1.770 81.490 2.770 ;
        RECT 79.850 1.120 80.360 1.770 ;
        RECT 80.610 1.440 80.840 1.770 ;
        RECT 80.560 1.120 80.890 1.440 ;
        RECT 81.090 1.180 81.490 1.770 ;
        RECT 81.630 2.800 81.930 3.960 ;
        RECT 82.640 3.570 82.870 4.570 ;
        RECT 86.550 4.440 86.910 4.580 ;
        RECT 86.680 3.570 86.910 4.440 ;
        RECT 88.450 4.260 88.740 4.270 ;
        RECT 89.480 4.260 89.650 4.990 ;
        RECT 90.080 4.750 90.410 5.030 ;
        RECT 94.260 4.580 94.400 6.330 ;
        RECT 97.060 6.260 97.360 9.240 ;
        RECT 101.380 9.050 103.210 9.070 ;
        RECT 101.380 8.910 103.420 9.050 ;
        RECT 98.610 8.420 98.930 8.740 ;
        RECT 101.380 8.720 101.520 8.910 ;
        RECT 101.380 8.450 101.710 8.720 ;
        RECT 102.240 8.410 102.580 8.730 ;
        RECT 98.170 7.840 98.490 8.160 ;
        RECT 101.790 7.830 102.130 8.170 ;
        RECT 102.990 8.050 103.420 8.910 ;
        RECT 103.620 8.750 103.950 9.090 ;
        RECT 103.670 8.050 103.900 8.750 ;
        RECT 104.150 8.050 104.630 9.050 ;
        RECT 102.990 7.050 103.240 8.050 ;
        RECT 103.400 7.560 103.690 7.890 ;
        RECT 103.960 7.190 104.250 7.500 ;
        RECT 104.400 7.050 104.630 8.050 ;
        RECT 101.190 6.800 101.510 7.000 ;
        RECT 102.070 6.800 102.390 7.000 ;
        RECT 101.220 6.660 102.390 6.800 ;
        RECT 102.990 6.470 103.500 7.050 ;
        RECT 103.750 6.720 103.980 7.050 ;
        RECT 95.760 5.950 97.360 6.260 ;
        RECT 97.190 5.130 97.360 5.950 ;
        RECT 94.560 4.990 97.360 5.130 ;
        RECT 101.970 6.400 103.500 6.470 ;
        RECT 103.700 6.400 104.030 6.720 ;
        RECT 104.230 6.460 104.630 7.050 ;
        RECT 104.230 6.400 104.460 6.460 ;
        RECT 101.970 6.330 103.240 6.400 ;
        RECT 94.560 4.760 94.890 4.990 ;
        RECT 88.450 4.120 89.650 4.260 ;
        RECT 88.450 3.960 89.640 4.120 ;
        RECT 87.760 3.750 87.990 3.770 ;
        RECT 82.370 3.120 82.700 3.400 ;
        RECT 86.850 3.100 87.180 3.390 ;
        RECT 83.980 2.800 84.270 2.970 ;
        RECT 81.630 2.630 84.270 2.800 ;
        RECT 87.560 2.770 87.990 3.750 ;
        RECT 88.190 3.470 88.520 3.810 ;
        RECT 88.240 2.770 88.470 3.470 ;
        RECT 88.720 2.770 89.200 3.770 ;
        RECT 81.090 1.120 81.320 1.180 ;
        RECT 81.630 0.980 81.930 2.630 ;
        RECT 87.560 2.500 87.810 2.770 ;
        RECT 82.160 2.090 82.540 2.410 ;
        RECT 87.460 2.170 87.810 2.500 ;
        RECT 87.970 2.280 88.260 2.610 ;
        RECT 87.560 1.770 87.810 2.170 ;
        RECT 88.530 1.910 88.820 2.220 ;
        RECT 88.970 1.770 89.200 2.770 ;
        RECT 87.560 1.120 88.070 1.770 ;
        RECT 88.320 1.440 88.550 1.770 ;
        RECT 88.270 1.120 88.600 1.440 ;
        RECT 88.800 1.180 89.200 1.770 ;
        RECT 89.340 2.800 89.640 3.960 ;
        RECT 90.350 3.570 90.580 4.570 ;
        RECT 94.260 4.440 94.620 4.580 ;
        RECT 94.390 3.570 94.620 4.440 ;
        RECT 96.160 4.260 96.450 4.270 ;
        RECT 97.190 4.260 97.360 4.990 ;
        RECT 97.790 4.750 98.120 5.030 ;
        RECT 101.970 4.580 102.110 6.330 ;
        RECT 104.770 6.260 105.070 9.240 ;
        RECT 109.090 9.050 110.920 9.070 ;
        RECT 109.090 8.910 111.130 9.050 ;
        RECT 106.320 8.420 106.640 8.740 ;
        RECT 109.090 8.720 109.230 8.910 ;
        RECT 109.090 8.450 109.420 8.720 ;
        RECT 109.950 8.410 110.290 8.730 ;
        RECT 105.880 7.840 106.200 8.160 ;
        RECT 109.500 7.830 109.840 8.170 ;
        RECT 110.700 8.050 111.130 8.910 ;
        RECT 111.330 8.750 111.660 9.090 ;
        RECT 111.380 8.050 111.610 8.750 ;
        RECT 111.860 8.050 112.340 9.050 ;
        RECT 110.700 7.050 110.950 8.050 ;
        RECT 111.110 7.560 111.400 7.890 ;
        RECT 111.670 7.190 111.960 7.500 ;
        RECT 112.110 7.050 112.340 8.050 ;
        RECT 108.900 6.800 109.220 7.000 ;
        RECT 109.780 6.800 110.100 7.000 ;
        RECT 108.930 6.660 110.100 6.800 ;
        RECT 110.700 6.470 111.210 7.050 ;
        RECT 111.460 6.720 111.690 7.050 ;
        RECT 103.470 5.950 105.070 6.260 ;
        RECT 104.900 5.130 105.070 5.950 ;
        RECT 102.270 4.990 105.070 5.130 ;
        RECT 109.680 6.400 111.210 6.470 ;
        RECT 111.410 6.400 111.740 6.720 ;
        RECT 111.940 6.460 112.340 7.050 ;
        RECT 111.940 6.400 112.170 6.460 ;
        RECT 109.680 6.330 110.950 6.400 ;
        RECT 102.270 4.760 102.600 4.990 ;
        RECT 96.160 4.120 97.360 4.260 ;
        RECT 96.160 3.960 97.350 4.120 ;
        RECT 95.470 3.750 95.700 3.770 ;
        RECT 90.080 3.120 90.410 3.400 ;
        RECT 94.560 3.100 94.890 3.390 ;
        RECT 91.690 2.800 91.980 2.970 ;
        RECT 89.340 2.630 91.980 2.800 ;
        RECT 95.270 2.770 95.700 3.750 ;
        RECT 95.900 3.470 96.230 3.810 ;
        RECT 95.950 2.770 96.180 3.470 ;
        RECT 96.430 2.770 96.910 3.770 ;
        RECT 88.800 1.120 89.030 1.180 ;
        RECT 89.340 0.980 89.640 2.630 ;
        RECT 95.270 2.500 95.520 2.770 ;
        RECT 89.870 2.090 90.250 2.410 ;
        RECT 95.170 2.170 95.520 2.500 ;
        RECT 95.680 2.280 95.970 2.610 ;
        RECT 95.270 1.770 95.520 2.170 ;
        RECT 96.240 1.910 96.530 2.220 ;
        RECT 96.680 1.770 96.910 2.770 ;
        RECT 95.270 1.120 95.780 1.770 ;
        RECT 96.030 1.440 96.260 1.770 ;
        RECT 95.980 1.120 96.310 1.440 ;
        RECT 96.510 1.180 96.910 1.770 ;
        RECT 97.050 2.800 97.350 3.960 ;
        RECT 98.060 3.570 98.290 4.570 ;
        RECT 101.970 4.440 102.330 4.580 ;
        RECT 102.100 3.570 102.330 4.440 ;
        RECT 103.870 4.260 104.160 4.270 ;
        RECT 104.900 4.260 105.070 4.990 ;
        RECT 105.500 4.750 105.830 5.030 ;
        RECT 109.680 4.580 109.820 6.330 ;
        RECT 112.480 6.260 112.780 9.240 ;
        RECT 116.800 9.050 118.630 9.070 ;
        RECT 116.800 8.910 118.840 9.050 ;
        RECT 114.030 8.420 114.350 8.740 ;
        RECT 116.800 8.720 116.940 8.910 ;
        RECT 116.800 8.450 117.130 8.720 ;
        RECT 117.660 8.410 118.000 8.730 ;
        RECT 113.590 7.840 113.910 8.160 ;
        RECT 117.210 7.830 117.550 8.170 ;
        RECT 118.410 8.050 118.840 8.910 ;
        RECT 119.040 8.750 119.370 9.090 ;
        RECT 119.090 8.050 119.320 8.750 ;
        RECT 119.570 8.050 120.050 9.050 ;
        RECT 118.410 7.050 118.660 8.050 ;
        RECT 118.820 7.560 119.110 7.890 ;
        RECT 119.380 7.190 119.670 7.500 ;
        RECT 119.820 7.050 120.050 8.050 ;
        RECT 116.610 6.800 116.930 7.000 ;
        RECT 117.490 6.800 117.810 7.000 ;
        RECT 116.640 6.660 117.810 6.800 ;
        RECT 118.410 6.470 118.920 7.050 ;
        RECT 119.170 6.720 119.400 7.050 ;
        RECT 111.180 5.950 112.780 6.260 ;
        RECT 112.610 5.130 112.780 5.950 ;
        RECT 109.980 4.990 112.780 5.130 ;
        RECT 117.390 6.400 118.920 6.470 ;
        RECT 119.120 6.400 119.450 6.720 ;
        RECT 119.650 6.460 120.050 7.050 ;
        RECT 119.650 6.400 119.880 6.460 ;
        RECT 117.390 6.330 118.660 6.400 ;
        RECT 109.980 4.760 110.310 4.990 ;
        RECT 103.870 4.120 105.070 4.260 ;
        RECT 103.870 3.960 105.060 4.120 ;
        RECT 103.180 3.750 103.410 3.770 ;
        RECT 97.790 3.120 98.120 3.400 ;
        RECT 102.270 3.100 102.600 3.390 ;
        RECT 99.400 2.800 99.690 2.970 ;
        RECT 97.050 2.630 99.690 2.800 ;
        RECT 102.980 2.770 103.410 3.750 ;
        RECT 103.610 3.470 103.940 3.810 ;
        RECT 103.660 2.770 103.890 3.470 ;
        RECT 104.140 2.770 104.620 3.770 ;
        RECT 96.510 1.120 96.740 1.180 ;
        RECT 97.050 0.980 97.350 2.630 ;
        RECT 102.980 2.500 103.230 2.770 ;
        RECT 97.580 2.090 97.960 2.410 ;
        RECT 102.880 2.170 103.230 2.500 ;
        RECT 103.390 2.280 103.680 2.610 ;
        RECT 102.980 1.770 103.230 2.170 ;
        RECT 103.950 1.910 104.240 2.220 ;
        RECT 104.390 1.770 104.620 2.770 ;
        RECT 102.980 1.120 103.490 1.770 ;
        RECT 103.740 1.440 103.970 1.770 ;
        RECT 103.690 1.120 104.020 1.440 ;
        RECT 104.220 1.180 104.620 1.770 ;
        RECT 104.760 2.800 105.060 3.960 ;
        RECT 105.770 3.570 106.000 4.570 ;
        RECT 109.680 4.440 110.040 4.580 ;
        RECT 109.810 3.570 110.040 4.440 ;
        RECT 111.580 4.260 111.870 4.270 ;
        RECT 112.610 4.260 112.780 4.990 ;
        RECT 113.210 4.750 113.540 5.030 ;
        RECT 117.390 4.580 117.530 6.330 ;
        RECT 120.190 6.260 120.490 9.240 ;
        RECT 121.740 8.420 122.060 8.740 ;
        RECT 121.300 7.840 121.620 8.160 ;
        RECT 118.890 5.950 120.490 6.260 ;
        RECT 120.320 5.130 120.490 5.950 ;
        RECT 117.690 4.990 120.490 5.130 ;
        RECT 117.690 4.760 118.020 4.990 ;
        RECT 111.580 4.120 112.780 4.260 ;
        RECT 111.580 3.960 112.770 4.120 ;
        RECT 110.890 3.750 111.120 3.770 ;
        RECT 105.500 3.120 105.830 3.400 ;
        RECT 109.980 3.100 110.310 3.390 ;
        RECT 107.110 2.800 107.400 2.970 ;
        RECT 104.760 2.630 107.400 2.800 ;
        RECT 110.690 2.770 111.120 3.750 ;
        RECT 111.320 3.470 111.650 3.810 ;
        RECT 111.370 2.770 111.600 3.470 ;
        RECT 111.850 2.770 112.330 3.770 ;
        RECT 104.220 1.120 104.450 1.180 ;
        RECT 104.760 0.980 105.060 2.630 ;
        RECT 110.690 2.500 110.940 2.770 ;
        RECT 105.290 2.090 105.670 2.410 ;
        RECT 110.590 2.170 110.940 2.500 ;
        RECT 111.100 2.280 111.390 2.610 ;
        RECT 110.690 1.770 110.940 2.170 ;
        RECT 111.660 1.910 111.950 2.220 ;
        RECT 112.100 1.770 112.330 2.770 ;
        RECT 110.690 1.120 111.200 1.770 ;
        RECT 111.450 1.440 111.680 1.770 ;
        RECT 111.400 1.120 111.730 1.440 ;
        RECT 111.930 1.180 112.330 1.770 ;
        RECT 112.470 2.800 112.770 3.960 ;
        RECT 113.480 3.570 113.710 4.570 ;
        RECT 117.390 4.440 117.750 4.580 ;
        RECT 117.520 3.570 117.750 4.440 ;
        RECT 119.290 4.260 119.580 4.270 ;
        RECT 120.320 4.260 120.490 4.990 ;
        RECT 120.920 4.750 121.250 5.030 ;
        RECT 119.290 4.120 120.490 4.260 ;
        RECT 119.290 3.960 120.480 4.120 ;
        RECT 118.600 3.750 118.830 3.770 ;
        RECT 113.210 3.120 113.540 3.400 ;
        RECT 117.690 3.100 118.020 3.390 ;
        RECT 114.820 2.800 115.110 2.970 ;
        RECT 112.470 2.630 115.110 2.800 ;
        RECT 118.400 2.770 118.830 3.750 ;
        RECT 119.030 3.470 119.360 3.810 ;
        RECT 119.080 2.770 119.310 3.470 ;
        RECT 119.560 2.770 120.040 3.770 ;
        RECT 111.930 1.120 112.160 1.180 ;
        RECT 112.470 0.980 112.770 2.630 ;
        RECT 118.400 2.500 118.650 2.770 ;
        RECT 113.000 2.090 113.380 2.410 ;
        RECT 118.300 2.170 118.650 2.500 ;
        RECT 118.810 2.280 119.100 2.610 ;
        RECT 118.400 1.770 118.650 2.170 ;
        RECT 119.370 1.910 119.660 2.220 ;
        RECT 119.810 1.770 120.040 2.770 ;
        RECT 118.400 1.120 118.910 1.770 ;
        RECT 119.160 1.440 119.390 1.770 ;
        RECT 119.110 1.120 119.440 1.440 ;
        RECT 119.640 1.180 120.040 1.770 ;
        RECT 120.180 2.800 120.480 3.960 ;
        RECT 121.190 3.570 121.420 4.570 ;
        RECT 120.920 3.120 121.250 3.400 ;
        RECT 122.530 2.800 122.820 2.970 ;
        RECT 120.180 2.630 122.820 2.800 ;
        RECT 119.640 1.120 119.870 1.180 ;
        RECT 120.180 0.980 120.480 2.630 ;
        RECT 120.710 2.090 121.090 2.410 ;
        RECT 3.230 0.670 4.830 0.980 ;
        RECT 10.940 0.670 12.540 0.980 ;
        RECT 18.650 0.670 20.250 0.980 ;
        RECT 26.360 0.670 27.960 0.980 ;
        RECT 34.070 0.670 35.670 0.980 ;
        RECT 41.780 0.670 43.380 0.980 ;
        RECT 49.490 0.670 51.090 0.980 ;
        RECT 57.200 0.670 58.800 0.980 ;
        RECT 64.910 0.670 66.510 0.980 ;
        RECT 72.620 0.670 74.220 0.980 ;
        RECT 80.330 0.670 81.930 0.980 ;
        RECT 88.040 0.670 89.640 0.980 ;
        RECT 95.750 0.670 97.350 0.980 ;
        RECT 103.460 0.670 105.060 0.980 ;
        RECT 111.170 0.670 112.770 0.980 ;
        RECT 118.880 0.670 120.480 0.980 ;
      LAYER via ;
        RECT 2.030 31.080 2.290 31.340 ;
        RECT 3.630 32.050 3.890 32.310 ;
        RECT 4.450 30.990 4.710 31.260 ;
        RECT 9.740 31.080 10.000 31.340 ;
        RECT 3.720 29.690 3.980 29.950 ;
        RECT 11.340 32.050 11.600 32.310 ;
        RECT 12.160 30.990 12.420 31.260 ;
        RECT 17.450 31.080 17.710 31.340 ;
        RECT 11.430 29.690 11.690 29.950 ;
        RECT 1.450 25.330 1.710 25.590 ;
        RECT 1.010 24.750 1.270 25.010 ;
        RECT 19.050 32.050 19.310 32.310 ;
        RECT 19.870 30.990 20.130 31.260 ;
        RECT 25.160 31.080 25.420 31.340 ;
        RECT 19.140 29.690 19.400 29.950 ;
        RECT 3.620 26.770 3.880 27.030 ;
        RECT 5.260 26.490 5.520 26.760 ;
        RECT 6.140 26.490 6.400 26.760 ;
        RECT 3.710 24.410 3.970 24.670 ;
        RECT 5.530 25.320 5.790 25.580 ;
        RECT 9.160 25.330 9.420 25.590 ;
        RECT 5.070 24.760 5.330 25.020 ;
        RECT 8.720 24.750 8.980 25.010 ;
        RECT 26.760 32.050 27.020 32.310 ;
        RECT 27.580 30.990 27.840 31.260 ;
        RECT 32.870 31.080 33.130 31.340 ;
        RECT 26.850 29.690 27.110 29.950 ;
        RECT 11.330 26.770 11.590 27.030 ;
        RECT 12.970 26.490 13.230 26.760 ;
        RECT 13.850 26.490 14.110 26.760 ;
        RECT 11.420 24.410 11.680 24.670 ;
        RECT 13.240 25.320 13.500 25.580 ;
        RECT 16.870 25.330 17.130 25.590 ;
        RECT 12.780 24.760 13.040 25.020 ;
        RECT 16.430 24.750 16.690 25.010 ;
        RECT 34.470 32.050 34.730 32.310 ;
        RECT 35.290 30.990 35.550 31.260 ;
        RECT 40.580 31.080 40.840 31.340 ;
        RECT 34.560 29.690 34.820 29.950 ;
        RECT 19.040 26.770 19.300 27.030 ;
        RECT 20.680 26.490 20.940 26.760 ;
        RECT 21.560 26.490 21.820 26.760 ;
        RECT 19.130 24.410 19.390 24.670 ;
        RECT 20.950 25.320 21.210 25.580 ;
        RECT 24.580 25.330 24.840 25.590 ;
        RECT 20.490 24.760 20.750 25.020 ;
        RECT 24.140 24.750 24.400 25.010 ;
        RECT 42.180 32.050 42.440 32.310 ;
        RECT 43.000 30.990 43.260 31.260 ;
        RECT 48.290 31.080 48.550 31.340 ;
        RECT 42.270 29.690 42.530 29.950 ;
        RECT 26.750 26.770 27.010 27.030 ;
        RECT 28.390 26.490 28.650 26.760 ;
        RECT 29.270 26.490 29.530 26.760 ;
        RECT 26.840 24.410 27.100 24.670 ;
        RECT 28.660 25.320 28.920 25.580 ;
        RECT 32.290 25.330 32.550 25.590 ;
        RECT 28.200 24.760 28.460 25.020 ;
        RECT 31.850 24.750 32.110 25.010 ;
        RECT 49.890 32.050 50.150 32.310 ;
        RECT 50.710 30.990 50.970 31.260 ;
        RECT 56.000 31.080 56.260 31.340 ;
        RECT 49.980 29.690 50.240 29.950 ;
        RECT 34.460 26.770 34.720 27.030 ;
        RECT 36.100 26.490 36.360 26.760 ;
        RECT 36.980 26.490 37.240 26.760 ;
        RECT 34.550 24.410 34.810 24.670 ;
        RECT 36.370 25.320 36.630 25.580 ;
        RECT 40.000 25.330 40.260 25.590 ;
        RECT 35.910 24.760 36.170 25.020 ;
        RECT 39.560 24.750 39.820 25.010 ;
        RECT 57.600 32.050 57.860 32.310 ;
        RECT 58.420 30.990 58.680 31.260 ;
        RECT 63.710 31.080 63.970 31.340 ;
        RECT 57.690 29.690 57.950 29.950 ;
        RECT 42.170 26.770 42.430 27.030 ;
        RECT 43.810 26.490 44.070 26.760 ;
        RECT 44.690 26.490 44.950 26.760 ;
        RECT 42.260 24.410 42.520 24.670 ;
        RECT 44.080 25.320 44.340 25.580 ;
        RECT 47.710 25.330 47.970 25.590 ;
        RECT 43.620 24.760 43.880 25.020 ;
        RECT 47.270 24.750 47.530 25.010 ;
        RECT 65.310 32.050 65.570 32.310 ;
        RECT 66.130 30.990 66.390 31.260 ;
        RECT 71.420 31.080 71.680 31.340 ;
        RECT 65.400 29.690 65.660 29.950 ;
        RECT 49.880 26.770 50.140 27.030 ;
        RECT 51.520 26.490 51.780 26.760 ;
        RECT 52.400 26.490 52.660 26.760 ;
        RECT 49.970 24.410 50.230 24.670 ;
        RECT 51.790 25.320 52.050 25.580 ;
        RECT 55.420 25.330 55.680 25.590 ;
        RECT 51.330 24.760 51.590 25.020 ;
        RECT 54.980 24.750 55.240 25.010 ;
        RECT 73.020 32.050 73.280 32.310 ;
        RECT 73.840 30.990 74.100 31.260 ;
        RECT 79.130 31.080 79.390 31.340 ;
        RECT 73.110 29.690 73.370 29.950 ;
        RECT 57.590 26.770 57.850 27.030 ;
        RECT 59.230 26.490 59.490 26.760 ;
        RECT 60.110 26.490 60.370 26.760 ;
        RECT 57.680 24.410 57.940 24.670 ;
        RECT 59.500 25.320 59.760 25.580 ;
        RECT 63.130 25.330 63.390 25.590 ;
        RECT 59.040 24.760 59.300 25.020 ;
        RECT 62.690 24.750 62.950 25.010 ;
        RECT 80.730 32.050 80.990 32.310 ;
        RECT 81.550 30.990 81.810 31.260 ;
        RECT 86.840 31.080 87.100 31.340 ;
        RECT 80.820 29.690 81.080 29.950 ;
        RECT 65.300 26.770 65.560 27.030 ;
        RECT 66.940 26.490 67.200 26.760 ;
        RECT 67.820 26.490 68.080 26.760 ;
        RECT 65.390 24.410 65.650 24.670 ;
        RECT 67.210 25.320 67.470 25.580 ;
        RECT 70.840 25.330 71.100 25.590 ;
        RECT 66.750 24.760 67.010 25.020 ;
        RECT 70.400 24.750 70.660 25.010 ;
        RECT 88.440 32.050 88.700 32.310 ;
        RECT 89.260 30.990 89.520 31.260 ;
        RECT 94.550 31.080 94.810 31.340 ;
        RECT 88.530 29.690 88.790 29.950 ;
        RECT 73.010 26.770 73.270 27.030 ;
        RECT 74.650 26.490 74.910 26.760 ;
        RECT 75.530 26.490 75.790 26.760 ;
        RECT 73.100 24.410 73.360 24.670 ;
        RECT 74.920 25.320 75.180 25.580 ;
        RECT 78.550 25.330 78.810 25.590 ;
        RECT 74.460 24.760 74.720 25.020 ;
        RECT 78.110 24.750 78.370 25.010 ;
        RECT 96.150 32.050 96.410 32.310 ;
        RECT 96.970 30.990 97.230 31.260 ;
        RECT 102.260 31.080 102.520 31.340 ;
        RECT 96.240 29.690 96.500 29.950 ;
        RECT 80.720 26.770 80.980 27.030 ;
        RECT 82.360 26.490 82.620 26.760 ;
        RECT 83.240 26.490 83.500 26.760 ;
        RECT 80.810 24.410 81.070 24.670 ;
        RECT 82.630 25.320 82.890 25.580 ;
        RECT 86.260 25.330 86.520 25.590 ;
        RECT 82.170 24.760 82.430 25.020 ;
        RECT 85.820 24.750 86.080 25.010 ;
        RECT 103.860 32.050 104.120 32.310 ;
        RECT 104.680 30.990 104.940 31.260 ;
        RECT 109.970 31.080 110.230 31.340 ;
        RECT 103.950 29.690 104.210 29.950 ;
        RECT 88.430 26.770 88.690 27.030 ;
        RECT 90.070 26.490 90.330 26.760 ;
        RECT 90.950 26.490 91.210 26.760 ;
        RECT 88.520 24.410 88.780 24.670 ;
        RECT 90.340 25.320 90.600 25.580 ;
        RECT 93.970 25.330 94.230 25.590 ;
        RECT 89.880 24.760 90.140 25.020 ;
        RECT 93.530 24.750 93.790 25.010 ;
        RECT 111.570 32.050 111.830 32.310 ;
        RECT 112.390 30.990 112.650 31.260 ;
        RECT 117.680 31.080 117.940 31.340 ;
        RECT 111.660 29.690 111.920 29.950 ;
        RECT 96.140 26.770 96.400 27.030 ;
        RECT 97.780 26.490 98.040 26.760 ;
        RECT 98.660 26.490 98.920 26.760 ;
        RECT 96.230 24.410 96.490 24.670 ;
        RECT 98.050 25.320 98.310 25.580 ;
        RECT 101.680 25.330 101.940 25.590 ;
        RECT 97.590 24.760 97.850 25.020 ;
        RECT 101.240 24.750 101.500 25.010 ;
        RECT 119.280 32.050 119.540 32.310 ;
        RECT 120.100 30.990 120.360 31.260 ;
        RECT 119.370 29.690 119.630 29.950 ;
        RECT 103.850 26.770 104.110 27.030 ;
        RECT 105.490 26.490 105.750 26.760 ;
        RECT 106.370 26.490 106.630 26.760 ;
        RECT 103.940 24.410 104.200 24.670 ;
        RECT 105.760 25.320 106.020 25.580 ;
        RECT 109.390 25.330 109.650 25.590 ;
        RECT 105.300 24.760 105.560 25.020 ;
        RECT 108.950 24.750 109.210 25.010 ;
        RECT 111.560 26.770 111.820 27.030 ;
        RECT 113.200 26.490 113.460 26.760 ;
        RECT 114.080 26.490 114.340 26.760 ;
        RECT 111.650 24.410 111.910 24.670 ;
        RECT 113.470 25.320 113.730 25.580 ;
        RECT 117.100 25.330 117.360 25.590 ;
        RECT 113.010 24.760 113.270 25.020 ;
        RECT 116.660 24.750 116.920 25.010 ;
        RECT 119.270 26.770 119.530 27.030 ;
        RECT 120.910 26.490 121.170 26.760 ;
        RECT 121.790 26.490 122.050 26.760 ;
        RECT 119.360 24.410 119.620 24.670 ;
        RECT 121.180 25.320 121.440 25.580 ;
        RECT 120.720 24.760 120.980 25.020 ;
        RECT 28.700 20.600 28.970 20.860 ;
        RECT 90.360 20.610 90.630 20.870 ;
        RECT 58.530 19.880 58.790 20.140 ;
        RECT 58.550 15.830 58.810 16.090 ;
        RECT 124.550 15.860 124.830 16.120 ;
        RECT 58.440 13.640 58.710 13.900 ;
        RECT 28.820 11.920 29.090 12.220 ;
        RECT 90.480 11.960 90.770 12.220 ;
        RECT 2.060 8.440 2.320 8.700 ;
        RECT 1.600 7.880 1.860 8.140 ;
        RECT 3.420 8.790 3.680 9.050 ;
        RECT 0.990 6.700 1.250 6.970 ;
        RECT 1.870 6.700 2.130 6.970 ;
        RECT 3.510 6.430 3.770 6.690 ;
        RECT 6.120 8.450 6.380 8.710 ;
        RECT 9.770 8.440 10.030 8.700 ;
        RECT 5.680 7.870 5.940 8.130 ;
        RECT 9.310 7.880 9.570 8.140 ;
        RECT 11.130 8.790 11.390 9.050 ;
        RECT 8.700 6.700 8.960 6.970 ;
        RECT 9.580 6.700 9.840 6.970 ;
        RECT 11.220 6.430 11.480 6.690 ;
        RECT 13.830 8.450 14.090 8.710 ;
        RECT 17.480 8.440 17.740 8.700 ;
        RECT 13.390 7.870 13.650 8.130 ;
        RECT 17.020 7.880 17.280 8.140 ;
        RECT 18.840 8.790 19.100 9.050 ;
        RECT 16.410 6.700 16.670 6.970 ;
        RECT 17.290 6.700 17.550 6.970 ;
        RECT 18.930 6.430 19.190 6.690 ;
        RECT 3.410 3.510 3.670 3.770 ;
        RECT 2.680 2.200 2.940 2.470 ;
        RECT 3.500 1.150 3.760 1.410 ;
        RECT 21.540 8.450 21.800 8.710 ;
        RECT 25.190 8.440 25.450 8.700 ;
        RECT 21.100 7.870 21.360 8.130 ;
        RECT 24.730 7.880 24.990 8.140 ;
        RECT 26.550 8.790 26.810 9.050 ;
        RECT 24.120 6.700 24.380 6.970 ;
        RECT 25.000 6.700 25.260 6.970 ;
        RECT 26.640 6.430 26.900 6.690 ;
        RECT 11.120 3.510 11.380 3.770 ;
        RECT 5.100 2.120 5.360 2.380 ;
        RECT 10.390 2.200 10.650 2.470 ;
        RECT 11.210 1.150 11.470 1.410 ;
        RECT 29.250 8.450 29.510 8.710 ;
        RECT 32.900 8.440 33.160 8.700 ;
        RECT 28.810 7.870 29.070 8.130 ;
        RECT 32.440 7.880 32.700 8.140 ;
        RECT 34.260 8.790 34.520 9.050 ;
        RECT 31.830 6.700 32.090 6.970 ;
        RECT 32.710 6.700 32.970 6.970 ;
        RECT 34.350 6.430 34.610 6.690 ;
        RECT 18.830 3.510 19.090 3.770 ;
        RECT 12.810 2.120 13.070 2.380 ;
        RECT 18.100 2.200 18.360 2.470 ;
        RECT 18.920 1.150 19.180 1.410 ;
        RECT 36.960 8.450 37.220 8.710 ;
        RECT 40.610 8.440 40.870 8.700 ;
        RECT 36.520 7.870 36.780 8.130 ;
        RECT 40.150 7.880 40.410 8.140 ;
        RECT 41.970 8.790 42.230 9.050 ;
        RECT 39.540 6.700 39.800 6.970 ;
        RECT 40.420 6.700 40.680 6.970 ;
        RECT 42.060 6.430 42.320 6.690 ;
        RECT 26.540 3.510 26.800 3.770 ;
        RECT 20.520 2.120 20.780 2.380 ;
        RECT 25.810 2.200 26.070 2.470 ;
        RECT 26.630 1.150 26.890 1.410 ;
        RECT 44.670 8.450 44.930 8.710 ;
        RECT 48.320 8.440 48.580 8.700 ;
        RECT 44.230 7.870 44.490 8.130 ;
        RECT 47.860 7.880 48.120 8.140 ;
        RECT 49.680 8.790 49.940 9.050 ;
        RECT 47.250 6.700 47.510 6.970 ;
        RECT 48.130 6.700 48.390 6.970 ;
        RECT 49.770 6.430 50.030 6.690 ;
        RECT 34.250 3.510 34.510 3.770 ;
        RECT 28.230 2.120 28.490 2.380 ;
        RECT 33.520 2.200 33.780 2.470 ;
        RECT 34.340 1.150 34.600 1.410 ;
        RECT 52.380 8.450 52.640 8.710 ;
        RECT 56.030 8.440 56.290 8.700 ;
        RECT 51.940 7.870 52.200 8.130 ;
        RECT 55.570 7.880 55.830 8.140 ;
        RECT 57.390 8.790 57.650 9.050 ;
        RECT 54.960 6.700 55.220 6.970 ;
        RECT 55.840 6.700 56.100 6.970 ;
        RECT 57.480 6.430 57.740 6.690 ;
        RECT 41.960 3.510 42.220 3.770 ;
        RECT 35.940 2.120 36.200 2.380 ;
        RECT 41.230 2.200 41.490 2.470 ;
        RECT 42.050 1.150 42.310 1.410 ;
        RECT 60.090 8.450 60.350 8.710 ;
        RECT 63.740 8.440 64.000 8.700 ;
        RECT 59.650 7.870 59.910 8.130 ;
        RECT 63.280 7.880 63.540 8.140 ;
        RECT 65.100 8.790 65.360 9.050 ;
        RECT 62.670 6.700 62.930 6.970 ;
        RECT 63.550 6.700 63.810 6.970 ;
        RECT 65.190 6.430 65.450 6.690 ;
        RECT 49.670 3.510 49.930 3.770 ;
        RECT 43.650 2.120 43.910 2.380 ;
        RECT 48.940 2.200 49.200 2.470 ;
        RECT 49.760 1.150 50.020 1.410 ;
        RECT 67.800 8.450 68.060 8.710 ;
        RECT 71.450 8.440 71.710 8.700 ;
        RECT 67.360 7.870 67.620 8.130 ;
        RECT 70.990 7.880 71.250 8.140 ;
        RECT 72.810 8.790 73.070 9.050 ;
        RECT 70.380 6.700 70.640 6.970 ;
        RECT 71.260 6.700 71.520 6.970 ;
        RECT 72.900 6.430 73.160 6.690 ;
        RECT 57.380 3.510 57.640 3.770 ;
        RECT 51.360 2.120 51.620 2.380 ;
        RECT 56.650 2.200 56.910 2.470 ;
        RECT 57.470 1.150 57.730 1.410 ;
        RECT 75.510 8.450 75.770 8.710 ;
        RECT 79.160 8.440 79.420 8.700 ;
        RECT 75.070 7.870 75.330 8.130 ;
        RECT 78.700 7.880 78.960 8.140 ;
        RECT 80.520 8.790 80.780 9.050 ;
        RECT 78.090 6.700 78.350 6.970 ;
        RECT 78.970 6.700 79.230 6.970 ;
        RECT 80.610 6.430 80.870 6.690 ;
        RECT 65.090 3.510 65.350 3.770 ;
        RECT 59.070 2.120 59.330 2.380 ;
        RECT 64.360 2.200 64.620 2.470 ;
        RECT 65.180 1.150 65.440 1.410 ;
        RECT 83.220 8.450 83.480 8.710 ;
        RECT 86.870 8.440 87.130 8.700 ;
        RECT 82.780 7.870 83.040 8.130 ;
        RECT 86.410 7.880 86.670 8.140 ;
        RECT 88.230 8.790 88.490 9.050 ;
        RECT 85.800 6.700 86.060 6.970 ;
        RECT 86.680 6.700 86.940 6.970 ;
        RECT 88.320 6.430 88.580 6.690 ;
        RECT 72.800 3.510 73.060 3.770 ;
        RECT 66.780 2.120 67.040 2.380 ;
        RECT 72.070 2.200 72.330 2.470 ;
        RECT 72.890 1.150 73.150 1.410 ;
        RECT 90.930 8.450 91.190 8.710 ;
        RECT 94.580 8.440 94.840 8.700 ;
        RECT 90.490 7.870 90.750 8.130 ;
        RECT 94.120 7.880 94.380 8.140 ;
        RECT 95.940 8.790 96.200 9.050 ;
        RECT 93.510 6.700 93.770 6.970 ;
        RECT 94.390 6.700 94.650 6.970 ;
        RECT 96.030 6.430 96.290 6.690 ;
        RECT 80.510 3.510 80.770 3.770 ;
        RECT 74.490 2.120 74.750 2.380 ;
        RECT 79.780 2.200 80.040 2.470 ;
        RECT 80.600 1.150 80.860 1.410 ;
        RECT 98.640 8.450 98.900 8.710 ;
        RECT 102.290 8.440 102.550 8.700 ;
        RECT 98.200 7.870 98.460 8.130 ;
        RECT 101.830 7.880 102.090 8.140 ;
        RECT 103.650 8.790 103.910 9.050 ;
        RECT 101.220 6.700 101.480 6.970 ;
        RECT 102.100 6.700 102.360 6.970 ;
        RECT 103.740 6.430 104.000 6.690 ;
        RECT 88.220 3.510 88.480 3.770 ;
        RECT 82.200 2.120 82.460 2.380 ;
        RECT 87.490 2.200 87.750 2.470 ;
        RECT 88.310 1.150 88.570 1.410 ;
        RECT 106.350 8.450 106.610 8.710 ;
        RECT 110.000 8.440 110.260 8.700 ;
        RECT 105.910 7.870 106.170 8.130 ;
        RECT 109.540 7.880 109.800 8.140 ;
        RECT 111.360 8.790 111.620 9.050 ;
        RECT 108.930 6.700 109.190 6.970 ;
        RECT 109.810 6.700 110.070 6.970 ;
        RECT 111.450 6.430 111.710 6.690 ;
        RECT 95.930 3.510 96.190 3.770 ;
        RECT 89.910 2.120 90.170 2.380 ;
        RECT 95.200 2.200 95.460 2.470 ;
        RECT 96.020 1.150 96.280 1.410 ;
        RECT 114.060 8.450 114.320 8.710 ;
        RECT 117.710 8.440 117.970 8.700 ;
        RECT 113.620 7.870 113.880 8.130 ;
        RECT 117.250 7.880 117.510 8.140 ;
        RECT 119.070 8.790 119.330 9.050 ;
        RECT 116.640 6.700 116.900 6.970 ;
        RECT 117.520 6.700 117.780 6.970 ;
        RECT 119.160 6.430 119.420 6.690 ;
        RECT 103.640 3.510 103.900 3.770 ;
        RECT 97.620 2.120 97.880 2.380 ;
        RECT 102.910 2.200 103.170 2.470 ;
        RECT 103.730 1.150 103.990 1.410 ;
        RECT 121.770 8.450 122.030 8.710 ;
        RECT 121.330 7.870 121.590 8.130 ;
        RECT 111.350 3.510 111.610 3.770 ;
        RECT 105.330 2.120 105.590 2.380 ;
        RECT 110.620 2.200 110.880 2.470 ;
        RECT 111.440 1.150 111.700 1.410 ;
        RECT 119.060 3.510 119.320 3.770 ;
        RECT 113.040 2.120 113.300 2.380 ;
        RECT 118.330 2.200 118.590 2.470 ;
        RECT 119.150 1.150 119.410 1.410 ;
        RECT 120.750 2.120 121.010 2.380 ;
      LAYER met2 ;
        RECT 3.600 32.300 3.930 32.340 ;
        RECT 11.310 32.300 11.640 32.340 ;
        RECT 19.020 32.300 19.350 32.340 ;
        RECT 26.730 32.300 27.060 32.340 ;
        RECT 34.440 32.300 34.770 32.340 ;
        RECT 42.150 32.300 42.480 32.340 ;
        RECT 49.860 32.300 50.190 32.340 ;
        RECT 57.570 32.300 57.900 32.340 ;
        RECT 65.280 32.300 65.610 32.340 ;
        RECT 72.990 32.300 73.320 32.340 ;
        RECT 80.700 32.300 81.030 32.340 ;
        RECT 88.410 32.300 88.740 32.340 ;
        RECT 96.120 32.300 96.450 32.340 ;
        RECT 103.830 32.300 104.160 32.340 ;
        RECT 111.540 32.300 111.870 32.340 ;
        RECT 119.250 32.300 119.580 32.340 ;
        RECT 0.490 32.160 3.930 32.300 ;
        RECT 0.490 26.830 0.630 32.160 ;
        RECT 3.600 32.020 3.930 32.160 ;
        RECT 1.950 31.350 2.330 31.370 ;
        RECT 1.950 31.210 2.790 31.350 ;
        RECT 1.950 31.050 2.330 31.210 ;
        RECT -0.740 26.650 0.630 26.830 ;
        RECT -0.740 22.470 -0.560 26.650 ;
        RECT 2.650 25.620 2.790 31.210 ;
        RECT 3.680 29.990 3.930 32.020 ;
        RECT 8.200 32.160 11.640 32.300 ;
        RECT 4.390 30.960 4.740 31.290 ;
        RECT 3.680 29.650 4.010 29.990 ;
        RECT 4.390 28.630 4.530 30.960 ;
        RECT 4.390 28.490 5.830 28.630 ;
        RECT 3.590 26.800 3.920 27.060 ;
        RECT 3.590 26.740 5.550 26.800 ;
        RECT 3.660 26.660 5.550 26.740 ;
        RECT 1.420 25.480 2.790 25.620 ;
        RECT 1.420 25.300 1.740 25.480 ;
        RECT 0.980 24.820 1.300 25.040 ;
        RECT 0.980 24.720 1.310 24.820 ;
        RECT 1.170 24.200 1.310 24.720 ;
        RECT 3.670 24.710 3.920 26.660 ;
        RECT 5.230 26.460 5.550 26.660 ;
        RECT 5.690 25.630 5.830 28.490 ;
        RECT 8.200 26.830 8.340 32.160 ;
        RECT 11.310 32.020 11.640 32.160 ;
        RECT 9.660 31.350 10.040 31.370 ;
        RECT 9.660 31.210 10.500 31.350 ;
        RECT 9.660 31.050 10.040 31.210 ;
        RECT 6.430 26.800 8.340 26.830 ;
        RECT 6.400 26.790 8.340 26.800 ;
        RECT 6.110 26.650 8.340 26.790 ;
        RECT 6.110 26.460 6.430 26.650 ;
        RECT 5.490 25.290 5.830 25.630 ;
        RECT 10.360 25.620 10.500 31.210 ;
        RECT 11.390 29.990 11.640 32.020 ;
        RECT 15.910 32.160 19.350 32.300 ;
        RECT 12.100 30.960 12.450 31.290 ;
        RECT 11.390 29.650 11.720 29.990 ;
        RECT 12.100 28.630 12.240 30.960 ;
        RECT 12.100 28.490 13.540 28.630 ;
        RECT 11.300 26.800 11.630 27.060 ;
        RECT 11.300 26.740 13.260 26.800 ;
        RECT 11.370 26.660 13.260 26.740 ;
        RECT 9.130 25.480 10.500 25.620 ;
        RECT 9.130 25.300 9.450 25.480 ;
        RECT 5.040 24.730 5.380 25.050 ;
        RECT 8.690 24.820 9.010 25.040 ;
        RECT 3.670 24.370 4.000 24.710 ;
        RECT 5.040 24.200 5.180 24.730 ;
        RECT 8.690 24.720 9.020 24.820 ;
        RECT 8.880 24.200 9.020 24.720 ;
        RECT 11.380 24.710 11.630 26.660 ;
        RECT 12.940 26.460 13.260 26.660 ;
        RECT 13.400 25.630 13.540 28.490 ;
        RECT 15.910 26.830 16.050 32.160 ;
        RECT 19.020 32.020 19.350 32.160 ;
        RECT 17.370 31.350 17.750 31.370 ;
        RECT 17.370 31.210 18.210 31.350 ;
        RECT 17.370 31.050 17.750 31.210 ;
        RECT 14.140 26.800 16.050 26.830 ;
        RECT 14.110 26.790 16.050 26.800 ;
        RECT 13.820 26.650 16.050 26.790 ;
        RECT 13.820 26.460 14.140 26.650 ;
        RECT 13.200 25.290 13.540 25.630 ;
        RECT 18.070 25.620 18.210 31.210 ;
        RECT 19.100 29.990 19.350 32.020 ;
        RECT 23.620 32.160 27.060 32.300 ;
        RECT 19.810 30.960 20.160 31.290 ;
        RECT 19.100 29.650 19.430 29.990 ;
        RECT 19.810 28.630 19.950 30.960 ;
        RECT 19.810 28.490 21.250 28.630 ;
        RECT 19.010 26.800 19.340 27.060 ;
        RECT 19.010 26.740 20.970 26.800 ;
        RECT 19.080 26.660 20.970 26.740 ;
        RECT 16.840 25.480 18.210 25.620 ;
        RECT 16.840 25.300 17.160 25.480 ;
        RECT 12.750 24.730 13.090 25.050 ;
        RECT 16.400 24.820 16.720 25.040 ;
        RECT 11.380 24.370 11.710 24.710 ;
        RECT 12.750 24.200 12.890 24.730 ;
        RECT 16.400 24.720 16.730 24.820 ;
        RECT 16.590 24.200 16.730 24.720 ;
        RECT 19.090 24.710 19.340 26.660 ;
        RECT 20.650 26.460 20.970 26.660 ;
        RECT 21.110 25.630 21.250 28.490 ;
        RECT 23.620 26.830 23.760 32.160 ;
        RECT 26.730 32.020 27.060 32.160 ;
        RECT 25.080 31.350 25.460 31.370 ;
        RECT 25.080 31.210 25.920 31.350 ;
        RECT 25.080 31.050 25.460 31.210 ;
        RECT 21.850 26.800 23.760 26.830 ;
        RECT 21.820 26.790 23.760 26.800 ;
        RECT 21.530 26.650 23.760 26.790 ;
        RECT 21.530 26.460 21.850 26.650 ;
        RECT 20.910 25.290 21.250 25.630 ;
        RECT 25.780 25.620 25.920 31.210 ;
        RECT 26.810 29.990 27.060 32.020 ;
        RECT 31.330 32.160 34.770 32.300 ;
        RECT 27.520 30.960 27.870 31.290 ;
        RECT 26.810 29.650 27.140 29.990 ;
        RECT 27.520 28.630 27.660 30.960 ;
        RECT 27.520 28.490 28.960 28.630 ;
        RECT 26.720 26.800 27.050 27.060 ;
        RECT 26.720 26.740 28.680 26.800 ;
        RECT 26.790 26.660 28.680 26.740 ;
        RECT 24.550 25.480 25.920 25.620 ;
        RECT 24.550 25.300 24.870 25.480 ;
        RECT 20.460 24.730 20.800 25.050 ;
        RECT 24.110 24.820 24.430 25.040 ;
        RECT 19.090 24.370 19.420 24.710 ;
        RECT 20.460 24.200 20.600 24.730 ;
        RECT 24.110 24.720 24.440 24.820 ;
        RECT 24.300 24.200 24.440 24.720 ;
        RECT 26.800 24.710 27.050 26.660 ;
        RECT 28.360 26.460 28.680 26.660 ;
        RECT 28.820 25.630 28.960 28.490 ;
        RECT 31.330 26.830 31.470 32.160 ;
        RECT 34.440 32.020 34.770 32.160 ;
        RECT 32.790 31.350 33.170 31.370 ;
        RECT 32.790 31.210 33.630 31.350 ;
        RECT 32.790 31.050 33.170 31.210 ;
        RECT 29.560 26.800 31.470 26.830 ;
        RECT 29.530 26.790 31.470 26.800 ;
        RECT 29.240 26.650 31.470 26.790 ;
        RECT 29.240 26.460 29.560 26.650 ;
        RECT 28.620 25.290 28.960 25.630 ;
        RECT 33.490 25.620 33.630 31.210 ;
        RECT 34.520 29.990 34.770 32.020 ;
        RECT 39.040 32.160 42.480 32.300 ;
        RECT 35.230 30.960 35.580 31.290 ;
        RECT 34.520 29.650 34.850 29.990 ;
        RECT 35.230 28.630 35.370 30.960 ;
        RECT 35.230 28.490 36.670 28.630 ;
        RECT 34.430 26.800 34.760 27.060 ;
        RECT 34.430 26.740 36.390 26.800 ;
        RECT 34.500 26.660 36.390 26.740 ;
        RECT 32.260 25.480 33.630 25.620 ;
        RECT 32.260 25.300 32.580 25.480 ;
        RECT 28.170 24.730 28.510 25.050 ;
        RECT 31.820 24.820 32.140 25.040 ;
        RECT 26.800 24.370 27.130 24.710 ;
        RECT 28.170 24.200 28.310 24.730 ;
        RECT 31.820 24.720 32.150 24.820 ;
        RECT 32.010 24.200 32.150 24.720 ;
        RECT 34.510 24.710 34.760 26.660 ;
        RECT 36.070 26.460 36.390 26.660 ;
        RECT 36.530 25.630 36.670 28.490 ;
        RECT 39.040 26.830 39.180 32.160 ;
        RECT 42.150 32.020 42.480 32.160 ;
        RECT 40.500 31.350 40.880 31.370 ;
        RECT 40.500 31.210 41.340 31.350 ;
        RECT 40.500 31.050 40.880 31.210 ;
        RECT 37.270 26.800 39.180 26.830 ;
        RECT 37.240 26.790 39.180 26.800 ;
        RECT 36.950 26.650 39.180 26.790 ;
        RECT 36.950 26.460 37.270 26.650 ;
        RECT 36.330 25.290 36.670 25.630 ;
        RECT 41.200 25.620 41.340 31.210 ;
        RECT 42.230 29.990 42.480 32.020 ;
        RECT 46.750 32.160 50.190 32.300 ;
        RECT 42.940 30.960 43.290 31.290 ;
        RECT 42.230 29.650 42.560 29.990 ;
        RECT 42.940 28.630 43.080 30.960 ;
        RECT 42.940 28.490 44.380 28.630 ;
        RECT 42.140 26.800 42.470 27.060 ;
        RECT 42.140 26.740 44.100 26.800 ;
        RECT 42.210 26.660 44.100 26.740 ;
        RECT 39.970 25.480 41.340 25.620 ;
        RECT 39.970 25.300 40.290 25.480 ;
        RECT 35.880 24.730 36.220 25.050 ;
        RECT 39.530 24.820 39.850 25.040 ;
        RECT 34.510 24.370 34.840 24.710 ;
        RECT 35.880 24.200 36.020 24.730 ;
        RECT 39.530 24.720 39.860 24.820 ;
        RECT 39.720 24.200 39.860 24.720 ;
        RECT 42.220 24.710 42.470 26.660 ;
        RECT 43.780 26.460 44.100 26.660 ;
        RECT 44.240 25.630 44.380 28.490 ;
        RECT 46.750 26.830 46.890 32.160 ;
        RECT 49.860 32.020 50.190 32.160 ;
        RECT 48.210 31.350 48.590 31.370 ;
        RECT 48.210 31.210 49.050 31.350 ;
        RECT 48.210 31.050 48.590 31.210 ;
        RECT 44.980 26.800 46.890 26.830 ;
        RECT 44.950 26.790 46.890 26.800 ;
        RECT 44.660 26.650 46.890 26.790 ;
        RECT 44.660 26.460 44.980 26.650 ;
        RECT 44.040 25.290 44.380 25.630 ;
        RECT 48.910 25.620 49.050 31.210 ;
        RECT 49.940 29.990 50.190 32.020 ;
        RECT 54.460 32.160 57.900 32.300 ;
        RECT 50.650 30.960 51.000 31.290 ;
        RECT 49.940 29.650 50.270 29.990 ;
        RECT 50.650 28.630 50.790 30.960 ;
        RECT 50.650 28.490 52.090 28.630 ;
        RECT 49.850 26.800 50.180 27.060 ;
        RECT 49.850 26.740 51.810 26.800 ;
        RECT 49.920 26.660 51.810 26.740 ;
        RECT 47.680 25.480 49.050 25.620 ;
        RECT 47.680 25.300 48.000 25.480 ;
        RECT 43.590 24.730 43.930 25.050 ;
        RECT 47.240 24.820 47.560 25.040 ;
        RECT 42.220 24.370 42.550 24.710 ;
        RECT 43.590 24.200 43.730 24.730 ;
        RECT 47.240 24.720 47.570 24.820 ;
        RECT 47.430 24.200 47.570 24.720 ;
        RECT 49.930 24.710 50.180 26.660 ;
        RECT 51.490 26.460 51.810 26.660 ;
        RECT 51.950 25.630 52.090 28.490 ;
        RECT 54.460 26.830 54.600 32.160 ;
        RECT 57.570 32.020 57.900 32.160 ;
        RECT 55.920 31.350 56.300 31.370 ;
        RECT 55.920 31.210 56.760 31.350 ;
        RECT 55.920 31.050 56.300 31.210 ;
        RECT 52.690 26.800 54.600 26.830 ;
        RECT 52.660 26.790 54.600 26.800 ;
        RECT 52.370 26.650 54.600 26.790 ;
        RECT 52.370 26.460 52.690 26.650 ;
        RECT 51.750 25.290 52.090 25.630 ;
        RECT 56.620 25.620 56.760 31.210 ;
        RECT 57.650 29.990 57.900 32.020 ;
        RECT 62.170 32.160 65.610 32.300 ;
        RECT 58.360 30.960 58.710 31.290 ;
        RECT 57.650 29.650 57.980 29.990 ;
        RECT 58.360 28.630 58.500 30.960 ;
        RECT 58.360 28.490 59.800 28.630 ;
        RECT 57.560 26.800 57.890 27.060 ;
        RECT 57.560 26.740 59.520 26.800 ;
        RECT 57.630 26.660 59.520 26.740 ;
        RECT 55.390 25.480 56.760 25.620 ;
        RECT 55.390 25.300 55.710 25.480 ;
        RECT 51.300 24.730 51.640 25.050 ;
        RECT 54.950 24.820 55.270 25.040 ;
        RECT 49.930 24.370 50.260 24.710 ;
        RECT 51.300 24.200 51.440 24.730 ;
        RECT 54.950 24.720 55.280 24.820 ;
        RECT 55.140 24.200 55.280 24.720 ;
        RECT 57.640 24.710 57.890 26.660 ;
        RECT 59.200 26.460 59.520 26.660 ;
        RECT 59.660 25.630 59.800 28.490 ;
        RECT 62.170 26.830 62.310 32.160 ;
        RECT 65.280 32.020 65.610 32.160 ;
        RECT 63.630 31.350 64.010 31.370 ;
        RECT 63.630 31.210 64.470 31.350 ;
        RECT 63.630 31.050 64.010 31.210 ;
        RECT 60.400 26.800 62.310 26.830 ;
        RECT 60.370 26.790 62.310 26.800 ;
        RECT 60.080 26.650 62.310 26.790 ;
        RECT 60.080 26.460 60.400 26.650 ;
        RECT 59.460 25.290 59.800 25.630 ;
        RECT 64.330 25.620 64.470 31.210 ;
        RECT 65.360 29.990 65.610 32.020 ;
        RECT 69.880 32.160 73.320 32.300 ;
        RECT 66.070 30.960 66.420 31.290 ;
        RECT 65.360 29.650 65.690 29.990 ;
        RECT 66.070 28.630 66.210 30.960 ;
        RECT 66.070 28.490 67.510 28.630 ;
        RECT 65.270 26.800 65.600 27.060 ;
        RECT 65.270 26.740 67.230 26.800 ;
        RECT 65.340 26.660 67.230 26.740 ;
        RECT 63.100 25.480 64.470 25.620 ;
        RECT 63.100 25.300 63.420 25.480 ;
        RECT 59.010 24.730 59.350 25.050 ;
        RECT 62.660 24.820 62.980 25.040 ;
        RECT 57.640 24.370 57.970 24.710 ;
        RECT 59.010 24.200 59.150 24.730 ;
        RECT 62.660 24.720 62.990 24.820 ;
        RECT 62.850 24.200 62.990 24.720 ;
        RECT 65.350 24.710 65.600 26.660 ;
        RECT 66.910 26.460 67.230 26.660 ;
        RECT 67.370 25.630 67.510 28.490 ;
        RECT 69.880 26.830 70.020 32.160 ;
        RECT 72.990 32.020 73.320 32.160 ;
        RECT 71.340 31.350 71.720 31.370 ;
        RECT 71.340 31.210 72.180 31.350 ;
        RECT 71.340 31.050 71.720 31.210 ;
        RECT 68.110 26.800 70.020 26.830 ;
        RECT 68.080 26.790 70.020 26.800 ;
        RECT 67.790 26.650 70.020 26.790 ;
        RECT 67.790 26.460 68.110 26.650 ;
        RECT 67.170 25.290 67.510 25.630 ;
        RECT 72.040 25.620 72.180 31.210 ;
        RECT 73.070 29.990 73.320 32.020 ;
        RECT 77.590 32.160 81.030 32.300 ;
        RECT 73.780 30.960 74.130 31.290 ;
        RECT 73.070 29.650 73.400 29.990 ;
        RECT 73.780 28.630 73.920 30.960 ;
        RECT 73.780 28.490 75.220 28.630 ;
        RECT 72.980 26.800 73.310 27.060 ;
        RECT 72.980 26.740 74.940 26.800 ;
        RECT 73.050 26.660 74.940 26.740 ;
        RECT 70.810 25.480 72.180 25.620 ;
        RECT 70.810 25.300 71.130 25.480 ;
        RECT 66.720 24.730 67.060 25.050 ;
        RECT 70.370 24.820 70.690 25.040 ;
        RECT 65.350 24.370 65.680 24.710 ;
        RECT 66.720 24.200 66.860 24.730 ;
        RECT 70.370 24.720 70.700 24.820 ;
        RECT 70.560 24.200 70.700 24.720 ;
        RECT 73.060 24.710 73.310 26.660 ;
        RECT 74.620 26.460 74.940 26.660 ;
        RECT 75.080 25.630 75.220 28.490 ;
        RECT 77.590 26.830 77.730 32.160 ;
        RECT 80.700 32.020 81.030 32.160 ;
        RECT 79.050 31.350 79.430 31.370 ;
        RECT 79.050 31.210 79.890 31.350 ;
        RECT 79.050 31.050 79.430 31.210 ;
        RECT 75.820 26.800 77.730 26.830 ;
        RECT 75.790 26.790 77.730 26.800 ;
        RECT 75.500 26.650 77.730 26.790 ;
        RECT 75.500 26.460 75.820 26.650 ;
        RECT 74.880 25.290 75.220 25.630 ;
        RECT 79.750 25.620 79.890 31.210 ;
        RECT 80.780 29.990 81.030 32.020 ;
        RECT 85.300 32.160 88.740 32.300 ;
        RECT 81.490 30.960 81.840 31.290 ;
        RECT 80.780 29.650 81.110 29.990 ;
        RECT 81.490 28.630 81.630 30.960 ;
        RECT 81.490 28.490 82.930 28.630 ;
        RECT 80.690 26.800 81.020 27.060 ;
        RECT 80.690 26.740 82.650 26.800 ;
        RECT 80.760 26.660 82.650 26.740 ;
        RECT 78.520 25.480 79.890 25.620 ;
        RECT 78.520 25.300 78.840 25.480 ;
        RECT 74.430 24.730 74.770 25.050 ;
        RECT 78.080 24.820 78.400 25.040 ;
        RECT 73.060 24.370 73.390 24.710 ;
        RECT 74.430 24.200 74.570 24.730 ;
        RECT 78.080 24.720 78.410 24.820 ;
        RECT 78.270 24.200 78.410 24.720 ;
        RECT 80.770 24.710 81.020 26.660 ;
        RECT 82.330 26.460 82.650 26.660 ;
        RECT 82.790 25.630 82.930 28.490 ;
        RECT 85.300 26.830 85.440 32.160 ;
        RECT 88.410 32.020 88.740 32.160 ;
        RECT 86.760 31.350 87.140 31.370 ;
        RECT 86.760 31.210 87.600 31.350 ;
        RECT 86.760 31.050 87.140 31.210 ;
        RECT 83.530 26.800 85.440 26.830 ;
        RECT 83.500 26.790 85.440 26.800 ;
        RECT 83.210 26.650 85.440 26.790 ;
        RECT 83.210 26.460 83.530 26.650 ;
        RECT 82.590 25.290 82.930 25.630 ;
        RECT 87.460 25.620 87.600 31.210 ;
        RECT 88.490 29.990 88.740 32.020 ;
        RECT 93.010 32.160 96.450 32.300 ;
        RECT 89.200 30.960 89.550 31.290 ;
        RECT 88.490 29.650 88.820 29.990 ;
        RECT 89.200 28.630 89.340 30.960 ;
        RECT 89.200 28.490 90.640 28.630 ;
        RECT 88.400 26.800 88.730 27.060 ;
        RECT 88.400 26.740 90.360 26.800 ;
        RECT 88.470 26.660 90.360 26.740 ;
        RECT 86.230 25.480 87.600 25.620 ;
        RECT 86.230 25.300 86.550 25.480 ;
        RECT 82.140 24.730 82.480 25.050 ;
        RECT 85.790 24.820 86.110 25.040 ;
        RECT 80.770 24.370 81.100 24.710 ;
        RECT 82.140 24.200 82.280 24.730 ;
        RECT 85.790 24.720 86.120 24.820 ;
        RECT 85.980 24.200 86.120 24.720 ;
        RECT 88.480 24.710 88.730 26.660 ;
        RECT 90.040 26.460 90.360 26.660 ;
        RECT 90.500 25.630 90.640 28.490 ;
        RECT 93.010 26.830 93.150 32.160 ;
        RECT 96.120 32.020 96.450 32.160 ;
        RECT 94.470 31.350 94.850 31.370 ;
        RECT 94.470 31.210 95.310 31.350 ;
        RECT 94.470 31.050 94.850 31.210 ;
        RECT 91.240 26.800 93.150 26.830 ;
        RECT 91.210 26.790 93.150 26.800 ;
        RECT 90.920 26.650 93.150 26.790 ;
        RECT 90.920 26.460 91.240 26.650 ;
        RECT 90.300 25.290 90.640 25.630 ;
        RECT 95.170 25.620 95.310 31.210 ;
        RECT 96.200 29.990 96.450 32.020 ;
        RECT 100.720 32.160 104.160 32.300 ;
        RECT 96.910 30.960 97.260 31.290 ;
        RECT 96.200 29.650 96.530 29.990 ;
        RECT 96.910 28.630 97.050 30.960 ;
        RECT 96.910 28.490 98.350 28.630 ;
        RECT 96.110 26.800 96.440 27.060 ;
        RECT 96.110 26.740 98.070 26.800 ;
        RECT 96.180 26.660 98.070 26.740 ;
        RECT 93.940 25.480 95.310 25.620 ;
        RECT 93.940 25.300 94.260 25.480 ;
        RECT 89.850 24.730 90.190 25.050 ;
        RECT 93.500 24.820 93.820 25.040 ;
        RECT 88.480 24.370 88.810 24.710 ;
        RECT 89.850 24.200 89.990 24.730 ;
        RECT 93.500 24.720 93.830 24.820 ;
        RECT 93.690 24.200 93.830 24.720 ;
        RECT 96.190 24.710 96.440 26.660 ;
        RECT 97.750 26.460 98.070 26.660 ;
        RECT 98.210 25.630 98.350 28.490 ;
        RECT 100.720 26.830 100.860 32.160 ;
        RECT 103.830 32.020 104.160 32.160 ;
        RECT 102.180 31.350 102.560 31.370 ;
        RECT 102.180 31.210 103.020 31.350 ;
        RECT 102.180 31.050 102.560 31.210 ;
        RECT 98.950 26.800 100.860 26.830 ;
        RECT 98.920 26.790 100.860 26.800 ;
        RECT 98.630 26.650 100.860 26.790 ;
        RECT 98.630 26.460 98.950 26.650 ;
        RECT 98.010 25.290 98.350 25.630 ;
        RECT 102.880 25.620 103.020 31.210 ;
        RECT 103.910 29.990 104.160 32.020 ;
        RECT 108.430 32.160 111.870 32.300 ;
        RECT 104.620 30.960 104.970 31.290 ;
        RECT 103.910 29.650 104.240 29.990 ;
        RECT 104.620 28.630 104.760 30.960 ;
        RECT 104.620 28.490 106.060 28.630 ;
        RECT 103.820 26.800 104.150 27.060 ;
        RECT 103.820 26.740 105.780 26.800 ;
        RECT 103.890 26.660 105.780 26.740 ;
        RECT 101.650 25.480 103.020 25.620 ;
        RECT 101.650 25.300 101.970 25.480 ;
        RECT 97.560 24.730 97.900 25.050 ;
        RECT 101.210 24.820 101.530 25.040 ;
        RECT 96.190 24.370 96.520 24.710 ;
        RECT 97.560 24.200 97.700 24.730 ;
        RECT 101.210 24.720 101.540 24.820 ;
        RECT 101.400 24.200 101.540 24.720 ;
        RECT 103.900 24.710 104.150 26.660 ;
        RECT 105.460 26.460 105.780 26.660 ;
        RECT 105.920 25.630 106.060 28.490 ;
        RECT 108.430 26.830 108.570 32.160 ;
        RECT 111.540 32.020 111.870 32.160 ;
        RECT 109.890 31.350 110.270 31.370 ;
        RECT 109.890 31.210 110.730 31.350 ;
        RECT 109.890 31.050 110.270 31.210 ;
        RECT 106.660 26.800 108.570 26.830 ;
        RECT 106.630 26.790 108.570 26.800 ;
        RECT 106.340 26.650 108.570 26.790 ;
        RECT 106.340 26.460 106.660 26.650 ;
        RECT 105.720 25.290 106.060 25.630 ;
        RECT 110.590 25.620 110.730 31.210 ;
        RECT 111.620 29.990 111.870 32.020 ;
        RECT 116.140 32.160 119.580 32.300 ;
        RECT 112.330 30.960 112.680 31.290 ;
        RECT 111.620 29.650 111.950 29.990 ;
        RECT 112.330 28.630 112.470 30.960 ;
        RECT 112.330 28.490 113.770 28.630 ;
        RECT 111.530 26.800 111.860 27.060 ;
        RECT 111.530 26.740 113.490 26.800 ;
        RECT 111.600 26.660 113.490 26.740 ;
        RECT 109.360 25.480 110.730 25.620 ;
        RECT 109.360 25.300 109.680 25.480 ;
        RECT 105.270 24.730 105.610 25.050 ;
        RECT 108.920 24.820 109.240 25.040 ;
        RECT 103.900 24.370 104.230 24.710 ;
        RECT 105.270 24.200 105.410 24.730 ;
        RECT 108.920 24.720 109.250 24.820 ;
        RECT 109.110 24.200 109.250 24.720 ;
        RECT 111.610 24.710 111.860 26.660 ;
        RECT 113.170 26.460 113.490 26.660 ;
        RECT 113.630 25.630 113.770 28.490 ;
        RECT 116.140 26.830 116.280 32.160 ;
        RECT 119.250 32.020 119.580 32.160 ;
        RECT 117.600 31.350 117.980 31.370 ;
        RECT 117.600 31.210 118.440 31.350 ;
        RECT 117.600 31.050 117.980 31.210 ;
        RECT 114.370 26.800 116.280 26.830 ;
        RECT 114.340 26.790 116.280 26.800 ;
        RECT 114.050 26.650 116.280 26.790 ;
        RECT 114.050 26.460 114.370 26.650 ;
        RECT 113.430 25.290 113.770 25.630 ;
        RECT 118.300 25.620 118.440 31.210 ;
        RECT 119.330 29.990 119.580 32.020 ;
        RECT 120.040 30.960 120.390 31.290 ;
        RECT 119.330 29.650 119.660 29.990 ;
        RECT 120.040 28.630 120.180 30.960 ;
        RECT 120.040 28.490 121.480 28.630 ;
        RECT 119.240 26.800 119.570 27.060 ;
        RECT 119.240 26.740 121.200 26.800 ;
        RECT 119.310 26.660 121.200 26.740 ;
        RECT 117.070 25.480 118.440 25.620 ;
        RECT 117.070 25.300 117.390 25.480 ;
        RECT 112.980 24.730 113.320 25.050 ;
        RECT 116.630 24.820 116.950 25.040 ;
        RECT 111.610 24.370 111.940 24.710 ;
        RECT 112.980 24.200 113.120 24.730 ;
        RECT 116.630 24.720 116.960 24.820 ;
        RECT 116.820 24.200 116.960 24.720 ;
        RECT 119.320 24.710 119.570 26.660 ;
        RECT 120.880 26.460 121.200 26.660 ;
        RECT 121.340 25.630 121.480 28.490 ;
        RECT 122.080 26.810 123.040 26.830 ;
        RECT 122.080 26.800 123.990 26.810 ;
        RECT 122.050 26.790 123.990 26.800 ;
        RECT 121.760 26.650 123.990 26.790 ;
        RECT 121.760 26.460 122.080 26.650 ;
        RECT 122.840 26.630 123.990 26.650 ;
        RECT 121.140 25.290 121.480 25.630 ;
        RECT 120.690 24.730 121.030 25.050 ;
        RECT 119.320 24.370 119.650 24.710 ;
        RECT 120.690 24.200 120.830 24.730 ;
        RECT -0.320 24.060 60.950 24.200 ;
        RECT 61.910 24.060 123.040 24.200 ;
        RECT -0.750 21.950 -0.560 22.470 ;
        RECT -0.750 6.810 -0.570 21.950 ;
        RECT 28.840 20.890 29.000 24.060 ;
        RECT 28.660 20.570 29.000 20.890 ;
        RECT 90.300 20.910 90.450 24.060 ;
        RECT 90.300 20.840 90.660 20.910 ;
        RECT 90.310 20.560 90.660 20.840 ;
        RECT 58.500 19.840 58.820 20.160 ;
        RECT 58.500 16.120 58.650 19.840 ;
        RECT 58.500 15.940 58.840 16.120 ;
        RECT 58.510 15.800 58.840 15.940 ;
        RECT 123.810 15.980 123.990 26.630 ;
        RECT 124.510 15.980 124.860 16.150 ;
        RECT 123.810 15.830 124.860 15.980 ;
        RECT 58.510 13.940 58.650 15.800 ;
        RECT 58.400 13.610 58.740 13.940 ;
        RECT 28.790 11.980 29.140 12.250 ;
        RECT 90.430 12.040 90.810 12.290 ;
        RECT 28.780 11.880 29.140 11.980 ;
        RECT 90.420 11.910 90.810 12.040 ;
        RECT 28.780 9.400 28.990 11.880 ;
        RECT 90.420 9.400 90.670 11.910 ;
        RECT 0.000 9.260 61.130 9.400 ;
        RECT 62.090 9.260 123.360 9.400 ;
        RECT 2.210 8.730 2.350 9.260 ;
        RECT 3.390 8.750 3.720 9.090 ;
        RECT 2.010 8.410 2.350 8.730 ;
        RECT 1.560 7.830 1.900 8.170 ;
        RECT 0.960 6.810 1.280 7.000 ;
        RECT -0.750 6.670 1.280 6.810 ;
        RECT -0.750 6.660 0.990 6.670 ;
        RECT -0.750 6.630 0.960 6.660 ;
        RECT 1.560 4.970 1.700 7.830 ;
        RECT 1.840 6.800 2.160 7.000 ;
        RECT 3.470 6.800 3.720 8.750 ;
        RECT 6.080 8.740 6.220 9.260 ;
        RECT 6.080 8.640 6.410 8.740 ;
        RECT 9.920 8.730 10.060 9.260 ;
        RECT 11.100 8.750 11.430 9.090 ;
        RECT 6.090 8.420 6.410 8.640 ;
        RECT 9.720 8.410 10.060 8.730 ;
        RECT 5.650 7.980 5.970 8.160 ;
        RECT 4.600 7.840 5.970 7.980 ;
        RECT 1.840 6.720 3.730 6.800 ;
        RECT 1.840 6.660 3.800 6.720 ;
        RECT 3.470 6.400 3.800 6.660 ;
        RECT 1.560 4.830 3.000 4.970 ;
        RECT 2.860 2.500 3.000 4.830 ;
        RECT 3.380 3.470 3.710 3.810 ;
        RECT 2.650 2.170 3.000 2.500 ;
        RECT 3.460 1.440 3.710 3.470 ;
        RECT 4.600 2.250 4.740 7.840 ;
        RECT 9.270 7.830 9.610 8.170 ;
        RECT 8.670 6.810 8.990 7.000 ;
        RECT 6.760 6.670 8.990 6.810 ;
        RECT 6.760 6.660 8.700 6.670 ;
        RECT 6.760 6.630 8.670 6.660 ;
        RECT 5.060 2.250 5.440 2.410 ;
        RECT 4.600 2.110 5.440 2.250 ;
        RECT 5.060 2.090 5.440 2.110 ;
        RECT 3.460 1.300 3.790 1.440 ;
        RECT 6.760 1.300 6.900 6.630 ;
        RECT 9.270 4.970 9.410 7.830 ;
        RECT 9.550 6.800 9.870 7.000 ;
        RECT 11.180 6.800 11.430 8.750 ;
        RECT 13.790 8.740 13.930 9.260 ;
        RECT 13.790 8.640 14.120 8.740 ;
        RECT 17.630 8.730 17.770 9.260 ;
        RECT 18.810 8.750 19.140 9.090 ;
        RECT 13.800 8.420 14.120 8.640 ;
        RECT 17.430 8.410 17.770 8.730 ;
        RECT 13.360 7.980 13.680 8.160 ;
        RECT 12.310 7.840 13.680 7.980 ;
        RECT 9.550 6.720 11.440 6.800 ;
        RECT 9.550 6.660 11.510 6.720 ;
        RECT 11.180 6.400 11.510 6.660 ;
        RECT 9.270 4.830 10.710 4.970 ;
        RECT 10.570 2.500 10.710 4.830 ;
        RECT 11.090 3.470 11.420 3.810 ;
        RECT 10.360 2.170 10.710 2.500 ;
        RECT 3.460 1.160 6.900 1.300 ;
        RECT 11.170 1.440 11.420 3.470 ;
        RECT 12.310 2.250 12.450 7.840 ;
        RECT 16.980 7.830 17.320 8.170 ;
        RECT 16.380 6.810 16.700 7.000 ;
        RECT 14.470 6.670 16.700 6.810 ;
        RECT 14.470 6.660 16.410 6.670 ;
        RECT 14.470 6.630 16.380 6.660 ;
        RECT 12.770 2.250 13.150 2.410 ;
        RECT 12.310 2.110 13.150 2.250 ;
        RECT 12.770 2.090 13.150 2.110 ;
        RECT 11.170 1.300 11.500 1.440 ;
        RECT 14.470 1.300 14.610 6.630 ;
        RECT 16.980 4.970 17.120 7.830 ;
        RECT 17.260 6.800 17.580 7.000 ;
        RECT 18.890 6.800 19.140 8.750 ;
        RECT 21.500 8.740 21.640 9.260 ;
        RECT 21.500 8.640 21.830 8.740 ;
        RECT 25.340 8.730 25.480 9.260 ;
        RECT 26.520 8.750 26.850 9.090 ;
        RECT 21.510 8.420 21.830 8.640 ;
        RECT 25.140 8.410 25.480 8.730 ;
        RECT 21.070 7.980 21.390 8.160 ;
        RECT 20.020 7.840 21.390 7.980 ;
        RECT 17.260 6.720 19.150 6.800 ;
        RECT 17.260 6.660 19.220 6.720 ;
        RECT 18.890 6.400 19.220 6.660 ;
        RECT 16.980 4.830 18.420 4.970 ;
        RECT 18.280 2.500 18.420 4.830 ;
        RECT 18.800 3.470 19.130 3.810 ;
        RECT 18.070 2.170 18.420 2.500 ;
        RECT 11.170 1.160 14.610 1.300 ;
        RECT 18.880 1.440 19.130 3.470 ;
        RECT 20.020 2.250 20.160 7.840 ;
        RECT 24.690 7.830 25.030 8.170 ;
        RECT 24.090 6.810 24.410 7.000 ;
        RECT 22.180 6.670 24.410 6.810 ;
        RECT 22.180 6.660 24.120 6.670 ;
        RECT 22.180 6.630 24.090 6.660 ;
        RECT 20.480 2.250 20.860 2.410 ;
        RECT 20.020 2.110 20.860 2.250 ;
        RECT 20.480 2.090 20.860 2.110 ;
        RECT 18.880 1.300 19.210 1.440 ;
        RECT 22.180 1.300 22.320 6.630 ;
        RECT 24.690 4.970 24.830 7.830 ;
        RECT 24.970 6.800 25.290 7.000 ;
        RECT 26.600 6.800 26.850 8.750 ;
        RECT 29.210 8.740 29.350 9.260 ;
        RECT 29.210 8.640 29.540 8.740 ;
        RECT 33.050 8.730 33.190 9.260 ;
        RECT 34.230 8.750 34.560 9.090 ;
        RECT 29.220 8.420 29.540 8.640 ;
        RECT 32.850 8.410 33.190 8.730 ;
        RECT 28.780 7.980 29.100 8.160 ;
        RECT 27.730 7.840 29.100 7.980 ;
        RECT 24.970 6.720 26.860 6.800 ;
        RECT 24.970 6.660 26.930 6.720 ;
        RECT 26.600 6.400 26.930 6.660 ;
        RECT 24.690 4.830 26.130 4.970 ;
        RECT 25.990 2.500 26.130 4.830 ;
        RECT 26.510 3.470 26.840 3.810 ;
        RECT 25.780 2.170 26.130 2.500 ;
        RECT 18.880 1.160 22.320 1.300 ;
        RECT 26.590 1.440 26.840 3.470 ;
        RECT 27.730 2.250 27.870 7.840 ;
        RECT 32.400 7.830 32.740 8.170 ;
        RECT 31.800 6.810 32.120 7.000 ;
        RECT 29.890 6.670 32.120 6.810 ;
        RECT 29.890 6.660 31.830 6.670 ;
        RECT 29.890 6.630 31.800 6.660 ;
        RECT 28.190 2.250 28.570 2.410 ;
        RECT 27.730 2.110 28.570 2.250 ;
        RECT 28.190 2.090 28.570 2.110 ;
        RECT 26.590 1.300 26.920 1.440 ;
        RECT 29.890 1.300 30.030 6.630 ;
        RECT 32.400 4.970 32.540 7.830 ;
        RECT 32.680 6.800 33.000 7.000 ;
        RECT 34.310 6.800 34.560 8.750 ;
        RECT 36.920 8.740 37.060 9.260 ;
        RECT 36.920 8.640 37.250 8.740 ;
        RECT 40.760 8.730 40.900 9.260 ;
        RECT 41.940 8.750 42.270 9.090 ;
        RECT 36.930 8.420 37.250 8.640 ;
        RECT 40.560 8.410 40.900 8.730 ;
        RECT 36.490 7.980 36.810 8.160 ;
        RECT 35.440 7.840 36.810 7.980 ;
        RECT 32.680 6.720 34.570 6.800 ;
        RECT 32.680 6.660 34.640 6.720 ;
        RECT 34.310 6.400 34.640 6.660 ;
        RECT 32.400 4.830 33.840 4.970 ;
        RECT 33.700 2.500 33.840 4.830 ;
        RECT 34.220 3.470 34.550 3.810 ;
        RECT 33.490 2.170 33.840 2.500 ;
        RECT 26.590 1.160 30.030 1.300 ;
        RECT 34.300 1.440 34.550 3.470 ;
        RECT 35.440 2.250 35.580 7.840 ;
        RECT 40.110 7.830 40.450 8.170 ;
        RECT 39.510 6.810 39.830 7.000 ;
        RECT 37.600 6.670 39.830 6.810 ;
        RECT 37.600 6.660 39.540 6.670 ;
        RECT 37.600 6.630 39.510 6.660 ;
        RECT 35.900 2.250 36.280 2.410 ;
        RECT 35.440 2.110 36.280 2.250 ;
        RECT 35.900 2.090 36.280 2.110 ;
        RECT 34.300 1.300 34.630 1.440 ;
        RECT 37.600 1.300 37.740 6.630 ;
        RECT 40.110 4.970 40.250 7.830 ;
        RECT 40.390 6.800 40.710 7.000 ;
        RECT 42.020 6.800 42.270 8.750 ;
        RECT 44.630 8.740 44.770 9.260 ;
        RECT 44.630 8.640 44.960 8.740 ;
        RECT 48.470 8.730 48.610 9.260 ;
        RECT 49.650 8.750 49.980 9.090 ;
        RECT 44.640 8.420 44.960 8.640 ;
        RECT 48.270 8.410 48.610 8.730 ;
        RECT 44.200 7.980 44.520 8.160 ;
        RECT 43.150 7.840 44.520 7.980 ;
        RECT 40.390 6.720 42.280 6.800 ;
        RECT 40.390 6.660 42.350 6.720 ;
        RECT 42.020 6.400 42.350 6.660 ;
        RECT 40.110 4.830 41.550 4.970 ;
        RECT 41.410 2.500 41.550 4.830 ;
        RECT 41.930 3.470 42.260 3.810 ;
        RECT 41.200 2.170 41.550 2.500 ;
        RECT 34.300 1.160 37.740 1.300 ;
        RECT 42.010 1.440 42.260 3.470 ;
        RECT 43.150 2.250 43.290 7.840 ;
        RECT 47.820 7.830 48.160 8.170 ;
        RECT 47.220 6.810 47.540 7.000 ;
        RECT 45.310 6.670 47.540 6.810 ;
        RECT 45.310 6.660 47.250 6.670 ;
        RECT 45.310 6.630 47.220 6.660 ;
        RECT 43.610 2.250 43.990 2.410 ;
        RECT 43.150 2.110 43.990 2.250 ;
        RECT 43.610 2.090 43.990 2.110 ;
        RECT 42.010 1.300 42.340 1.440 ;
        RECT 45.310 1.300 45.450 6.630 ;
        RECT 47.820 4.970 47.960 7.830 ;
        RECT 48.100 6.800 48.420 7.000 ;
        RECT 49.730 6.800 49.980 8.750 ;
        RECT 52.340 8.740 52.480 9.260 ;
        RECT 52.340 8.640 52.670 8.740 ;
        RECT 56.180 8.730 56.320 9.260 ;
        RECT 57.360 8.750 57.690 9.090 ;
        RECT 52.350 8.420 52.670 8.640 ;
        RECT 55.980 8.410 56.320 8.730 ;
        RECT 51.910 7.980 52.230 8.160 ;
        RECT 50.860 7.840 52.230 7.980 ;
        RECT 48.100 6.720 49.990 6.800 ;
        RECT 48.100 6.660 50.060 6.720 ;
        RECT 49.730 6.400 50.060 6.660 ;
        RECT 47.820 4.830 49.260 4.970 ;
        RECT 49.120 2.500 49.260 4.830 ;
        RECT 49.640 3.470 49.970 3.810 ;
        RECT 48.910 2.170 49.260 2.500 ;
        RECT 42.010 1.160 45.450 1.300 ;
        RECT 49.720 1.440 49.970 3.470 ;
        RECT 50.860 2.250 51.000 7.840 ;
        RECT 55.530 7.830 55.870 8.170 ;
        RECT 54.930 6.810 55.250 7.000 ;
        RECT 53.020 6.670 55.250 6.810 ;
        RECT 53.020 6.660 54.960 6.670 ;
        RECT 53.020 6.630 54.930 6.660 ;
        RECT 51.320 2.250 51.700 2.410 ;
        RECT 50.860 2.110 51.700 2.250 ;
        RECT 51.320 2.090 51.700 2.110 ;
        RECT 49.720 1.300 50.050 1.440 ;
        RECT 53.020 1.300 53.160 6.630 ;
        RECT 55.530 4.970 55.670 7.830 ;
        RECT 55.810 6.800 56.130 7.000 ;
        RECT 57.440 6.800 57.690 8.750 ;
        RECT 60.050 8.740 60.190 9.260 ;
        RECT 60.050 8.640 60.380 8.740 ;
        RECT 63.890 8.730 64.030 9.260 ;
        RECT 65.070 8.750 65.400 9.090 ;
        RECT 60.060 8.420 60.380 8.640 ;
        RECT 63.690 8.410 64.030 8.730 ;
        RECT 59.620 7.980 59.940 8.160 ;
        RECT 58.570 7.840 59.940 7.980 ;
        RECT 55.810 6.720 57.700 6.800 ;
        RECT 55.810 6.660 57.770 6.720 ;
        RECT 57.440 6.400 57.770 6.660 ;
        RECT 55.530 4.830 56.970 4.970 ;
        RECT 56.830 2.500 56.970 4.830 ;
        RECT 57.350 3.470 57.680 3.810 ;
        RECT 56.620 2.170 56.970 2.500 ;
        RECT 49.720 1.160 53.160 1.300 ;
        RECT 57.430 1.440 57.680 3.470 ;
        RECT 58.570 2.250 58.710 7.840 ;
        RECT 63.240 7.830 63.580 8.170 ;
        RECT 62.640 6.810 62.960 7.000 ;
        RECT 60.730 6.670 62.960 6.810 ;
        RECT 60.730 6.660 62.670 6.670 ;
        RECT 60.730 6.630 62.640 6.660 ;
        RECT 59.030 2.250 59.410 2.410 ;
        RECT 58.570 2.110 59.410 2.250 ;
        RECT 59.030 2.090 59.410 2.110 ;
        RECT 57.430 1.300 57.760 1.440 ;
        RECT 60.730 1.300 60.870 6.630 ;
        RECT 63.240 4.970 63.380 7.830 ;
        RECT 63.520 6.800 63.840 7.000 ;
        RECT 65.150 6.800 65.400 8.750 ;
        RECT 67.760 8.740 67.900 9.260 ;
        RECT 67.760 8.640 68.090 8.740 ;
        RECT 71.600 8.730 71.740 9.260 ;
        RECT 72.780 8.750 73.110 9.090 ;
        RECT 67.770 8.420 68.090 8.640 ;
        RECT 71.400 8.410 71.740 8.730 ;
        RECT 67.330 7.980 67.650 8.160 ;
        RECT 66.280 7.840 67.650 7.980 ;
        RECT 63.520 6.720 65.410 6.800 ;
        RECT 63.520 6.660 65.480 6.720 ;
        RECT 65.150 6.400 65.480 6.660 ;
        RECT 63.240 4.830 64.680 4.970 ;
        RECT 64.540 2.500 64.680 4.830 ;
        RECT 65.060 3.470 65.390 3.810 ;
        RECT 64.330 2.170 64.680 2.500 ;
        RECT 57.430 1.160 60.870 1.300 ;
        RECT 65.140 1.440 65.390 3.470 ;
        RECT 66.280 2.250 66.420 7.840 ;
        RECT 70.950 7.830 71.290 8.170 ;
        RECT 70.350 6.810 70.670 7.000 ;
        RECT 68.440 6.670 70.670 6.810 ;
        RECT 68.440 6.660 70.380 6.670 ;
        RECT 68.440 6.630 70.350 6.660 ;
        RECT 66.740 2.250 67.120 2.410 ;
        RECT 66.280 2.110 67.120 2.250 ;
        RECT 66.740 2.090 67.120 2.110 ;
        RECT 65.140 1.300 65.470 1.440 ;
        RECT 68.440 1.300 68.580 6.630 ;
        RECT 70.950 4.970 71.090 7.830 ;
        RECT 71.230 6.800 71.550 7.000 ;
        RECT 72.860 6.800 73.110 8.750 ;
        RECT 75.470 8.740 75.610 9.260 ;
        RECT 75.470 8.640 75.800 8.740 ;
        RECT 79.310 8.730 79.450 9.260 ;
        RECT 80.490 8.750 80.820 9.090 ;
        RECT 75.480 8.420 75.800 8.640 ;
        RECT 79.110 8.410 79.450 8.730 ;
        RECT 75.040 7.980 75.360 8.160 ;
        RECT 73.990 7.840 75.360 7.980 ;
        RECT 71.230 6.720 73.120 6.800 ;
        RECT 71.230 6.660 73.190 6.720 ;
        RECT 72.860 6.400 73.190 6.660 ;
        RECT 70.950 4.830 72.390 4.970 ;
        RECT 72.250 2.500 72.390 4.830 ;
        RECT 72.770 3.470 73.100 3.810 ;
        RECT 72.040 2.170 72.390 2.500 ;
        RECT 65.140 1.160 68.580 1.300 ;
        RECT 72.850 1.440 73.100 3.470 ;
        RECT 73.990 2.250 74.130 7.840 ;
        RECT 78.660 7.830 79.000 8.170 ;
        RECT 78.060 6.810 78.380 7.000 ;
        RECT 76.150 6.670 78.380 6.810 ;
        RECT 76.150 6.660 78.090 6.670 ;
        RECT 76.150 6.630 78.060 6.660 ;
        RECT 74.450 2.250 74.830 2.410 ;
        RECT 73.990 2.110 74.830 2.250 ;
        RECT 74.450 2.090 74.830 2.110 ;
        RECT 72.850 1.300 73.180 1.440 ;
        RECT 76.150 1.300 76.290 6.630 ;
        RECT 78.660 4.970 78.800 7.830 ;
        RECT 78.940 6.800 79.260 7.000 ;
        RECT 80.570 6.800 80.820 8.750 ;
        RECT 83.180 8.740 83.320 9.260 ;
        RECT 83.180 8.640 83.510 8.740 ;
        RECT 87.020 8.730 87.160 9.260 ;
        RECT 88.200 8.750 88.530 9.090 ;
        RECT 83.190 8.420 83.510 8.640 ;
        RECT 86.820 8.410 87.160 8.730 ;
        RECT 82.750 7.980 83.070 8.160 ;
        RECT 81.700 7.840 83.070 7.980 ;
        RECT 78.940 6.720 80.830 6.800 ;
        RECT 78.940 6.660 80.900 6.720 ;
        RECT 80.570 6.400 80.900 6.660 ;
        RECT 78.660 4.830 80.100 4.970 ;
        RECT 79.960 2.500 80.100 4.830 ;
        RECT 80.480 3.470 80.810 3.810 ;
        RECT 79.750 2.170 80.100 2.500 ;
        RECT 72.850 1.160 76.290 1.300 ;
        RECT 80.560 1.440 80.810 3.470 ;
        RECT 81.700 2.250 81.840 7.840 ;
        RECT 86.370 7.830 86.710 8.170 ;
        RECT 85.770 6.810 86.090 7.000 ;
        RECT 83.860 6.670 86.090 6.810 ;
        RECT 83.860 6.660 85.800 6.670 ;
        RECT 83.860 6.630 85.770 6.660 ;
        RECT 82.160 2.250 82.540 2.410 ;
        RECT 81.700 2.110 82.540 2.250 ;
        RECT 82.160 2.090 82.540 2.110 ;
        RECT 80.560 1.300 80.890 1.440 ;
        RECT 83.860 1.300 84.000 6.630 ;
        RECT 86.370 4.970 86.510 7.830 ;
        RECT 86.650 6.800 86.970 7.000 ;
        RECT 88.280 6.800 88.530 8.750 ;
        RECT 90.890 8.740 91.030 9.260 ;
        RECT 90.890 8.640 91.220 8.740 ;
        RECT 94.730 8.730 94.870 9.260 ;
        RECT 95.910 8.750 96.240 9.090 ;
        RECT 90.900 8.420 91.220 8.640 ;
        RECT 94.530 8.410 94.870 8.730 ;
        RECT 90.460 7.980 90.780 8.160 ;
        RECT 89.410 7.840 90.780 7.980 ;
        RECT 86.650 6.720 88.540 6.800 ;
        RECT 86.650 6.660 88.610 6.720 ;
        RECT 88.280 6.400 88.610 6.660 ;
        RECT 86.370 4.830 87.810 4.970 ;
        RECT 87.670 2.500 87.810 4.830 ;
        RECT 88.190 3.470 88.520 3.810 ;
        RECT 87.460 2.170 87.810 2.500 ;
        RECT 80.560 1.160 84.000 1.300 ;
        RECT 88.270 1.440 88.520 3.470 ;
        RECT 89.410 2.250 89.550 7.840 ;
        RECT 94.080 7.830 94.420 8.170 ;
        RECT 93.480 6.810 93.800 7.000 ;
        RECT 91.570 6.670 93.800 6.810 ;
        RECT 91.570 6.660 93.510 6.670 ;
        RECT 91.570 6.630 93.480 6.660 ;
        RECT 89.870 2.250 90.250 2.410 ;
        RECT 89.410 2.110 90.250 2.250 ;
        RECT 89.870 2.090 90.250 2.110 ;
        RECT 88.270 1.300 88.600 1.440 ;
        RECT 91.570 1.300 91.710 6.630 ;
        RECT 94.080 4.970 94.220 7.830 ;
        RECT 94.360 6.800 94.680 7.000 ;
        RECT 95.990 6.800 96.240 8.750 ;
        RECT 98.600 8.740 98.740 9.260 ;
        RECT 98.600 8.640 98.930 8.740 ;
        RECT 102.440 8.730 102.580 9.260 ;
        RECT 103.620 8.750 103.950 9.090 ;
        RECT 98.610 8.420 98.930 8.640 ;
        RECT 102.240 8.410 102.580 8.730 ;
        RECT 98.170 7.980 98.490 8.160 ;
        RECT 97.120 7.840 98.490 7.980 ;
        RECT 94.360 6.720 96.250 6.800 ;
        RECT 94.360 6.660 96.320 6.720 ;
        RECT 95.990 6.400 96.320 6.660 ;
        RECT 94.080 4.830 95.520 4.970 ;
        RECT 95.380 2.500 95.520 4.830 ;
        RECT 95.900 3.470 96.230 3.810 ;
        RECT 95.170 2.170 95.520 2.500 ;
        RECT 88.270 1.160 91.710 1.300 ;
        RECT 95.980 1.440 96.230 3.470 ;
        RECT 97.120 2.250 97.260 7.840 ;
        RECT 101.790 7.830 102.130 8.170 ;
        RECT 101.190 6.810 101.510 7.000 ;
        RECT 99.280 6.670 101.510 6.810 ;
        RECT 99.280 6.660 101.220 6.670 ;
        RECT 99.280 6.630 101.190 6.660 ;
        RECT 97.580 2.250 97.960 2.410 ;
        RECT 97.120 2.110 97.960 2.250 ;
        RECT 97.580 2.090 97.960 2.110 ;
        RECT 95.980 1.300 96.310 1.440 ;
        RECT 99.280 1.300 99.420 6.630 ;
        RECT 101.790 4.970 101.930 7.830 ;
        RECT 102.070 6.800 102.390 7.000 ;
        RECT 103.700 6.800 103.950 8.750 ;
        RECT 106.310 8.740 106.450 9.260 ;
        RECT 106.310 8.640 106.640 8.740 ;
        RECT 110.150 8.730 110.290 9.260 ;
        RECT 111.330 8.750 111.660 9.090 ;
        RECT 106.320 8.420 106.640 8.640 ;
        RECT 109.950 8.410 110.290 8.730 ;
        RECT 105.880 7.980 106.200 8.160 ;
        RECT 104.830 7.840 106.200 7.980 ;
        RECT 102.070 6.720 103.960 6.800 ;
        RECT 102.070 6.660 104.030 6.720 ;
        RECT 103.700 6.400 104.030 6.660 ;
        RECT 101.790 4.830 103.230 4.970 ;
        RECT 103.090 2.500 103.230 4.830 ;
        RECT 103.610 3.470 103.940 3.810 ;
        RECT 102.880 2.170 103.230 2.500 ;
        RECT 95.980 1.160 99.420 1.300 ;
        RECT 103.690 1.440 103.940 3.470 ;
        RECT 104.830 2.250 104.970 7.840 ;
        RECT 109.500 7.830 109.840 8.170 ;
        RECT 108.900 6.810 109.220 7.000 ;
        RECT 106.990 6.670 109.220 6.810 ;
        RECT 106.990 6.660 108.930 6.670 ;
        RECT 106.990 6.630 108.900 6.660 ;
        RECT 105.290 2.250 105.670 2.410 ;
        RECT 104.830 2.110 105.670 2.250 ;
        RECT 105.290 2.090 105.670 2.110 ;
        RECT 103.690 1.300 104.020 1.440 ;
        RECT 106.990 1.300 107.130 6.630 ;
        RECT 109.500 4.970 109.640 7.830 ;
        RECT 109.780 6.800 110.100 7.000 ;
        RECT 111.410 6.800 111.660 8.750 ;
        RECT 114.020 8.740 114.160 9.260 ;
        RECT 114.020 8.640 114.350 8.740 ;
        RECT 117.860 8.730 118.000 9.260 ;
        RECT 119.040 8.750 119.370 9.090 ;
        RECT 114.030 8.420 114.350 8.640 ;
        RECT 117.660 8.410 118.000 8.730 ;
        RECT 113.590 7.980 113.910 8.160 ;
        RECT 112.540 7.840 113.910 7.980 ;
        RECT 109.780 6.720 111.670 6.800 ;
        RECT 109.780 6.660 111.740 6.720 ;
        RECT 111.410 6.400 111.740 6.660 ;
        RECT 109.500 4.830 110.940 4.970 ;
        RECT 110.800 2.500 110.940 4.830 ;
        RECT 111.320 3.470 111.650 3.810 ;
        RECT 110.590 2.170 110.940 2.500 ;
        RECT 103.690 1.160 107.130 1.300 ;
        RECT 111.400 1.440 111.650 3.470 ;
        RECT 112.540 2.250 112.680 7.840 ;
        RECT 117.210 7.830 117.550 8.170 ;
        RECT 116.610 6.810 116.930 7.000 ;
        RECT 114.700 6.670 116.930 6.810 ;
        RECT 114.700 6.660 116.640 6.670 ;
        RECT 114.700 6.630 116.610 6.660 ;
        RECT 113.000 2.250 113.380 2.410 ;
        RECT 112.540 2.110 113.380 2.250 ;
        RECT 113.000 2.090 113.380 2.110 ;
        RECT 111.400 1.300 111.730 1.440 ;
        RECT 114.700 1.300 114.840 6.630 ;
        RECT 117.210 4.970 117.350 7.830 ;
        RECT 117.490 6.800 117.810 7.000 ;
        RECT 119.120 6.800 119.370 8.750 ;
        RECT 121.730 8.740 121.870 9.260 ;
        RECT 121.730 8.640 122.060 8.740 ;
        RECT 121.740 8.420 122.060 8.640 ;
        RECT 121.300 7.980 121.620 8.160 ;
        RECT 120.250 7.840 121.620 7.980 ;
        RECT 117.490 6.720 119.380 6.800 ;
        RECT 117.490 6.660 119.450 6.720 ;
        RECT 119.120 6.400 119.450 6.660 ;
        RECT 117.210 4.830 118.650 4.970 ;
        RECT 118.510 2.500 118.650 4.830 ;
        RECT 119.030 3.470 119.360 3.810 ;
        RECT 118.300 2.170 118.650 2.500 ;
        RECT 111.400 1.160 114.840 1.300 ;
        RECT 119.110 1.440 119.360 3.470 ;
        RECT 120.250 2.250 120.390 7.840 ;
        RECT 123.810 6.810 123.990 15.830 ;
        RECT 122.410 6.630 123.990 6.810 ;
        RECT 120.710 2.250 121.090 2.410 ;
        RECT 120.250 2.110 121.090 2.250 ;
        RECT 120.710 2.090 121.090 2.110 ;
        RECT 119.110 1.300 119.440 1.440 ;
        RECT 122.410 1.300 122.550 6.630 ;
        RECT 119.110 1.160 122.550 1.300 ;
        RECT 3.460 1.120 3.790 1.160 ;
        RECT 11.170 1.120 11.500 1.160 ;
        RECT 18.880 1.120 19.210 1.160 ;
        RECT 26.590 1.120 26.920 1.160 ;
        RECT 34.300 1.120 34.630 1.160 ;
        RECT 42.010 1.120 42.340 1.160 ;
        RECT 49.720 1.120 50.050 1.160 ;
        RECT 57.430 1.120 57.760 1.160 ;
        RECT 65.140 1.120 65.470 1.160 ;
        RECT 72.850 1.120 73.180 1.160 ;
        RECT 80.560 1.120 80.890 1.160 ;
        RECT 88.270 1.120 88.600 1.160 ;
        RECT 95.980 1.120 96.310 1.160 ;
        RECT 103.690 1.120 104.020 1.160 ;
        RECT 111.400 1.120 111.730 1.160 ;
        RECT 119.110 1.120 119.440 1.160 ;
  END
END 32BR
END LIBRARY

