magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 42 21 228 203
rect 42 17 63 21
rect 29 -17 63 17
<< locali >>
rect 144 297 210 493
rect 64 215 130 263
rect 164 177 210 297
rect 144 51 210 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 68 299 110 527
rect 64 17 110 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel locali s 64 215 130 263 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 276 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 42 17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 42 21 228 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 314 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 276 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 144 51 210 177 6 Y
port 6 nsew signal output
rlabel locali s 164 177 210 297 6 Y
port 6 nsew signal output
rlabel locali s 144 297 210 493 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 276 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2228044
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2224550
<< end >>
