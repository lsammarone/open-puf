magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 3835 6565 6265 6671
rect 6295 5999 6467 7237
rect 3900 4537 5249 5153
rect 3900 4431 6254 4537
rect 3900 4400 5264 4431
rect 3900 3857 5249 4400
rect 6325 3857 6467 5111
<< pwell >>
rect 3845 7556 6259 7642
rect 3842 5594 6280 5680
rect 5298 5447 6280 5594
rect 5088 3452 6291 3538
rect 5088 3358 5174 3452
<< mvpsubdiff >>
rect 3871 7582 3895 7616
rect 3929 7582 3963 7616
rect 3997 7582 4031 7616
rect 4065 7582 4099 7616
rect 4133 7582 4167 7616
rect 4201 7582 4235 7616
rect 4269 7582 4303 7616
rect 4337 7582 4371 7616
rect 4405 7582 4439 7616
rect 4473 7582 4507 7616
rect 4541 7582 4575 7616
rect 4609 7582 4643 7616
rect 4677 7582 4711 7616
rect 4745 7582 4779 7616
rect 4813 7582 4847 7616
rect 4881 7582 4915 7616
rect 4949 7582 4983 7616
rect 5017 7582 5051 7616
rect 5085 7582 5119 7616
rect 5153 7582 5187 7616
rect 5221 7582 5255 7616
rect 5289 7582 5323 7616
rect 5357 7582 5391 7616
rect 5425 7582 5459 7616
rect 5493 7582 5527 7616
rect 5561 7582 5595 7616
rect 5629 7582 5663 7616
rect 5697 7582 5731 7616
rect 5765 7582 5799 7616
rect 5833 7582 5867 7616
rect 5901 7582 5935 7616
rect 5969 7582 6003 7616
rect 6037 7582 6071 7616
rect 6105 7582 6139 7616
rect 6173 7582 6233 7616
rect 3868 5620 3892 5654
rect 3926 5620 3960 5654
rect 3994 5620 4028 5654
rect 4062 5620 4096 5654
rect 4130 5620 4164 5654
rect 4198 5620 4232 5654
rect 4266 5620 4300 5654
rect 4334 5620 4368 5654
rect 4402 5620 4436 5654
rect 4470 5620 4504 5654
rect 4538 5620 4572 5654
rect 4606 5620 4640 5654
rect 4674 5620 4708 5654
rect 4742 5620 4776 5654
rect 4810 5620 4844 5654
rect 4878 5620 4912 5654
rect 4946 5620 4980 5654
rect 5014 5620 5048 5654
rect 5082 5620 5116 5654
rect 5150 5620 5184 5654
rect 5218 5620 5252 5654
rect 5286 5620 5320 5654
rect 5354 5620 5388 5654
rect 5422 5620 5456 5654
rect 5490 5620 5524 5654
rect 5558 5620 5592 5654
rect 5626 5620 5660 5654
rect 5694 5620 5728 5654
rect 5762 5620 5796 5654
rect 5830 5620 5864 5654
rect 5898 5620 5932 5654
rect 5966 5620 6000 5654
rect 6034 5620 6068 5654
rect 6102 5620 6136 5654
rect 6170 5620 6254 5654
rect 5324 5581 6254 5620
rect 5324 5547 5348 5581
rect 5382 5547 5416 5581
rect 5450 5547 5484 5581
rect 5518 5547 5552 5581
rect 5586 5547 5620 5581
rect 5654 5547 5688 5581
rect 5722 5547 5756 5581
rect 5790 5547 5824 5581
rect 5858 5547 5892 5581
rect 5926 5547 5960 5581
rect 5994 5547 6028 5581
rect 6062 5547 6096 5581
rect 6130 5547 6164 5581
rect 6198 5547 6254 5581
rect 5324 5507 6254 5547
rect 5324 5473 5348 5507
rect 5382 5473 5416 5507
rect 5450 5473 5484 5507
rect 5518 5473 5552 5507
rect 5586 5473 5620 5507
rect 5654 5473 5688 5507
rect 5722 5473 5756 5507
rect 5790 5473 5824 5507
rect 5858 5473 5892 5507
rect 5926 5473 5960 5507
rect 5994 5473 6028 5507
rect 6062 5473 6096 5507
rect 6130 5473 6164 5507
rect 6198 5473 6254 5507
rect 5114 3478 5138 3512
rect 5172 3478 5206 3512
rect 5240 3478 5274 3512
rect 5308 3478 5342 3512
rect 5376 3478 5410 3512
rect 5444 3478 5478 3512
rect 5512 3478 5546 3512
rect 5580 3478 5614 3512
rect 5648 3478 5682 3512
rect 5716 3478 5750 3512
rect 5784 3478 5818 3512
rect 5852 3478 5886 3512
rect 5920 3478 5954 3512
rect 5988 3478 6022 3512
rect 6056 3478 6090 3512
rect 6124 3478 6158 3512
rect 6192 3478 6265 3512
rect 5114 3444 5148 3478
rect 5114 3384 5148 3410
<< mvnsubdiff >>
rect 3871 6601 3895 6635
rect 3929 6601 3963 6635
rect 3997 6601 4031 6635
rect 4065 6601 4099 6635
rect 4133 6601 4167 6635
rect 4201 6601 4235 6635
rect 4269 6601 4303 6635
rect 4337 6601 4371 6635
rect 4405 6601 4439 6635
rect 4473 6601 4507 6635
rect 4541 6601 4575 6635
rect 4609 6601 4643 6635
rect 4677 6601 4711 6635
rect 4745 6601 4779 6635
rect 4813 6601 4847 6635
rect 4881 6601 4915 6635
rect 4949 6601 4983 6635
rect 5017 6601 5051 6635
rect 5085 6601 5119 6635
rect 5153 6601 5187 6635
rect 5221 6601 5255 6635
rect 5289 6601 5323 6635
rect 5357 6601 5391 6635
rect 5425 6601 5459 6635
rect 5493 6601 5527 6635
rect 5561 6601 5595 6635
rect 5629 6601 5663 6635
rect 5697 6601 5731 6635
rect 5765 6601 5799 6635
rect 5833 6601 5867 6635
rect 5901 6601 5935 6635
rect 5969 6601 6003 6635
rect 6037 6601 6071 6635
rect 6105 6601 6139 6635
rect 6173 6601 6229 6635
rect 5194 4470 5230 4501
rect 3996 4436 4035 4470
rect 4069 4436 4103 4470
rect 4137 4436 4171 4470
rect 4205 4436 4239 4470
rect 4273 4436 4307 4470
rect 4341 4436 4375 4470
rect 4409 4436 4443 4470
rect 4477 4436 4511 4470
rect 4545 4436 4579 4470
rect 4613 4436 4647 4470
rect 4681 4436 4715 4470
rect 4749 4436 4783 4470
rect 4817 4436 4851 4470
rect 4885 4436 4919 4470
rect 4953 4436 4987 4470
rect 5021 4436 5055 4470
rect 5089 4436 5123 4470
rect 5157 4467 5230 4470
rect 5264 4467 5298 4501
rect 5332 4467 5366 4501
rect 5400 4467 5434 4501
rect 5468 4467 5502 4501
rect 5536 4467 5570 4501
rect 5604 4467 5638 4501
rect 5672 4467 5706 4501
rect 5740 4467 5774 4501
rect 5808 4467 5842 4501
rect 5876 4467 5910 4501
rect 5944 4467 5978 4501
rect 6012 4467 6046 4501
rect 6080 4467 6114 4501
rect 6148 4467 6218 4501
rect 5157 4436 5228 4467
<< mvpsubdiffcont >>
rect 3895 7582 3929 7616
rect 3963 7582 3997 7616
rect 4031 7582 4065 7616
rect 4099 7582 4133 7616
rect 4167 7582 4201 7616
rect 4235 7582 4269 7616
rect 4303 7582 4337 7616
rect 4371 7582 4405 7616
rect 4439 7582 4473 7616
rect 4507 7582 4541 7616
rect 4575 7582 4609 7616
rect 4643 7582 4677 7616
rect 4711 7582 4745 7616
rect 4779 7582 4813 7616
rect 4847 7582 4881 7616
rect 4915 7582 4949 7616
rect 4983 7582 5017 7616
rect 5051 7582 5085 7616
rect 5119 7582 5153 7616
rect 5187 7582 5221 7616
rect 5255 7582 5289 7616
rect 5323 7582 5357 7616
rect 5391 7582 5425 7616
rect 5459 7582 5493 7616
rect 5527 7582 5561 7616
rect 5595 7582 5629 7616
rect 5663 7582 5697 7616
rect 5731 7582 5765 7616
rect 5799 7582 5833 7616
rect 5867 7582 5901 7616
rect 5935 7582 5969 7616
rect 6003 7582 6037 7616
rect 6071 7582 6105 7616
rect 6139 7582 6173 7616
rect 3892 5620 3926 5654
rect 3960 5620 3994 5654
rect 4028 5620 4062 5654
rect 4096 5620 4130 5654
rect 4164 5620 4198 5654
rect 4232 5620 4266 5654
rect 4300 5620 4334 5654
rect 4368 5620 4402 5654
rect 4436 5620 4470 5654
rect 4504 5620 4538 5654
rect 4572 5620 4606 5654
rect 4640 5620 4674 5654
rect 4708 5620 4742 5654
rect 4776 5620 4810 5654
rect 4844 5620 4878 5654
rect 4912 5620 4946 5654
rect 4980 5620 5014 5654
rect 5048 5620 5082 5654
rect 5116 5620 5150 5654
rect 5184 5620 5218 5654
rect 5252 5620 5286 5654
rect 5320 5620 5354 5654
rect 5388 5620 5422 5654
rect 5456 5620 5490 5654
rect 5524 5620 5558 5654
rect 5592 5620 5626 5654
rect 5660 5620 5694 5654
rect 5728 5620 5762 5654
rect 5796 5620 5830 5654
rect 5864 5620 5898 5654
rect 5932 5620 5966 5654
rect 6000 5620 6034 5654
rect 6068 5620 6102 5654
rect 6136 5620 6170 5654
rect 5348 5547 5382 5581
rect 5416 5547 5450 5581
rect 5484 5547 5518 5581
rect 5552 5547 5586 5581
rect 5620 5547 5654 5581
rect 5688 5547 5722 5581
rect 5756 5547 5790 5581
rect 5824 5547 5858 5581
rect 5892 5547 5926 5581
rect 5960 5547 5994 5581
rect 6028 5547 6062 5581
rect 6096 5547 6130 5581
rect 6164 5547 6198 5581
rect 5348 5473 5382 5507
rect 5416 5473 5450 5507
rect 5484 5473 5518 5507
rect 5552 5473 5586 5507
rect 5620 5473 5654 5507
rect 5688 5473 5722 5507
rect 5756 5473 5790 5507
rect 5824 5473 5858 5507
rect 5892 5473 5926 5507
rect 5960 5473 5994 5507
rect 6028 5473 6062 5507
rect 6096 5473 6130 5507
rect 6164 5473 6198 5507
rect 5138 3478 5172 3512
rect 5206 3478 5240 3512
rect 5274 3478 5308 3512
rect 5342 3478 5376 3512
rect 5410 3478 5444 3512
rect 5478 3478 5512 3512
rect 5546 3478 5580 3512
rect 5614 3478 5648 3512
rect 5682 3478 5716 3512
rect 5750 3478 5784 3512
rect 5818 3478 5852 3512
rect 5886 3478 5920 3512
rect 5954 3478 5988 3512
rect 6022 3478 6056 3512
rect 6090 3478 6124 3512
rect 6158 3478 6192 3512
rect 5114 3410 5148 3444
<< mvnsubdiffcont >>
rect 3895 6601 3929 6635
rect 3963 6601 3997 6635
rect 4031 6601 4065 6635
rect 4099 6601 4133 6635
rect 4167 6601 4201 6635
rect 4235 6601 4269 6635
rect 4303 6601 4337 6635
rect 4371 6601 4405 6635
rect 4439 6601 4473 6635
rect 4507 6601 4541 6635
rect 4575 6601 4609 6635
rect 4643 6601 4677 6635
rect 4711 6601 4745 6635
rect 4779 6601 4813 6635
rect 4847 6601 4881 6635
rect 4915 6601 4949 6635
rect 4983 6601 5017 6635
rect 5051 6601 5085 6635
rect 5119 6601 5153 6635
rect 5187 6601 5221 6635
rect 5255 6601 5289 6635
rect 5323 6601 5357 6635
rect 5391 6601 5425 6635
rect 5459 6601 5493 6635
rect 5527 6601 5561 6635
rect 5595 6601 5629 6635
rect 5663 6601 5697 6635
rect 5731 6601 5765 6635
rect 5799 6601 5833 6635
rect 5867 6601 5901 6635
rect 5935 6601 5969 6635
rect 6003 6601 6037 6635
rect 6071 6601 6105 6635
rect 6139 6601 6173 6635
rect 4035 4436 4069 4470
rect 4103 4436 4137 4470
rect 4171 4436 4205 4470
rect 4239 4436 4273 4470
rect 4307 4436 4341 4470
rect 4375 4436 4409 4470
rect 4443 4436 4477 4470
rect 4511 4436 4545 4470
rect 4579 4436 4613 4470
rect 4647 4436 4681 4470
rect 4715 4436 4749 4470
rect 4783 4436 4817 4470
rect 4851 4436 4885 4470
rect 4919 4436 4953 4470
rect 4987 4436 5021 4470
rect 5055 4436 5089 4470
rect 5123 4436 5157 4470
rect 5230 4467 5264 4501
rect 5298 4467 5332 4501
rect 5366 4467 5400 4501
rect 5434 4467 5468 4501
rect 5502 4467 5536 4501
rect 5570 4467 5604 4501
rect 5638 4467 5672 4501
rect 5706 4467 5740 4501
rect 5774 4467 5808 4501
rect 5842 4467 5876 4501
rect 5910 4467 5944 4501
rect 5978 4467 6012 4501
rect 6046 4467 6080 4501
rect 6114 4467 6148 4501
<< locali >>
rect 3871 7582 3883 7616
rect 3929 7582 3955 7616
rect 3997 7582 4027 7616
rect 4065 7582 4099 7616
rect 4133 7582 4167 7616
rect 4205 7582 4235 7616
rect 4277 7582 4303 7616
rect 4349 7582 4371 7616
rect 4421 7582 4439 7616
rect 4493 7582 4507 7616
rect 4565 7582 4575 7616
rect 4637 7582 4643 7616
rect 4709 7582 4711 7616
rect 4745 7582 4747 7616
rect 4813 7582 4819 7616
rect 4881 7582 4891 7616
rect 4949 7582 4963 7616
rect 5017 7582 5035 7616
rect 5085 7582 5107 7616
rect 5153 7582 5179 7616
rect 5221 7582 5251 7616
rect 5289 7582 5323 7616
rect 5357 7582 5391 7616
rect 5429 7582 5459 7616
rect 5501 7582 5527 7616
rect 5573 7582 5595 7616
rect 5645 7582 5663 7616
rect 5717 7582 5731 7616
rect 5789 7582 5799 7616
rect 5861 7582 5867 7616
rect 5933 7582 5935 7616
rect 5969 7582 5971 7616
rect 6037 7582 6043 7616
rect 6105 7582 6115 7616
rect 6173 7582 6187 7616
rect 6221 7582 6233 7616
rect 3971 7230 4005 7268
rect 4443 7233 4477 7271
rect 4055 6982 4089 7020
rect 4124 6939 4190 7218
rect 4429 7199 4443 7218
rect 4612 7233 4646 7271
rect 4477 7199 4495 7218
rect 4600 7199 4612 7218
rect 4795 7237 4829 7275
rect 4646 7199 4666 7218
rect 4968 7237 5002 7275
rect 5445 7237 5479 7275
rect 4530 7085 4564 7123
rect 5257 7025 5323 7218
rect 5659 7095 5693 7133
rect 5730 7034 5796 7218
rect 5904 7167 5968 7218
rect 5904 7133 5917 7167
rect 5951 7133 5968 7167
rect 5904 7095 5968 7133
rect 5904 7061 5917 7095
rect 5951 7061 5968 7095
rect 5904 7043 5968 7061
rect 6089 7167 6151 7218
rect 6089 7133 6111 7167
rect 6145 7133 6151 7167
rect 6089 7095 6151 7133
rect 6089 7061 6111 7095
rect 6145 7061 6151 7095
rect 6089 7043 6151 7061
rect 4124 6905 4144 6939
rect 4178 6905 4190 6939
rect 4883 6953 4917 6991
rect 5257 6991 5267 7025
rect 5301 6991 5323 7025
rect 5257 6953 5323 6991
rect 5257 6921 5267 6953
rect 5301 6921 5323 6953
rect 5359 6955 5393 6993
rect 5730 7000 5743 7034
rect 5777 7000 5796 7034
rect 5730 6962 5796 7000
rect 5730 6928 5743 6962
rect 5777 6928 5796 6962
rect 4124 6867 4190 6905
rect 6011 6910 6045 6948
rect 4124 6833 4144 6867
rect 4178 6833 4190 6867
rect 4124 6831 4190 6833
rect 3871 6601 3883 6635
rect 3929 6601 3955 6635
rect 3997 6601 4027 6635
rect 4065 6601 4099 6635
rect 4133 6601 4167 6635
rect 4205 6601 4235 6635
rect 4277 6601 4303 6635
rect 4349 6601 4371 6635
rect 4421 6601 4439 6635
rect 4493 6601 4507 6635
rect 4565 6601 4575 6635
rect 4637 6601 4643 6635
rect 4709 6601 4711 6635
rect 4745 6601 4747 6635
rect 4813 6601 4819 6635
rect 4881 6601 4891 6635
rect 4949 6601 4963 6635
rect 5017 6601 5035 6635
rect 5085 6601 5107 6635
rect 5153 6601 5179 6635
rect 5221 6601 5251 6635
rect 5289 6601 5323 6635
rect 5357 6601 5391 6635
rect 5429 6601 5459 6635
rect 5501 6601 5527 6635
rect 5573 6601 5595 6635
rect 5645 6601 5663 6635
rect 5717 6601 5731 6635
rect 5789 6601 5799 6635
rect 5861 6601 5867 6635
rect 5933 6601 5935 6635
rect 5969 6601 5971 6635
rect 6037 6601 6043 6635
rect 6105 6601 6115 6635
rect 6173 6601 6229 6635
rect 4127 6337 4193 6341
rect 4127 6303 4140 6337
rect 4174 6303 4193 6337
rect 4127 6265 4193 6303
rect 4127 6231 4140 6265
rect 4174 6231 4193 6265
rect 5258 6330 5324 6348
rect 5258 6296 5274 6330
rect 5308 6296 5324 6330
rect 5258 6258 5324 6296
rect 6011 6308 6045 6346
rect 4055 6030 4089 6068
rect 4127 6018 4193 6231
rect 4430 6212 4439 6238
rect 4473 6212 4496 6238
rect 5258 6224 5274 6258
rect 5308 6224 5324 6258
rect 4430 6174 4496 6212
rect 4430 6140 4439 6174
rect 4473 6140 4496 6174
rect 4430 6018 4496 6140
rect 5007 6149 5041 6187
rect 5076 6109 5093 6143
rect 5127 6109 5142 6143
rect 5076 6071 5142 6109
rect 5076 6037 5093 6071
rect 5127 6037 5142 6071
rect 5076 6017 5142 6037
rect 5258 6018 5324 6224
rect 5903 6175 5968 6193
rect 5359 6071 5393 6109
rect 5659 6103 5693 6141
rect 5903 6141 5917 6175
rect 5951 6141 5968 6175
rect 5903 6103 5968 6141
rect 5903 6069 5917 6103
rect 5951 6069 5968 6103
rect 3962 5945 3996 5983
rect 3949 5911 3962 5917
rect 3996 5911 4015 5917
rect 3949 5898 4015 5911
rect 4615 5913 4649 5951
rect 4741 5956 4779 5990
rect 4813 5956 4865 5990
rect 4899 5956 4937 5990
rect 5903 6018 5968 6069
rect 6089 6175 6152 6193
rect 6089 6141 6111 6175
rect 6145 6141 6152 6175
rect 6089 6103 6152 6141
rect 6089 6069 6111 6103
rect 6145 6069 6152 6103
rect 6089 6018 6152 6069
rect 4707 5859 4741 5956
rect 5446 5915 5480 5953
rect 5737 5950 5771 5988
rect 3868 5620 3880 5654
rect 3926 5620 3952 5654
rect 3994 5620 4024 5654
rect 4062 5620 4096 5654
rect 4130 5620 4164 5654
rect 4202 5620 4232 5654
rect 4274 5620 4300 5654
rect 4346 5620 4368 5654
rect 4418 5620 4436 5654
rect 4490 5620 4504 5654
rect 4562 5620 4572 5654
rect 4634 5620 4640 5654
rect 4706 5620 4708 5654
rect 4742 5620 4744 5654
rect 4810 5620 4816 5654
rect 4878 5620 4888 5654
rect 4946 5620 4960 5654
rect 5014 5620 5032 5654
rect 5082 5620 5104 5654
rect 5150 5620 5176 5654
rect 5218 5620 5248 5654
rect 5286 5620 5320 5654
rect 5354 5620 5388 5654
rect 5426 5620 5456 5654
rect 5498 5620 5524 5654
rect 5570 5620 5592 5654
rect 5642 5620 5660 5654
rect 5714 5620 5728 5654
rect 5786 5620 5796 5654
rect 5858 5620 5864 5654
rect 5930 5620 5932 5654
rect 5966 5620 5968 5654
rect 6034 5620 6040 5654
rect 6102 5620 6112 5654
rect 6170 5620 6184 5654
rect 6218 5620 6254 5654
rect 5324 5581 6254 5620
rect 5324 5547 5336 5581
rect 5382 5547 5408 5581
rect 5450 5547 5480 5581
rect 5518 5547 5552 5581
rect 5586 5547 5620 5581
rect 5658 5547 5688 5581
rect 5730 5547 5756 5581
rect 5802 5547 5824 5581
rect 5874 5547 5892 5581
rect 5946 5547 5960 5581
rect 6018 5547 6028 5581
rect 6090 5547 6096 5581
rect 6162 5547 6164 5581
rect 6198 5547 6200 5581
rect 6234 5547 6254 5581
rect 5324 5507 6254 5547
rect 5324 5473 5336 5507
rect 5382 5473 5408 5507
rect 5450 5473 5480 5507
rect 5518 5473 5552 5507
rect 5586 5473 5620 5507
rect 5658 5473 5688 5507
rect 5730 5473 5756 5507
rect 5802 5473 5824 5507
rect 5874 5473 5892 5507
rect 5946 5473 5960 5507
rect 6018 5473 6028 5507
rect 6090 5473 6096 5507
rect 6162 5473 6164 5507
rect 6198 5473 6200 5507
rect 6234 5473 6254 5507
rect 4233 5283 4271 5317
rect 5421 5045 5487 5092
rect 5524 5084 5558 5122
rect 6088 5132 6122 5170
rect 5421 5011 5435 5045
rect 5469 5011 5487 5045
rect 4766 4905 4800 4943
rect 5421 4973 5487 5011
rect 5421 4939 5435 4973
rect 5469 4939 5487 4973
rect 5716 5041 5781 5092
rect 5716 5007 5725 5041
rect 5759 5007 5781 5041
rect 5716 4969 5781 5007
rect 5716 4935 5725 4969
rect 5759 4935 5781 4969
rect 5716 4917 5781 4935
rect 5902 5041 5966 5092
rect 5902 5007 5919 5041
rect 5953 5007 5966 5041
rect 5902 4969 5966 5007
rect 5902 4935 5919 4969
rect 5953 4935 5966 4969
rect 6177 4969 6211 5007
rect 5902 4917 5966 4935
rect 4463 4802 4501 4836
rect 5823 4762 5857 4800
rect 5194 4470 5230 4501
rect 3996 4436 4035 4470
rect 4089 4436 4103 4470
rect 4161 4436 4171 4470
rect 4233 4436 4239 4470
rect 4305 4436 4307 4470
rect 4341 4436 4343 4470
rect 4409 4436 4415 4470
rect 4477 4436 4487 4470
rect 4545 4436 4559 4470
rect 4613 4436 4631 4470
rect 4681 4436 4703 4470
rect 4749 4436 4775 4470
rect 4817 4436 4847 4470
rect 4885 4436 4919 4470
rect 4953 4436 4987 4470
rect 5025 4436 5055 4470
rect 5097 4436 5123 4470
rect 5169 4467 5230 4470
rect 5264 4467 5298 4501
rect 5336 4467 5366 4501
rect 5408 4467 5434 4501
rect 5480 4467 5502 4501
rect 5552 4467 5570 4501
rect 5624 4467 5638 4501
rect 5696 4467 5706 4501
rect 5768 4467 5774 4501
rect 5840 4467 5842 4501
rect 5876 4467 5878 4501
rect 5944 4467 5950 4501
rect 6012 4467 6022 4501
rect 6080 4467 6094 4501
rect 6148 4467 6218 4501
rect 5169 4436 5228 4467
rect 5323 4174 5357 4212
rect 6100 4212 6116 4246
rect 6150 4212 6166 4246
rect 6100 4174 6166 4212
rect 6100 4140 6116 4174
rect 6150 4140 6166 4174
rect 5744 4033 5808 4049
rect 5744 3999 5752 4033
rect 5786 3999 5808 4033
rect 4429 3935 4467 3969
rect 5744 3961 5808 3999
rect 4199 3884 4233 3922
rect 5744 3927 5752 3961
rect 5786 3927 5808 3961
rect 4736 3797 4770 3835
rect 5409 3805 5443 3843
rect 5744 3874 5808 3927
rect 5929 4031 5992 4049
rect 5929 3997 5946 4031
rect 5980 3997 5992 4031
rect 5929 3959 5992 3997
rect 5929 3925 5946 3959
rect 5980 3925 5992 3959
rect 5588 3804 5622 3842
rect 5929 3874 5992 3925
rect 6100 3876 6166 4140
rect 6204 3959 6238 3997
rect 5850 3813 5884 3851
rect 5114 3478 5126 3512
rect 5172 3478 5198 3512
rect 5240 3478 5270 3512
rect 5308 3478 5342 3512
rect 5376 3478 5410 3512
rect 5448 3478 5478 3512
rect 5520 3478 5546 3512
rect 5592 3478 5614 3512
rect 5664 3478 5682 3512
rect 5736 3478 5750 3512
rect 5808 3478 5818 3512
rect 5880 3478 5886 3512
rect 5952 3478 5954 3512
rect 5988 3478 5990 3512
rect 6056 3478 6062 3512
rect 6124 3478 6134 3512
rect 6192 3478 6206 3512
rect 6240 3478 6265 3512
rect 5114 3444 5148 3478
rect 5114 3384 5148 3410
rect -9024 2453 -9006 2487
rect -8972 2453 -8958 2487
rect -9024 2415 -8958 2453
rect -9024 2381 -9006 2415
rect -8972 2381 -8958 2415
rect -9202 2336 -9180 2343
rect -9146 2336 -9136 2343
rect -9024 2336 -8958 2381
rect -8845 2453 -8827 2487
rect -8793 2453 -8779 2487
rect -8845 2415 -8779 2453
rect -8744 2461 -8710 2499
rect -8845 2381 -8827 2415
rect -8793 2381 -8779 2415
rect -8845 2336 -8779 2381
rect -9180 2271 -9146 2309
rect -9096 2264 -9062 2302
rect -8649 2264 -8615 2302
<< viali >>
rect 3883 7582 3895 7616
rect 3895 7582 3917 7616
rect 3955 7582 3963 7616
rect 3963 7582 3989 7616
rect 4027 7582 4031 7616
rect 4031 7582 4061 7616
rect 4099 7582 4133 7616
rect 4171 7582 4201 7616
rect 4201 7582 4205 7616
rect 4243 7582 4269 7616
rect 4269 7582 4277 7616
rect 4315 7582 4337 7616
rect 4337 7582 4349 7616
rect 4387 7582 4405 7616
rect 4405 7582 4421 7616
rect 4459 7582 4473 7616
rect 4473 7582 4493 7616
rect 4531 7582 4541 7616
rect 4541 7582 4565 7616
rect 4603 7582 4609 7616
rect 4609 7582 4637 7616
rect 4675 7582 4677 7616
rect 4677 7582 4709 7616
rect 4747 7582 4779 7616
rect 4779 7582 4781 7616
rect 4819 7582 4847 7616
rect 4847 7582 4853 7616
rect 4891 7582 4915 7616
rect 4915 7582 4925 7616
rect 4963 7582 4983 7616
rect 4983 7582 4997 7616
rect 5035 7582 5051 7616
rect 5051 7582 5069 7616
rect 5107 7582 5119 7616
rect 5119 7582 5141 7616
rect 5179 7582 5187 7616
rect 5187 7582 5213 7616
rect 5251 7582 5255 7616
rect 5255 7582 5285 7616
rect 5323 7582 5357 7616
rect 5395 7582 5425 7616
rect 5425 7582 5429 7616
rect 5467 7582 5493 7616
rect 5493 7582 5501 7616
rect 5539 7582 5561 7616
rect 5561 7582 5573 7616
rect 5611 7582 5629 7616
rect 5629 7582 5645 7616
rect 5683 7582 5697 7616
rect 5697 7582 5717 7616
rect 5755 7582 5765 7616
rect 5765 7582 5789 7616
rect 5827 7582 5833 7616
rect 5833 7582 5861 7616
rect 5899 7582 5901 7616
rect 5901 7582 5933 7616
rect 5971 7582 6003 7616
rect 6003 7582 6005 7616
rect 6043 7582 6071 7616
rect 6071 7582 6077 7616
rect 6115 7582 6139 7616
rect 6139 7582 6149 7616
rect 6187 7582 6221 7616
rect 3971 7268 4005 7302
rect 3971 7196 4005 7230
rect 4443 7271 4477 7305
rect 4055 7020 4089 7054
rect 4055 6948 4089 6982
rect 4443 7199 4477 7233
rect 4612 7271 4646 7305
rect 4612 7199 4646 7233
rect 4795 7275 4829 7309
rect 4795 7203 4829 7237
rect 4968 7275 5002 7309
rect 4968 7203 5002 7237
rect 5445 7275 5479 7309
rect 4530 7123 4564 7157
rect 4530 7051 4564 7085
rect 5445 7203 5479 7237
rect 5659 7133 5693 7167
rect 5659 7061 5693 7095
rect 5917 7133 5951 7167
rect 5917 7061 5951 7095
rect 6111 7133 6145 7167
rect 6111 7061 6145 7095
rect 4144 6905 4178 6939
rect 4883 6991 4917 7025
rect 4883 6919 4917 6953
rect 5267 6991 5301 7025
rect 5267 6919 5301 6953
rect 5359 6993 5393 7027
rect 5359 6921 5393 6955
rect 5743 7000 5777 7034
rect 5743 6928 5777 6962
rect 6011 6948 6045 6982
rect 6011 6876 6045 6910
rect 4144 6833 4178 6867
rect 3883 6601 3895 6635
rect 3895 6601 3917 6635
rect 3955 6601 3963 6635
rect 3963 6601 3989 6635
rect 4027 6601 4031 6635
rect 4031 6601 4061 6635
rect 4099 6601 4133 6635
rect 4171 6601 4201 6635
rect 4201 6601 4205 6635
rect 4243 6601 4269 6635
rect 4269 6601 4277 6635
rect 4315 6601 4337 6635
rect 4337 6601 4349 6635
rect 4387 6601 4405 6635
rect 4405 6601 4421 6635
rect 4459 6601 4473 6635
rect 4473 6601 4493 6635
rect 4531 6601 4541 6635
rect 4541 6601 4565 6635
rect 4603 6601 4609 6635
rect 4609 6601 4637 6635
rect 4675 6601 4677 6635
rect 4677 6601 4709 6635
rect 4747 6601 4779 6635
rect 4779 6601 4781 6635
rect 4819 6601 4847 6635
rect 4847 6601 4853 6635
rect 4891 6601 4915 6635
rect 4915 6601 4925 6635
rect 4963 6601 4983 6635
rect 4983 6601 4997 6635
rect 5035 6601 5051 6635
rect 5051 6601 5069 6635
rect 5107 6601 5119 6635
rect 5119 6601 5141 6635
rect 5179 6601 5187 6635
rect 5187 6601 5213 6635
rect 5251 6601 5255 6635
rect 5255 6601 5285 6635
rect 5323 6601 5357 6635
rect 5395 6601 5425 6635
rect 5425 6601 5429 6635
rect 5467 6601 5493 6635
rect 5493 6601 5501 6635
rect 5539 6601 5561 6635
rect 5561 6601 5573 6635
rect 5611 6601 5629 6635
rect 5629 6601 5645 6635
rect 5683 6601 5697 6635
rect 5697 6601 5717 6635
rect 5755 6601 5765 6635
rect 5765 6601 5789 6635
rect 5827 6601 5833 6635
rect 5833 6601 5861 6635
rect 5899 6601 5901 6635
rect 5901 6601 5933 6635
rect 5971 6601 6003 6635
rect 6003 6601 6005 6635
rect 6043 6601 6071 6635
rect 6071 6601 6077 6635
rect 6115 6601 6139 6635
rect 6139 6601 6149 6635
rect 4140 6303 4174 6337
rect 4140 6231 4174 6265
rect 5274 6296 5308 6330
rect 6011 6346 6045 6380
rect 6011 6274 6045 6308
rect 4055 6068 4089 6102
rect 3962 5983 3996 6017
rect 4055 5996 4089 6030
rect 4439 6212 4473 6246
rect 5274 6224 5308 6258
rect 4439 6140 4473 6174
rect 5007 6187 5041 6221
rect 5007 6115 5041 6149
rect 5093 6109 5127 6143
rect 5093 6037 5127 6071
rect 5359 6109 5393 6143
rect 5359 6037 5393 6071
rect 5659 6141 5693 6175
rect 5659 6069 5693 6103
rect 5917 6141 5951 6175
rect 5917 6069 5951 6103
rect 3962 5911 3996 5945
rect 4615 5951 4649 5985
rect 4615 5879 4649 5913
rect 4707 5956 4741 5990
rect 4779 5956 4813 5990
rect 4865 5956 4899 5990
rect 4937 5956 4971 5990
rect 5737 5988 5771 6022
rect 6111 6141 6145 6175
rect 6111 6069 6145 6103
rect 5446 5953 5480 5987
rect 5737 5916 5771 5950
rect 5446 5881 5480 5915
rect 3880 5620 3892 5654
rect 3892 5620 3914 5654
rect 3952 5620 3960 5654
rect 3960 5620 3986 5654
rect 4024 5620 4028 5654
rect 4028 5620 4058 5654
rect 4096 5620 4130 5654
rect 4168 5620 4198 5654
rect 4198 5620 4202 5654
rect 4240 5620 4266 5654
rect 4266 5620 4274 5654
rect 4312 5620 4334 5654
rect 4334 5620 4346 5654
rect 4384 5620 4402 5654
rect 4402 5620 4418 5654
rect 4456 5620 4470 5654
rect 4470 5620 4490 5654
rect 4528 5620 4538 5654
rect 4538 5620 4562 5654
rect 4600 5620 4606 5654
rect 4606 5620 4634 5654
rect 4672 5620 4674 5654
rect 4674 5620 4706 5654
rect 4744 5620 4776 5654
rect 4776 5620 4778 5654
rect 4816 5620 4844 5654
rect 4844 5620 4850 5654
rect 4888 5620 4912 5654
rect 4912 5620 4922 5654
rect 4960 5620 4980 5654
rect 4980 5620 4994 5654
rect 5032 5620 5048 5654
rect 5048 5620 5066 5654
rect 5104 5620 5116 5654
rect 5116 5620 5138 5654
rect 5176 5620 5184 5654
rect 5184 5620 5210 5654
rect 5248 5620 5252 5654
rect 5252 5620 5282 5654
rect 5320 5620 5354 5654
rect 5392 5620 5422 5654
rect 5422 5620 5426 5654
rect 5464 5620 5490 5654
rect 5490 5620 5498 5654
rect 5536 5620 5558 5654
rect 5558 5620 5570 5654
rect 5608 5620 5626 5654
rect 5626 5620 5642 5654
rect 5680 5620 5694 5654
rect 5694 5620 5714 5654
rect 5752 5620 5762 5654
rect 5762 5620 5786 5654
rect 5824 5620 5830 5654
rect 5830 5620 5858 5654
rect 5896 5620 5898 5654
rect 5898 5620 5930 5654
rect 5968 5620 6000 5654
rect 6000 5620 6002 5654
rect 6040 5620 6068 5654
rect 6068 5620 6074 5654
rect 6112 5620 6136 5654
rect 6136 5620 6146 5654
rect 6184 5620 6218 5654
rect 5336 5547 5348 5581
rect 5348 5547 5370 5581
rect 5408 5547 5416 5581
rect 5416 5547 5442 5581
rect 5480 5547 5484 5581
rect 5484 5547 5514 5581
rect 5552 5547 5586 5581
rect 5624 5547 5654 5581
rect 5654 5547 5658 5581
rect 5696 5547 5722 5581
rect 5722 5547 5730 5581
rect 5768 5547 5790 5581
rect 5790 5547 5802 5581
rect 5840 5547 5858 5581
rect 5858 5547 5874 5581
rect 5912 5547 5926 5581
rect 5926 5547 5946 5581
rect 5984 5547 5994 5581
rect 5994 5547 6018 5581
rect 6056 5547 6062 5581
rect 6062 5547 6090 5581
rect 6128 5547 6130 5581
rect 6130 5547 6162 5581
rect 6200 5547 6234 5581
rect 5336 5473 5348 5507
rect 5348 5473 5370 5507
rect 5408 5473 5416 5507
rect 5416 5473 5442 5507
rect 5480 5473 5484 5507
rect 5484 5473 5514 5507
rect 5552 5473 5586 5507
rect 5624 5473 5654 5507
rect 5654 5473 5658 5507
rect 5696 5473 5722 5507
rect 5722 5473 5730 5507
rect 5768 5473 5790 5507
rect 5790 5473 5802 5507
rect 5840 5473 5858 5507
rect 5858 5473 5874 5507
rect 5912 5473 5926 5507
rect 5926 5473 5946 5507
rect 5984 5473 5994 5507
rect 5994 5473 6018 5507
rect 6056 5473 6062 5507
rect 6062 5473 6090 5507
rect 6128 5473 6130 5507
rect 6130 5473 6162 5507
rect 6200 5473 6234 5507
rect 4199 5283 4233 5317
rect 4271 5283 4305 5317
rect 6088 5170 6122 5204
rect 5524 5122 5558 5156
rect 6088 5098 6122 5132
rect 5524 5050 5558 5084
rect 5435 5011 5469 5045
rect 4766 4943 4800 4977
rect 5435 4939 5469 4973
rect 5725 5007 5759 5041
rect 5725 4935 5759 4969
rect 5919 5007 5953 5041
rect 5919 4935 5953 4969
rect 6177 5007 6211 5041
rect 6177 4935 6211 4969
rect 4766 4871 4800 4905
rect 4429 4802 4463 4836
rect 4501 4802 4535 4836
rect 5823 4800 5857 4834
rect 5823 4728 5857 4762
rect 4055 4436 4069 4470
rect 4069 4436 4089 4470
rect 4127 4436 4137 4470
rect 4137 4436 4161 4470
rect 4199 4436 4205 4470
rect 4205 4436 4233 4470
rect 4271 4436 4273 4470
rect 4273 4436 4305 4470
rect 4343 4436 4375 4470
rect 4375 4436 4377 4470
rect 4415 4436 4443 4470
rect 4443 4436 4449 4470
rect 4487 4436 4511 4470
rect 4511 4436 4521 4470
rect 4559 4436 4579 4470
rect 4579 4436 4593 4470
rect 4631 4436 4647 4470
rect 4647 4436 4665 4470
rect 4703 4436 4715 4470
rect 4715 4436 4737 4470
rect 4775 4436 4783 4470
rect 4783 4436 4809 4470
rect 4847 4436 4851 4470
rect 4851 4436 4881 4470
rect 4919 4436 4953 4470
rect 4991 4436 5021 4470
rect 5021 4436 5025 4470
rect 5063 4436 5089 4470
rect 5089 4436 5097 4470
rect 5135 4436 5157 4470
rect 5157 4436 5169 4470
rect 5230 4467 5264 4501
rect 5302 4467 5332 4501
rect 5332 4467 5336 4501
rect 5374 4467 5400 4501
rect 5400 4467 5408 4501
rect 5446 4467 5468 4501
rect 5468 4467 5480 4501
rect 5518 4467 5536 4501
rect 5536 4467 5552 4501
rect 5590 4467 5604 4501
rect 5604 4467 5624 4501
rect 5662 4467 5672 4501
rect 5672 4467 5696 4501
rect 5734 4467 5740 4501
rect 5740 4467 5768 4501
rect 5806 4467 5808 4501
rect 5808 4467 5840 4501
rect 5878 4467 5910 4501
rect 5910 4467 5912 4501
rect 5950 4467 5978 4501
rect 5978 4467 5984 4501
rect 6022 4467 6046 4501
rect 6046 4467 6056 4501
rect 6094 4467 6114 4501
rect 6114 4467 6128 4501
rect 5323 4212 5357 4246
rect 5323 4140 5357 4174
rect 6116 4212 6150 4246
rect 6116 4140 6150 4174
rect 5752 3999 5786 4033
rect 4199 3922 4233 3956
rect 4395 3935 4429 3969
rect 4467 3935 4501 3969
rect 4199 3850 4233 3884
rect 5752 3927 5786 3961
rect 4736 3835 4770 3869
rect 4736 3763 4770 3797
rect 5409 3843 5443 3877
rect 5409 3771 5443 3805
rect 5588 3842 5622 3876
rect 5946 3997 5980 4031
rect 5946 3925 5980 3959
rect 5588 3770 5622 3804
rect 5850 3851 5884 3885
rect 6204 3997 6238 4031
rect 6204 3925 6238 3959
rect 5850 3779 5884 3813
rect 5126 3478 5138 3512
rect 5138 3478 5160 3512
rect 5198 3478 5206 3512
rect 5206 3478 5232 3512
rect 5270 3478 5274 3512
rect 5274 3478 5304 3512
rect 5342 3478 5376 3512
rect 5414 3478 5444 3512
rect 5444 3478 5448 3512
rect 5486 3478 5512 3512
rect 5512 3478 5520 3512
rect 5558 3478 5580 3512
rect 5580 3478 5592 3512
rect 5630 3478 5648 3512
rect 5648 3478 5664 3512
rect 5702 3478 5716 3512
rect 5716 3478 5736 3512
rect 5774 3478 5784 3512
rect 5784 3478 5808 3512
rect 5846 3478 5852 3512
rect 5852 3478 5880 3512
rect 5918 3478 5920 3512
rect 5920 3478 5952 3512
rect 5990 3478 6022 3512
rect 6022 3478 6024 3512
rect 6062 3478 6090 3512
rect 6090 3478 6096 3512
rect 6134 3478 6158 3512
rect 6158 3478 6168 3512
rect 6206 3478 6240 3512
rect -8744 2499 -8710 2533
rect -9006 2453 -8972 2487
rect -9006 2381 -8972 2415
rect -9180 2309 -9146 2343
rect -8827 2453 -8793 2487
rect -8744 2427 -8710 2461
rect -8827 2381 -8793 2415
rect -9180 2237 -9146 2271
rect -9096 2302 -9062 2336
rect -9096 2230 -9062 2264
rect -8649 2302 -8615 2336
rect -8649 2230 -8615 2264
<< metal1 >>
rect 3836 7623 6233 7628
rect 3836 7616 5099 7623
rect 3836 7582 3883 7616
rect 3917 7582 3955 7616
rect 3989 7582 4027 7616
rect 4061 7582 4099 7616
rect 4133 7582 4171 7616
rect 4205 7582 4243 7616
rect 4277 7582 4315 7616
rect 4349 7582 4387 7616
rect 4421 7582 4459 7616
rect 4493 7582 4531 7616
rect 4565 7582 4603 7616
rect 4637 7582 4675 7616
rect 4709 7582 4747 7616
rect 4781 7582 4819 7616
rect 4853 7582 4891 7616
rect 4925 7582 4963 7616
rect 4997 7582 5035 7616
rect 5069 7582 5099 7616
rect 3836 7571 5099 7582
rect 5151 7571 5178 7623
rect 5230 7616 5256 7623
rect 5308 7616 6233 7623
rect 5230 7582 5251 7616
rect 5308 7582 5323 7616
rect 5357 7582 5395 7616
rect 5429 7582 5467 7616
rect 5501 7582 5539 7616
rect 5573 7582 5611 7616
rect 5645 7582 5683 7616
rect 5717 7582 5755 7616
rect 5789 7582 5827 7616
rect 5861 7582 5899 7616
rect 5933 7582 5971 7616
rect 6005 7582 6043 7616
rect 6077 7582 6115 7616
rect 6149 7582 6187 7616
rect 6221 7582 6233 7616
rect 5230 7571 5256 7582
rect 5308 7571 6233 7582
rect 3836 7544 6233 7571
rect 3836 7492 5099 7544
rect 5151 7492 5178 7544
rect 5230 7492 5256 7544
rect 5308 7492 6233 7544
rect 3836 7465 6233 7492
rect 3836 7413 5099 7465
rect 5151 7413 5178 7465
rect 5230 7413 5256 7465
rect 5308 7413 6233 7465
rect 3836 7412 6233 7413
rect 3965 7302 4011 7314
rect 3965 7268 3971 7302
rect 4005 7268 4011 7302
rect 3965 7230 4011 7268
rect 3965 7196 3971 7230
rect 4005 7196 4011 7230
rect 3965 7184 4011 7196
rect 4434 7312 4486 7318
rect 4434 7245 4486 7260
rect 4434 7187 4486 7193
rect 4603 7312 4655 7318
rect 4603 7245 4655 7260
rect 4603 7187 4655 7193
rect 4786 7316 4838 7322
rect 4786 7249 4838 7264
rect 4786 7191 4838 7197
rect 4959 7316 5011 7322
rect 4959 7249 5011 7264
rect 4959 7191 5011 7197
rect 5436 7316 5488 7322
rect 5436 7249 5488 7264
rect 5436 7191 5488 7197
rect 5579 7246 5659 7298
rect 5711 7246 5723 7298
rect 5775 7246 5781 7298
tri 5575 7187 5579 7191 se
rect 5579 7187 5613 7246
tri 5613 7212 5647 7246 nw
tri 5572 7184 5575 7187 se
rect 5575 7184 5613 7187
tri 5567 7179 5572 7184 se
rect 5572 7179 5613 7184
tri 5557 7169 5567 7179 se
rect 5567 7169 5613 7179
rect 4524 7167 4570 7169
tri 4570 7167 4572 7169 sw
tri 5555 7167 5557 7169 se
rect 5557 7167 5613 7169
rect 4524 7157 4572 7167
tri 4572 7157 4582 7167 sw
tri 5545 7157 5555 7167 se
rect 5555 7157 5613 7167
rect 4524 7123 4530 7157
rect 4564 7123 5613 7157
rect 5653 7167 5699 7179
tri 5699 7167 5706 7174 sw
tri 5904 7167 5911 7174 se
rect 5911 7167 5957 7179
tri 5957 7167 5964 7174 sw
tri 6098 7167 6105 7174 se
rect 6105 7167 6151 7179
rect 5653 7133 5659 7167
rect 5693 7140 5706 7167
tri 5706 7140 5733 7167 sw
tri 5877 7140 5904 7167 se
rect 5904 7140 5917 7167
rect 5693 7133 5917 7140
rect 5951 7140 5964 7167
tri 5964 7140 5991 7167 sw
tri 6071 7140 6098 7167 se
rect 6098 7140 6111 7167
rect 5951 7133 6111 7140
rect 6145 7133 6151 7167
rect 4524 7095 4576 7123
tri 4576 7095 4604 7123 nw
rect 5653 7095 6151 7133
rect 4524 7085 4570 7095
tri 4570 7089 4576 7095 nw
rect 4049 7054 4095 7066
rect 4049 7020 4055 7054
rect 4089 7039 4095 7054
rect 4524 7051 4530 7085
rect 4564 7051 4570 7085
tri 4095 7039 4106 7050 sw
rect 4524 7039 4570 7051
rect 4794 7067 5442 7095
rect 4794 7061 4856 7067
tri 4856 7061 4862 7067 nw
tri 5412 7061 5418 7067 ne
rect 5418 7061 5442 7067
rect 4794 7045 4840 7061
tri 4840 7045 4856 7061 nw
tri 5418 7045 5434 7061 ne
rect 5434 7045 5442 7061
tri 4792 7043 4794 7045 se
rect 4794 7043 4838 7045
tri 4838 7043 4840 7045 nw
tri 5434 7043 5436 7045 ne
rect 5436 7043 5442 7045
rect 5494 7043 5506 7095
rect 5558 7043 5564 7095
rect 5653 7061 5659 7095
rect 5693 7076 5917 7095
rect 5693 7061 5711 7076
tri 5711 7061 5726 7076 nw
tri 5884 7061 5899 7076 ne
rect 5899 7061 5917 7076
rect 5951 7076 6111 7095
rect 5951 7061 5969 7076
tri 5969 7061 5984 7076 nw
tri 6078 7061 6093 7076 ne
rect 6093 7061 6111 7076
rect 6145 7061 6151 7095
rect 5653 7049 5699 7061
tri 5699 7049 5711 7061 nw
tri 5899 7049 5911 7061 ne
rect 5911 7049 5957 7061
tri 5957 7049 5969 7061 nw
tri 6093 7049 6105 7061 ne
rect 6105 7049 6151 7061
tri 4788 7039 4792 7043 se
rect 4792 7039 4834 7043
tri 4834 7039 4838 7043 nw
rect 4089 7037 4106 7039
tri 4106 7037 4108 7039 sw
tri 4786 7037 4788 7039 se
rect 4788 7037 4832 7039
tri 4832 7037 4834 7039 nw
rect 4089 7034 4108 7037
tri 4108 7034 4111 7037 sw
tri 4783 7034 4786 7037 se
rect 4786 7034 4829 7037
tri 4829 7034 4832 7037 nw
rect 4089 7027 4111 7034
tri 4111 7027 4118 7034 sw
tri 4776 7027 4783 7034 se
rect 4783 7027 4828 7034
tri 4828 7033 4829 7034 nw
rect 4089 7025 4118 7027
tri 4118 7025 4120 7027 sw
tri 4774 7025 4776 7027 se
rect 4776 7025 4828 7027
rect 4089 7020 4120 7025
rect 4049 7016 4120 7020
tri 4120 7016 4129 7025 sw
tri 4765 7016 4774 7025 se
rect 4774 7016 4828 7025
rect 4049 7011 4414 7016
tri 4414 7011 4419 7016 sw
tri 4760 7011 4765 7016 se
rect 4765 7011 4828 7016
rect 4049 6982 4828 7011
rect 4049 6948 4055 6982
rect 4089 6962 4107 6982
tri 4107 6962 4127 6982 nw
tri 4358 6977 4363 6982 ne
rect 4363 6977 4828 6982
rect 4877 7025 5307 7037
rect 4877 6991 4883 7025
rect 4917 6992 5267 7025
rect 4917 6991 4957 6992
tri 4957 6991 4958 6992 nw
tri 5226 6991 5227 6992 ne
rect 5227 6991 5267 6992
rect 5301 6991 5307 7025
rect 4877 6982 4948 6991
tri 4948 6982 4957 6991 nw
tri 5227 6982 5236 6991 ne
rect 5236 6982 5307 6991
rect 4877 6962 4928 6982
tri 4928 6962 4948 6982 nw
tri 5236 6964 5254 6982 ne
rect 5254 6964 5307 6982
rect 4089 6955 4100 6962
tri 4100 6955 4107 6962 nw
rect 4089 6953 4098 6955
tri 4098 6953 4100 6955 nw
rect 4877 6953 4923 6962
tri 4923 6957 4928 6962 nw
rect 5002 6958 5054 6964
tri 5254 6962 5256 6964 ne
rect 5256 6962 5307 6964
rect 4089 6951 4096 6953
tri 4096 6951 4098 6953 nw
rect 4089 6948 4095 6951
tri 4095 6950 4096 6951 nw
rect 4049 6936 4095 6948
rect 4138 6939 4184 6951
rect 4138 6905 4144 6939
rect 4178 6910 4184 6939
rect 4877 6919 4883 6953
rect 4917 6919 4923 6953
tri 4184 6910 4187 6913 sw
rect 4178 6907 4187 6910
tri 4187 6907 4190 6910 sw
rect 4877 6907 4923 6919
tri 4999 6910 5002 6913 se
tri 4996 6907 4999 6910 se
rect 4999 6907 5002 6910
rect 4178 6905 4190 6907
rect 4138 6879 4190 6905
tri 4190 6879 4218 6907 sw
tri 4968 6879 4996 6907 se
rect 4996 6906 5002 6907
tri 5256 6957 5261 6962 ne
rect 5261 6953 5307 6962
rect 5261 6919 5267 6953
rect 5301 6919 5307 6953
rect 5261 6907 5307 6919
rect 5353 7034 5399 7039
tri 5399 7034 5403 7038 sw
tri 5733 7034 5737 7038 se
rect 5737 7034 5783 7046
rect 5353 7027 5403 7034
rect 5353 6993 5359 7027
rect 5393 7004 5403 7027
tri 5403 7004 5433 7034 sw
tri 5703 7004 5733 7034 se
rect 5733 7004 5743 7034
rect 5393 7000 5743 7004
rect 5777 7000 5783 7034
rect 5393 6993 5783 7000
rect 5353 6962 5783 6993
rect 5353 6958 5743 6962
rect 5353 6955 5403 6958
rect 5353 6921 5359 6955
rect 5393 6928 5403 6955
tri 5403 6928 5433 6958 nw
tri 5695 6928 5725 6958 ne
rect 5725 6928 5743 6958
rect 5777 6928 5783 6962
rect 5393 6921 5399 6928
tri 5399 6924 5403 6928 nw
tri 5725 6924 5729 6928 ne
rect 5729 6924 5783 6928
rect 5353 6909 5399 6921
tri 5729 6916 5737 6924 ne
rect 5737 6916 5783 6924
rect 6005 6982 6051 6994
rect 6005 6948 6011 6982
rect 6045 6948 6051 6982
rect 6005 6910 6051 6948
rect 4996 6894 5054 6906
rect 4996 6879 5002 6894
rect 4138 6867 5002 6879
rect 4138 6833 4144 6867
rect 4178 6842 5002 6867
rect 6005 6876 6011 6910
rect 6045 6876 6051 6910
rect 6005 6864 6051 6876
rect 4178 6836 5054 6842
rect 4178 6833 4184 6836
rect 4138 6821 4184 6833
tri 4184 6821 4199 6836 nw
rect 4277 6647 6233 6793
rect 3871 6635 6233 6647
rect 3871 6601 3883 6635
rect 3917 6601 3955 6635
rect 3989 6601 4027 6635
rect 4061 6601 4099 6635
rect 4133 6601 4171 6635
rect 4205 6601 4243 6635
rect 4277 6601 4315 6635
rect 4349 6601 4387 6635
rect 4421 6601 4459 6635
rect 4493 6601 4531 6635
rect 4565 6601 4603 6635
rect 4637 6601 4675 6635
rect 4709 6601 4747 6635
rect 4781 6601 4819 6635
rect 4853 6601 4891 6635
rect 4925 6601 4963 6635
rect 4997 6601 5035 6635
rect 5069 6601 5107 6635
rect 5141 6601 5179 6635
rect 5213 6601 5251 6635
rect 5285 6601 5323 6635
rect 5357 6601 5395 6635
rect 5429 6601 5467 6635
rect 5501 6601 5539 6635
rect 5573 6601 5611 6635
rect 5645 6601 5683 6635
rect 5717 6601 5755 6635
rect 5789 6601 5827 6635
rect 5861 6601 5899 6635
rect 5933 6601 5971 6635
rect 6005 6601 6043 6635
rect 6077 6601 6115 6635
rect 6149 6601 6233 6635
tri 3836 6559 3867 6590 ne
rect 3871 6589 6233 6601
rect 4277 6443 6233 6589
rect 6005 6380 6051 6392
rect 4134 6346 4180 6349
tri 4180 6346 4183 6349 sw
rect 6005 6346 6011 6380
rect 6045 6346 6051 6380
rect 4134 6340 4183 6346
tri 4183 6340 4189 6346 sw
tri 5266 6340 5268 6342 se
rect 5268 6340 5314 6342
rect 4134 6337 4564 6340
rect 4134 6303 4140 6337
rect 4174 6303 4564 6337
tri 5262 6336 5266 6340 se
rect 5266 6336 5314 6340
rect 4134 6294 4564 6303
rect 4134 6274 4194 6294
tri 4194 6274 4214 6294 nw
tri 4484 6274 4504 6294 ne
rect 4504 6274 4564 6294
rect 4134 6265 4182 6274
rect 4134 6231 4140 6265
rect 4174 6262 4182 6265
tri 4182 6262 4194 6274 nw
tri 4504 6262 4516 6274 ne
rect 4516 6262 4564 6274
rect 4174 6231 4180 6262
tri 4180 6260 4182 6262 nw
tri 4516 6260 4518 6262 ne
rect 4134 6219 4180 6231
rect 4433 6246 4479 6258
rect 4433 6212 4439 6246
rect 4473 6212 4479 6246
tri 4412 6187 4433 6208 se
rect 4433 6187 4479 6212
tri 4400 6175 4412 6187 se
rect 4412 6175 4479 6187
tri 4399 6174 4400 6175 se
rect 4400 6174 4479 6175
rect 4049 6140 4439 6174
rect 4473 6140 4479 6174
rect 4049 6128 4479 6140
rect 4518 6208 4564 6262
rect 4695 6330 5314 6336
rect 4747 6296 5274 6330
rect 5308 6296 5314 6330
rect 4747 6284 5314 6296
rect 4747 6278 4771 6284
rect 4695 6274 4771 6278
tri 4771 6274 4781 6284 nw
tri 5234 6274 5244 6284 ne
rect 5244 6274 5314 6284
rect 4695 6266 4759 6274
rect 4747 6262 4759 6266
tri 4759 6262 4771 6274 nw
tri 5244 6262 5256 6274 ne
rect 5256 6262 5314 6274
rect 6005 6308 6051 6346
rect 6005 6274 6011 6308
rect 6045 6274 6051 6308
rect 6005 6262 6051 6274
rect 4747 6258 4755 6262
tri 4755 6258 4759 6262 nw
tri 5256 6258 5260 6262 ne
rect 5260 6258 5314 6262
tri 4747 6250 4755 6258 nw
tri 5260 6250 5268 6258 ne
tri 4564 6208 4570 6214 sw
rect 4695 6208 4747 6214
rect 4786 6240 4838 6246
rect 4518 6206 4570 6208
tri 4570 6206 4572 6208 sw
rect 4518 6187 4572 6206
tri 4572 6187 4591 6206 sw
tri 4767 6187 4786 6206 se
rect 4786 6187 4838 6188
rect 4518 6180 4591 6187
tri 4591 6180 4598 6187 sw
tri 4760 6180 4767 6187 se
rect 4767 6180 4838 6187
rect 4518 6176 4838 6180
rect 4518 6134 4786 6176
tri 4770 6128 4776 6134 ne
rect 4776 6128 4786 6134
rect 4049 6115 4116 6128
tri 4116 6115 4129 6128 nw
tri 4776 6118 4786 6128 ne
rect 4786 6118 4838 6124
rect 5001 6227 5054 6233
rect 5001 6175 5002 6227
rect 5268 6224 5274 6258
rect 5308 6224 5314 6258
rect 5268 6212 5314 6224
rect 5001 6161 5054 6175
rect 4049 6109 4110 6115
tri 4110 6109 4116 6115 nw
rect 5001 6109 5002 6161
rect 5653 6175 5699 6187
tri 5699 6175 5711 6187 sw
tri 5899 6175 5911 6187 se
rect 5911 6175 5957 6187
tri 5957 6175 5969 6187 sw
tri 6093 6175 6105 6187 se
rect 6105 6175 6151 6187
rect 4049 6103 4104 6109
tri 4104 6103 4110 6109 nw
rect 5001 6103 5054 6109
rect 5087 6143 5133 6155
tri 5133 6143 5137 6147 sw
tri 5349 6143 5353 6147 se
rect 5353 6143 5399 6155
rect 5087 6109 5093 6143
rect 5127 6113 5137 6143
tri 5137 6113 5167 6143 sw
tri 5319 6113 5349 6143 se
rect 5349 6113 5359 6143
rect 5127 6109 5359 6113
rect 5393 6109 5399 6143
rect 4049 6102 4095 6103
rect 4049 6068 4055 6102
rect 4089 6068 4095 6102
tri 4095 6094 4104 6103 nw
rect 4049 6030 4095 6068
rect 3956 6017 4002 6029
rect 3956 5983 3962 6017
rect 3996 5983 4002 6017
rect 4049 5996 4055 6030
rect 4089 5996 4095 6030
rect 4049 5984 4095 5996
rect 4176 6030 4821 6076
rect 4176 6022 4261 6030
tri 4261 6022 4269 6030 nw
tri 4791 6024 4797 6030 ne
rect 4797 6024 4821 6030
rect 4873 6024 4885 6076
rect 4937 6024 4943 6076
rect 5087 6071 5399 6109
rect 5087 6037 5093 6071
rect 5127 6067 5359 6071
rect 5127 6037 5137 6067
tri 5137 6037 5167 6067 nw
tri 5319 6037 5349 6067 ne
rect 5349 6037 5359 6067
rect 5393 6037 5399 6071
rect 5653 6141 5659 6175
rect 5693 6160 5711 6175
tri 5711 6160 5726 6175 sw
tri 5884 6160 5899 6175 se
rect 5899 6160 5917 6175
rect 5693 6141 5917 6160
rect 5951 6160 5969 6175
tri 5969 6160 5984 6175 sw
tri 6078 6160 6093 6175 se
rect 6093 6160 6111 6175
rect 5951 6141 6111 6160
rect 6145 6141 6151 6175
rect 5653 6103 6151 6141
rect 5653 6069 5659 6103
rect 5693 6096 5917 6103
rect 5693 6069 5706 6096
tri 5706 6069 5733 6096 nw
tri 5877 6069 5904 6096 ne
rect 5904 6069 5917 6096
rect 5951 6096 6111 6103
rect 5951 6069 5964 6096
tri 5964 6069 5991 6096 nw
tri 6071 6069 6098 6096 ne
rect 6098 6069 6111 6096
rect 6145 6069 6151 6103
rect 5653 6057 5699 6069
tri 5699 6062 5706 6069 nw
tri 5904 6062 5911 6069 ne
rect 5911 6057 5957 6069
tri 5957 6062 5964 6069 nw
tri 6098 6062 6105 6069 ne
rect 6105 6057 6151 6069
rect 5087 6025 5133 6037
tri 5133 6033 5137 6037 nw
tri 5349 6033 5353 6037 ne
rect 5353 6025 5399 6037
rect 5729 6033 5781 6039
rect 4176 5997 4236 6022
tri 4236 5997 4261 6022 nw
rect 3956 5951 4002 5983
tri 4002 5951 4030 5979 sw
tri 4148 5951 4176 5979 se
rect 4176 5951 4235 5997
tri 4235 5996 4236 5997 nw
rect 3956 5950 4030 5951
tri 4030 5950 4031 5951 sw
tri 4147 5950 4148 5951 se
rect 4148 5950 4235 5951
rect 3956 5945 4031 5950
tri 4031 5945 4036 5950 sw
tri 4142 5945 4147 5950 se
rect 4147 5945 4235 5950
rect 3956 5911 3962 5945
rect 3996 5911 4235 5945
rect 3956 5899 4235 5911
rect 4519 5991 4655 5997
rect 4571 5985 4655 5991
rect 4571 5951 4615 5985
rect 4649 5951 4655 5985
rect 4571 5939 4655 5951
rect 4695 5990 4983 5996
rect 4695 5956 4707 5990
rect 4741 5956 4779 5990
rect 4813 5956 4865 5990
rect 4899 5956 4937 5990
rect 4971 5956 4983 5990
rect 5440 5993 5572 5999
rect 5440 5987 5520 5993
rect 5356 5976 5408 5982
rect 4695 5950 4983 5956
tri 5347 5953 5356 5962 se
tri 5344 5950 5347 5953 se
rect 5347 5950 5356 5953
rect 4519 5925 4655 5939
rect 4571 5922 4655 5925
tri 4655 5922 4683 5950 sw
tri 5316 5922 5344 5950 se
rect 5344 5924 5356 5950
rect 5344 5922 5408 5924
rect 4571 5913 5408 5922
rect 4571 5879 4615 5913
rect 4649 5912 5408 5913
rect 4649 5879 5356 5912
rect 4571 5876 5356 5879
rect 4571 5873 4659 5876
rect 4519 5871 4659 5873
tri 4659 5871 4664 5876 nw
tri 5334 5871 5339 5876 ne
rect 5339 5871 5356 5876
rect 4519 5867 4655 5871
tri 4655 5867 4659 5871 nw
tri 5339 5867 5343 5871 ne
rect 5343 5867 5356 5871
tri 5343 5854 5356 5867 ne
rect 5440 5953 5446 5987
rect 5480 5953 5520 5987
rect 5440 5941 5520 5953
rect 5440 5929 5572 5941
rect 5440 5915 5520 5929
rect 5440 5881 5446 5915
rect 5480 5881 5520 5915
rect 5440 5877 5520 5881
rect 5729 5962 5781 5981
rect 5729 5904 5781 5910
rect 5440 5865 5572 5877
rect 5356 5854 5408 5860
rect 3867 5819 6265 5825
rect 3867 5767 5095 5819
rect 5147 5767 5178 5819
rect 5230 5767 5261 5819
rect 5313 5767 6265 5819
rect 3867 5753 6265 5767
rect 3867 5701 5095 5753
rect 5147 5701 5178 5753
rect 5230 5701 5261 5753
rect 5313 5701 6265 5753
rect 3867 5687 6265 5701
rect 3867 5654 5095 5687
rect 5147 5654 5178 5687
rect 5230 5654 5261 5687
rect 5313 5654 6265 5687
rect 3867 5620 3880 5654
rect 3914 5620 3952 5654
rect 3986 5620 4024 5654
rect 4058 5620 4096 5654
rect 4130 5620 4168 5654
rect 4202 5620 4240 5654
rect 4274 5620 4312 5654
rect 4346 5620 4384 5654
rect 4418 5620 4456 5654
rect 4490 5620 4528 5654
rect 4562 5620 4600 5654
rect 4634 5620 4672 5654
rect 4706 5620 4744 5654
rect 4778 5620 4816 5654
rect 4850 5620 4888 5654
rect 4922 5620 4960 5654
rect 4994 5620 5032 5654
rect 5066 5635 5095 5654
rect 5147 5635 5176 5654
rect 5230 5635 5248 5654
rect 5313 5635 5320 5654
rect 5066 5621 5104 5635
rect 5138 5621 5176 5635
rect 5210 5621 5248 5635
rect 5282 5621 5320 5635
rect 5066 5620 5095 5621
rect 5147 5620 5176 5621
rect 5230 5620 5248 5621
rect 5313 5620 5320 5621
rect 5354 5620 5392 5654
rect 5426 5620 5464 5654
rect 5498 5620 5536 5654
rect 5570 5620 5608 5654
rect 5642 5620 5680 5654
rect 5714 5620 5752 5654
rect 5786 5620 5824 5654
rect 5858 5620 5896 5654
rect 5930 5620 5968 5654
rect 6002 5620 6040 5654
rect 6074 5620 6112 5654
rect 6146 5620 6184 5654
rect 6218 5620 6265 5654
rect 3867 5569 5095 5620
rect 5147 5569 5178 5620
rect 5230 5569 5261 5620
rect 5313 5581 6265 5620
rect 5313 5569 5336 5581
rect 3867 5555 5336 5569
rect 3867 5503 5095 5555
rect 5147 5503 5178 5555
rect 5230 5503 5261 5555
rect 5313 5547 5336 5555
rect 5370 5547 5408 5581
rect 5442 5547 5480 5581
rect 5514 5547 5552 5581
rect 5586 5547 5624 5581
rect 5658 5547 5696 5581
rect 5730 5547 5768 5581
rect 5802 5547 5840 5581
rect 5874 5547 5912 5581
rect 5946 5547 5984 5581
rect 6018 5547 6056 5581
rect 6090 5547 6128 5581
rect 6162 5547 6200 5581
rect 6234 5547 6265 5581
rect 5313 5507 6265 5547
rect 5313 5503 5336 5507
rect 3867 5489 5336 5503
rect 3867 5437 5095 5489
rect 5147 5437 5178 5489
rect 5230 5437 5261 5489
rect 5313 5473 5336 5489
rect 5370 5473 5408 5507
rect 5442 5473 5480 5507
rect 5514 5473 5552 5507
rect 5586 5473 5624 5507
rect 5658 5473 5696 5507
rect 5730 5473 5768 5507
rect 5802 5473 5840 5507
rect 5874 5473 5912 5507
rect 5946 5473 5984 5507
rect 6018 5473 6056 5507
rect 6090 5473 6128 5507
rect 6162 5473 6200 5507
rect 6234 5473 6265 5507
rect 5313 5437 6265 5473
rect 3867 5424 6265 5437
rect 3867 5372 5095 5424
rect 5147 5372 5178 5424
rect 5230 5372 5261 5424
rect 5313 5372 6265 5424
rect 3867 5351 6265 5372
tri 5218 5323 5246 5351 ne
rect 5246 5323 6265 5351
rect 3816 5271 3822 5323
rect 3874 5271 3886 5323
rect 3938 5317 4317 5323
rect 3938 5283 4199 5317
rect 4233 5283 4271 5317
rect 4305 5283 4317 5317
tri 5246 5287 5282 5323 ne
rect 5282 5287 6265 5323
rect 3938 5277 4317 5283
rect 3938 5271 3962 5277
tri 3962 5271 3968 5277 nw
rect 6082 5204 6128 5216
tri 6068 5170 6082 5184 se
rect 6082 5170 6088 5204
rect 6122 5170 6128 5204
tri 6066 5168 6068 5170 se
rect 6068 5168 6128 5170
rect 5518 5156 5564 5168
rect 5518 5122 5524 5156
rect 5558 5154 5564 5156
tri 5564 5154 5578 5168 sw
tri 6052 5154 6066 5168 se
rect 6066 5154 6128 5168
rect 5558 5132 6128 5154
rect 5558 5122 6088 5132
rect 5518 5120 6088 5122
rect 4434 5098 4486 5104
tri 4486 5098 4492 5104 sw
rect 5518 5098 5576 5120
tri 5576 5098 5598 5120 nw
tri 6048 5098 6070 5120 ne
rect 6070 5098 6088 5120
rect 6122 5098 6128 5132
rect 4486 5084 4492 5098
tri 4492 5084 4506 5098 sw
rect 5518 5084 5564 5098
tri 5564 5086 5576 5098 nw
tri 6070 5086 6082 5098 ne
rect 6082 5086 6128 5098
rect 4486 5069 4506 5084
tri 4506 5069 4521 5084 sw
rect 4486 5046 5225 5069
rect 4434 5034 5225 5046
rect 4486 5017 5225 5034
rect 4486 5011 4510 5017
tri 4510 5011 4516 5017 nw
tri 5097 5011 5103 5017 ne
rect 5103 5011 5225 5017
rect 4486 5007 4506 5011
tri 4506 5007 4510 5011 nw
tri 5103 5007 5107 5011 ne
rect 5107 5007 5225 5011
rect 4486 4989 4488 5007
tri 4488 4989 4506 5007 nw
tri 5107 4989 5125 5007 ne
rect 5125 4989 5225 5007
tri 4486 4987 4488 4989 nw
rect 4434 4976 4486 4982
rect 4528 4937 4534 4989
rect 4586 4937 4598 4989
rect 4650 4977 4806 4989
rect 4650 4943 4766 4977
rect 4800 4943 4806 4977
tri 5125 4973 5141 4989 ne
rect 5141 4973 5225 4989
rect 4650 4937 4806 4943
tri 5141 4941 5173 4973 ne
tri 4726 4935 4728 4937 ne
rect 4728 4935 4806 4937
tri 4728 4923 4740 4935 ne
rect 4740 4923 4806 4935
tri 4740 4905 4758 4923 ne
rect 4758 4905 4806 4923
tri 4758 4903 4760 4905 ne
rect 4760 4871 4766 4905
rect 4800 4871 4806 4905
rect 4760 4859 4806 4871
rect 5173 4903 5225 4973
rect 5429 5051 5488 5057
rect 5429 5045 5436 5051
rect 5429 5011 5435 5045
rect 5518 5050 5524 5084
rect 5558 5050 5564 5084
rect 5518 5038 5564 5050
rect 5719 5041 5765 5053
tri 5912 5047 5913 5048 se
rect 5913 5047 5959 5053
tri 5765 5041 5771 5047 sw
tri 5906 5041 5912 5047 se
rect 5912 5041 5959 5047
tri 5959 5041 5966 5048 sw
tri 6164 5041 6171 5048 se
rect 6171 5041 6217 5053
rect 5429 4999 5436 5011
rect 5429 4985 5488 4999
rect 5429 4973 5436 4985
rect 5429 4939 5435 4973
rect 5429 4933 5436 4939
rect 5429 4927 5488 4933
rect 5719 5007 5725 5041
rect 5759 5014 5771 5041
tri 5771 5014 5798 5041 sw
tri 5879 5014 5906 5041 se
rect 5906 5014 5919 5041
rect 5759 5007 5919 5014
rect 5953 5014 5966 5041
tri 5966 5014 5993 5041 sw
tri 6137 5014 6164 5041 se
rect 6164 5014 6177 5041
rect 5953 5007 6177 5014
rect 6211 5007 6217 5041
rect 5719 4969 6217 5007
rect 5719 4935 5725 4969
rect 5759 4950 5919 4969
rect 5759 4935 5777 4950
tri 5777 4935 5792 4950 nw
tri 5886 4935 5901 4950 ne
rect 5901 4935 5919 4950
rect 5953 4950 6177 4969
rect 5953 4935 5971 4950
tri 5971 4935 5986 4950 nw
tri 6144 4935 6159 4950 ne
rect 6159 4935 6177 4950
rect 6211 4935 6217 4969
rect 5719 4923 5765 4935
tri 5765 4923 5777 4935 nw
tri 5901 4923 5913 4935 ne
rect 5913 4923 5959 4935
tri 5959 4923 5971 4935 nw
tri 6159 4923 6171 4935 ne
rect 6171 4923 6217 4935
tri 5225 4903 5239 4917 sw
rect 5520 4912 5572 4918
rect 5173 4869 5239 4903
tri 5239 4869 5273 4903 sw
tri 5486 4869 5520 4903 se
rect 5173 4860 5520 4869
rect 5173 4848 5572 4860
tri 4547 4842 4553 4848 se
rect 4553 4842 4565 4848
rect 4417 4836 4565 4842
rect 4417 4802 4429 4836
rect 4463 4802 4501 4836
rect 4535 4802 4565 4836
rect 4417 4796 4565 4802
rect 4617 4796 4629 4848
rect 4681 4796 4687 4848
rect 5173 4799 5520 4848
tri 5511 4796 5514 4799 ne
rect 5514 4796 5520 4799
tri 5514 4790 5520 4796 ne
rect 5520 4790 5572 4796
rect 5733 4840 5863 4846
rect 5785 4834 5863 4840
rect 5785 4800 5823 4834
rect 5857 4800 5863 4834
rect 5785 4788 5863 4800
rect 5733 4774 5863 4788
tri 4123 4728 4144 4749 se
tri 4062 4667 4123 4728 se
rect 4123 4667 4144 4728
tri 4044 4649 4062 4667 se
rect 4062 4649 4144 4667
tri 4894 4728 4915 4749 sw
rect 4894 4667 4915 4728
tri 4915 4667 4976 4728 sw
rect 5785 4762 5863 4774
rect 5785 4728 5823 4762
rect 5857 4728 5863 4762
rect 5785 4722 5863 4728
rect 5733 4716 5863 4722
rect 4894 4649 5336 4667
rect 3868 4513 5336 4649
rect 5571 4513 5642 4667
rect 5876 4513 6187 4619
rect 3868 4501 6218 4513
rect 6265 4504 6292 4667
rect 3868 4470 5230 4501
rect 3868 4436 4055 4470
rect 4089 4436 4127 4470
rect 4161 4436 4199 4470
rect 4233 4436 4271 4470
rect 4305 4436 4343 4470
rect 4377 4436 4415 4470
rect 4449 4436 4487 4470
rect 4521 4436 4559 4470
rect 4593 4436 4631 4470
rect 4665 4436 4703 4470
rect 4737 4436 4775 4470
rect 4809 4436 4847 4470
rect 4881 4436 4919 4470
rect 4953 4436 4991 4470
rect 5025 4436 5063 4470
rect 5097 4436 5135 4470
rect 5169 4467 5230 4470
rect 5264 4467 5302 4501
rect 5336 4467 5374 4501
rect 5408 4467 5446 4501
rect 5480 4467 5518 4501
rect 5552 4467 5590 4501
rect 5624 4467 5662 4501
rect 5696 4467 5734 4501
rect 5768 4467 5806 4501
rect 5840 4467 5878 4501
rect 5912 4467 5950 4501
rect 5984 4467 6022 4501
rect 6056 4467 6094 4501
rect 6128 4467 6218 4501
rect 5169 4455 6218 4467
rect 5169 4447 5336 4455
rect 5169 4436 5311 4447
rect 3868 4303 5311 4436
rect 5876 4387 6187 4455
tri 3995 4258 4040 4303 ne
rect 4040 4301 5311 4303
rect 4040 4284 4965 4301
rect 4040 4258 4144 4284
tri 4040 4246 4052 4258 ne
rect 4052 4246 4144 4258
tri 4052 4212 4086 4246 ne
rect 4086 4212 4144 4246
tri 4086 4174 4124 4212 ne
rect 4124 4174 4144 4212
tri 4124 4154 4144 4174 ne
rect 4861 4258 4965 4284
tri 4965 4258 5008 4301 nw
rect 4861 4246 4953 4258
tri 4953 4246 4965 4258 nw
rect 5317 4246 5363 4258
rect 6109 4252 6161 4258
tri 5363 4246 5367 4250 sw
tri 6105 4246 6109 4250 se
rect 4861 4212 4919 4246
tri 4919 4212 4953 4246 nw
rect 5317 4212 5323 4246
rect 5357 4216 5367 4246
tri 5367 4216 5397 4246 sw
tri 6075 4216 6105 4246 se
rect 6105 4216 6109 4246
rect 5357 4212 6109 4216
rect 4861 4174 4881 4212
tri 4881 4174 4919 4212 nw
rect 5317 4200 6109 4212
rect 5317 4183 6161 4200
rect 5317 4174 6109 4183
tri 4861 4154 4881 4174 nw
rect 5317 4140 5323 4174
rect 5357 4170 6109 4174
rect 5357 4140 5367 4170
tri 5367 4140 5397 4170 nw
tri 6075 4140 6105 4170 ne
rect 6105 4140 6109 4170
rect 5317 4128 5363 4140
tri 5363 4136 5367 4140 nw
tri 6105 4136 6109 4140 ne
rect 6109 4125 6161 4131
rect 5746 4033 5792 4045
tri 5939 4042 5940 4043 se
rect 5940 4042 5986 4043
rect 5746 3999 5752 4033
rect 5786 4031 5792 4033
tri 5792 4031 5803 4042 sw
tri 5928 4031 5939 4042 se
rect 5939 4031 5986 4042
tri 5986 4031 5998 4043 sw
tri 6186 4031 6198 4043 se
rect 6198 4031 6244 4043
rect 5786 4016 5803 4031
tri 5803 4016 5818 4031 sw
tri 5913 4016 5928 4031 se
rect 5928 4016 5946 4031
rect 5786 3999 5946 4016
rect 5746 3997 5946 3999
rect 5980 4016 5998 4031
tri 5998 4016 6013 4031 sw
tri 6171 4016 6186 4031 se
rect 6186 4016 6204 4031
rect 5980 3997 6204 4016
rect 6238 3997 6244 4031
rect 4383 3969 5628 3975
rect 3952 3962 4004 3968
tri 4181 3956 4193 3968 se
rect 4193 3956 4239 3968
tri 4172 3947 4181 3956 se
rect 4181 3947 4199 3956
tri 4004 3922 4029 3947 sw
tri 4147 3922 4172 3947 se
rect 4172 3922 4199 3947
rect 4233 3922 4239 3956
rect 4383 3935 4395 3969
rect 4429 3935 4467 3969
rect 4501 3935 5628 3969
rect 4383 3929 5628 3935
tri 5548 3927 5550 3929 ne
rect 5550 3927 5628 3929
tri 5550 3925 5552 3927 ne
rect 5552 3925 5628 3927
rect 4004 3913 4029 3922
tri 4029 3913 4038 3922 sw
tri 4138 3913 4147 3922 se
rect 4147 3913 4239 3922
tri 5552 3915 5562 3925 ne
rect 5562 3915 5628 3925
rect 5746 3961 6244 3997
rect 5746 3927 5752 3961
rect 5786 3959 6244 3961
rect 5786 3952 5946 3959
rect 5786 3927 5799 3952
rect 5746 3925 5799 3927
tri 5799 3925 5826 3952 nw
tri 5901 3925 5928 3952 ne
rect 5928 3925 5946 3952
rect 5980 3952 6204 3959
rect 5980 3925 5998 3952
tri 5998 3925 6025 3952 nw
tri 6165 3925 6192 3952 ne
rect 6192 3925 6204 3952
rect 6238 3925 6244 3959
rect 5746 3915 5792 3925
tri 5792 3918 5799 3925 nw
tri 5928 3918 5935 3925 ne
rect 5935 3918 5986 3925
tri 5935 3915 5938 3918 ne
rect 5938 3915 5986 3918
tri 5562 3913 5564 3915 ne
rect 5564 3913 5628 3915
tri 5938 3913 5940 3915 ne
rect 5940 3913 5986 3915
tri 5986 3913 5998 3925 nw
tri 6192 3919 6198 3925 ne
rect 6198 3913 6244 3925
rect 4004 3910 4239 3913
rect 3952 3898 4239 3910
rect 4004 3884 4239 3898
tri 5564 3897 5580 3913 ne
rect 5580 3897 5628 3913
tri 5580 3895 5582 3897 ne
rect 4004 3861 4199 3884
rect 4004 3850 4014 3861
tri 4014 3850 4025 3861 nw
tri 4170 3850 4181 3861 ne
rect 4181 3850 4199 3861
rect 4233 3850 4239 3884
rect 3952 3840 4004 3846
tri 4004 3840 4014 3850 nw
tri 4181 3840 4191 3850 ne
rect 4191 3840 4239 3850
tri 4191 3838 4193 3840 ne
rect 4193 3838 4239 3840
rect 4358 3829 4364 3881
rect 4416 3829 4428 3881
rect 4480 3869 4776 3881
rect 4480 3835 4736 3869
rect 4770 3835 4776 3869
rect 4480 3829 4776 3835
tri 4696 3813 4712 3829 ne
rect 4712 3813 4776 3829
tri 4712 3805 4720 3813 ne
rect 4720 3805 4776 3813
tri 4720 3797 4728 3805 ne
rect 4728 3797 4776 3805
tri 4728 3795 4730 3797 ne
rect 4730 3763 4736 3797
rect 4770 3763 4776 3797
rect 4730 3751 4776 3763
rect 4891 3877 4943 3882
tri 4943 3877 4947 3881 sw
rect 5403 3877 5449 3889
rect 4891 3876 4947 3877
rect 4943 3871 4947 3876
tri 4947 3871 4953 3877 sw
rect 4943 3843 4953 3871
tri 4953 3843 4981 3871 sw
tri 5375 3843 5403 3871 se
rect 5403 3843 5409 3877
rect 5443 3843 5449 3877
rect 4943 3842 4981 3843
tri 4981 3842 4982 3843 sw
tri 5374 3842 5375 3843 se
rect 5375 3842 5449 3843
rect 4943 3837 4982 3842
tri 4982 3837 4987 3842 sw
tri 5369 3837 5374 3842 se
rect 5374 3837 5449 3842
rect 4943 3824 5449 3837
rect 4891 3812 5449 3824
rect 4943 3805 5449 3812
rect 4943 3799 5409 3805
rect 4943 3795 4964 3799
tri 4964 3795 4968 3799 nw
tri 5369 3795 5373 3799 ne
rect 5373 3795 5409 3799
tri 4943 3774 4964 3795 nw
tri 5373 3774 5394 3795 ne
rect 5394 3774 5409 3795
tri 5394 3771 5397 3774 ne
rect 5397 3771 5409 3774
rect 5443 3771 5449 3805
tri 5397 3770 5398 3771 ne
rect 5398 3770 5449 3771
tri 5398 3765 5403 3770 ne
rect 4891 3754 4943 3760
rect 5403 3759 5449 3770
rect 5582 3876 5628 3897
rect 5582 3842 5588 3876
rect 5622 3842 5628 3876
rect 5582 3804 5628 3842
rect 5582 3770 5588 3804
rect 5622 3770 5628 3804
rect 5582 3758 5628 3770
rect 5814 3891 5890 3897
rect 5866 3885 5890 3891
rect 5884 3851 5890 3885
rect 5866 3839 5890 3851
rect 5814 3825 5890 3839
rect 5866 3813 5890 3825
rect 5884 3779 5890 3813
rect 5866 3773 5890 3779
rect 5814 3767 5890 3773
tri 5109 3553 5237 3681 se
rect 5237 3675 5458 3681
rect 5237 3623 5238 3675
rect 5290 3623 5322 3675
rect 5374 3623 5406 3675
rect 5237 3599 5458 3623
rect 5237 3553 5238 3599
rect -8872 3542 -8635 3548
rect -8872 3490 -8687 3542
rect -8872 3476 -8635 3490
rect -8872 3424 -8687 3476
rect -8872 3418 -8635 3424
rect 4057 3547 5238 3553
rect 5290 3547 5322 3599
rect 5374 3547 5406 3599
rect 6046 3553 6213 3609
rect 5458 3547 6292 3553
rect 4057 3523 6292 3547
rect 4057 3512 5238 3523
rect 5290 3512 5322 3523
rect 5374 3512 5406 3523
rect 5458 3512 6292 3523
rect 4057 3478 5126 3512
rect 5160 3478 5198 3512
rect 5232 3478 5238 3512
rect 5304 3478 5322 3512
rect 5376 3478 5406 3512
rect 5458 3478 5486 3512
rect 5520 3478 5558 3512
rect 5592 3478 5630 3512
rect 5664 3478 5702 3512
rect 5736 3478 5774 3512
rect 5808 3478 5846 3512
rect 5880 3478 5918 3512
rect 5952 3478 5990 3512
rect 6024 3478 6062 3512
rect 6096 3478 6134 3512
rect 6168 3478 6206 3512
rect 6240 3478 6292 3512
rect 4057 3471 5238 3478
rect 5290 3471 5322 3478
rect 5374 3471 5406 3478
rect 5458 3471 6292 3478
rect 4057 3448 6292 3471
rect 4057 3396 5238 3448
rect 5290 3396 5322 3448
rect 5374 3396 5406 3448
rect 5458 3396 6292 3448
rect 4057 3390 6292 3396
tri -8913 3102 -8856 3159 se
rect -8856 3102 -8473 3159
rect -9329 2761 -9284 2963
rect -8491 2848 -8429 2957
tri -8429 2848 -8320 2957 nw
rect 4430 2899 4741 3074
tri -8491 2786 -8429 2848 nw
rect 6040 2842 6168 2848
rect 6092 2790 6116 2842
rect 6040 2776 6168 2790
rect 6092 2724 6116 2776
rect 6040 2718 6168 2724
rect -8750 2539 -8635 2545
rect -8750 2533 -8687 2539
rect -8750 2499 -8744 2533
rect -8710 2499 -8687 2533
rect -9012 2487 -8966 2499
rect -9012 2453 -9006 2487
rect -8972 2453 -8966 2487
rect -9012 2415 -8966 2453
rect -9012 2381 -9006 2415
rect -8972 2381 -8966 2415
rect -9012 2369 -8966 2381
rect -8833 2487 -8787 2499
rect -8833 2453 -8827 2487
rect -8793 2453 -8787 2487
rect -8833 2415 -8787 2453
rect -8750 2487 -8687 2499
rect 4316 2518 4387 2555
rect 5657 2525 5698 2569
rect 6220 2490 6294 2525
rect -8750 2473 -8635 2487
rect -8750 2461 -8687 2473
rect -8750 2427 -8744 2461
rect -8710 2427 -8687 2461
rect -8750 2421 -8687 2427
rect -8750 2415 -8635 2421
rect -8833 2381 -8827 2415
rect -8793 2381 -8787 2415
rect -8833 2369 -8787 2381
rect -9186 2343 -9140 2355
rect -9186 2309 -9180 2343
rect -9146 2309 -9140 2343
rect -9186 2271 -9140 2309
rect -9186 2237 -9180 2271
rect -9146 2237 -9140 2271
rect -9186 2225 -9140 2237
rect -9102 2336 -9056 2348
rect -9102 2302 -9096 2336
rect -9062 2302 -9056 2336
rect -8655 2336 -8609 2348
tri -9056 2302 -9052 2306 sw
rect -8655 2302 -8649 2336
rect -8615 2302 -8609 2336
rect -9102 2300 -9052 2302
tri -9052 2300 -9050 2302 sw
rect -9102 2264 -9050 2300
tri -9050 2264 -9014 2300 sw
tri -8691 2264 -8655 2300 se
rect -8655 2264 -8609 2302
rect -9102 2230 -9096 2264
rect -9062 2230 -8649 2264
rect -8615 2230 -8609 2264
rect -9102 2218 -8609 2230
rect 4310 2196 4377 2240
rect -8496 2079 -8491 2141
tri -8491 2079 -8429 2141 sw
rect -8496 2010 -8429 2079
tri -8429 2010 -8360 2079 sw
rect 5343 2073 5459 2079
rect 4346 1898 4513 2054
rect 5395 2021 5407 2073
rect 5343 2006 5459 2021
rect 5395 1954 5407 2006
rect 5343 1940 5459 1954
rect 5395 1888 5407 1940
rect 5343 1882 5459 1888
tri 6162 1847 6196 1881 ne
rect 6196 1744 6248 1881
tri 6248 1855 6274 1881 nw
rect 6003 1703 6045 1741
rect 6033 1340 6168 1457
<< via1 >>
rect 5099 7616 5151 7623
rect 5099 7582 5107 7616
rect 5107 7582 5141 7616
rect 5141 7582 5151 7616
rect 5099 7571 5151 7582
rect 5178 7616 5230 7623
rect 5256 7616 5308 7623
rect 5178 7582 5179 7616
rect 5179 7582 5213 7616
rect 5213 7582 5230 7616
rect 5256 7582 5285 7616
rect 5285 7582 5308 7616
rect 5178 7571 5230 7582
rect 5256 7571 5308 7582
rect 5099 7492 5151 7544
rect 5178 7492 5230 7544
rect 5256 7492 5308 7544
rect 5099 7413 5151 7465
rect 5178 7413 5230 7465
rect 5256 7413 5308 7465
rect 4434 7305 4486 7312
rect 4434 7271 4443 7305
rect 4443 7271 4477 7305
rect 4477 7271 4486 7305
rect 4434 7260 4486 7271
rect 4434 7233 4486 7245
rect 4434 7199 4443 7233
rect 4443 7199 4477 7233
rect 4477 7199 4486 7233
rect 4434 7193 4486 7199
rect 4603 7305 4655 7312
rect 4603 7271 4612 7305
rect 4612 7271 4646 7305
rect 4646 7271 4655 7305
rect 4603 7260 4655 7271
rect 4603 7233 4655 7245
rect 4603 7199 4612 7233
rect 4612 7199 4646 7233
rect 4646 7199 4655 7233
rect 4603 7193 4655 7199
rect 4786 7309 4838 7316
rect 4786 7275 4795 7309
rect 4795 7275 4829 7309
rect 4829 7275 4838 7309
rect 4786 7264 4838 7275
rect 4786 7237 4838 7249
rect 4786 7203 4795 7237
rect 4795 7203 4829 7237
rect 4829 7203 4838 7237
rect 4786 7197 4838 7203
rect 4959 7309 5011 7316
rect 4959 7275 4968 7309
rect 4968 7275 5002 7309
rect 5002 7275 5011 7309
rect 4959 7264 5011 7275
rect 4959 7237 5011 7249
rect 4959 7203 4968 7237
rect 4968 7203 5002 7237
rect 5002 7203 5011 7237
rect 4959 7197 5011 7203
rect 5436 7309 5488 7316
rect 5436 7275 5445 7309
rect 5445 7275 5479 7309
rect 5479 7275 5488 7309
rect 5436 7264 5488 7275
rect 5436 7237 5488 7249
rect 5436 7203 5445 7237
rect 5445 7203 5479 7237
rect 5479 7203 5488 7237
rect 5436 7197 5488 7203
rect 5659 7246 5711 7298
rect 5723 7246 5775 7298
rect 5442 7043 5494 7095
rect 5506 7043 5558 7095
rect 5002 6906 5054 6958
rect 5002 6842 5054 6894
rect 4695 6278 4747 6330
rect 4695 6214 4747 6266
rect 4786 6188 4838 6240
rect 4786 6124 4838 6176
rect 5002 6221 5054 6227
rect 5002 6187 5007 6221
rect 5007 6187 5041 6221
rect 5041 6187 5054 6221
rect 5002 6175 5054 6187
rect 5002 6149 5054 6161
rect 5002 6115 5007 6149
rect 5007 6115 5041 6149
rect 5041 6115 5054 6149
rect 5002 6109 5054 6115
rect 4821 6024 4873 6076
rect 4885 6024 4937 6076
rect 5729 6022 5781 6033
rect 4519 5939 4571 5991
rect 4519 5873 4571 5925
rect 5356 5924 5408 5976
rect 5356 5860 5408 5912
rect 5520 5941 5572 5993
rect 5520 5877 5572 5929
rect 5729 5988 5737 6022
rect 5737 5988 5771 6022
rect 5771 5988 5781 6022
rect 5729 5981 5781 5988
rect 5729 5950 5781 5962
rect 5729 5916 5737 5950
rect 5737 5916 5771 5950
rect 5771 5916 5781 5950
rect 5729 5910 5781 5916
rect 5095 5767 5147 5819
rect 5178 5767 5230 5819
rect 5261 5767 5313 5819
rect 5095 5701 5147 5753
rect 5178 5701 5230 5753
rect 5261 5701 5313 5753
rect 5095 5654 5147 5687
rect 5178 5654 5230 5687
rect 5261 5654 5313 5687
rect 5095 5635 5104 5654
rect 5104 5635 5138 5654
rect 5138 5635 5147 5654
rect 5178 5635 5210 5654
rect 5210 5635 5230 5654
rect 5261 5635 5282 5654
rect 5282 5635 5313 5654
rect 5095 5620 5104 5621
rect 5104 5620 5138 5621
rect 5138 5620 5147 5621
rect 5178 5620 5210 5621
rect 5210 5620 5230 5621
rect 5261 5620 5282 5621
rect 5282 5620 5313 5621
rect 5095 5569 5147 5620
rect 5178 5569 5230 5620
rect 5261 5569 5313 5620
rect 5095 5503 5147 5555
rect 5178 5503 5230 5555
rect 5261 5503 5313 5555
rect 5095 5437 5147 5489
rect 5178 5437 5230 5489
rect 5261 5437 5313 5489
rect 5095 5372 5147 5424
rect 5178 5372 5230 5424
rect 5261 5372 5313 5424
rect 3822 5271 3874 5323
rect 3886 5271 3938 5323
rect 4434 5046 4486 5098
rect 4434 4982 4486 5034
rect 4534 4937 4586 4989
rect 4598 4937 4650 4989
rect 5436 5045 5488 5051
rect 5436 5011 5469 5045
rect 5469 5011 5488 5045
rect 5436 4999 5488 5011
rect 5436 4973 5488 4985
rect 5436 4939 5469 4973
rect 5469 4939 5488 4973
rect 5436 4933 5488 4939
rect 5520 4860 5572 4912
rect 4565 4796 4617 4848
rect 4629 4796 4681 4848
rect 5520 4796 5572 4848
rect 5733 4788 5785 4840
rect 5733 4722 5785 4774
rect 6109 4246 6161 4252
rect 6109 4212 6116 4246
rect 6116 4212 6150 4246
rect 6150 4212 6161 4246
rect 6109 4200 6161 4212
rect 6109 4174 6161 4183
rect 6109 4140 6116 4174
rect 6116 4140 6150 4174
rect 6150 4140 6161 4174
rect 6109 4131 6161 4140
rect 3952 3910 4004 3962
rect 3952 3846 4004 3898
rect 4364 3829 4416 3881
rect 4428 3829 4480 3881
rect 4891 3824 4943 3876
rect 4891 3760 4943 3812
rect 5814 3885 5866 3891
rect 5814 3851 5850 3885
rect 5850 3851 5866 3885
rect 5814 3839 5866 3851
rect 5814 3813 5866 3825
rect 5814 3779 5850 3813
rect 5850 3779 5866 3813
rect 5814 3773 5866 3779
rect 5238 3623 5290 3675
rect 5322 3623 5374 3675
rect 5406 3623 5458 3675
rect -8687 3490 -8635 3542
rect -8687 3424 -8635 3476
rect 5238 3547 5290 3599
rect 5322 3547 5374 3599
rect 5406 3547 5458 3599
rect 5238 3512 5290 3523
rect 5322 3512 5374 3523
rect 5406 3512 5458 3523
rect 5238 3478 5270 3512
rect 5270 3478 5290 3512
rect 5322 3478 5342 3512
rect 5342 3478 5374 3512
rect 5406 3478 5414 3512
rect 5414 3478 5448 3512
rect 5448 3478 5458 3512
rect 5238 3471 5290 3478
rect 5322 3471 5374 3478
rect 5406 3471 5458 3478
rect 5238 3396 5290 3448
rect 5322 3396 5374 3448
rect 5406 3396 5458 3448
rect 6040 2790 6092 2842
rect 6116 2790 6168 2842
rect 6040 2724 6092 2776
rect 6116 2724 6168 2776
rect -8687 2487 -8635 2539
rect -8687 2421 -8635 2473
rect 5343 2021 5395 2073
rect 5407 2021 5459 2073
rect 5343 1954 5395 2006
rect 5407 1954 5459 2006
rect 5343 1888 5395 1940
rect 5407 1888 5459 1940
<< metal2 >>
rect 5093 7623 5314 7624
rect 5093 7571 5099 7623
rect 5151 7571 5178 7623
rect 5230 7571 5256 7623
rect 5308 7571 5314 7623
rect 5093 7544 5314 7571
rect 5093 7492 5099 7544
rect 5151 7492 5178 7544
rect 5230 7492 5256 7544
rect 5308 7492 5314 7544
tri 3907 5372 3952 5417 se
rect 3952 5372 4004 7362
tri 3858 5323 3907 5372 se
rect 3907 5323 4004 5372
rect 3816 5271 3822 5323
rect 3874 5271 3886 5323
rect 3938 5271 4004 5323
tri 3858 5177 3952 5271 ne
rect 3952 3962 4004 5271
rect 4434 7312 4486 7432
rect 4434 7245 4486 7260
rect 4434 5098 4486 7193
rect 4519 5991 4571 7453
rect 4519 5925 4571 5939
rect 4519 5867 4571 5873
rect 4603 7312 4655 7425
rect 4603 7245 4655 7260
tri 4590 5051 4603 5064 se
rect 4603 5051 4655 7193
rect 4786 7316 4838 7473
rect 4786 7249 4838 7264
rect 4959 7316 5011 7473
rect 4959 7249 5011 7264
tri 4925 7209 4959 7243 se
rect 4434 5034 4486 5046
tri 4538 4999 4590 5051 se
rect 4590 4999 4655 5051
rect 3952 3898 4004 3910
tri 4385 3891 4434 3940 se
rect 4434 3891 4486 4982
tri 4528 4989 4538 4999 se
rect 4538 4989 4655 4999
rect 4695 6330 4747 6336
rect 4695 6266 4747 6278
tri 4655 4989 4656 4990 sw
rect 4528 4937 4534 4989
rect 4586 4937 4598 4989
rect 4650 4937 4656 4989
tri 4655 4860 4695 4900 se
rect 4695 4860 4747 6214
rect 4786 6240 4838 7197
rect 4786 6176 4838 6188
rect 4786 6118 4838 6124
rect 4891 7197 4959 7209
rect 4891 7157 5011 7197
rect 5093 7465 5314 7492
rect 5093 7413 5099 7465
rect 5151 7413 5178 7465
rect 5230 7413 5256 7465
rect 5308 7413 5314 7465
tri 4890 6109 4891 6110 se
rect 4891 6109 4943 7157
tri 4943 7123 4977 7157 nw
tri 4857 6076 4890 6109 se
rect 4890 6076 4943 6109
rect 5002 6958 5054 6964
rect 5002 6894 5054 6906
rect 5002 6227 5054 6842
rect 5002 6161 5054 6175
rect 5002 6103 5054 6109
rect 4815 6024 4821 6076
rect 4873 6024 4885 6076
rect 4937 6024 4943 6076
tri 4857 5993 4888 6024 ne
rect 4888 5993 4943 6024
tri 4888 5990 4891 5993 ne
tri 4643 4848 4655 4860 se
rect 4655 4848 4747 4860
rect 4559 4796 4565 4848
rect 4617 4796 4629 4848
rect 4681 4796 4747 4848
tri 4376 3882 4385 3891 se
rect 4385 3882 4486 3891
tri 4375 3881 4376 3882 se
rect 4376 3881 4486 3882
rect 3952 3840 4004 3846
rect 4358 3829 4364 3881
rect 4416 3829 4428 3881
rect 4480 3829 4486 3881
rect 4891 3876 4943 5993
rect 4891 3812 4943 3824
rect 4891 3754 4943 3760
rect 5093 5819 5314 7413
rect 5436 7316 5488 7473
tri 5414 7264 5436 7286 se
tri 5399 7249 5414 7264 se
rect 5414 7249 5488 7264
tri 5380 7230 5399 7249 se
rect 5399 7230 5436 7249
rect 5356 7197 5436 7230
rect 5653 7246 5659 7298
rect 5711 7246 5723 7298
rect 5775 7246 5781 7298
tri 5695 7212 5729 7246 ne
rect 5356 7191 5488 7197
rect 5356 7157 5443 7191
tri 5443 7157 5477 7191 nw
rect 5356 7123 5409 7157
tri 5409 7123 5443 7157 nw
rect 5356 5976 5408 7123
tri 5408 7122 5409 7123 nw
rect 5356 5912 5408 5924
rect 5356 5854 5408 5860
rect 5436 7043 5442 7095
rect 5494 7043 5506 7095
rect 5558 7043 5564 7095
rect 5093 5767 5095 5819
rect 5147 5767 5178 5819
rect 5230 5767 5261 5819
rect 5313 5767 5314 5819
rect 5093 5753 5314 5767
rect 5093 5701 5095 5753
rect 5147 5701 5178 5753
rect 5230 5701 5261 5753
rect 5313 5701 5314 5753
rect 5093 5687 5314 5701
rect 5093 5635 5095 5687
rect 5147 5635 5178 5687
rect 5230 5635 5261 5687
rect 5313 5635 5314 5687
rect 5093 5621 5314 5635
rect 5093 5569 5095 5621
rect 5147 5569 5178 5621
rect 5230 5569 5261 5621
rect 5313 5569 5314 5621
rect 5093 5555 5314 5569
rect 5093 5503 5095 5555
rect 5147 5503 5178 5555
rect 5230 5503 5261 5555
rect 5313 5503 5314 5555
rect 5093 5489 5314 5503
rect 5093 5437 5095 5489
rect 5147 5437 5178 5489
rect 5230 5437 5261 5489
rect 5313 5437 5314 5489
rect 5093 5424 5314 5437
rect 5093 5372 5095 5424
rect 5147 5372 5178 5424
rect 5230 5372 5261 5424
rect 5313 5372 5314 5424
rect 5093 3897 5314 5372
rect 5436 5051 5488 7043
tri 5488 7009 5522 7043 nw
rect 5729 6033 5781 7246
rect 5436 4985 5488 4999
rect 5436 4927 5488 4933
rect 5520 5993 5572 5999
rect 5520 5929 5572 5941
rect 5729 5962 5781 5981
rect 5729 5904 5781 5910
rect 5520 4912 5572 5877
rect 5520 4848 5572 4860
rect 5520 4790 5572 4796
rect 5733 4840 5785 4846
rect 5733 4774 5785 4788
rect 5733 4716 5785 4722
rect 6109 4252 6161 4258
rect 6109 4183 6161 4200
rect 6109 4125 6161 4131
tri 5314 3897 5399 3982 sw
rect 5093 3891 5399 3897
tri 5399 3891 5405 3897 sw
rect 5814 3891 5866 3897
rect 5093 3839 5405 3891
tri 5405 3839 5457 3891 sw
rect 5093 3837 5457 3839
tri 5457 3837 5459 3839 sw
rect 5093 3675 5459 3837
rect 5814 3825 5866 3839
rect 5814 3767 5866 3773
rect 5093 3623 5238 3675
rect 5290 3623 5322 3675
rect 5374 3623 5406 3675
rect 5458 3623 5459 3675
rect 5093 3599 5459 3623
rect -8687 3542 -8635 3548
rect -8687 3476 -8635 3490
rect -8687 2539 -8635 3424
rect 5093 3547 5238 3599
rect 5290 3547 5322 3599
rect 5374 3547 5406 3599
rect 5458 3547 5459 3599
rect 5093 3523 5459 3547
rect 5093 3471 5238 3523
rect 5290 3471 5322 3523
rect 5374 3471 5406 3523
rect 5458 3471 5459 3523
rect 5093 3448 5459 3471
rect 5093 3396 5238 3448
rect 5290 3396 5322 3448
rect 5374 3396 5406 3448
rect 5458 3396 5459 3448
rect 5093 3310 5459 3396
tri 5093 3201 5202 3310 ne
rect 5202 3107 5459 3310
rect -8687 2473 -8635 2487
rect -8687 2415 -8635 2421
rect 5237 2073 5459 3107
rect 6040 2842 6168 2848
rect 6092 2790 6116 2842
rect 6040 2776 6168 2790
rect 6092 2724 6116 2776
rect 6040 2688 6168 2724
tri 5755 2254 5789 2288 se
rect 5237 2021 5343 2073
rect 5395 2021 5407 2073
rect 5237 2006 5459 2021
rect 5237 1954 5343 2006
rect 5395 1954 5407 2006
rect 5237 1940 5459 1954
rect 5237 1888 5343 1940
rect 5395 1888 5407 1940
rect 5237 1878 5459 1888
use sky130_fd_io__com_ctl_ls_octl  sky130_fd_io__com_ctl_ls_octl_0
timestamp 1648127584
transform 1 0 4281 0 -1 3202
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1648127584
transform -1 0 5943 0 1 5584
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1648127584
transform 1 0 5926 0 -1 5526
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1648127584
transform -1 0 5943 0 -1 7652
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_3
timestamp 1648127584
transform 1 0 5274 0 -1 5526
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_4
timestamp 1648127584
transform 1 0 5953 0 1 3442
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1648127584
transform -1 0 6295 0 1 5584
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_1
timestamp 1648127584
transform 1 0 5761 0 -1 7652
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_2
timestamp 1648127584
transform 1 0 5601 0 1 3442
box 0 24 534 1116
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_3
timestamp 1648127584
transform 1 0 5574 0 -1 5526
box 0 24 534 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1648127584
transform 1 0 -8994 0 1 1902
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1648127584
transform -1 0 5291 0 1 5584
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1648127584
transform 1 0 5109 0 1 5584
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1648127584
transform 1 0 4281 0 1 5584
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_4
timestamp 1648127584
transform -1 0 4339 0 -1 7652
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_5
timestamp 1648127584
transform 1 0 4633 0 -1 7652
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_6
timestamp 1648127584
transform -1 0 5643 0 -1 7652
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_7
timestamp 1648127584
transform -1 0 4815 0 -1 7652
box -42 24 569 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1648127584
transform -1 0 -8812 0 1 1902
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1648127584
transform -1 0 4339 0 1 5584
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_2
timestamp 1648127584
transform -1 0 5783 0 1 3442
box 0 24 534 1116
use sky130_fd_io__hvsbt_xor  sky130_fd_io__hvsbt_xor_0
timestamp 1648127584
transform 1 0 3805 0 -1 5656
box 95 75 1333 1135
use sky130_fd_io__hvsbt_xorv2  sky130_fd_io__hvsbt_xorv2_0
timestamp 1648127584
transform 1 0 3772 0 1 3247
box 95 75 1333 1135
<< labels >>
flabel metal2 s 4436 7368 4485 7431 3 FreeSans 520 270 0 0 DM_H[0]
port 1 nsew
flabel metal2 s 3965 7295 3991 7344 3 FreeSans 520 270 0 0 DM_H[2]
port 2 nsew
flabel metal2 s 5442 7419 5486 7468 3 FreeSans 520 270 0 0 DM_H_N[0]
port 3 nsew
flabel metal2 s 4968 7412 5002 7461 3 FreeSans 520 270 0 0 DM_H_N[1]
port 4 nsew
flabel metal2 s 4796 7417 4831 7462 3 FreeSans 520 270 0 0 DM_H_N[2]
port 5 nsew
flabel metal2 s 5020 6773 5051 6867 3 FreeSans 520 0 0 0 PUEN_2OR1_H
port 6 nsew
flabel metal2 s 4604 7370 4653 7423 3 FreeSans 520 270 0 0 DM_H[1]
port 7 nsew
flabel comment s 5456 7513 5456 7513 0 FreeSans 440 90 0 0 DM_H_N<0>
flabel comment s 4980 7575 4980 7575 0 FreeSans 440 270 0 0 DM_H_N<1>
flabel comment s 4804 7579 4804 7579 0 FreeSans 440 270 0 0 DM_H_N<2>
flabel comment s 4452 6892 4452 6892 0 FreeSans 440 90 0 0 DM_H<0>
flabel comment s 4630 6909 4630 6909 0 FreeSans 440 90 0 0 DM_H<1>
flabel comment s 3971 6510 3971 6510 0 FreeSans 440 270 0 0 DM_H<2>
flabel metal1 s 6014 6884 6044 6944 3 FreeSans 520 0 0 0 PDEN_H_N[1]
port 8 nsew
flabel metal1 s 6012 6289 6046 6353 3 FreeSans 520 0 0 0 PDEN_H_N[0]
port 9 nsew
flabel metal1 s 6003 1703 6045 1741 3 FreeSans 520 180 0 0 OD_H
port 10 nsew
flabel metal1 s 6220 2490 6294 2525 3 FreeSans 520 180 0 0 SLOW
port 11 nsew
flabel metal1 s 4316 2518 4387 2555 3 FreeSans 520 180 0 0 SLOW_H
port 12 nsew
flabel metal1 s 4310 2196 4377 2240 3 FreeSans 520 180 0 0 SLOW_H_N
port 13 nsew
flabel metal1 s 5657 2525 5698 2569 3 FreeSans 520 180 0 0 HLD_I_H_N
port 14 nsew
flabel metal1 s 5876 6498 6187 6730 3 FreeSans 520 0 0 0 VCC_IO
port 15 nsew
flabel metal1 s 6019 7436 6186 7606 3 FreeSans 520 0 0 0 VGND
port 16 nsew
flabel metal1 s 6033 1340 6168 1457 3 FreeSans 520 180 0 0 VPWR
port 17 nsew
flabel metal1 s 5876 4387 6187 4619 3 FreeSans 520 0 0 0 VCC_IO
port 15 nsew
flabel metal1 s 6019 5485 6186 5641 3 FreeSans 520 0 0 0 VGND
port 16 nsew
flabel metal1 s 6046 3453 6213 3609 3 FreeSans 520 0 0 0 VGND
port 16 nsew
flabel metal1 s 4346 1898 4513 2054 3 FreeSans 520 180 0 0 VGND
port 16 nsew
flabel metal1 s 4430 2899 4741 3074 3 FreeSans 520 180 0 0 VCC_IO
port 15 nsew
<< properties >>
string GDS_END 6893798
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6828852
<< end >>
