magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 1951 203
rect 30 -17 64 21
<< locali >>
rect 607 323 673 493
rect 775 323 841 493
rect 943 323 1009 493
rect 1111 323 1177 493
rect 1279 323 1345 493
rect 1447 323 1513 493
rect 1615 323 1681 493
rect 1783 323 1849 493
rect 1952 323 2007 472
rect 607 289 2007 323
rect 17 215 497 255
rect 1931 181 2007 289
rect 607 147 2007 181
rect 607 52 673 147
rect 607 51 657 52
rect 775 52 841 147
rect 791 51 825 52
rect 943 52 1009 147
rect 959 51 993 52
rect 1111 52 1177 147
rect 1279 52 1345 147
rect 1447 52 1513 147
rect 1615 52 1681 147
rect 1783 52 1849 147
rect 1952 73 2007 147
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 35 289 69 527
rect 103 323 169 493
rect 203 367 237 527
rect 271 323 337 493
rect 371 367 405 527
rect 439 323 505 493
rect 539 367 573 527
rect 707 367 741 527
rect 875 367 909 527
rect 1043 367 1077 527
rect 1211 367 1245 527
rect 1379 367 1413 527
rect 1547 367 1581 527
rect 1715 367 1749 527
rect 1883 367 1917 527
rect 103 289 573 323
rect 538 255 573 289
rect 538 215 1882 255
rect 538 181 573 215
rect 35 17 69 181
rect 103 147 573 181
rect 103 52 169 147
rect 203 17 237 113
rect 271 52 337 147
rect 371 17 405 113
rect 439 52 505 147
rect 539 17 573 113
rect 707 17 741 113
rect 875 17 909 113
rect 1043 17 1077 113
rect 1211 17 1245 113
rect 1379 17 1413 113
rect 1547 17 1581 113
rect 1715 17 1749 113
rect 1883 17 1917 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
rlabel locali s 17 215 497 255 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 1951 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 959 51 993 52 6 X
port 6 nsew signal output
rlabel locali s 791 51 825 52 6 X
port 6 nsew signal output
rlabel locali s 607 51 657 52 6 X
port 6 nsew signal output
rlabel locali s 1952 73 2007 147 6 X
port 6 nsew signal output
rlabel locali s 1783 52 1849 147 6 X
port 6 nsew signal output
rlabel locali s 1615 52 1681 147 6 X
port 6 nsew signal output
rlabel locali s 1447 52 1513 147 6 X
port 6 nsew signal output
rlabel locali s 1279 52 1345 147 6 X
port 6 nsew signal output
rlabel locali s 1111 52 1177 147 6 X
port 6 nsew signal output
rlabel locali s 943 52 1009 147 6 X
port 6 nsew signal output
rlabel locali s 775 52 841 147 6 X
port 6 nsew signal output
rlabel locali s 607 52 673 147 6 X
port 6 nsew signal output
rlabel locali s 607 147 2007 181 6 X
port 6 nsew signal output
rlabel locali s 1931 181 2007 289 6 X
port 6 nsew signal output
rlabel locali s 607 289 2007 323 6 X
port 6 nsew signal output
rlabel locali s 1952 323 2007 472 6 X
port 6 nsew signal output
rlabel locali s 1783 323 1849 493 6 X
port 6 nsew signal output
rlabel locali s 1615 323 1681 493 6 X
port 6 nsew signal output
rlabel locali s 1447 323 1513 493 6 X
port 6 nsew signal output
rlabel locali s 1279 323 1345 493 6 X
port 6 nsew signal output
rlabel locali s 1111 323 1177 493 6 X
port 6 nsew signal output
rlabel locali s 943 323 1009 493 6 X
port 6 nsew signal output
rlabel locali s 775 323 841 493 6 X
port 6 nsew signal output
rlabel locali s 607 323 673 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3140136
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3124628
<< end >>
