magic
tech sky130A
magscale 1 2
timestamp 1654664132
<< nwell >>
rect 30591 9642 30703 9963
rect 30870 9642 30959 9963
<< viali >>
rect 27864 9722 27898 9756
rect 29381 9735 29415 9769
rect 29549 9735 29583 9769
rect 29717 9735 29751 9769
rect 29885 9735 29919 9769
rect 30053 9735 30087 9769
rect 30221 9735 30255 9769
rect 30389 9735 30423 9769
rect 31129 9734 31163 9768
rect 31297 9734 31331 9768
rect 31465 9734 31499 9768
rect 31633 9734 31667 9768
rect 31801 9734 31835 9768
rect 31969 9734 32003 9768
rect 32137 9734 32171 9768
rect 27678 9596 27712 9630
rect 28353 9602 28387 9636
rect 28435 9602 28469 9636
rect 28526 9602 28560 9636
rect 28620 9602 28654 9636
rect 28940 9595 28974 9629
rect 29141 9600 29175 9634
rect 29260 9600 29294 9634
rect 29379 9600 29413 9634
rect 29498 9600 29532 9634
rect 29617 9600 29651 9634
rect 29736 9600 29770 9634
rect 29855 9600 29889 9634
rect 31065 9602 31099 9636
rect 31184 9602 31218 9636
rect 31303 9602 31337 9636
rect 31422 9602 31456 9636
rect 31541 9602 31575 9636
rect 31660 9602 31694 9636
rect 31779 9602 31813 9636
<< metal1 >>
rect 427 13891 785 13911
rect 427 13890 727 13891
rect 427 13838 451 13890
rect 503 13839 727 13890
rect 779 13839 785 13891
rect 503 13838 785 13839
rect 427 13814 785 13838
rect 61150 13149 61394 13227
rect 0 12219 29210 12224
rect 0 12167 29120 12219
rect 29172 12167 29210 12219
rect 0 12163 29210 12167
rect 30969 12216 61648 12221
rect 30969 12164 31007 12216
rect 31059 12164 61648 12216
rect 30969 12160 61648 12164
rect 0 12077 27302 12082
rect 0 12025 27232 12077
rect 27284 12025 27302 12077
rect 0 12021 27302 12025
rect 32877 12074 61648 12079
rect 32877 12022 32895 12074
rect 32947 12022 61648 12074
rect 32877 12018 61648 12022
rect 0 11936 25444 11940
rect 0 11884 25345 11936
rect 25397 11884 25444 11936
rect 0 11879 25444 11884
rect 34735 11933 61648 11937
rect 34735 11881 34782 11933
rect 34834 11881 61648 11933
rect 34735 11876 61648 11881
rect 0 11795 23520 11798
rect 0 11743 23456 11795
rect 23508 11743 23520 11795
rect 0 11737 23520 11743
rect 36659 11792 61648 11795
rect 36659 11740 36671 11792
rect 36723 11740 61648 11792
rect 36659 11734 61648 11740
rect 0 11652 21644 11656
rect 0 11600 21568 11652
rect 21620 11600 21644 11652
rect 0 11595 21644 11600
rect 38535 11649 61648 11653
rect 38535 11597 38559 11649
rect 38611 11597 61648 11649
rect 38535 11592 61648 11597
rect 0 11509 19762 11514
rect 0 11457 19678 11509
rect 19730 11457 19762 11509
rect 0 11453 19762 11457
rect 40417 11506 61648 11511
rect 40417 11454 40449 11506
rect 40501 11454 61648 11506
rect 40417 11450 61648 11454
rect 0 11368 17854 11372
rect 0 11316 17792 11368
rect 17844 11316 17854 11368
rect 0 11311 17854 11316
rect 42325 11365 61648 11369
rect 42325 11313 42335 11365
rect 42387 11313 61648 11365
rect 42325 11308 61648 11313
rect 0 11225 15978 11230
rect 0 11173 15904 11225
rect 15956 11173 15978 11225
rect 0 11169 15978 11173
rect 44201 11222 61648 11227
rect 44201 11170 44223 11222
rect 44275 11170 61648 11222
rect 44201 11166 61648 11170
rect 0 11083 14108 11088
rect 0 11031 14023 11083
rect 14075 11031 14108 11083
rect 0 11027 14108 11031
rect 46071 11080 61648 11085
rect 46071 11028 46104 11080
rect 46156 11028 61648 11080
rect 46071 11024 61648 11028
rect 0 10940 12236 10946
rect 0 10888 12135 10940
rect 12187 10888 12236 10940
rect 0 10885 12236 10888
rect 47943 10937 61648 10943
rect 47943 10885 47992 10937
rect 48044 10885 61648 10937
rect 47943 10882 61648 10885
rect 0 10798 10350 10804
rect 0 10746 10247 10798
rect 10299 10746 10350 10798
rect 0 10743 10350 10746
rect 49829 10800 59808 10801
rect 61176 10800 61648 10801
rect 49829 10795 61648 10800
rect 49829 10743 49880 10795
rect 49932 10743 61648 10795
rect 49829 10740 61648 10743
rect 59711 10739 61648 10740
rect 0 10656 8439 10662
rect 0 10604 8360 10656
rect 8412 10604 8439 10656
rect 0 10601 8439 10604
rect 51740 10653 61648 10659
rect 51740 10601 51767 10653
rect 51819 10601 61648 10653
rect 51740 10598 61648 10601
rect 0 10515 6563 10520
rect 0 10463 6470 10515
rect 6522 10463 6563 10515
rect 0 10459 6563 10463
rect 53616 10512 61648 10517
rect 53616 10460 53657 10512
rect 53709 10460 61648 10512
rect 53616 10456 61648 10460
rect 0 10373 4666 10378
rect 0 10321 4583 10373
rect 4635 10321 4666 10373
rect 0 10317 4666 10321
rect 55513 10370 61648 10375
rect 55513 10318 55544 10370
rect 55596 10318 61648 10370
rect 55513 10314 61648 10318
rect 0 10230 2794 10236
rect 0 10178 2694 10230
rect 2746 10178 2794 10230
rect 0 10175 2794 10178
rect 57385 10227 61648 10233
rect 57385 10175 57433 10227
rect 57485 10175 61648 10227
rect 57385 10172 61648 10175
rect 0 10089 935 10094
rect 0 10037 806 10089
rect 858 10037 935 10089
rect 0 10033 935 10037
rect 59244 10086 61648 10091
rect 59244 10034 59321 10086
rect 59373 10034 61648 10086
rect 59244 10030 61648 10034
rect 0 9947 1157 9952
rect 0 9895 1033 9947
rect 1085 9895 1157 9947
rect 0 9891 1157 9895
rect 28101 9877 28177 9973
rect 29005 9877 29081 9973
rect 30553 9877 30740 9973
rect 30832 9877 31019 9973
rect 59479 9944 61648 9949
rect 59479 9892 59551 9944
rect 59603 9892 61648 9944
rect 59479 9888 61648 9892
rect 0 9808 3016 9810
rect 0 9756 2920 9808
rect 2972 9756 3016 9808
rect 57620 9805 61648 9807
rect 0 9749 3016 9756
rect 27854 9756 27907 9773
rect 27854 9722 27864 9756
rect 27898 9722 27907 9756
rect 0 9663 4927 9668
rect 0 9611 4809 9663
rect 4861 9611 4927 9663
rect 0 9607 4927 9611
rect 7162 9652 7509 9674
rect 7162 9640 27730 9652
rect 7162 9588 7251 9640
rect 7303 9588 7349 9640
rect 7401 9630 27730 9640
rect 7401 9596 27678 9630
rect 27712 9596 27730 9630
rect 7401 9588 27730 9596
rect 27854 9651 27907 9722
rect 29369 9769 32186 9794
rect 29369 9735 29381 9769
rect 29415 9735 29549 9769
rect 29583 9735 29717 9769
rect 29751 9735 29885 9769
rect 29919 9735 30053 9769
rect 30087 9735 30221 9769
rect 30255 9735 30389 9769
rect 30423 9768 32186 9769
rect 30423 9760 31129 9768
rect 30423 9735 30601 9760
rect 29369 9708 30601 9735
rect 30653 9708 30704 9760
rect 30756 9708 30807 9760
rect 30859 9708 30910 9760
rect 30962 9734 31129 9760
rect 31163 9734 31297 9768
rect 31331 9734 31465 9768
rect 31499 9734 31633 9768
rect 31667 9734 31801 9768
rect 31835 9734 31969 9768
rect 32003 9734 32137 9768
rect 32171 9734 32186 9768
rect 57620 9753 57664 9805
rect 57716 9753 61648 9805
rect 57620 9746 61648 9753
rect 30962 9708 32186 9734
rect 29369 9686 32186 9708
rect 55709 9660 61648 9665
rect 27854 9636 28699 9651
rect 27854 9602 28353 9636
rect 28387 9602 28435 9636
rect 28469 9602 28526 9636
rect 28560 9602 28620 9636
rect 28654 9602 28699 9636
rect 27854 9590 28699 9602
rect 28918 9636 32109 9645
rect 28918 9634 31065 9636
rect 28918 9629 29141 9634
rect 28918 9595 28940 9629
rect 28974 9600 29141 9629
rect 29175 9600 29260 9634
rect 29294 9600 29379 9634
rect 29413 9600 29498 9634
rect 29532 9600 29617 9634
rect 29651 9600 29736 9634
rect 29770 9600 29855 9634
rect 29889 9602 31065 9634
rect 31099 9602 31184 9636
rect 31218 9602 31303 9636
rect 31337 9602 31422 9636
rect 31456 9602 31541 9636
rect 31575 9602 31660 9636
rect 31694 9602 31779 9636
rect 31813 9602 32109 9636
rect 55709 9608 55775 9660
rect 55827 9608 61648 9660
rect 55709 9604 61648 9608
rect 29889 9600 32109 9602
rect 28974 9595 32109 9600
rect 28918 9588 32109 9595
rect 7162 9578 27730 9588
rect 7162 9550 7509 9578
rect 0 9522 6773 9526
rect 0 9470 6698 9522
rect 6750 9470 6773 9522
rect 0 9465 6773 9470
rect 53863 9519 61648 9523
rect 53863 9467 53886 9519
rect 53938 9467 61648 9519
rect 53863 9462 61648 9467
rect 0 9378 8664 9384
rect 0 9326 8585 9378
rect 8637 9326 8664 9378
rect 28101 9333 28177 9429
rect 29005 9332 29081 9428
rect 30553 9333 30740 9429
rect 30832 9333 31019 9429
rect 51972 9375 61648 9381
rect 0 9323 8664 9326
rect 51972 9323 51999 9375
rect 52051 9323 61648 9375
rect 51972 9320 61648 9323
rect 0 9237 10552 9242
rect 0 9185 10473 9237
rect 10525 9185 10552 9237
rect 0 9181 10552 9185
rect 50084 9234 61648 9239
rect 50084 9182 50111 9234
rect 50163 9182 61648 9234
rect 50084 9178 61648 9182
rect 0 9095 12453 9100
rect 0 9043 12362 9095
rect 12414 9043 12453 9095
rect 0 9039 12453 9043
rect 48183 9092 61648 9097
rect 48183 9040 48222 9092
rect 48274 9040 61648 9092
rect 48183 9036 61648 9040
rect 0 8950 14328 8958
rect 0 8898 14250 8950
rect 14302 8898 14328 8950
rect 0 8897 14328 8898
rect 46308 8947 61648 8955
rect 46308 8895 46334 8947
rect 46386 8895 61648 8947
rect 46308 8894 61648 8895
rect 0 8811 16239 8816
rect 0 8759 16128 8811
rect 16180 8759 16239 8811
rect 0 8755 16239 8759
rect 44397 8808 61648 8813
rect 44397 8756 44456 8808
rect 44508 8756 61648 8808
rect 44397 8752 61648 8756
rect 0 8670 18137 8674
rect 0 8618 18019 8670
rect 18071 8618 18137 8670
rect 0 8613 18137 8618
rect 42499 8667 61648 8671
rect 42499 8615 42565 8667
rect 42617 8615 61648 8667
rect 42499 8610 61648 8615
rect 0 8529 20044 8532
rect 0 8477 19904 8529
rect 19956 8477 20044 8529
rect 0 8471 20044 8477
rect 40592 8526 61648 8529
rect 40592 8474 40680 8526
rect 40732 8474 61648 8526
rect 40592 8468 61648 8474
rect 0 8386 21894 8390
rect 0 8334 21795 8386
rect 21847 8334 21894 8386
rect 0 8329 21894 8334
rect 38742 8383 61648 8387
rect 38742 8331 38789 8383
rect 38841 8331 61648 8383
rect 38742 8326 61648 8331
rect 0 8243 23769 8248
rect 0 8191 23685 8243
rect 23737 8191 23769 8243
rect 0 8187 23769 8191
rect 36867 8240 61648 8245
rect 36867 8188 36899 8240
rect 36951 8188 61648 8240
rect 36867 8184 61648 8188
rect 0 8099 25666 8106
rect 0 8047 25568 8099
rect 25620 8047 25666 8099
rect 0 8045 25666 8047
rect 34970 8096 61648 8103
rect 34970 8044 35016 8096
rect 35068 8044 61648 8096
rect 34970 8042 61648 8044
rect 0 7957 27596 7964
rect 0 7905 27458 7957
rect 27510 7905 27596 7957
rect 0 7903 27596 7905
rect 33040 7954 61648 7961
rect 33040 7902 33126 7954
rect 33178 7902 61648 7954
rect 33040 7900 61648 7902
rect 0 7817 29446 7822
rect 0 7765 29350 7817
rect 29402 7765 29446 7817
rect 0 7761 29446 7765
rect 31190 7814 61648 7819
rect 31190 7762 31234 7814
rect 31286 7762 61648 7814
rect 31190 7758 61648 7762
rect 174 6112 955 6127
rect 174 6104 896 6112
rect 174 6052 191 6104
rect 243 6060 896 6104
rect 948 6060 955 6112
rect 243 6052 955 6060
rect 174 6034 955 6052
<< via1 >>
rect 30637 15452 30689 15504
rect 30754 15452 30806 15504
rect 30871 15452 30923 15504
rect 451 13838 503 13890
rect 727 13839 779 13891
rect 29120 12167 29172 12219
rect 31007 12164 31059 12216
rect 27232 12025 27284 12077
rect 32895 12022 32947 12074
rect 25345 11884 25397 11936
rect 34782 11881 34834 11933
rect 23456 11743 23508 11795
rect 36671 11740 36723 11792
rect 21568 11600 21620 11652
rect 38559 11597 38611 11649
rect 19678 11457 19730 11509
rect 40449 11454 40501 11506
rect 17792 11316 17844 11368
rect 42335 11313 42387 11365
rect 15904 11173 15956 11225
rect 44223 11170 44275 11222
rect 14023 11031 14075 11083
rect 46104 11028 46156 11080
rect 12135 10888 12187 10940
rect 47992 10885 48044 10937
rect 10247 10746 10299 10798
rect 49880 10743 49932 10795
rect 8360 10604 8412 10656
rect 51767 10601 51819 10653
rect 6470 10463 6522 10515
rect 53657 10460 53709 10512
rect 4583 10321 4635 10373
rect 55544 10318 55596 10370
rect 2694 10178 2746 10230
rect 57433 10175 57485 10227
rect 806 10037 858 10089
rect 59321 10034 59373 10086
rect 1033 9895 1085 9947
rect 31704 9891 31756 9943
rect 31834 9891 31886 9943
rect 31964 9891 32016 9943
rect 59551 9892 59603 9944
rect 2920 9756 2972 9808
rect 4809 9611 4861 9663
rect 7251 9588 7303 9640
rect 7349 9588 7401 9640
rect 30601 9708 30653 9760
rect 30704 9708 30756 9760
rect 30807 9708 30859 9760
rect 30910 9708 30962 9760
rect 57664 9753 57716 9805
rect 55775 9608 55827 9660
rect 6698 9470 6750 9522
rect 53886 9467 53938 9519
rect 8585 9326 8637 9378
rect 31694 9361 31746 9413
rect 31807 9361 31859 9413
rect 31920 9361 31972 9413
rect 32033 9361 32085 9413
rect 32146 9361 32198 9413
rect 51999 9323 52051 9375
rect 10473 9185 10525 9237
rect 50111 9182 50163 9234
rect 12362 9043 12414 9095
rect 48222 9040 48274 9092
rect 14250 8898 14302 8950
rect 46334 8895 46386 8947
rect 16128 8759 16180 8811
rect 44456 8756 44508 8808
rect 18019 8618 18071 8670
rect 42565 8615 42617 8667
rect 19904 8477 19956 8529
rect 40680 8474 40732 8526
rect 21795 8334 21847 8386
rect 38789 8331 38841 8383
rect 23685 8191 23737 8243
rect 36899 8188 36951 8240
rect 25568 8047 25620 8099
rect 35016 8044 35068 8096
rect 27458 7905 27510 7957
rect 33126 7902 33178 7954
rect 29350 7765 29402 7817
rect 31234 7762 31286 7814
rect 31694 7472 31746 7524
rect 31807 7472 31859 7524
rect 31920 7472 31972 7524
rect 32033 7472 32085 7524
rect 32146 7472 32198 7524
rect 31694 7367 31746 7419
rect 31807 7367 31859 7419
rect 31920 7367 31972 7419
rect 32033 7367 32085 7419
rect 32146 7367 32198 7419
rect 191 6052 243 6104
rect 896 6060 948 6112
rect 30626 3223 30678 3275
rect 30709 3223 30761 3275
rect 30792 3223 30844 3275
rect 30875 3223 30927 3275
<< metal2 >>
rect 2180 19017 2224 20184
rect 4068 19017 4112 19992
rect 5956 19017 6000 19992
rect 7844 19017 7888 19992
rect 9732 19017 9776 19992
rect 11620 19017 11664 19992
rect 13508 19017 13552 19992
rect 15396 19017 15440 19992
rect 17284 19017 17328 19992
rect 19172 19017 19216 19992
rect 21060 19017 21104 19992
rect 22948 19017 22992 19992
rect 24836 19017 24880 19992
rect 26724 19017 26768 19992
rect 28612 19017 28656 19992
rect 30500 19017 30544 19992
rect 32388 19017 32432 19992
rect 34276 19017 34320 19992
rect 36164 19017 36208 19992
rect 38052 19017 38096 19992
rect 39940 19017 39984 19992
rect 41828 19017 41872 19992
rect 43716 19017 43760 19992
rect 45604 19017 45648 19992
rect 47492 19017 47536 19992
rect 49380 19017 49424 20151
rect 51268 19017 51312 19992
rect 53156 19017 53200 19992
rect 55044 19017 55088 19992
rect 56932 19017 56976 19992
rect 58820 19017 58864 19992
rect 60708 19017 60752 19992
rect 61283 18335 61319 18368
rect 182 18299 896 18335
rect 60572 18299 61319 18335
rect 182 6127 218 18299
rect 30573 15559 30969 15588
rect 30573 15503 30604 15559
rect 30660 15504 30713 15559
rect 30769 15504 30822 15559
rect 30878 15504 30969 15559
rect 30689 15503 30713 15504
rect 30806 15503 30822 15504
rect 30573 15457 30637 15503
rect 30689 15457 30754 15503
rect 30806 15457 30871 15503
rect 30573 15401 30604 15457
rect 30689 15452 30713 15457
rect 30806 15452 30822 15457
rect 30923 15452 30969 15504
rect 30660 15401 30713 15452
rect 30769 15401 30822 15452
rect 30878 15401 30969 15452
rect 30573 15380 30969 15401
rect 416 13890 514 13917
rect 416 13838 451 13890
rect 503 13838 514 13890
rect 416 13798 514 13838
rect 714 13891 818 13914
rect 714 13839 727 13891
rect 779 13879 818 13891
rect 61283 13879 61319 18299
rect 779 13843 990 13879
rect 60666 13843 61319 13879
rect 779 13839 818 13843
rect 714 13814 818 13839
rect 181 6104 292 6127
rect 181 6052 191 6104
rect 243 6052 292 6104
rect 181 6012 292 6052
rect 448 1648 484 13798
rect 810 10099 854 13161
rect 2698 10242 2742 13161
rect 4586 10382 4630 13161
rect 6474 10526 6518 13161
rect 8362 10666 8406 13161
rect 10250 10808 10294 12753
rect 12138 10950 12182 12773
rect 14026 11092 14070 12763
rect 15908 11233 15952 12770
rect 17796 11374 17840 12823
rect 19684 11519 19728 12763
rect 21572 11662 21616 12743
rect 23460 11804 23504 12743
rect 25348 11945 25392 12703
rect 27236 12088 27280 12747
rect 29124 12234 29168 12757
rect 29101 12219 29195 12234
rect 31011 12231 31055 12596
rect 29101 12167 29120 12219
rect 29172 12167 29195 12219
rect 29101 12153 29195 12167
rect 30984 12216 31078 12231
rect 30984 12164 31007 12216
rect 31059 12164 31078 12216
rect 29124 12109 29168 12153
rect 30984 12150 31078 12164
rect 31011 12106 31055 12150
rect 27221 12077 27298 12088
rect 32899 12085 32943 12617
rect 27221 12025 27232 12077
rect 27284 12025 27298 12077
rect 27221 12015 27298 12025
rect 32881 12074 32958 12085
rect 32881 12022 32895 12074
rect 32947 12022 32958 12074
rect 27236 11972 27280 12015
rect 32881 12012 32958 12022
rect 32899 11969 32943 12012
rect 25332 11936 25409 11945
rect 34787 11942 34831 12673
rect 25332 11884 25345 11936
rect 25397 11884 25409 11936
rect 25332 11872 25409 11884
rect 34770 11933 34847 11942
rect 34770 11881 34782 11933
rect 34834 11881 34847 11933
rect 25348 11842 25392 11872
rect 34770 11869 34847 11881
rect 34787 11839 34831 11869
rect 23445 11795 23522 11804
rect 36675 11801 36719 12598
rect 23445 11743 23456 11795
rect 23508 11743 23522 11795
rect 23445 11731 23522 11743
rect 36657 11792 36734 11801
rect 36657 11740 36671 11792
rect 36723 11740 36734 11792
rect 23460 11695 23504 11731
rect 36657 11728 36734 11740
rect 36675 11692 36719 11728
rect 21556 11652 21633 11662
rect 38563 11659 38607 12608
rect 21556 11600 21568 11652
rect 21620 11600 21633 11652
rect 21556 11589 21633 11600
rect 38546 11649 38623 11659
rect 38546 11597 38559 11649
rect 38611 11597 38623 11649
rect 21572 11555 21616 11589
rect 38546 11586 38623 11597
rect 38563 11552 38607 11586
rect 19670 11509 19747 11519
rect 40451 11516 40495 12636
rect 19670 11457 19678 11509
rect 19730 11457 19747 11509
rect 19670 11446 19747 11457
rect 40432 11506 40509 11516
rect 40432 11454 40449 11506
rect 40501 11454 40509 11506
rect 19684 11404 19728 11446
rect 40432 11443 40509 11454
rect 40451 11401 40495 11443
rect 17779 11368 17856 11374
rect 42339 11371 42383 12629
rect 17779 11316 17792 11368
rect 17844 11316 17856 11368
rect 17779 11301 17856 11316
rect 42323 11365 42400 11371
rect 42323 11313 42335 11365
rect 42387 11313 42400 11365
rect 17796 11258 17840 11301
rect 42323 11298 42400 11313
rect 42339 11255 42383 11298
rect 15892 11225 15969 11233
rect 44227 11230 44271 12627
rect 15892 11173 15904 11225
rect 15956 11173 15969 11225
rect 15892 11160 15969 11173
rect 44210 11222 44287 11230
rect 44210 11170 44223 11222
rect 44275 11170 44287 11222
rect 15908 11131 15952 11160
rect 44210 11157 44287 11170
rect 44227 11128 44271 11157
rect 14011 11083 14088 11092
rect 46109 11089 46153 12595
rect 14011 11031 14023 11083
rect 14075 11031 14088 11083
rect 14011 11019 14088 11031
rect 46091 11080 46168 11089
rect 46091 11028 46104 11080
rect 46156 11028 46168 11080
rect 14026 10991 14070 11019
rect 46091 11016 46168 11028
rect 46109 10988 46153 11016
rect 12123 10940 12200 10950
rect 47997 10947 48041 12633
rect 12123 10888 12135 10940
rect 12187 10888 12200 10940
rect 12123 10877 12200 10888
rect 47979 10937 48056 10947
rect 47979 10885 47992 10937
rect 48044 10885 48056 10937
rect 12138 10854 12182 10877
rect 47979 10874 48056 10885
rect 47997 10851 48041 10874
rect 10234 10798 10311 10808
rect 49885 10805 49929 12618
rect 10234 10746 10247 10798
rect 10299 10746 10311 10798
rect 10234 10735 10311 10746
rect 49868 10795 49945 10805
rect 49868 10743 49880 10795
rect 49932 10743 49945 10795
rect 10250 10697 10294 10735
rect 49868 10732 49945 10743
rect 49885 10694 49929 10732
rect 8348 10656 8425 10666
rect 51773 10663 51817 12618
rect 8348 10604 8360 10656
rect 8412 10604 8425 10656
rect 8348 10593 8425 10604
rect 51754 10653 51831 10663
rect 51754 10601 51767 10653
rect 51819 10601 51831 10653
rect 8362 10560 8406 10593
rect 51754 10590 51831 10601
rect 51773 10557 51817 10590
rect 6460 10515 6537 10526
rect 53661 10523 53705 12631
rect 6460 10463 6470 10515
rect 6522 10463 6537 10515
rect 6460 10453 6537 10463
rect 53642 10512 53719 10523
rect 53642 10460 53657 10512
rect 53709 10460 53719 10512
rect 6474 10417 6518 10453
rect 53642 10450 53719 10460
rect 4570 10373 4647 10382
rect 4570 10321 4583 10373
rect 4635 10321 4647 10373
rect 4570 10309 4647 10321
rect 30574 10377 30971 10416
rect 53661 10414 53705 10450
rect 55549 10379 55593 12648
rect 30574 10321 30597 10377
rect 30653 10321 30701 10377
rect 30757 10321 30805 10377
rect 30861 10321 30909 10377
rect 30965 10321 30971 10377
rect 4586 10270 4630 10309
rect 30574 10278 30971 10321
rect 55532 10370 55609 10379
rect 55532 10318 55544 10370
rect 55596 10318 55609 10370
rect 55532 10306 55609 10318
rect 2686 10230 2763 10242
rect 2686 10178 2694 10230
rect 2746 10178 2763 10230
rect 2686 10169 2763 10178
rect 30574 10222 30597 10278
rect 30653 10222 30701 10278
rect 30757 10222 30805 10278
rect 30861 10222 30909 10278
rect 30965 10222 30971 10278
rect 55549 10267 55593 10306
rect 57437 10239 57481 12646
rect 2698 10133 2742 10169
rect 793 10089 870 10099
rect 793 10037 806 10089
rect 858 10037 870 10089
rect 793 10026 870 10037
rect 810 10003 854 10026
rect 1039 9958 1083 9988
rect 1022 9947 1101 9958
rect 1022 9895 1033 9947
rect 1085 9895 1101 9947
rect 1022 9882 1101 9895
rect 1039 7250 1083 9882
rect 2927 9817 2971 9861
rect 2908 9808 2987 9817
rect 2908 9756 2920 9808
rect 2972 9756 2987 9808
rect 2908 9741 2987 9756
rect 30574 9760 30971 10222
rect 57416 10227 57493 10239
rect 57416 10175 57433 10227
rect 57485 10175 57493 10227
rect 57416 10166 57493 10175
rect 57437 10130 57481 10166
rect 59325 10096 59369 12644
rect 59309 10086 59386 10096
rect 59309 10034 59321 10086
rect 59373 10034 59386 10086
rect 59309 10023 59386 10034
rect 59325 10000 59369 10023
rect 31665 9947 32066 9972
rect 59553 9955 59597 9985
rect 31665 9891 31704 9947
rect 31760 9891 31833 9947
rect 31889 9891 31962 9947
rect 32018 9891 32066 9947
rect 31665 9878 32066 9891
rect 59535 9944 59614 9955
rect 59535 9892 59551 9944
rect 59603 9892 59614 9944
rect 59535 9879 59614 9892
rect 57665 9814 57709 9858
rect 2927 7204 2971 9741
rect 4815 9671 4859 9744
rect 30574 9708 30601 9760
rect 30653 9708 30704 9760
rect 30756 9708 30807 9760
rect 30859 9708 30910 9760
rect 30962 9708 30971 9760
rect 57649 9805 57728 9814
rect 57649 9753 57664 9805
rect 57716 9753 57728 9805
rect 4790 9663 4869 9671
rect 4790 9611 4809 9663
rect 4861 9611 4869 9663
rect 4790 9595 4869 9611
rect 7162 9644 7509 9674
rect 7162 9640 7252 9644
rect 4815 7167 4859 9595
rect 6703 9530 6747 9604
rect 7162 9588 7251 9640
rect 7308 9588 7349 9644
rect 7405 9588 7509 9644
rect 7162 9550 7509 9588
rect 6685 9522 6764 9530
rect 6685 9470 6698 9522
rect 6750 9470 6764 9522
rect 6685 9454 6764 9470
rect 6703 7216 6747 9454
rect 8591 9389 8635 9438
rect 8574 9378 8653 9389
rect 8574 9326 8585 9378
rect 8637 9326 8653 9378
rect 8574 9313 8653 9326
rect 8591 7253 8635 9313
rect 10479 9247 10523 9292
rect 10462 9237 10541 9247
rect 10462 9185 10473 9237
rect 10525 9185 10541 9237
rect 10462 9171 10541 9185
rect 10479 7216 10523 9171
rect 12367 9104 12411 9145
rect 12351 9095 12430 9104
rect 12351 9043 12362 9095
rect 12414 9043 12430 9095
rect 12351 9028 12430 9043
rect 30574 9048 30971 9708
rect 55777 9668 55821 9741
rect 57649 9738 57728 9753
rect 55767 9660 55846 9668
rect 55767 9608 55775 9660
rect 55827 9608 55846 9660
rect 53889 9527 53933 9601
rect 55767 9592 55846 9608
rect 53872 9519 53951 9527
rect 53872 9467 53886 9519
rect 53938 9467 53951 9519
rect 53872 9451 53951 9467
rect 12367 7192 12411 9028
rect 30574 8992 30610 9048
rect 30666 8992 30698 9048
rect 30754 8992 30786 9048
rect 30842 8992 30874 9048
rect 30930 8992 30971 9048
rect 14255 8959 14299 8986
rect 14239 8950 14318 8959
rect 14239 8898 14250 8950
rect 14302 8898 14318 8950
rect 14239 8883 14318 8898
rect 30574 8953 30971 8992
rect 30574 8897 30610 8953
rect 30666 8897 30698 8953
rect 30754 8897 30786 8953
rect 30842 8897 30874 8953
rect 30930 8897 30971 8953
rect 14255 7216 14299 8883
rect 30574 8866 30971 8897
rect 31639 9413 32306 9430
rect 31639 9361 31694 9413
rect 31746 9361 31807 9413
rect 31859 9361 31920 9413
rect 31972 9361 32033 9413
rect 32085 9361 32146 9413
rect 32198 9361 32306 9413
rect 52001 9386 52045 9435
rect 16137 8821 16181 8863
rect 16117 8811 16196 8821
rect 16117 8759 16128 8811
rect 16180 8759 16196 8811
rect 16117 8745 16196 8759
rect 16137 7161 16181 8745
rect 18025 8679 18069 8735
rect 18007 8670 18086 8679
rect 18007 8618 18019 8670
rect 18071 8618 18086 8670
rect 18007 8603 18086 8618
rect 18025 7192 18069 8603
rect 19913 8538 19957 8594
rect 19893 8529 19972 8538
rect 19893 8477 19904 8529
rect 19956 8477 19972 8529
rect 19893 8462 19972 8477
rect 19913 7234 19957 8462
rect 21801 8396 21845 8453
rect 21783 8386 21862 8396
rect 21783 8334 21795 8386
rect 21847 8334 21862 8386
rect 21783 8320 21862 8334
rect 21801 7210 21845 8320
rect 23689 8253 23733 8319
rect 23673 8243 23752 8253
rect 23673 8191 23685 8243
rect 23737 8191 23752 8243
rect 23673 8177 23752 8191
rect 23689 7161 23733 8177
rect 25577 8112 25621 8166
rect 25555 8099 25634 8112
rect 25555 8047 25568 8099
rect 25620 8047 25634 8099
rect 25555 8036 25634 8047
rect 25577 7192 25621 8036
rect 27465 7970 27509 8007
rect 27449 7957 27528 7970
rect 27449 7905 27458 7957
rect 27510 7905 27528 7957
rect 27449 7894 27528 7905
rect 27465 7192 27509 7894
rect 29353 7828 29397 7903
rect 29339 7817 29418 7828
rect 31239 7825 31283 7900
rect 29339 7765 29350 7817
rect 29402 7765 29418 7817
rect 29339 7752 29418 7765
rect 31218 7814 31297 7825
rect 31218 7762 31234 7814
rect 31286 7762 31297 7814
rect 29353 7198 29397 7752
rect 31218 7749 31297 7762
rect 31239 7293 31283 7749
rect 31639 7524 32306 9361
rect 51983 9375 52062 9386
rect 51983 9323 51999 9375
rect 52051 9323 52062 9375
rect 51983 9310 52062 9323
rect 50113 9244 50157 9289
rect 50095 9234 50174 9244
rect 50095 9182 50111 9234
rect 50163 9182 50174 9234
rect 50095 9168 50174 9182
rect 48225 9101 48269 9142
rect 48206 9092 48285 9101
rect 48206 9040 48222 9092
rect 48274 9040 48285 9092
rect 48206 9025 48285 9040
rect 46337 8956 46381 8983
rect 46318 8947 46397 8956
rect 46318 8895 46334 8947
rect 46386 8895 46397 8947
rect 46318 8880 46397 8895
rect 44455 8818 44499 8860
rect 44440 8808 44519 8818
rect 44440 8756 44456 8808
rect 44508 8756 44519 8808
rect 44440 8742 44519 8756
rect 42567 8676 42611 8732
rect 42550 8667 42629 8676
rect 42550 8615 42565 8667
rect 42617 8615 42629 8667
rect 42550 8600 42629 8615
rect 40679 8535 40723 8591
rect 40664 8526 40743 8535
rect 40664 8474 40680 8526
rect 40732 8474 40743 8526
rect 40664 8459 40743 8474
rect 38791 8393 38835 8450
rect 38774 8383 38853 8393
rect 38774 8331 38789 8383
rect 38841 8331 38853 8383
rect 38774 8317 38853 8331
rect 36903 8250 36947 8316
rect 36884 8240 36963 8250
rect 36884 8188 36899 8240
rect 36951 8188 36963 8240
rect 36884 8174 36963 8188
rect 35015 8109 35059 8163
rect 35002 8096 35081 8109
rect 35002 8044 35016 8096
rect 35068 8044 35081 8096
rect 35002 8033 35081 8044
rect 33127 7967 33171 8004
rect 33108 7954 33187 7967
rect 33108 7902 33126 7954
rect 33178 7902 33187 7954
rect 33108 7891 33187 7902
rect 31639 7472 31694 7524
rect 31746 7472 31807 7524
rect 31859 7472 31920 7524
rect 31972 7472 32033 7524
rect 32085 7472 32146 7524
rect 32198 7472 32306 7524
rect 31639 7419 32306 7472
rect 31639 7367 31694 7419
rect 31746 7367 31807 7419
rect 31859 7367 31920 7419
rect 31972 7367 32033 7419
rect 32085 7367 32146 7419
rect 32198 7367 32306 7419
rect 31639 7319 32306 7367
rect 33127 7340 33171 7891
rect 35015 7302 35059 8033
rect 36903 7299 36947 8174
rect 38791 7293 38835 8317
rect 40679 7319 40723 8459
rect 42567 7244 42611 8600
rect 44455 7287 44499 8742
rect 46337 7306 46381 8880
rect 48225 7270 48269 9025
rect 50113 7259 50157 9168
rect 52001 7285 52045 9310
rect 53889 7310 53933 9451
rect 55777 7268 55821 9592
rect 57665 7329 57709 9738
rect 59553 7299 59597 9879
rect 889 6112 959 6133
rect 889 6060 896 6112
rect 948 6104 959 6112
rect 948 6068 1219 6104
rect 60895 6068 61620 6104
rect 948 6060 959 6068
rect 889 6029 959 6060
rect 30574 3324 30971 3357
rect 30574 3268 30615 3324
rect 30671 3275 30707 3324
rect 30763 3275 30799 3324
rect 30855 3275 30891 3324
rect 30678 3268 30707 3275
rect 30763 3268 30792 3275
rect 30855 3268 30875 3275
rect 30947 3268 30971 3324
rect 30574 3233 30626 3268
rect 30678 3233 30709 3268
rect 30761 3233 30792 3268
rect 30844 3233 30875 3268
rect 30927 3233 30971 3268
rect 30574 3177 30615 3233
rect 30678 3223 30707 3233
rect 30763 3223 30792 3233
rect 30855 3223 30875 3233
rect 30671 3177 30707 3223
rect 30763 3177 30799 3223
rect 30855 3177 30891 3223
rect 30947 3177 30971 3233
rect 30574 3151 30971 3177
rect 61584 1648 61620 6068
rect 448 1612 1125 1648
rect 60801 1612 61620 1648
rect 61584 1601 61620 1612
rect 2409 0 2465 930
rect 4297 0 4353 930
rect 6185 0 6241 930
rect 8073 0 8129 930
rect 9961 0 10017 930
rect 11849 0 11905 930
rect 13737 0 13793 930
rect 15625 0 15681 930
rect 17513 0 17569 930
rect 19401 0 19457 930
rect 21289 0 21345 930
rect 23177 0 23233 930
rect 25065 0 25121 930
rect 26953 0 27009 930
rect 28841 0 28897 930
rect 30729 0 30785 930
rect 32617 0 32673 930
rect 34505 0 34561 930
rect 36393 0 36449 930
rect 38281 0 38337 930
rect 40169 0 40225 930
rect 42057 0 42113 930
rect 43945 0 44001 930
rect 45833 0 45889 930
rect 47721 0 47777 930
rect 49609 0 49665 930
rect 51497 0 51553 930
rect 53385 0 53441 930
rect 55273 0 55329 930
rect 57161 0 57217 930
rect 59049 0 59105 930
rect 60937 0 60993 930
<< via2 >>
rect 30604 15504 30660 15559
rect 30713 15504 30769 15559
rect 30822 15504 30878 15559
rect 30604 15503 30637 15504
rect 30637 15503 30660 15504
rect 30713 15503 30754 15504
rect 30754 15503 30769 15504
rect 30822 15503 30871 15504
rect 30871 15503 30878 15504
rect 30604 15452 30637 15457
rect 30637 15452 30660 15457
rect 30713 15452 30754 15457
rect 30754 15452 30769 15457
rect 30822 15452 30871 15457
rect 30871 15452 30878 15457
rect 30604 15401 30660 15452
rect 30713 15401 30769 15452
rect 30822 15401 30878 15452
rect 30597 10321 30653 10377
rect 30701 10321 30757 10377
rect 30805 10321 30861 10377
rect 30909 10321 30965 10377
rect 30597 10222 30653 10278
rect 30701 10222 30757 10278
rect 30805 10222 30861 10278
rect 30909 10222 30965 10278
rect 31704 9943 31760 9947
rect 31704 9891 31756 9943
rect 31756 9891 31760 9943
rect 31833 9943 31889 9947
rect 31833 9891 31834 9943
rect 31834 9891 31886 9943
rect 31886 9891 31889 9943
rect 31962 9943 32018 9947
rect 31962 9891 31964 9943
rect 31964 9891 32016 9943
rect 32016 9891 32018 9943
rect 7252 9640 7308 9644
rect 7252 9588 7303 9640
rect 7303 9588 7308 9640
rect 7349 9640 7405 9644
rect 7349 9588 7401 9640
rect 7401 9588 7405 9640
rect 30610 8992 30666 9048
rect 30698 8992 30754 9048
rect 30786 8992 30842 9048
rect 30874 8992 30930 9048
rect 30610 8897 30666 8953
rect 30698 8897 30754 8953
rect 30786 8897 30842 8953
rect 30874 8897 30930 8953
rect 30615 3275 30671 3324
rect 30707 3275 30763 3324
rect 30799 3275 30855 3324
rect 30891 3275 30947 3324
rect 30615 3268 30626 3275
rect 30626 3268 30671 3275
rect 30707 3268 30709 3275
rect 30709 3268 30761 3275
rect 30761 3268 30763 3275
rect 30799 3268 30844 3275
rect 30844 3268 30855 3275
rect 30891 3268 30927 3275
rect 30927 3268 30947 3275
rect 30615 3223 30626 3233
rect 30626 3223 30671 3233
rect 30707 3223 30709 3233
rect 30709 3223 30761 3233
rect 30761 3223 30763 3233
rect 30799 3223 30844 3233
rect 30844 3223 30855 3233
rect 30891 3223 30927 3233
rect 30927 3223 30947 3233
rect 30615 3177 30671 3223
rect 30707 3177 30763 3223
rect 30799 3177 30855 3223
rect 30891 3177 30947 3223
<< metal3 >>
rect 30573 15559 30968 15588
rect 30573 15503 30604 15559
rect 30660 15536 30713 15559
rect 30769 15503 30822 15559
rect 30878 15503 30968 15559
rect 30573 15457 30647 15503
rect 30743 15457 30968 15503
rect 30573 15401 30604 15457
rect 30660 15401 30713 15428
rect 30769 15401 30822 15457
rect 30878 15401 30968 15457
rect 30573 15380 30968 15401
rect 30573 10377 30970 10419
rect 30573 10321 30597 10377
rect 30653 10352 30701 10377
rect 30757 10321 30805 10377
rect 30861 10352 30909 10377
rect 30965 10321 30970 10377
rect 30573 10278 30638 10321
rect 30734 10278 30820 10321
rect 30916 10278 30970 10321
rect 30573 10222 30597 10278
rect 30653 10222 30701 10244
rect 30757 10222 30805 10278
rect 30861 10222 30909 10244
rect 30965 10222 30970 10278
rect 30573 10195 30970 10222
rect 31665 9961 32066 9972
rect 31665 9947 31786 9961
rect 31960 9947 32066 9961
rect 31665 9891 31704 9947
rect 31760 9897 31786 9947
rect 31960 9897 31962 9947
rect 31760 9891 31833 9897
rect 31889 9891 31962 9897
rect 32018 9891 32066 9947
rect 31665 9878 32066 9891
rect 7162 9660 7509 9674
rect 61 9644 7509 9660
rect 61 9588 7252 9644
rect 7308 9588 7349 9644
rect 7405 9588 7509 9644
rect 61 9570 7509 9588
rect 7162 9550 7509 9570
rect 30574 9048 30971 9106
rect 30574 8992 30610 9048
rect 30666 9029 30698 9048
rect 30754 8992 30786 9048
rect 30842 9029 30874 9048
rect 30930 8992 30971 9048
rect 30574 8953 30630 8992
rect 30726 8953 30820 8992
rect 30916 8953 30971 8992
rect 30574 8897 30610 8953
rect 30666 8897 30698 8921
rect 30754 8897 30786 8953
rect 30842 8897 30874 8921
rect 30930 8897 30971 8953
rect 30574 8866 30971 8897
rect 30574 3324 30971 3357
rect 30574 3268 30615 3324
rect 30671 3300 30707 3324
rect 30763 3268 30799 3324
rect 30855 3301 30891 3324
rect 30947 3268 30971 3324
rect 30574 3233 30642 3268
rect 30738 3233 30816 3268
rect 30912 3233 30971 3268
rect 30574 3177 30615 3233
rect 30671 3177 30707 3192
rect 30763 3177 30799 3233
rect 30855 3177 30891 3193
rect 30947 3177 30971 3233
rect 30574 3151 30971 3177
<< via3 >>
rect 20135 19603 20241 19781
rect 20309 19603 20415 19781
rect 20483 19603 20589 19781
rect 35110 19580 35216 19758
rect 35293 19580 35399 19758
rect 35476 19580 35582 19758
rect 50608 19593 50714 19771
rect 50791 19593 50897 19771
rect 50974 19593 51080 19771
rect 18612 17459 18718 17637
rect 18786 17459 18892 17637
rect 18960 17459 19066 17637
rect 33589 17464 33695 17642
rect 33772 17464 33878 17642
rect 33955 17464 34061 17642
rect 49083 17455 49189 17633
rect 49266 17455 49372 17633
rect 49449 17455 49555 17633
rect 30647 15503 30660 15536
rect 30660 15503 30713 15536
rect 30713 15503 30743 15536
rect 30647 15457 30743 15503
rect 30647 15428 30660 15457
rect 30660 15428 30713 15457
rect 30713 15428 30743 15457
rect 18625 14531 18731 14709
rect 18799 14531 18905 14709
rect 18973 14531 19079 14709
rect 31710 14534 31834 14700
rect 31909 14534 32033 14700
rect 33575 14529 33681 14707
rect 33758 14529 33864 14707
rect 33941 14529 34047 14707
rect 49114 14526 49220 14704
rect 49297 14526 49403 14704
rect 49480 14526 49586 14704
rect 20135 12395 20241 12573
rect 20309 12395 20415 12573
rect 20483 12395 20589 12573
rect 35125 12406 35231 12584
rect 35308 12406 35414 12584
rect 35491 12406 35597 12584
rect 50583 12397 50689 12575
rect 50766 12397 50872 12575
rect 50949 12397 51055 12575
rect 30638 10321 30653 10352
rect 30653 10321 30701 10352
rect 30701 10321 30734 10352
rect 30820 10321 30861 10352
rect 30861 10321 30909 10352
rect 30909 10321 30916 10352
rect 30638 10278 30734 10321
rect 30820 10278 30916 10321
rect 30638 10244 30653 10278
rect 30653 10244 30701 10278
rect 30701 10244 30734 10278
rect 30820 10244 30861 10278
rect 30861 10244 30909 10278
rect 30909 10244 30916 10278
rect 31786 9947 31960 9961
rect 31786 9897 31833 9947
rect 31833 9897 31889 9947
rect 31889 9897 31960 9947
rect 30630 8992 30666 9029
rect 30666 8992 30698 9029
rect 30698 8992 30726 9029
rect 30820 8992 30842 9029
rect 30842 8992 30874 9029
rect 30874 8992 30916 9029
rect 30630 8953 30726 8992
rect 30820 8953 30916 8992
rect 30630 8921 30666 8953
rect 30666 8921 30698 8953
rect 30698 8921 30726 8953
rect 30820 8921 30842 8953
rect 30842 8921 30874 8953
rect 30874 8921 30916 8953
rect 3333 7354 3439 7532
rect 3584 7354 3690 7532
rect 3835 7354 3941 7532
rect 20113 7357 20219 7535
rect 20287 7357 20393 7535
rect 20461 7357 20567 7535
rect 35080 7364 35186 7542
rect 35263 7364 35369 7542
rect 35446 7364 35552 7542
rect 50585 7356 50691 7534
rect 50768 7356 50874 7534
rect 50951 7356 51057 7534
rect 2108 5225 2214 5403
rect 2284 5225 2390 5403
rect 2460 5225 2566 5403
rect 18611 5231 18717 5409
rect 18785 5231 18891 5409
rect 18959 5231 19065 5409
rect 33587 5232 33693 5410
rect 33770 5232 33876 5410
rect 33953 5232 34059 5410
rect 49082 5228 49188 5406
rect 49265 5228 49371 5406
rect 49448 5228 49554 5406
rect 30642 3268 30671 3300
rect 30671 3268 30707 3300
rect 30707 3268 30738 3300
rect 30816 3268 30855 3301
rect 30855 3268 30891 3301
rect 30891 3268 30912 3301
rect 30642 3233 30738 3268
rect 30816 3233 30912 3268
rect 30642 3192 30671 3233
rect 30671 3192 30707 3233
rect 30707 3192 30738 3233
rect 30816 3193 30855 3233
rect 30855 3193 30891 3233
rect 30891 3193 30912 3233
rect 2104 2292 2210 2470
rect 2280 2292 2386 2470
rect 2456 2292 2562 2470
rect 18608 2295 18714 2473
rect 18782 2295 18888 2473
rect 18956 2295 19062 2473
rect 33599 2291 33705 2469
rect 33782 2291 33888 2469
rect 33965 2291 34071 2469
rect 49090 2295 49196 2473
rect 49273 2295 49379 2473
rect 49456 2295 49562 2473
rect 3367 170 3473 348
rect 3618 170 3724 348
rect 3869 170 3975 348
rect 20117 173 20223 351
rect 20291 173 20397 351
rect 20465 173 20571 351
rect 35126 184 35232 362
rect 35309 184 35415 362
rect 35492 184 35598 362
rect 50626 176 50732 354
rect 50809 176 50915 354
rect 50992 176 51098 354
<< metal4 >>
rect 2024 5403 2642 20087
rect 2024 5225 2108 5403
rect 2214 5225 2284 5403
rect 2390 5225 2460 5403
rect 2566 5225 2642 5403
rect 2024 2470 2642 5225
rect 2024 2292 2104 2470
rect 2210 2292 2280 2470
rect 2386 2292 2456 2470
rect 2562 2292 2642 2470
rect 2024 38 2642 2292
rect 3257 7532 4041 20087
rect 3257 7354 3333 7532
rect 3439 7354 3584 7532
rect 3690 7354 3835 7532
rect 3941 7354 4041 7532
rect 3257 348 4041 7354
rect 3257 170 3367 348
rect 3473 170 3618 348
rect 3724 170 3869 348
rect 3975 170 4041 348
rect 3257 74 4041 170
rect 18524 17637 19142 20087
rect 18524 17459 18612 17637
rect 18718 17459 18786 17637
rect 18892 17459 18960 17637
rect 19066 17459 19142 17637
rect 18524 14709 19142 17459
rect 18524 14531 18625 14709
rect 18731 14531 18799 14709
rect 18905 14531 18973 14709
rect 19079 14531 19142 14709
rect 18524 5409 19142 14531
rect 18524 5231 18611 5409
rect 18717 5231 18785 5409
rect 18891 5231 18959 5409
rect 19065 5231 19142 5409
rect 18524 2473 19142 5231
rect 18524 2295 18608 2473
rect 18714 2295 18782 2473
rect 18888 2295 18956 2473
rect 19062 2295 19142 2473
rect 18524 38 19142 2295
rect 20024 19781 20642 20087
rect 20024 19603 20135 19781
rect 20241 19603 20309 19781
rect 20415 19603 20483 19781
rect 20589 19603 20642 19781
rect 20024 12573 20642 19603
rect 33524 17642 34142 20087
rect 33524 17464 33589 17642
rect 33695 17464 33772 17642
rect 33878 17464 33955 17642
rect 34061 17464 34142 17642
rect 20024 12395 20135 12573
rect 20241 12395 20309 12573
rect 20415 12395 20483 12573
rect 20589 12395 20642 12573
rect 20024 7535 20642 12395
rect 30573 15536 30970 15648
rect 30573 15428 30647 15536
rect 30743 15428 30970 15536
rect 30573 10856 30970 15428
rect 30572 10495 30970 10856
rect 30573 10352 30970 10495
rect 30573 10244 30638 10352
rect 30734 10244 30820 10352
rect 30916 10244 30970 10352
rect 30573 10195 30970 10244
rect 31658 14700 32062 14819
rect 31658 14534 31710 14700
rect 31834 14534 31909 14700
rect 32033 14534 32062 14700
rect 31658 9989 32062 14534
rect 33524 14707 34142 17464
rect 33524 14529 33575 14707
rect 33681 14529 33758 14707
rect 33864 14529 33941 14707
rect 34047 14529 34142 14707
rect 31658 9967 32066 9989
rect 31665 9961 32066 9967
rect 31665 9897 31786 9961
rect 31960 9897 32066 9961
rect 31665 9878 32066 9897
rect 20024 7357 20113 7535
rect 20219 7357 20287 7535
rect 20393 7357 20461 7535
rect 20567 7357 20642 7535
rect 20024 351 20642 7357
rect 30575 9029 30971 9105
rect 30575 8921 30630 9029
rect 30726 8921 30820 9029
rect 30916 8921 30971 9029
rect 30575 3301 30971 8921
rect 30575 3300 30816 3301
rect 30575 3192 30642 3300
rect 30738 3193 30816 3300
rect 30912 3193 30971 3301
rect 30738 3192 30971 3193
rect 30575 3089 30971 3192
rect 33524 5410 34142 14529
rect 33524 5232 33587 5410
rect 33693 5232 33770 5410
rect 33876 5232 33953 5410
rect 34059 5232 34142 5410
rect 20024 173 20117 351
rect 20223 173 20291 351
rect 20397 173 20465 351
rect 20571 173 20642 351
rect 20024 38 20642 173
rect 33524 2469 34142 5232
rect 33524 2291 33599 2469
rect 33705 2291 33782 2469
rect 33888 2291 33965 2469
rect 34071 2291 34142 2469
rect 33524 38 34142 2291
rect 35024 19758 35642 20087
rect 35024 19580 35110 19758
rect 35216 19580 35293 19758
rect 35399 19580 35476 19758
rect 35582 19580 35642 19758
rect 35024 12584 35642 19580
rect 35024 12406 35125 12584
rect 35231 12406 35308 12584
rect 35414 12406 35491 12584
rect 35597 12406 35642 12584
rect 35024 7542 35642 12406
rect 35024 7364 35080 7542
rect 35186 7364 35263 7542
rect 35369 7364 35446 7542
rect 35552 7364 35642 7542
rect 35024 362 35642 7364
rect 35024 184 35126 362
rect 35232 184 35309 362
rect 35415 184 35492 362
rect 35598 184 35642 362
rect 35024 38 35642 184
rect 49024 17633 49642 20087
rect 49024 17455 49083 17633
rect 49189 17455 49266 17633
rect 49372 17455 49449 17633
rect 49555 17455 49642 17633
rect 49024 14704 49642 17455
rect 49024 14526 49114 14704
rect 49220 14526 49297 14704
rect 49403 14526 49480 14704
rect 49586 14526 49642 14704
rect 49024 5406 49642 14526
rect 49024 5228 49082 5406
rect 49188 5228 49265 5406
rect 49371 5228 49448 5406
rect 49554 5228 49642 5406
rect 49024 2473 49642 5228
rect 49024 2295 49090 2473
rect 49196 2295 49273 2473
rect 49379 2295 49456 2473
rect 49562 2295 49642 2473
rect 49024 38 49642 2295
rect 50524 19771 51142 20087
rect 50524 19593 50608 19771
rect 50714 19593 50791 19771
rect 50897 19593 50974 19771
rect 51080 19593 51142 19771
rect 50524 12575 51142 19593
rect 50524 12397 50583 12575
rect 50689 12397 50766 12575
rect 50872 12397 50949 12575
rect 51055 12397 51142 12575
rect 50524 7534 51142 12397
rect 50524 7356 50585 7534
rect 50691 7356 50768 7534
rect 50874 7356 50951 7534
rect 51057 7356 51142 7534
rect 50524 354 51142 7356
rect 50524 176 50626 354
rect 50732 176 50809 354
rect 50915 176 50992 354
rect 51098 176 51142 354
rect 50524 38 51142 176
use BR128half  BR128half_0
timestamp 1654664110
transform 1 0 790 0 1 12369
box -430 -58 60604 7443
use BR128half  BR128half_1
timestamp 1654664110
transform -1 0 61001 0 1 138
box -430 -58 60604 7443
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 27641 0 1 9381
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1654402208
transform 1 0 28177 0 1 9381
box -38 -48 866 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654402208
transform 1 0 29081 0 1 9381
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654402208
transform 1 0 30997 0 1 9381
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 30740 0 1 9381
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1650294714
transform 1 0 28009 0 1 9381
box -38 -48 130 592
<< labels >>
flabel metal1 61150 13149 61394 13227 1 FreeSans 800 0 0 0 OUT
port 3 n
flabel metal1 61176 12160 61648 12221 1 FreeSans 800 0 0 0 C[112]
port 19 n
flabel metal1 61176 12018 61648 12079 1 FreeSans 800 0 0 0 C[113]
port 18 n
flabel metal1 61176 11876 61648 11937 1 FreeSans 800 0 0 0 C[114]
port 17 n
flabel metal1 61176 11734 61648 11795 1 FreeSans 800 0 0 0 C[115]
port 16 n
flabel metal1 61176 11592 61648 11653 1 FreeSans 800 0 0 0 C[116]
port 15 n
flabel metal1 61176 11450 61648 11511 1 FreeSans 800 0 0 0 C[117]
port 14 n
flabel metal1 61176 11308 61648 11369 1 FreeSans 800 0 0 0 C[118]
port 13 n
flabel metal1 61176 11166 61648 11227 1 FreeSans 800 0 0 0 C[119]
port 12 n
flabel metal1 61176 11024 61648 11085 1 FreeSans 800 0 0 0 C[120]
port 11 n
flabel metal1 61176 10882 61648 10943 1 FreeSans 800 0 0 0 C[121]
port 10 n
flabel metal1 61176 10740 61648 10801 1 FreeSans 800 0 0 0 C[122]
port 9 n
flabel metal1 61176 10598 61648 10659 1 FreeSans 800 0 0 0 C[123]
port 8 n
flabel metal1 61176 10456 61648 10517 1 FreeSans 800 0 0 0 C[124]
port 7 n
flabel metal1 61176 10314 61648 10375 1 FreeSans 800 0 0 0 C[125]
port 6 n
flabel metal1 61176 10172 61648 10233 1 FreeSans 800 0 0 0 C[126]
port 5 n
flabel metal1 61176 10030 61648 10091 1 FreeSans 800 0 0 0 C[127]
port 4 n
flabel metal1 61176 9888 61648 9949 1 FreeSans 800 0 0 0 C[63]
port 68 n
flabel metal1 61176 9746 61648 9807 1 FreeSans 800 0 0 0 C[62]
port 69 n
flabel metal1 61176 9604 61648 9665 1 FreeSans 800 0 0 0 C[61]
port 70 n
flabel metal1 61176 9462 61648 9523 1 FreeSans 800 0 0 0 C[60]
port 71 n
flabel metal1 61176 9320 61648 9381 1 FreeSans 800 0 0 0 C[59]
port 72 n
flabel metal1 61176 9178 61648 9239 1 FreeSans 800 0 0 0 C[58]
port 73 n
flabel metal1 61176 9036 61648 9097 1 FreeSans 800 0 0 0 C[57]
port 74 n
flabel metal1 61176 8894 61648 8955 1 FreeSans 800 0 0 0 C[56]
port 75 n
flabel metal1 61176 8752 61648 8813 1 FreeSans 800 0 0 0 C[55]
port 76 n
flabel metal1 61176 8610 61648 8671 1 FreeSans 800 0 0 0 C[54]
port 77 n
flabel metal1 61176 8468 61648 8529 1 FreeSans 800 0 0 0 C[53]
port 78 n
flabel metal1 61176 8326 61648 8387 1 FreeSans 800 0 0 0 C[52]
port 79 n
flabel metal1 61176 8184 61648 8245 1 FreeSans 800 0 0 0 C[51]
port 80 n
flabel metal1 61176 8042 61648 8103 1 FreeSans 800 0 0 0 C[50]
port 81 n
flabel metal1 61176 7900 61648 7961 1 FreeSans 800 0 0 0 C[49]
port 82 n
flabel metal1 61176 7758 61648 7819 1 FreeSans 800 0 0 0 C[48]
port 83 n
flabel metal3 61 9570 307 9660 1 FreeSans 400 0 0 0 RESET
port 132 n
flabel metal4 2024 38 2642 20087 1 FreeSans 1600 0 0 0 VDD
port 133 n
flabel metal4 3257 74 4041 20087 1 FreeSans 1600 0 0 0 VSS
port 134 n
flabel metal4 18524 38 19142 20087 1 FreeSans 1600 0 0 0 VDD
port 133 n
flabel metal4 20024 38 20642 20087 1 FreeSans 1600 0 0 0 VSS
port 134 n
flabel metal4 33524 38 34142 20087 1 FreeSans 1600 0 0 0 VDD
port 133 n
flabel metal4 35024 38 35642 20087 1 FreeSans 1600 0 0 0 VSS
port 134 n
flabel metal4 49024 38 49642 20087 1 FreeSans 1600 0 0 0 VDD
port 133 n
flabel metal4 50524 38 51142 20087 1 FreeSans 1600 0 0 0 VSS
port 134 n
flabel metal1 0 12163 460 12224 1 FreeSans 1200 0 0 0 C[111]
port 135 n
flabel metal1 0 12021 460 12082 1 FreeSans 1200 0 0 0 C[110]
port 136 n
flabel metal1 0 11879 460 11940 1 FreeSans 1200 0 0 0 C[109]
port 137 n
flabel metal1 0 11737 460 11798 1 FreeSans 1200 0 0 0 C[108]
port 138 n
flabel metal1 0 11595 460 11656 1 FreeSans 1200 0 0 0 C[107]
port 139 n
flabel metal1 0 11453 460 11514 1 FreeSans 1200 0 0 0 C[106]
port 140 n
flabel metal1 0 11311 460 11372 1 FreeSans 1200 0 0 0 C[105]
port 141 n
flabel metal1 0 11169 460 11230 1 FreeSans 1200 0 0 0 C[104]
port 142 n
flabel metal1 0 11027 460 11088 1 FreeSans 1200 0 0 0 C[103]
port 143 n
flabel metal1 0 10885 460 10946 1 FreeSans 1200 0 0 0 C[102]
port 144 n
flabel metal1 0 10743 460 10804 1 FreeSans 1200 0 0 0 C[101]
port 145 n
flabel metal1 0 10601 460 10662 1 FreeSans 1200 0 0 0 C[100]
port 146 n
flabel metal1 0 10459 460 10520 1 FreeSans 1200 0 0 0 C[99]
port 147 n
flabel metal1 0 10317 460 10378 1 FreeSans 1200 0 0 0 C[98]
port 148 n
flabel metal1 0 10175 460 10236 1 FreeSans 1200 0 0 0 C[97]
port 149 n
flabel metal1 0 10033 460 10094 1 FreeSans 1200 0 0 0 C[96]
port 150 n
flabel metal1 0 9891 460 9952 1 FreeSans 1200 0 0 0 C[32]
port 151 n
flabel metal1 0 9749 460 9810 1 FreeSans 1200 0 0 0 C[33]
port 152 n
flabel metal1 0 9607 460 9668 1 FreeSans 1200 0 0 0 C[34]
port 153 n
flabel metal1 0 9465 460 9526 1 FreeSans 1200 0 0 0 C[35]
port 154 n
flabel metal1 0 9323 460 9384 1 FreeSans 1200 0 0 0 C[36]
port 155 n
flabel metal1 0 9181 460 9242 1 FreeSans 1200 0 0 0 C[37]
port 156 n
flabel metal1 0 9039 460 9100 1 FreeSans 1200 0 0 0 C[38]
port 157 n
flabel metal1 0 8897 460 8958 1 FreeSans 1200 0 0 0 C[39]
port 158 n
flabel metal1 0 8755 460 8816 1 FreeSans 1200 0 0 0 C[40]
port 159 n
flabel metal1 0 8613 460 8674 1 FreeSans 1200 0 0 0 C[41]
port 160 n
flabel metal1 0 8471 460 8532 1 FreeSans 1200 0 0 0 C[42]
port 161 n
flabel metal1 0 8329 460 8390 1 FreeSans 1200 0 0 0 C[43]
port 162 n
flabel metal1 0 8187 460 8248 1 FreeSans 1200 0 0 0 C[44]
port 163 n
flabel metal1 0 8045 460 8106 1 FreeSans 1200 0 0 0 C[45]
port 164 n
flabel metal1 0 7903 460 7964 1 FreeSans 1200 0 0 0 C[46]
port 165 n
flabel metal1 0 7761 460 7822 1 FreeSans 1200 0 0 0 C[47]
port 166 n
flabel metal2 60708 19017 60752 19992 1 FreeSans 1600 0 0 0 C[0]
port 167 n
flabel metal2 58820 19017 58864 19992 1 FreeSans 1600 0 0 0 C[1]
port 168 n
flabel metal2 56932 19017 56976 19992 1 FreeSans 1600 0 0 0 C[2]
port 169 n
flabel metal2 55044 19017 55088 19992 1 FreeSans 1600 0 0 0 C[3]
port 170 n
flabel metal2 53156 19017 53200 19992 1 FreeSans 1600 0 0 0 C[4]
port 171 n
flabel metal2 51268 19017 51312 19992 1 FreeSans 1600 0 0 0 C[5]
port 172 n
flabel metal2 47492 19017 47536 19992 1 FreeSans 1600 0 0 0 C[7]
port 174 n
flabel metal2 45604 19017 45648 19992 1 FreeSans 1600 0 0 0 C[8]
port 175 n
flabel metal2 43716 19017 43760 19992 1 FreeSans 1600 0 0 0 C[9]
port 176 n
flabel metal2 41828 19017 41872 19992 1 FreeSans 1600 0 0 0 C[10]
port 177 n
flabel metal2 39940 19017 39984 19992 1 FreeSans 1600 0 0 0 C[11]
port 178 n
flabel metal2 38052 19017 38096 19992 1 FreeSans 1600 0 0 0 C[12]
port 179 n
flabel metal2 36164 19017 36208 19992 1 FreeSans 1600 0 0 0 C[13]
port 180 n
flabel metal2 34276 19017 34320 19992 1 FreeSans 1600 0 0 0 C[14]
port 181 n
flabel metal2 32388 19017 32432 19992 1 FreeSans 1600 0 0 0 C[15]
port 182 n
flabel metal2 30500 19017 30544 19992 1 FreeSans 1600 0 0 0 C[16]
port 183 n
flabel metal2 28612 19017 28656 19992 1 FreeSans 1600 0 0 0 C[17]
port 184 n
flabel metal2 26724 19017 26768 19992 1 FreeSans 1600 0 0 0 C[18]
port 185 n
flabel metal2 24836 19017 24880 19992 1 FreeSans 1600 0 0 0 C[19]
port 186 n
flabel metal2 22948 19017 22992 19992 1 FreeSans 1600 0 0 0 C[20]
port 187 n
flabel metal2 21060 19017 21104 19992 1 FreeSans 1600 0 0 0 C[21]
port 188 n
flabel metal2 19172 19017 19216 19992 1 FreeSans 1600 0 0 0 C[22]
port 189 n
flabel metal2 17284 19017 17328 19992 1 FreeSans 1600 0 0 0 C[23]
port 190 n
flabel metal2 15396 19017 15440 19992 1 FreeSans 1600 0 0 0 C[24]
port 191 n
flabel metal2 13508 19017 13552 19992 1 FreeSans 1600 0 0 0 C[25]
port 192 n
flabel metal2 11620 19017 11664 19992 1 FreeSans 1600 0 0 0 C[26]
port 193 n
flabel metal2 9732 19017 9776 19992 1 FreeSans 1600 0 0 0 C[27]
port 194 n
flabel metal2 7844 19017 7888 19992 1 FreeSans 1600 0 0 0 C[28]
port 195 n
flabel metal2 5956 19017 6000 19992 1 FreeSans 1600 0 0 0 C[29]
port 196 n
flabel metal2 4068 19017 4112 19992 1 FreeSans 1600 0 0 0 C[30]
port 197 n
flabel metal2 49380 19017 49424 20151 1 FreeSans 800 0 0 0 C[6]
port 199 n
flabel metal2 2180 19017 2224 20184 1 FreeSans 1600 0 0 0 C[31]
port 200 n
flabel metal2 2409 0 2465 930 1 FreeSans 1600 0 0 0 C[95]
port 201 n
flabel metal2 4297 0 4353 930 1 FreeSans 1600 0 0 0 C[94]
port 202 n
flabel metal2 6185 0 6241 930 1 FreeSans 1600 0 0 0 C[93]
port 203 n
flabel metal2 8073 0 8129 930 1 FreeSans 1600 0 0 0 C[92]
port 204 n
flabel metal2 9961 0 10017 930 1 FreeSans 1600 0 0 0 C[91]
port 205 n
flabel metal2 11849 0 11905 930 1 FreeSans 1600 0 0 0 C[90]
port 206 n
flabel metal2 13737 0 13793 930 1 FreeSans 1600 0 0 0 C[89]
port 207 n
flabel metal2 15625 0 15681 930 1 FreeSans 1600 0 0 0 C[88]
port 208 n
flabel metal2 17513 0 17569 930 1 FreeSans 1600 0 0 0 C[87]
port 209 n
flabel metal2 19401 0 19457 930 1 FreeSans 1600 0 0 0 C[86]
port 210 n
flabel metal2 21289 0 21345 930 1 FreeSans 1600 0 0 0 C[85]
port 211 n
flabel metal2 23177 0 23233 930 1 FreeSans 1600 0 0 0 C[84]
port 212 n
flabel metal2 25065 0 25121 930 1 FreeSans 1600 0 0 0 C[83]
port 213 n
flabel metal2 26953 0 27009 930 1 FreeSans 1600 0 0 0 C[82]
port 214 n
flabel metal2 28841 0 28897 930 1 FreeSans 1600 0 0 0 C[81]
port 215 n
flabel metal2 30729 0 30785 930 1 FreeSans 1600 0 0 0 C[80]
port 216 n
flabel metal2 32617 0 32673 930 1 FreeSans 1600 0 0 0 C[79]
port 217 n
flabel metal2 34505 0 34561 930 1 FreeSans 1600 0 0 0 C[78]
port 218 n
flabel metal2 36393 0 36449 930 1 FreeSans 1600 0 0 0 C[77]
port 219 n
flabel metal2 38281 0 38337 930 1 FreeSans 1600 0 0 0 C[76]
port 220 n
flabel metal2 40169 0 40225 930 1 FreeSans 1600 0 0 0 C[75]
port 221 n
flabel metal2 42057 0 42113 930 1 FreeSans 1600 0 0 0 C[74]
port 222 n
flabel metal2 43945 0 44001 930 1 FreeSans 1600 0 0 0 C[73]
port 223 n
flabel metal2 45833 0 45889 930 1 FreeSans 1600 0 0 0 C[72]
port 224 n
flabel metal2 47721 0 47777 930 1 FreeSans 1600 0 0 0 C[71]
port 225 n
flabel metal2 49609 0 49665 930 1 FreeSans 1600 0 0 0 C[70]
port 226 n
flabel metal2 51497 0 51553 930 1 FreeSans 1600 0 0 0 C[69]
port 227 n
flabel metal2 53385 0 53441 930 1 FreeSans 1600 0 0 0 C[68]
port 228 n
flabel metal2 55273 0 55329 930 1 FreeSans 1600 0 0 0 C[67]
port 229 n
flabel metal2 57161 0 57217 930 1 FreeSans 1600 0 0 0 C[66]
port 230 n
flabel metal2 59049 0 59105 930 1 FreeSans 1600 0 0 0 C[65]
port 231 n
flabel metal2 60937 0 60993 930 1 FreeSans 1600 0 0 0 C[64]
port 232 n
<< end >>
