magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< pwell >>
rect 76 211 90 226
<< obsli1 >>
rect 137 285 679 301
rect 137 251 139 285
rect 173 251 211 285
rect 245 251 283 285
rect 317 251 355 285
rect 389 251 427 285
rect 461 251 499 285
rect 533 251 571 285
rect 605 251 643 285
rect 677 251 679 285
rect 137 235 679 251
rect 47 173 81 189
rect 47 101 81 139
rect 47 51 81 67
rect 133 51 167 189
rect 219 173 253 189
rect 219 101 253 139
rect 219 51 253 67
rect 305 51 339 189
rect 391 173 425 189
rect 391 101 425 139
rect 391 51 425 67
rect 477 51 511 189
rect 563 173 597 189
rect 563 101 597 139
rect 563 51 597 67
rect 649 51 683 189
rect 735 173 769 189
rect 735 101 769 139
rect 735 51 769 67
<< obsli1c >>
rect 139 251 173 285
rect 211 251 245 285
rect 283 251 317 285
rect 355 251 389 285
rect 427 251 461 285
rect 499 251 533 285
rect 571 251 605 285
rect 643 251 677 285
rect 47 139 81 173
rect 47 67 81 101
rect 219 139 253 173
rect 219 67 253 101
rect 391 139 425 173
rect 391 67 425 101
rect 563 139 597 173
rect 563 67 597 101
rect 735 139 769 173
rect 735 67 769 101
<< metal1 >>
rect 127 285 689 297
rect 127 251 139 285
rect 173 251 211 285
rect 245 251 283 285
rect 317 251 355 285
rect 389 251 427 285
rect 461 251 499 285
rect 533 251 571 285
rect 605 251 643 285
rect 677 251 689 285
rect 127 239 689 251
rect 41 173 87 189
rect 41 139 47 173
rect 81 139 87 173
rect 41 101 87 139
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 213 173 259 189
rect 213 139 219 173
rect 253 139 259 173
rect 213 101 259 139
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 385 173 431 189
rect 385 139 391 173
rect 425 139 431 173
rect 385 101 431 139
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 557 173 603 189
rect 557 139 563 173
rect 597 139 603 173
rect 557 101 603 139
rect 557 67 563 101
rect 597 67 603 101
rect 557 -29 603 67
rect 729 173 775 189
rect 729 139 735 173
rect 769 139 775 173
rect 729 101 775 139
rect 729 67 735 101
rect 769 67 775 101
rect 729 -29 775 67
rect 41 -89 775 -29
<< obsm1 >>
rect 124 51 176 189
rect 296 51 348 189
rect 468 51 520 189
rect 640 51 692 189
<< obsm2 >>
rect 117 41 183 195
rect 289 41 355 195
rect 461 41 527 195
rect 633 41 699 195
<< metal3 >>
rect 117 129 699 195
rect 117 41 183 129
rect 289 41 355 129
rect 461 41 527 129
rect 633 41 699 129
<< labels >>
rlabel metal3 s 633 41 699 129 6 DRAIN
port 1 nsew
rlabel metal3 s 461 41 527 129 6 DRAIN
port 1 nsew
rlabel metal3 s 289 41 355 129 6 DRAIN
port 1 nsew
rlabel metal3 s 117 129 699 195 6 DRAIN
port 1 nsew
rlabel metal3 s 117 41 183 129 6 DRAIN
port 1 nsew
rlabel metal1 s 127 239 689 297 6 GATE
port 2 nsew
rlabel metal1 s 729 -29 775 189 6 SOURCE
port 3 nsew
rlabel metal1 s 557 -29 603 189 6 SOURCE
port 3 nsew
rlabel metal1 s 385 -29 431 189 6 SOURCE
port 3 nsew
rlabel metal1 s 213 -29 259 189 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -29 87 189 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -89 775 -29 8 SOURCE
port 3 nsew
rlabel pwell s 76 211 90 226 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 36 -89 780 301
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5942266
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5929644
<< end >>
