magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -66 377 6786 897
<< pwell >>
rect 4 43 6706 317
rect -26 -43 6746 43
<< mvnmos >>
rect 83 141 183 291
rect 239 141 339 291
rect 395 141 495 291
rect 551 141 651 291
rect 707 141 807 291
rect 863 141 963 291
rect 1019 141 1119 291
rect 1175 141 1275 291
rect 1331 141 1431 291
rect 1487 141 1587 291
rect 1691 141 1791 291
rect 1847 141 1947 291
rect 2003 141 2103 291
rect 2159 141 2259 291
rect 2315 141 2415 291
rect 2471 141 2571 291
rect 2627 141 2727 291
rect 2783 141 2883 291
rect 2939 141 3039 291
rect 3095 141 3195 291
rect 3251 141 3351 291
rect 3407 141 3507 291
rect 3563 141 3663 291
rect 3719 141 3819 291
rect 3875 141 3975 291
rect 4031 141 4131 291
rect 4187 141 4287 291
rect 4343 141 4443 291
rect 4499 141 4599 291
rect 4655 141 4755 291
rect 4811 141 4911 291
rect 4967 141 5067 291
rect 5123 141 5223 291
rect 5279 141 5379 291
rect 5435 141 5535 291
rect 5591 141 5691 291
rect 5747 141 5847 291
rect 5903 141 6003 291
rect 6059 141 6159 291
rect 6215 141 6315 291
rect 6371 141 6471 291
rect 6527 141 6627 291
<< mvpmos >>
rect 83 443 183 743
rect 239 443 339 743
rect 395 443 495 743
rect 551 443 651 743
rect 707 443 807 743
rect 863 443 963 743
rect 1019 443 1119 743
rect 1175 443 1275 743
rect 1331 443 1431 743
rect 1487 443 1587 743
rect 1691 443 1791 743
rect 1847 443 1947 743
rect 2003 443 2103 743
rect 2159 443 2259 743
rect 2315 443 2415 743
rect 2471 443 2571 743
rect 2627 443 2727 743
rect 2783 443 2883 743
rect 2939 443 3039 743
rect 3095 443 3195 743
rect 3251 443 3351 743
rect 3407 443 3507 743
rect 3563 443 3663 743
rect 3719 443 3819 743
rect 3875 443 3975 743
rect 4031 443 4131 743
rect 4187 443 4287 743
rect 4343 443 4443 743
rect 4499 443 4599 743
rect 4655 443 4755 743
rect 4811 443 4911 743
rect 4967 443 5067 743
rect 5123 443 5223 743
rect 5279 443 5379 743
rect 5435 443 5535 743
rect 5591 443 5691 743
rect 5747 443 5847 743
rect 5903 443 6003 743
rect 6059 443 6159 743
rect 6215 443 6315 743
rect 6371 443 6471 743
rect 6527 443 6627 743
<< mvndiff >>
rect 30 273 83 291
rect 30 239 38 273
rect 72 239 83 273
rect 30 205 83 239
rect 30 171 38 205
rect 72 171 83 205
rect 30 141 83 171
rect 183 269 239 291
rect 183 235 194 269
rect 228 235 239 269
rect 183 201 239 235
rect 183 167 194 201
rect 228 167 239 201
rect 183 141 239 167
rect 339 205 395 291
rect 339 171 350 205
rect 384 171 395 205
rect 339 141 395 171
rect 495 264 551 291
rect 495 230 506 264
rect 540 230 551 264
rect 495 196 551 230
rect 495 162 506 196
rect 540 162 551 196
rect 495 141 551 162
rect 651 205 707 291
rect 651 171 662 205
rect 696 171 707 205
rect 651 141 707 171
rect 807 264 863 291
rect 807 230 818 264
rect 852 230 863 264
rect 807 196 863 230
rect 807 162 818 196
rect 852 162 863 196
rect 807 141 863 162
rect 963 201 1019 291
rect 963 167 974 201
rect 1008 167 1019 201
rect 963 141 1019 167
rect 1119 264 1175 291
rect 1119 230 1130 264
rect 1164 230 1175 264
rect 1119 196 1175 230
rect 1119 162 1130 196
rect 1164 162 1175 196
rect 1119 141 1175 162
rect 1275 205 1331 291
rect 1275 171 1286 205
rect 1320 171 1331 205
rect 1275 141 1331 171
rect 1431 264 1487 291
rect 1431 230 1442 264
rect 1476 230 1487 264
rect 1431 196 1487 230
rect 1431 162 1442 196
rect 1476 162 1487 196
rect 1431 141 1487 162
rect 1587 269 1691 291
rect 1587 235 1646 269
rect 1680 235 1691 269
rect 1587 201 1691 235
rect 1587 167 1598 201
rect 1632 167 1691 201
rect 1587 141 1691 167
rect 1791 283 1847 291
rect 1791 249 1802 283
rect 1836 249 1847 283
rect 1791 208 1847 249
rect 1791 174 1802 208
rect 1836 174 1847 208
rect 1791 141 1847 174
rect 1947 269 2003 291
rect 1947 235 1958 269
rect 1992 235 2003 269
rect 1947 201 2003 235
rect 1947 167 1958 201
rect 1992 167 2003 201
rect 1947 141 2003 167
rect 2103 283 2159 291
rect 2103 249 2114 283
rect 2148 249 2159 283
rect 2103 208 2159 249
rect 2103 174 2114 208
rect 2148 174 2159 208
rect 2103 141 2159 174
rect 2259 269 2315 291
rect 2259 235 2270 269
rect 2304 235 2315 269
rect 2259 201 2315 235
rect 2259 167 2270 201
rect 2304 167 2315 201
rect 2259 141 2315 167
rect 2415 283 2471 291
rect 2415 249 2426 283
rect 2460 249 2471 283
rect 2415 208 2471 249
rect 2415 174 2426 208
rect 2460 174 2471 208
rect 2415 141 2471 174
rect 2571 269 2627 291
rect 2571 235 2582 269
rect 2616 235 2627 269
rect 2571 201 2627 235
rect 2571 167 2582 201
rect 2616 167 2627 201
rect 2571 141 2627 167
rect 2727 283 2783 291
rect 2727 249 2738 283
rect 2772 249 2783 283
rect 2727 208 2783 249
rect 2727 174 2738 208
rect 2772 174 2783 208
rect 2727 141 2783 174
rect 2883 269 2939 291
rect 2883 235 2894 269
rect 2928 235 2939 269
rect 2883 201 2939 235
rect 2883 167 2894 201
rect 2928 167 2939 201
rect 2883 141 2939 167
rect 3039 283 3095 291
rect 3039 249 3050 283
rect 3084 249 3095 283
rect 3039 208 3095 249
rect 3039 174 3050 208
rect 3084 174 3095 208
rect 3039 141 3095 174
rect 3195 269 3251 291
rect 3195 235 3206 269
rect 3240 235 3251 269
rect 3195 201 3251 235
rect 3195 167 3206 201
rect 3240 167 3251 201
rect 3195 141 3251 167
rect 3351 283 3407 291
rect 3351 249 3362 283
rect 3396 249 3407 283
rect 3351 208 3407 249
rect 3351 174 3362 208
rect 3396 174 3407 208
rect 3351 141 3407 174
rect 3507 269 3563 291
rect 3507 235 3518 269
rect 3552 235 3563 269
rect 3507 201 3563 235
rect 3507 167 3518 201
rect 3552 167 3563 201
rect 3507 141 3563 167
rect 3663 283 3719 291
rect 3663 249 3674 283
rect 3708 249 3719 283
rect 3663 208 3719 249
rect 3663 174 3674 208
rect 3708 174 3719 208
rect 3663 141 3719 174
rect 3819 269 3875 291
rect 3819 235 3830 269
rect 3864 235 3875 269
rect 3819 201 3875 235
rect 3819 167 3830 201
rect 3864 167 3875 201
rect 3819 141 3875 167
rect 3975 283 4031 291
rect 3975 249 3986 283
rect 4020 249 4031 283
rect 3975 208 4031 249
rect 3975 174 3986 208
rect 4020 174 4031 208
rect 3975 141 4031 174
rect 4131 269 4187 291
rect 4131 235 4142 269
rect 4176 235 4187 269
rect 4131 198 4187 235
rect 4131 164 4142 198
rect 4176 164 4187 198
rect 4131 141 4187 164
rect 4287 283 4343 291
rect 4287 249 4298 283
rect 4332 249 4343 283
rect 4287 208 4343 249
rect 4287 174 4298 208
rect 4332 174 4343 208
rect 4287 141 4343 174
rect 4443 269 4499 291
rect 4443 235 4454 269
rect 4488 235 4499 269
rect 4443 201 4499 235
rect 4443 167 4454 201
rect 4488 167 4499 201
rect 4443 141 4499 167
rect 4599 283 4655 291
rect 4599 249 4610 283
rect 4644 249 4655 283
rect 4599 208 4655 249
rect 4599 174 4610 208
rect 4644 174 4655 208
rect 4599 141 4655 174
rect 4755 269 4811 291
rect 4755 235 4766 269
rect 4800 235 4811 269
rect 4755 201 4811 235
rect 4755 167 4766 201
rect 4800 167 4811 201
rect 4755 141 4811 167
rect 4911 283 4967 291
rect 4911 249 4922 283
rect 4956 249 4967 283
rect 4911 208 4967 249
rect 4911 174 4922 208
rect 4956 174 4967 208
rect 4911 141 4967 174
rect 5067 269 5123 291
rect 5067 235 5078 269
rect 5112 235 5123 269
rect 5067 201 5123 235
rect 5067 167 5078 201
rect 5112 167 5123 201
rect 5067 141 5123 167
rect 5223 283 5279 291
rect 5223 249 5234 283
rect 5268 249 5279 283
rect 5223 208 5279 249
rect 5223 174 5234 208
rect 5268 174 5279 208
rect 5223 141 5279 174
rect 5379 269 5435 291
rect 5379 235 5390 269
rect 5424 235 5435 269
rect 5379 201 5435 235
rect 5379 167 5390 201
rect 5424 167 5435 201
rect 5379 141 5435 167
rect 5535 283 5591 291
rect 5535 249 5546 283
rect 5580 249 5591 283
rect 5535 208 5591 249
rect 5535 174 5546 208
rect 5580 174 5591 208
rect 5535 141 5591 174
rect 5691 269 5747 291
rect 5691 235 5702 269
rect 5736 235 5747 269
rect 5691 201 5747 235
rect 5691 167 5702 201
rect 5736 167 5747 201
rect 5691 141 5747 167
rect 5847 283 5903 291
rect 5847 249 5858 283
rect 5892 249 5903 283
rect 5847 208 5903 249
rect 5847 174 5858 208
rect 5892 174 5903 208
rect 5847 141 5903 174
rect 6003 269 6059 291
rect 6003 235 6014 269
rect 6048 235 6059 269
rect 6003 201 6059 235
rect 6003 167 6014 201
rect 6048 167 6059 201
rect 6003 141 6059 167
rect 6159 283 6215 291
rect 6159 249 6170 283
rect 6204 249 6215 283
rect 6159 208 6215 249
rect 6159 174 6170 208
rect 6204 174 6215 208
rect 6159 141 6215 174
rect 6315 269 6371 291
rect 6315 235 6326 269
rect 6360 235 6371 269
rect 6315 201 6371 235
rect 6315 167 6326 201
rect 6360 167 6371 201
rect 6315 141 6371 167
rect 6471 283 6527 291
rect 6471 249 6482 283
rect 6516 249 6527 283
rect 6471 208 6527 249
rect 6471 174 6482 208
rect 6516 174 6527 208
rect 6471 141 6527 174
rect 6627 279 6680 291
rect 6627 245 6638 279
rect 6672 245 6680 279
rect 6627 208 6680 245
rect 6627 174 6638 208
rect 6672 174 6680 208
rect 6627 141 6680 174
<< mvpdiff >>
rect 30 731 83 743
rect 30 697 38 731
rect 72 697 83 731
rect 30 642 83 697
rect 30 608 38 642
rect 72 608 83 642
rect 30 562 83 608
rect 30 528 38 562
rect 72 528 83 562
rect 30 489 83 528
rect 30 455 38 489
rect 72 455 83 489
rect 30 443 83 455
rect 183 735 239 743
rect 183 701 194 735
rect 228 701 239 735
rect 183 642 239 701
rect 183 608 194 642
rect 228 608 239 642
rect 183 558 239 608
rect 183 524 194 558
rect 228 524 239 558
rect 183 485 239 524
rect 183 451 194 485
rect 228 451 239 485
rect 183 443 239 451
rect 339 731 395 743
rect 339 697 350 731
rect 384 697 395 731
rect 339 663 395 697
rect 339 629 350 663
rect 384 629 395 663
rect 339 595 395 629
rect 339 561 350 595
rect 384 561 395 595
rect 339 527 395 561
rect 339 493 350 527
rect 384 493 395 527
rect 339 443 395 493
rect 495 735 551 743
rect 495 701 506 735
rect 540 701 551 735
rect 495 642 551 701
rect 495 608 506 642
rect 540 608 551 642
rect 495 558 551 608
rect 495 524 506 558
rect 540 524 551 558
rect 495 485 551 524
rect 495 451 506 485
rect 540 451 551 485
rect 495 443 551 451
rect 651 731 707 743
rect 651 697 662 731
rect 696 697 707 731
rect 651 663 707 697
rect 651 629 662 663
rect 696 629 707 663
rect 651 595 707 629
rect 651 561 662 595
rect 696 561 707 595
rect 651 527 707 561
rect 651 493 662 527
rect 696 493 707 527
rect 651 443 707 493
rect 807 735 863 743
rect 807 701 818 735
rect 852 701 863 735
rect 807 642 863 701
rect 807 608 818 642
rect 852 608 863 642
rect 807 558 863 608
rect 807 524 818 558
rect 852 524 863 558
rect 807 485 863 524
rect 807 451 818 485
rect 852 451 863 485
rect 807 443 863 451
rect 963 731 1019 743
rect 963 697 974 731
rect 1008 697 1019 731
rect 963 663 1019 697
rect 963 629 974 663
rect 1008 629 1019 663
rect 963 595 1019 629
rect 963 561 974 595
rect 1008 561 1019 595
rect 963 527 1019 561
rect 963 493 974 527
rect 1008 493 1019 527
rect 963 443 1019 493
rect 1119 735 1175 743
rect 1119 701 1130 735
rect 1164 701 1175 735
rect 1119 642 1175 701
rect 1119 608 1130 642
rect 1164 608 1175 642
rect 1119 558 1175 608
rect 1119 524 1130 558
rect 1164 524 1175 558
rect 1119 485 1175 524
rect 1119 451 1130 485
rect 1164 451 1175 485
rect 1119 443 1175 451
rect 1275 731 1331 743
rect 1275 697 1286 731
rect 1320 697 1331 731
rect 1275 663 1331 697
rect 1275 629 1286 663
rect 1320 629 1331 663
rect 1275 595 1331 629
rect 1275 561 1286 595
rect 1320 561 1331 595
rect 1275 527 1331 561
rect 1275 493 1286 527
rect 1320 493 1331 527
rect 1275 443 1331 493
rect 1431 735 1487 743
rect 1431 701 1442 735
rect 1476 701 1487 735
rect 1431 642 1487 701
rect 1431 608 1442 642
rect 1476 608 1487 642
rect 1431 558 1487 608
rect 1431 524 1442 558
rect 1476 524 1487 558
rect 1431 485 1487 524
rect 1431 451 1442 485
rect 1476 451 1487 485
rect 1431 443 1487 451
rect 1587 731 1691 743
rect 1587 697 1598 731
rect 1632 697 1691 731
rect 1587 663 1691 697
rect 1587 629 1646 663
rect 1680 629 1691 663
rect 1587 553 1691 629
rect 1587 519 1598 553
rect 1632 519 1691 553
rect 1587 485 1691 519
rect 1587 451 1646 485
rect 1680 451 1691 485
rect 1587 443 1691 451
rect 1791 735 1847 743
rect 1791 701 1802 735
rect 1836 701 1847 735
rect 1791 656 1847 701
rect 1791 622 1802 656
rect 1836 622 1847 656
rect 1791 576 1847 622
rect 1791 542 1802 576
rect 1836 542 1847 576
rect 1791 485 1847 542
rect 1791 451 1802 485
rect 1836 451 1847 485
rect 1791 443 1847 451
rect 1947 735 2003 743
rect 1947 701 1958 735
rect 1992 701 2003 735
rect 1947 656 2003 701
rect 1947 622 1958 656
rect 1992 622 2003 656
rect 1947 576 2003 622
rect 1947 542 1958 576
rect 1992 542 2003 576
rect 1947 485 2003 542
rect 1947 451 1958 485
rect 1992 451 2003 485
rect 1947 443 2003 451
rect 2103 735 2159 743
rect 2103 701 2114 735
rect 2148 701 2159 735
rect 2103 656 2159 701
rect 2103 622 2114 656
rect 2148 622 2159 656
rect 2103 576 2159 622
rect 2103 542 2114 576
rect 2148 542 2159 576
rect 2103 485 2159 542
rect 2103 451 2114 485
rect 2148 451 2159 485
rect 2103 443 2159 451
rect 2259 735 2315 743
rect 2259 701 2270 735
rect 2304 701 2315 735
rect 2259 656 2315 701
rect 2259 622 2270 656
rect 2304 622 2315 656
rect 2259 576 2315 622
rect 2259 542 2270 576
rect 2304 542 2315 576
rect 2259 485 2315 542
rect 2259 451 2270 485
rect 2304 451 2315 485
rect 2259 443 2315 451
rect 2415 735 2471 743
rect 2415 701 2426 735
rect 2460 701 2471 735
rect 2415 656 2471 701
rect 2415 622 2426 656
rect 2460 622 2471 656
rect 2415 576 2471 622
rect 2415 542 2426 576
rect 2460 542 2471 576
rect 2415 485 2471 542
rect 2415 451 2426 485
rect 2460 451 2471 485
rect 2415 443 2471 451
rect 2571 735 2627 743
rect 2571 701 2582 735
rect 2616 701 2627 735
rect 2571 656 2627 701
rect 2571 622 2582 656
rect 2616 622 2627 656
rect 2571 576 2627 622
rect 2571 542 2582 576
rect 2616 542 2627 576
rect 2571 485 2627 542
rect 2571 451 2582 485
rect 2616 451 2627 485
rect 2571 443 2627 451
rect 2727 735 2783 743
rect 2727 701 2738 735
rect 2772 701 2783 735
rect 2727 656 2783 701
rect 2727 622 2738 656
rect 2772 622 2783 656
rect 2727 576 2783 622
rect 2727 542 2738 576
rect 2772 542 2783 576
rect 2727 485 2783 542
rect 2727 451 2738 485
rect 2772 451 2783 485
rect 2727 443 2783 451
rect 2883 735 2939 743
rect 2883 701 2894 735
rect 2928 701 2939 735
rect 2883 656 2939 701
rect 2883 622 2894 656
rect 2928 622 2939 656
rect 2883 576 2939 622
rect 2883 542 2894 576
rect 2928 542 2939 576
rect 2883 485 2939 542
rect 2883 451 2894 485
rect 2928 451 2939 485
rect 2883 443 2939 451
rect 3039 735 3095 743
rect 3039 701 3050 735
rect 3084 701 3095 735
rect 3039 656 3095 701
rect 3039 622 3050 656
rect 3084 622 3095 656
rect 3039 576 3095 622
rect 3039 542 3050 576
rect 3084 542 3095 576
rect 3039 485 3095 542
rect 3039 451 3050 485
rect 3084 451 3095 485
rect 3039 443 3095 451
rect 3195 735 3251 743
rect 3195 701 3206 735
rect 3240 701 3251 735
rect 3195 656 3251 701
rect 3195 622 3206 656
rect 3240 622 3251 656
rect 3195 576 3251 622
rect 3195 542 3206 576
rect 3240 542 3251 576
rect 3195 485 3251 542
rect 3195 451 3206 485
rect 3240 451 3251 485
rect 3195 443 3251 451
rect 3351 735 3407 743
rect 3351 701 3362 735
rect 3396 701 3407 735
rect 3351 656 3407 701
rect 3351 622 3362 656
rect 3396 622 3407 656
rect 3351 576 3407 622
rect 3351 542 3362 576
rect 3396 542 3407 576
rect 3351 485 3407 542
rect 3351 451 3362 485
rect 3396 451 3407 485
rect 3351 443 3407 451
rect 3507 735 3563 743
rect 3507 701 3518 735
rect 3552 701 3563 735
rect 3507 656 3563 701
rect 3507 622 3518 656
rect 3552 622 3563 656
rect 3507 576 3563 622
rect 3507 542 3518 576
rect 3552 542 3563 576
rect 3507 485 3563 542
rect 3507 451 3518 485
rect 3552 451 3563 485
rect 3507 443 3563 451
rect 3663 735 3719 743
rect 3663 701 3674 735
rect 3708 701 3719 735
rect 3663 656 3719 701
rect 3663 622 3674 656
rect 3708 622 3719 656
rect 3663 576 3719 622
rect 3663 542 3674 576
rect 3708 542 3719 576
rect 3663 485 3719 542
rect 3663 451 3674 485
rect 3708 451 3719 485
rect 3663 443 3719 451
rect 3819 735 3875 743
rect 3819 701 3830 735
rect 3864 701 3875 735
rect 3819 656 3875 701
rect 3819 622 3830 656
rect 3864 622 3875 656
rect 3819 576 3875 622
rect 3819 542 3830 576
rect 3864 542 3875 576
rect 3819 485 3875 542
rect 3819 451 3830 485
rect 3864 451 3875 485
rect 3819 443 3875 451
rect 3975 735 4031 743
rect 3975 701 3986 735
rect 4020 701 4031 735
rect 3975 656 4031 701
rect 3975 622 3986 656
rect 4020 622 4031 656
rect 3975 576 4031 622
rect 3975 542 3986 576
rect 4020 542 4031 576
rect 3975 485 4031 542
rect 3975 451 3986 485
rect 4020 451 4031 485
rect 3975 443 4031 451
rect 4131 731 4187 743
rect 4131 697 4142 731
rect 4176 697 4187 731
rect 4131 656 4187 697
rect 4131 622 4142 656
rect 4176 622 4187 656
rect 4131 576 4187 622
rect 4131 542 4142 576
rect 4176 542 4187 576
rect 4131 489 4187 542
rect 4131 455 4142 489
rect 4176 455 4187 489
rect 4131 443 4187 455
rect 4287 735 4343 743
rect 4287 701 4298 735
rect 4332 701 4343 735
rect 4287 656 4343 701
rect 4287 622 4298 656
rect 4332 622 4343 656
rect 4287 576 4343 622
rect 4287 542 4298 576
rect 4332 542 4343 576
rect 4287 485 4343 542
rect 4287 451 4298 485
rect 4332 451 4343 485
rect 4287 443 4343 451
rect 4443 735 4499 743
rect 4443 701 4454 735
rect 4488 701 4499 735
rect 4443 656 4499 701
rect 4443 622 4454 656
rect 4488 622 4499 656
rect 4443 576 4499 622
rect 4443 542 4454 576
rect 4488 542 4499 576
rect 4443 485 4499 542
rect 4443 451 4454 485
rect 4488 451 4499 485
rect 4443 443 4499 451
rect 4599 735 4655 743
rect 4599 701 4610 735
rect 4644 701 4655 735
rect 4599 656 4655 701
rect 4599 622 4610 656
rect 4644 622 4655 656
rect 4599 576 4655 622
rect 4599 542 4610 576
rect 4644 542 4655 576
rect 4599 485 4655 542
rect 4599 451 4610 485
rect 4644 451 4655 485
rect 4599 443 4655 451
rect 4755 735 4811 743
rect 4755 701 4766 735
rect 4800 701 4811 735
rect 4755 656 4811 701
rect 4755 622 4766 656
rect 4800 622 4811 656
rect 4755 576 4811 622
rect 4755 542 4766 576
rect 4800 542 4811 576
rect 4755 485 4811 542
rect 4755 451 4766 485
rect 4800 451 4811 485
rect 4755 443 4811 451
rect 4911 735 4967 743
rect 4911 701 4922 735
rect 4956 701 4967 735
rect 4911 656 4967 701
rect 4911 622 4922 656
rect 4956 622 4967 656
rect 4911 576 4967 622
rect 4911 542 4922 576
rect 4956 542 4967 576
rect 4911 485 4967 542
rect 4911 451 4922 485
rect 4956 451 4967 485
rect 4911 443 4967 451
rect 5067 735 5123 743
rect 5067 701 5078 735
rect 5112 701 5123 735
rect 5067 656 5123 701
rect 5067 622 5078 656
rect 5112 622 5123 656
rect 5067 576 5123 622
rect 5067 542 5078 576
rect 5112 542 5123 576
rect 5067 485 5123 542
rect 5067 451 5078 485
rect 5112 451 5123 485
rect 5067 443 5123 451
rect 5223 735 5279 743
rect 5223 701 5234 735
rect 5268 701 5279 735
rect 5223 656 5279 701
rect 5223 622 5234 656
rect 5268 622 5279 656
rect 5223 576 5279 622
rect 5223 542 5234 576
rect 5268 542 5279 576
rect 5223 485 5279 542
rect 5223 451 5234 485
rect 5268 451 5279 485
rect 5223 443 5279 451
rect 5379 735 5435 743
rect 5379 701 5390 735
rect 5424 701 5435 735
rect 5379 656 5435 701
rect 5379 622 5390 656
rect 5424 622 5435 656
rect 5379 576 5435 622
rect 5379 542 5390 576
rect 5424 542 5435 576
rect 5379 485 5435 542
rect 5379 451 5390 485
rect 5424 451 5435 485
rect 5379 443 5435 451
rect 5535 735 5591 743
rect 5535 701 5546 735
rect 5580 701 5591 735
rect 5535 656 5591 701
rect 5535 622 5546 656
rect 5580 622 5591 656
rect 5535 576 5591 622
rect 5535 542 5546 576
rect 5580 542 5591 576
rect 5535 485 5591 542
rect 5535 451 5546 485
rect 5580 451 5591 485
rect 5535 443 5591 451
rect 5691 735 5747 743
rect 5691 701 5702 735
rect 5736 701 5747 735
rect 5691 656 5747 701
rect 5691 622 5702 656
rect 5736 622 5747 656
rect 5691 576 5747 622
rect 5691 542 5702 576
rect 5736 542 5747 576
rect 5691 485 5747 542
rect 5691 451 5702 485
rect 5736 451 5747 485
rect 5691 443 5747 451
rect 5847 735 5903 743
rect 5847 701 5858 735
rect 5892 701 5903 735
rect 5847 656 5903 701
rect 5847 622 5858 656
rect 5892 622 5903 656
rect 5847 576 5903 622
rect 5847 542 5858 576
rect 5892 542 5903 576
rect 5847 485 5903 542
rect 5847 451 5858 485
rect 5892 451 5903 485
rect 5847 443 5903 451
rect 6003 735 6059 743
rect 6003 701 6014 735
rect 6048 701 6059 735
rect 6003 656 6059 701
rect 6003 622 6014 656
rect 6048 622 6059 656
rect 6003 576 6059 622
rect 6003 542 6014 576
rect 6048 542 6059 576
rect 6003 485 6059 542
rect 6003 451 6014 485
rect 6048 451 6059 485
rect 6003 443 6059 451
rect 6159 735 6215 743
rect 6159 701 6170 735
rect 6204 701 6215 735
rect 6159 656 6215 701
rect 6159 622 6170 656
rect 6204 622 6215 656
rect 6159 576 6215 622
rect 6159 542 6170 576
rect 6204 542 6215 576
rect 6159 485 6215 542
rect 6159 451 6170 485
rect 6204 451 6215 485
rect 6159 443 6215 451
rect 6315 735 6371 743
rect 6315 701 6326 735
rect 6360 701 6371 735
rect 6315 656 6371 701
rect 6315 622 6326 656
rect 6360 622 6371 656
rect 6315 576 6371 622
rect 6315 542 6326 576
rect 6360 542 6371 576
rect 6315 485 6371 542
rect 6315 451 6326 485
rect 6360 451 6371 485
rect 6315 443 6371 451
rect 6471 735 6527 743
rect 6471 701 6482 735
rect 6516 701 6527 735
rect 6471 656 6527 701
rect 6471 622 6482 656
rect 6516 622 6527 656
rect 6471 576 6527 622
rect 6471 542 6482 576
rect 6516 542 6527 576
rect 6471 485 6527 542
rect 6471 451 6482 485
rect 6516 451 6527 485
rect 6471 443 6527 451
rect 6627 731 6680 743
rect 6627 697 6638 731
rect 6672 697 6680 731
rect 6627 656 6680 697
rect 6627 622 6638 656
rect 6672 622 6680 656
rect 6627 576 6680 622
rect 6627 542 6638 576
rect 6672 542 6680 576
rect 6627 489 6680 542
rect 6627 455 6638 489
rect 6672 455 6680 489
rect 6627 443 6680 455
<< mvndiffc >>
rect 38 239 72 273
rect 38 171 72 205
rect 194 235 228 269
rect 194 167 228 201
rect 350 171 384 205
rect 506 230 540 264
rect 506 162 540 196
rect 662 171 696 205
rect 818 230 852 264
rect 818 162 852 196
rect 974 167 1008 201
rect 1130 230 1164 264
rect 1130 162 1164 196
rect 1286 171 1320 205
rect 1442 230 1476 264
rect 1442 162 1476 196
rect 1646 235 1680 269
rect 1598 167 1632 201
rect 1802 249 1836 283
rect 1802 174 1836 208
rect 1958 235 1992 269
rect 1958 167 1992 201
rect 2114 249 2148 283
rect 2114 174 2148 208
rect 2270 235 2304 269
rect 2270 167 2304 201
rect 2426 249 2460 283
rect 2426 174 2460 208
rect 2582 235 2616 269
rect 2582 167 2616 201
rect 2738 249 2772 283
rect 2738 174 2772 208
rect 2894 235 2928 269
rect 2894 167 2928 201
rect 3050 249 3084 283
rect 3050 174 3084 208
rect 3206 235 3240 269
rect 3206 167 3240 201
rect 3362 249 3396 283
rect 3362 174 3396 208
rect 3518 235 3552 269
rect 3518 167 3552 201
rect 3674 249 3708 283
rect 3674 174 3708 208
rect 3830 235 3864 269
rect 3830 167 3864 201
rect 3986 249 4020 283
rect 3986 174 4020 208
rect 4142 235 4176 269
rect 4142 164 4176 198
rect 4298 249 4332 283
rect 4298 174 4332 208
rect 4454 235 4488 269
rect 4454 167 4488 201
rect 4610 249 4644 283
rect 4610 174 4644 208
rect 4766 235 4800 269
rect 4766 167 4800 201
rect 4922 249 4956 283
rect 4922 174 4956 208
rect 5078 235 5112 269
rect 5078 167 5112 201
rect 5234 249 5268 283
rect 5234 174 5268 208
rect 5390 235 5424 269
rect 5390 167 5424 201
rect 5546 249 5580 283
rect 5546 174 5580 208
rect 5702 235 5736 269
rect 5702 167 5736 201
rect 5858 249 5892 283
rect 5858 174 5892 208
rect 6014 235 6048 269
rect 6014 167 6048 201
rect 6170 249 6204 283
rect 6170 174 6204 208
rect 6326 235 6360 269
rect 6326 167 6360 201
rect 6482 249 6516 283
rect 6482 174 6516 208
rect 6638 245 6672 279
rect 6638 174 6672 208
<< mvpdiffc >>
rect 38 697 72 731
rect 38 608 72 642
rect 38 528 72 562
rect 38 455 72 489
rect 194 701 228 735
rect 194 608 228 642
rect 194 524 228 558
rect 194 451 228 485
rect 350 697 384 731
rect 350 629 384 663
rect 350 561 384 595
rect 350 493 384 527
rect 506 701 540 735
rect 506 608 540 642
rect 506 524 540 558
rect 506 451 540 485
rect 662 697 696 731
rect 662 629 696 663
rect 662 561 696 595
rect 662 493 696 527
rect 818 701 852 735
rect 818 608 852 642
rect 818 524 852 558
rect 818 451 852 485
rect 974 697 1008 731
rect 974 629 1008 663
rect 974 561 1008 595
rect 974 493 1008 527
rect 1130 701 1164 735
rect 1130 608 1164 642
rect 1130 524 1164 558
rect 1130 451 1164 485
rect 1286 697 1320 731
rect 1286 629 1320 663
rect 1286 561 1320 595
rect 1286 493 1320 527
rect 1442 701 1476 735
rect 1442 608 1476 642
rect 1442 524 1476 558
rect 1442 451 1476 485
rect 1598 697 1632 731
rect 1646 629 1680 663
rect 1598 519 1632 553
rect 1646 451 1680 485
rect 1802 701 1836 735
rect 1802 622 1836 656
rect 1802 542 1836 576
rect 1802 451 1836 485
rect 1958 701 1992 735
rect 1958 622 1992 656
rect 1958 542 1992 576
rect 1958 451 1992 485
rect 2114 701 2148 735
rect 2114 622 2148 656
rect 2114 542 2148 576
rect 2114 451 2148 485
rect 2270 701 2304 735
rect 2270 622 2304 656
rect 2270 542 2304 576
rect 2270 451 2304 485
rect 2426 701 2460 735
rect 2426 622 2460 656
rect 2426 542 2460 576
rect 2426 451 2460 485
rect 2582 701 2616 735
rect 2582 622 2616 656
rect 2582 542 2616 576
rect 2582 451 2616 485
rect 2738 701 2772 735
rect 2738 622 2772 656
rect 2738 542 2772 576
rect 2738 451 2772 485
rect 2894 701 2928 735
rect 2894 622 2928 656
rect 2894 542 2928 576
rect 2894 451 2928 485
rect 3050 701 3084 735
rect 3050 622 3084 656
rect 3050 542 3084 576
rect 3050 451 3084 485
rect 3206 701 3240 735
rect 3206 622 3240 656
rect 3206 542 3240 576
rect 3206 451 3240 485
rect 3362 701 3396 735
rect 3362 622 3396 656
rect 3362 542 3396 576
rect 3362 451 3396 485
rect 3518 701 3552 735
rect 3518 622 3552 656
rect 3518 542 3552 576
rect 3518 451 3552 485
rect 3674 701 3708 735
rect 3674 622 3708 656
rect 3674 542 3708 576
rect 3674 451 3708 485
rect 3830 701 3864 735
rect 3830 622 3864 656
rect 3830 542 3864 576
rect 3830 451 3864 485
rect 3986 701 4020 735
rect 3986 622 4020 656
rect 3986 542 4020 576
rect 3986 451 4020 485
rect 4142 697 4176 731
rect 4142 622 4176 656
rect 4142 542 4176 576
rect 4142 455 4176 489
rect 4298 701 4332 735
rect 4298 622 4332 656
rect 4298 542 4332 576
rect 4298 451 4332 485
rect 4454 701 4488 735
rect 4454 622 4488 656
rect 4454 542 4488 576
rect 4454 451 4488 485
rect 4610 701 4644 735
rect 4610 622 4644 656
rect 4610 542 4644 576
rect 4610 451 4644 485
rect 4766 701 4800 735
rect 4766 622 4800 656
rect 4766 542 4800 576
rect 4766 451 4800 485
rect 4922 701 4956 735
rect 4922 622 4956 656
rect 4922 542 4956 576
rect 4922 451 4956 485
rect 5078 701 5112 735
rect 5078 622 5112 656
rect 5078 542 5112 576
rect 5078 451 5112 485
rect 5234 701 5268 735
rect 5234 622 5268 656
rect 5234 542 5268 576
rect 5234 451 5268 485
rect 5390 701 5424 735
rect 5390 622 5424 656
rect 5390 542 5424 576
rect 5390 451 5424 485
rect 5546 701 5580 735
rect 5546 622 5580 656
rect 5546 542 5580 576
rect 5546 451 5580 485
rect 5702 701 5736 735
rect 5702 622 5736 656
rect 5702 542 5736 576
rect 5702 451 5736 485
rect 5858 701 5892 735
rect 5858 622 5892 656
rect 5858 542 5892 576
rect 5858 451 5892 485
rect 6014 701 6048 735
rect 6014 622 6048 656
rect 6014 542 6048 576
rect 6014 451 6048 485
rect 6170 701 6204 735
rect 6170 622 6204 656
rect 6170 542 6204 576
rect 6170 451 6204 485
rect 6326 701 6360 735
rect 6326 622 6360 656
rect 6326 542 6360 576
rect 6326 451 6360 485
rect 6482 701 6516 735
rect 6482 622 6516 656
rect 6482 542 6516 576
rect 6482 451 6516 485
rect 6638 697 6672 731
rect 6638 622 6672 656
rect 6638 542 6672 576
rect 6638 455 6672 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 5023 17
rect 5057 -17 5119 17
rect 5153 -17 5215 17
rect 5249 -17 5311 17
rect 5345 -17 5407 17
rect 5441 -17 5503 17
rect 5537 -17 5599 17
rect 5633 -17 5695 17
rect 5729 -17 5791 17
rect 5825 -17 5887 17
rect 5921 -17 5983 17
rect 6017 -17 6079 17
rect 6113 -17 6175 17
rect 6209 -17 6271 17
rect 6305 -17 6367 17
rect 6401 -17 6463 17
rect 6497 -17 6559 17
rect 6593 -17 6655 17
rect 6689 -17 6720 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4063 831
rect 4097 797 4159 831
rect 4193 797 4255 831
rect 4289 797 4351 831
rect 4385 797 4447 831
rect 4481 797 4543 831
rect 4577 797 4639 831
rect 4673 797 4735 831
rect 4769 797 4831 831
rect 4865 797 4927 831
rect 4961 797 5023 831
rect 5057 797 5119 831
rect 5153 797 5215 831
rect 5249 797 5311 831
rect 5345 797 5407 831
rect 5441 797 5503 831
rect 5537 797 5599 831
rect 5633 797 5695 831
rect 5729 797 5791 831
rect 5825 797 5887 831
rect 5921 797 5983 831
rect 6017 797 6079 831
rect 6113 797 6175 831
rect 6209 797 6271 831
rect 6305 797 6367 831
rect 6401 797 6463 831
rect 6497 797 6559 831
rect 6593 797 6655 831
rect 6689 797 6720 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect 4927 -17 4961 17
rect 5023 -17 5057 17
rect 5119 -17 5153 17
rect 5215 -17 5249 17
rect 5311 -17 5345 17
rect 5407 -17 5441 17
rect 5503 -17 5537 17
rect 5599 -17 5633 17
rect 5695 -17 5729 17
rect 5791 -17 5825 17
rect 5887 -17 5921 17
rect 5983 -17 6017 17
rect 6079 -17 6113 17
rect 6175 -17 6209 17
rect 6271 -17 6305 17
rect 6367 -17 6401 17
rect 6463 -17 6497 17
rect 6559 -17 6593 17
rect 6655 -17 6689 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
rect 4063 797 4097 831
rect 4159 797 4193 831
rect 4255 797 4289 831
rect 4351 797 4385 831
rect 4447 797 4481 831
rect 4543 797 4577 831
rect 4639 797 4673 831
rect 4735 797 4769 831
rect 4831 797 4865 831
rect 4927 797 4961 831
rect 5023 797 5057 831
rect 5119 797 5153 831
rect 5215 797 5249 831
rect 5311 797 5345 831
rect 5407 797 5441 831
rect 5503 797 5537 831
rect 5599 797 5633 831
rect 5695 797 5729 831
rect 5791 797 5825 831
rect 5887 797 5921 831
rect 5983 797 6017 831
rect 6079 797 6113 831
rect 6175 797 6209 831
rect 6271 797 6305 831
rect 6367 797 6401 831
rect 6463 797 6497 831
rect 6559 797 6593 831
rect 6655 797 6689 831
<< poly >>
rect 83 743 183 769
rect 239 743 339 769
rect 395 743 495 769
rect 551 743 651 769
rect 707 743 807 769
rect 863 743 963 769
rect 1019 743 1119 769
rect 1175 743 1275 769
rect 1331 743 1431 769
rect 1487 743 1587 769
rect 1691 743 1791 769
rect 1847 743 1947 769
rect 2003 743 2103 769
rect 2159 743 2259 769
rect 2315 743 2415 769
rect 2471 743 2571 769
rect 2627 743 2727 769
rect 2783 743 2883 769
rect 2939 743 3039 769
rect 3095 743 3195 769
rect 3251 743 3351 769
rect 3407 743 3507 769
rect 3563 743 3663 769
rect 3719 743 3819 769
rect 3875 743 3975 769
rect 4031 743 4131 769
rect 4187 743 4287 769
rect 4343 743 4443 769
rect 4499 743 4599 769
rect 4655 743 4755 769
rect 4811 743 4911 769
rect 4967 743 5067 769
rect 5123 743 5223 769
rect 5279 743 5379 769
rect 5435 743 5535 769
rect 5591 743 5691 769
rect 5747 743 5847 769
rect 5903 743 6003 769
rect 6059 743 6159 769
rect 6215 743 6315 769
rect 6371 743 6471 769
rect 6527 743 6627 769
rect 83 413 183 443
rect 239 413 339 443
rect 395 413 495 443
rect 551 413 651 443
rect 707 413 807 443
rect 863 413 963 443
rect 1019 413 1119 443
rect 1175 413 1275 443
rect 1331 413 1431 443
rect 1487 413 1587 443
rect 44 363 1587 413
rect 44 329 60 363
rect 94 329 128 363
rect 162 329 196 363
rect 230 329 264 363
rect 298 329 332 363
rect 366 329 400 363
rect 434 329 468 363
rect 502 329 536 363
rect 570 329 604 363
rect 638 329 672 363
rect 706 329 740 363
rect 774 329 808 363
rect 842 329 876 363
rect 910 329 1587 363
rect 44 313 1587 329
rect 83 291 183 313
rect 239 291 339 313
rect 395 291 495 313
rect 551 291 651 313
rect 707 291 807 313
rect 863 291 963 313
rect 1019 291 1119 313
rect 1175 291 1275 313
rect 1331 291 1431 313
rect 1487 291 1587 313
rect 1691 401 1791 443
rect 1847 401 1947 443
rect 2003 401 2103 443
rect 2159 401 2259 443
rect 2315 401 2415 443
rect 2471 401 2571 443
rect 2627 401 2727 443
rect 2783 401 2883 443
rect 2939 401 3039 443
rect 3095 401 3195 443
rect 3251 401 3351 443
rect 3407 401 3507 443
rect 3563 401 3663 443
rect 3719 401 3819 443
rect 3875 401 3975 443
rect 4031 401 4131 443
rect 4187 401 4287 443
rect 4343 401 4443 443
rect 4499 401 4599 443
rect 4655 401 4755 443
rect 4811 401 4911 443
rect 4967 401 5067 443
rect 5123 401 5223 443
rect 5279 401 5379 443
rect 5435 401 5535 443
rect 5591 401 5691 443
rect 5747 401 5847 443
rect 5903 401 6003 443
rect 6059 401 6159 443
rect 6215 401 6315 443
rect 6371 401 6471 443
rect 6527 401 6627 443
rect 1691 363 6627 401
rect 1691 329 1920 363
rect 1954 329 1988 363
rect 2022 329 2232 363
rect 2266 329 2300 363
rect 2334 329 2544 363
rect 2578 329 2612 363
rect 2646 329 2856 363
rect 2890 329 2924 363
rect 2958 329 3168 363
rect 3202 329 3236 363
rect 3270 329 3480 363
rect 3514 329 3548 363
rect 3582 329 3792 363
rect 3826 329 3860 363
rect 3894 329 4102 363
rect 4136 329 4170 363
rect 4204 329 4416 363
rect 4450 329 4484 363
rect 4518 329 4728 363
rect 4762 329 4796 363
rect 4830 329 5040 363
rect 5074 329 5108 363
rect 5142 329 5352 363
rect 5386 329 5420 363
rect 5454 329 5664 363
rect 5698 329 5732 363
rect 5766 329 5976 363
rect 6010 329 6044 363
rect 6078 329 6288 363
rect 6322 329 6356 363
rect 6390 329 6627 363
rect 1691 313 6627 329
rect 1691 291 1791 313
rect 1847 291 1947 313
rect 2003 291 2103 313
rect 2159 291 2259 313
rect 2315 291 2415 313
rect 2471 291 2571 313
rect 2627 291 2727 313
rect 2783 291 2883 313
rect 2939 291 3039 313
rect 3095 291 3195 313
rect 3251 291 3351 313
rect 3407 291 3507 313
rect 3563 291 3663 313
rect 3719 291 3819 313
rect 3875 291 3975 313
rect 4031 291 4131 313
rect 4187 291 4287 313
rect 4343 291 4443 313
rect 4499 291 4599 313
rect 4655 291 4755 313
rect 4811 291 4911 313
rect 4967 291 5067 313
rect 5123 291 5223 313
rect 5279 291 5379 313
rect 5435 291 5535 313
rect 5591 291 5691 313
rect 5747 291 5847 313
rect 5903 291 6003 313
rect 6059 291 6159 313
rect 6215 291 6315 313
rect 6371 291 6471 313
rect 6527 291 6627 313
rect 83 115 183 141
rect 239 115 339 141
rect 395 115 495 141
rect 551 115 651 141
rect 707 115 807 141
rect 863 115 963 141
rect 1019 115 1119 141
rect 1175 115 1275 141
rect 1331 115 1431 141
rect 1487 115 1587 141
rect 1691 115 1791 141
rect 1847 115 1947 141
rect 2003 115 2103 141
rect 2159 115 2259 141
rect 2315 115 2415 141
rect 2471 115 2571 141
rect 2627 115 2727 141
rect 2783 115 2883 141
rect 2939 115 3039 141
rect 3095 115 3195 141
rect 3251 115 3351 141
rect 3407 115 3507 141
rect 3563 115 3663 141
rect 3719 115 3819 141
rect 3875 115 3975 141
rect 4031 115 4131 141
rect 4187 115 4287 141
rect 4343 115 4443 141
rect 4499 115 4599 141
rect 4655 115 4755 141
rect 4811 115 4911 141
rect 4967 115 5067 141
rect 5123 115 5223 141
rect 5279 115 5379 141
rect 5435 115 5535 141
rect 5591 115 5691 141
rect 5747 115 5847 141
rect 5903 115 6003 141
rect 6059 115 6159 141
rect 6215 115 6315 141
rect 6371 115 6471 141
rect 6527 115 6627 141
<< polycont >>
rect 60 329 94 363
rect 128 329 162 363
rect 196 329 230 363
rect 264 329 298 363
rect 332 329 366 363
rect 400 329 434 363
rect 468 329 502 363
rect 536 329 570 363
rect 604 329 638 363
rect 672 329 706 363
rect 740 329 774 363
rect 808 329 842 363
rect 876 329 910 363
rect 1920 329 1954 363
rect 1988 329 2022 363
rect 2232 329 2266 363
rect 2300 329 2334 363
rect 2544 329 2578 363
rect 2612 329 2646 363
rect 2856 329 2890 363
rect 2924 329 2958 363
rect 3168 329 3202 363
rect 3236 329 3270 363
rect 3480 329 3514 363
rect 3548 329 3582 363
rect 3792 329 3826 363
rect 3860 329 3894 363
rect 4102 329 4136 363
rect 4170 329 4204 363
rect 4416 329 4450 363
rect 4484 329 4518 363
rect 4728 329 4762 363
rect 4796 329 4830 363
rect 5040 329 5074 363
rect 5108 329 5142 363
rect 5352 329 5386 363
rect 5420 329 5454 363
rect 5664 329 5698 363
rect 5732 329 5766 363
rect 5976 329 6010 363
rect 6044 329 6078 363
rect 6288 329 6322 363
rect 6356 329 6390 363
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4063 831
rect 4097 797 4159 831
rect 4193 797 4255 831
rect 4289 797 4351 831
rect 4385 797 4447 831
rect 4481 797 4543 831
rect 4577 797 4639 831
rect 4673 797 4735 831
rect 4769 797 4831 831
rect 4865 797 4927 831
rect 4961 797 5023 831
rect 5057 797 5119 831
rect 5153 797 5215 831
rect 5249 797 5311 831
rect 5345 797 5407 831
rect 5441 797 5503 831
rect 5537 797 5599 831
rect 5633 797 5695 831
rect 5729 797 5791 831
rect 5825 797 5887 831
rect 5921 797 5983 831
rect 6017 797 6079 831
rect 6113 797 6175 831
rect 6209 797 6271 831
rect 6305 797 6367 831
rect 6401 797 6463 831
rect 6497 797 6559 831
rect 6593 797 6655 831
rect 6689 797 6720 831
rect 22 731 136 751
rect 22 729 38 731
rect 72 729 136 731
rect 22 695 30 729
rect 72 697 102 729
rect 64 695 102 697
rect 22 642 136 695
rect 22 608 38 642
rect 72 608 136 642
rect 22 562 136 608
rect 22 528 38 562
rect 72 528 136 562
rect 22 489 136 528
rect 22 455 38 489
rect 72 455 136 489
rect 22 435 136 455
rect 170 735 232 751
rect 480 735 542 751
rect 788 735 858 751
rect 1104 735 1166 751
rect 1412 735 1482 751
rect 1786 735 1852 751
rect 170 701 194 735
rect 228 701 232 735
rect 170 642 232 701
rect 170 608 194 642
rect 228 608 232 642
rect 170 558 232 608
rect 170 524 194 558
rect 228 524 232 558
rect 170 485 232 524
rect 268 731 446 735
rect 268 729 350 731
rect 384 729 446 731
rect 302 695 340 729
rect 384 697 412 729
rect 374 695 412 697
rect 268 663 446 695
rect 268 629 350 663
rect 384 629 446 663
rect 268 595 446 629
rect 268 561 350 595
rect 384 561 446 595
rect 268 527 446 561
rect 268 493 350 527
rect 384 493 446 527
rect 268 489 446 493
rect 480 701 506 735
rect 540 701 542 735
rect 480 642 542 701
rect 480 608 506 642
rect 540 608 542 642
rect 480 558 542 608
rect 480 524 506 558
rect 540 524 542 558
rect 170 451 194 485
rect 228 453 232 485
rect 480 485 542 524
rect 576 731 754 735
rect 576 729 662 731
rect 696 729 754 731
rect 610 695 648 729
rect 696 697 720 729
rect 682 695 720 697
rect 576 663 754 695
rect 576 629 662 663
rect 696 629 754 663
rect 576 595 754 629
rect 576 561 662 595
rect 696 561 754 595
rect 576 527 754 561
rect 576 493 662 527
rect 696 493 754 527
rect 576 489 754 493
rect 788 701 818 735
rect 852 701 858 735
rect 788 642 858 701
rect 788 608 818 642
rect 852 608 858 642
rect 788 558 858 608
rect 788 524 818 558
rect 852 524 858 558
rect 480 453 506 485
rect 228 451 506 453
rect 540 453 542 485
rect 788 485 858 524
rect 892 731 1070 735
rect 892 729 974 731
rect 1008 729 1070 731
rect 926 695 964 729
rect 1008 697 1036 729
rect 998 695 1036 697
rect 892 663 1070 695
rect 892 629 974 663
rect 1008 629 1070 663
rect 892 595 1070 629
rect 892 561 974 595
rect 1008 561 1070 595
rect 892 527 1070 561
rect 892 493 974 527
rect 1008 493 1070 527
rect 892 489 1070 493
rect 1104 701 1130 735
rect 1164 701 1166 735
rect 1104 642 1166 701
rect 1104 608 1130 642
rect 1164 608 1166 642
rect 1104 558 1166 608
rect 1104 524 1130 558
rect 1164 524 1166 558
rect 788 453 818 485
rect 540 451 818 453
rect 852 453 858 485
rect 1104 485 1166 524
rect 1200 731 1378 735
rect 1200 729 1286 731
rect 1320 729 1378 731
rect 1234 695 1272 729
rect 1320 697 1344 729
rect 1306 695 1344 697
rect 1200 663 1378 695
rect 1200 629 1286 663
rect 1320 629 1378 663
rect 1200 595 1378 629
rect 1200 561 1286 595
rect 1320 561 1378 595
rect 1200 527 1378 561
rect 1200 493 1286 527
rect 1320 493 1378 527
rect 1200 489 1378 493
rect 1412 701 1442 735
rect 1476 701 1482 735
rect 1412 642 1482 701
rect 1412 608 1442 642
rect 1476 608 1482 642
rect 1412 558 1482 608
rect 1412 524 1442 558
rect 1476 524 1482 558
rect 1104 453 1130 485
rect 852 451 1130 453
rect 1164 453 1166 485
rect 1412 485 1482 524
rect 1412 453 1442 485
rect 1164 451 1442 453
rect 1476 451 1482 485
rect 170 397 1482 451
rect 1516 731 1696 735
rect 1516 729 1598 731
rect 1632 729 1696 731
rect 1550 695 1588 729
rect 1632 697 1660 729
rect 1622 695 1660 697
rect 1694 695 1696 729
rect 1516 663 1696 695
rect 1516 629 1646 663
rect 1680 629 1696 663
rect 1516 553 1696 629
rect 1516 519 1598 553
rect 1632 519 1696 553
rect 1516 485 1696 519
rect 1516 451 1646 485
rect 1680 451 1696 485
rect 1516 447 1696 451
rect 1786 701 1802 735
rect 1836 701 1852 735
rect 1786 656 1852 701
rect 1786 622 1802 656
rect 1836 622 1852 656
rect 1786 576 1852 622
rect 1786 542 1802 576
rect 1836 542 1852 576
rect 1786 498 1852 542
rect 1786 451 1802 498
rect 1836 451 1852 498
rect 44 329 60 363
rect 94 329 128 363
rect 162 329 196 363
rect 230 329 264 363
rect 298 329 332 363
rect 366 329 400 363
rect 434 329 468 363
rect 502 329 536 363
rect 570 329 604 363
rect 638 329 672 363
rect 706 329 740 363
rect 774 329 808 363
rect 842 329 876 363
rect 910 329 926 363
rect 44 316 926 329
rect 960 350 1482 397
rect 960 316 1004 350
rect 1038 316 1076 350
rect 1110 316 1148 350
rect 1182 316 1220 350
rect 1254 316 1292 350
rect 1326 316 1364 350
rect 1398 316 1436 350
rect 1470 316 1482 350
rect 960 282 1482 316
rect 22 273 129 282
rect 22 239 38 273
rect 72 239 129 273
rect 22 205 129 239
rect 22 171 38 205
rect 72 171 129 205
rect 22 119 129 171
rect 163 269 1482 282
rect 1786 283 1852 451
rect 1886 735 2064 751
rect 1886 729 1958 735
rect 1992 729 2064 735
rect 1920 695 1958 729
rect 1992 695 2030 729
rect 1886 656 2064 695
rect 1886 622 1958 656
rect 1992 622 2064 656
rect 1886 576 2064 622
rect 1886 542 1958 576
rect 1992 542 2064 576
rect 1886 485 2064 542
rect 1886 451 1958 485
rect 1992 451 2064 485
rect 1886 435 2064 451
rect 2098 735 2164 751
rect 2098 701 2114 735
rect 2148 701 2164 735
rect 2098 656 2164 701
rect 2098 622 2114 656
rect 2148 622 2164 656
rect 2098 576 2164 622
rect 2098 542 2114 576
rect 2148 542 2164 576
rect 2098 498 2164 542
rect 2098 451 2114 498
rect 2148 451 2164 498
rect 1904 363 2038 379
rect 1904 350 1920 363
rect 1904 316 1918 350
rect 1954 329 1988 363
rect 2022 350 2038 363
rect 1952 316 1990 329
rect 2024 316 2038 350
rect 1904 313 2038 316
rect 163 235 194 269
rect 228 264 1482 269
rect 228 239 506 264
rect 228 235 234 239
rect 163 201 234 235
rect 480 230 506 239
rect 540 239 818 264
rect 540 230 558 239
rect 163 167 194 201
rect 228 167 234 201
rect 163 151 234 167
rect 268 171 350 205
rect 384 171 446 205
rect 22 85 23 119
rect 57 85 95 119
rect 268 119 446 171
rect 480 196 558 230
rect 805 230 818 239
rect 852 239 1130 264
rect 852 230 854 239
rect 480 162 506 196
rect 540 162 558 196
rect 480 146 558 162
rect 592 171 662 205
rect 696 171 771 205
rect 302 85 340 119
rect 374 85 412 119
rect 592 119 771 171
rect 805 196 854 230
rect 1104 230 1130 239
rect 1164 239 1442 264
rect 1164 230 1182 239
rect 805 162 818 196
rect 852 162 854 196
rect 805 146 854 162
rect 888 201 1066 205
rect 888 167 974 201
rect 1008 167 1066 201
rect 626 85 664 119
rect 698 85 736 119
rect 770 85 771 119
rect 888 119 1066 167
rect 1104 196 1182 230
rect 1429 230 1442 239
rect 1476 239 1482 264
rect 1516 269 1696 279
rect 1476 230 1478 239
rect 1104 162 1130 196
rect 1164 162 1182 196
rect 1104 146 1182 162
rect 1216 171 1286 205
rect 1320 171 1395 205
rect 922 85 960 119
rect 994 85 1032 119
rect 1216 119 1395 171
rect 1429 196 1478 230
rect 1516 235 1646 269
rect 1680 235 1696 269
rect 1516 205 1696 235
rect 1429 162 1442 196
rect 1476 162 1478 196
rect 1429 146 1478 162
rect 1512 201 1696 205
rect 1512 167 1598 201
rect 1632 167 1696 201
rect 1250 85 1288 119
rect 1322 85 1360 119
rect 1394 85 1395 119
rect 1512 119 1696 167
rect 1786 249 1802 283
rect 1836 249 1852 283
rect 2098 283 2164 451
rect 2198 735 2376 751
rect 2198 729 2270 735
rect 2304 729 2376 735
rect 2232 695 2270 729
rect 2304 695 2342 729
rect 2198 656 2376 695
rect 2198 622 2270 656
rect 2304 622 2376 656
rect 2198 576 2376 622
rect 2198 542 2270 576
rect 2304 542 2376 576
rect 2198 485 2376 542
rect 2198 451 2270 485
rect 2304 451 2376 485
rect 2198 435 2376 451
rect 2410 735 2476 751
rect 2410 701 2426 735
rect 2460 701 2476 735
rect 2410 656 2476 701
rect 2410 622 2426 656
rect 2460 622 2476 656
rect 2410 576 2476 622
rect 2410 542 2426 576
rect 2460 542 2476 576
rect 2410 498 2476 542
rect 2410 451 2426 498
rect 2460 451 2476 498
rect 2216 363 2350 379
rect 2216 350 2232 363
rect 2216 316 2230 350
rect 2266 329 2300 363
rect 2334 350 2350 363
rect 2264 316 2302 329
rect 2336 316 2350 350
rect 2216 313 2350 316
rect 1786 208 1852 249
rect 1786 174 1802 208
rect 1836 174 1852 208
rect 1786 158 1852 174
rect 1886 269 2064 279
rect 1886 235 1958 269
rect 1992 235 2064 269
rect 1886 201 2064 235
rect 1886 167 1958 201
rect 1992 167 2064 201
rect 1546 85 1584 119
rect 1618 85 1656 119
rect 1690 85 1696 119
rect 1886 119 2064 167
rect 2098 249 2114 283
rect 2148 249 2164 283
rect 2410 283 2476 451
rect 2510 735 2688 751
rect 2510 729 2582 735
rect 2616 729 2688 735
rect 2544 695 2582 729
rect 2616 695 2654 729
rect 2510 656 2688 695
rect 2510 622 2582 656
rect 2616 622 2688 656
rect 2510 576 2688 622
rect 2510 542 2582 576
rect 2616 542 2688 576
rect 2510 485 2688 542
rect 2510 451 2582 485
rect 2616 451 2688 485
rect 2510 435 2688 451
rect 2722 735 2788 751
rect 2722 701 2738 735
rect 2772 701 2788 735
rect 2722 656 2788 701
rect 2722 622 2738 656
rect 2772 622 2788 656
rect 2722 576 2788 622
rect 2722 542 2738 576
rect 2772 542 2788 576
rect 2722 498 2788 542
rect 2722 451 2738 498
rect 2772 451 2788 498
rect 2528 363 2662 379
rect 2528 350 2544 363
rect 2528 316 2542 350
rect 2578 329 2612 363
rect 2646 350 2662 363
rect 2576 316 2614 329
rect 2648 316 2662 350
rect 2528 313 2662 316
rect 2098 208 2164 249
rect 2098 174 2114 208
rect 2148 174 2164 208
rect 2098 158 2164 174
rect 2198 269 2376 279
rect 2198 235 2270 269
rect 2304 235 2376 269
rect 2198 201 2376 235
rect 2198 167 2270 201
rect 2304 167 2376 201
rect 1920 85 1958 119
rect 1992 85 2030 119
rect 2198 119 2376 167
rect 2410 249 2426 283
rect 2460 249 2476 283
rect 2722 283 2788 451
rect 2822 735 3000 751
rect 2822 729 2894 735
rect 2928 729 3000 735
rect 2856 695 2894 729
rect 2928 695 2966 729
rect 2822 656 3000 695
rect 2822 622 2894 656
rect 2928 622 3000 656
rect 2822 576 3000 622
rect 2822 542 2894 576
rect 2928 542 3000 576
rect 2822 485 3000 542
rect 2822 451 2894 485
rect 2928 451 3000 485
rect 2822 435 3000 451
rect 3034 735 3100 751
rect 3034 701 3050 735
rect 3084 701 3100 735
rect 3034 656 3100 701
rect 3034 622 3050 656
rect 3084 622 3100 656
rect 3034 576 3100 622
rect 3034 542 3050 576
rect 3084 542 3100 576
rect 3034 498 3100 542
rect 3034 451 3050 498
rect 3084 451 3100 498
rect 2840 363 2974 379
rect 2840 350 2856 363
rect 2840 316 2854 350
rect 2890 329 2924 363
rect 2958 350 2974 363
rect 2888 316 2926 329
rect 2960 316 2974 350
rect 2840 313 2974 316
rect 2410 208 2476 249
rect 2410 174 2426 208
rect 2460 174 2476 208
rect 2410 158 2476 174
rect 2510 269 2688 279
rect 2510 235 2582 269
rect 2616 235 2688 269
rect 2510 201 2688 235
rect 2510 167 2582 201
rect 2616 167 2688 201
rect 2232 85 2270 119
rect 2304 85 2342 119
rect 2510 119 2688 167
rect 2722 249 2738 283
rect 2772 249 2788 283
rect 3034 283 3100 451
rect 3134 735 3312 751
rect 3134 729 3206 735
rect 3240 729 3312 735
rect 3168 695 3206 729
rect 3240 695 3278 729
rect 3134 656 3312 695
rect 3134 622 3206 656
rect 3240 622 3312 656
rect 3134 576 3312 622
rect 3134 542 3206 576
rect 3240 542 3312 576
rect 3134 485 3312 542
rect 3134 451 3206 485
rect 3240 451 3312 485
rect 3134 435 3312 451
rect 3346 735 3412 751
rect 3346 701 3362 735
rect 3396 701 3412 735
rect 3346 656 3412 701
rect 3346 622 3362 656
rect 3396 622 3412 656
rect 3346 576 3412 622
rect 3346 542 3362 576
rect 3396 542 3412 576
rect 3346 498 3412 542
rect 3346 451 3362 498
rect 3396 451 3412 498
rect 3152 363 3286 379
rect 3152 350 3168 363
rect 3152 316 3166 350
rect 3202 329 3236 363
rect 3270 350 3286 363
rect 3200 316 3238 329
rect 3272 316 3286 350
rect 3152 313 3286 316
rect 2722 208 2788 249
rect 2722 174 2738 208
rect 2772 174 2788 208
rect 2722 158 2788 174
rect 2822 269 3000 279
rect 2822 235 2894 269
rect 2928 235 3000 269
rect 2822 201 3000 235
rect 2822 167 2894 201
rect 2928 167 3000 201
rect 2544 85 2582 119
rect 2616 85 2654 119
rect 2822 119 3000 167
rect 3034 249 3050 283
rect 3084 249 3100 283
rect 3346 283 3412 451
rect 3446 735 3624 751
rect 3446 729 3518 735
rect 3552 729 3624 735
rect 3480 695 3518 729
rect 3552 695 3590 729
rect 3446 656 3624 695
rect 3446 622 3518 656
rect 3552 622 3624 656
rect 3446 576 3624 622
rect 3446 542 3518 576
rect 3552 542 3624 576
rect 3446 485 3624 542
rect 3446 451 3518 485
rect 3552 451 3624 485
rect 3446 435 3624 451
rect 3658 735 3724 751
rect 3658 701 3674 735
rect 3708 701 3724 735
rect 3658 656 3724 701
rect 3658 622 3674 656
rect 3708 622 3724 656
rect 3658 576 3724 622
rect 3658 542 3674 576
rect 3708 542 3724 576
rect 3658 498 3724 542
rect 3658 451 3674 498
rect 3708 451 3724 498
rect 3464 363 3598 379
rect 3464 350 3480 363
rect 3464 316 3478 350
rect 3514 329 3548 363
rect 3582 350 3598 363
rect 3512 316 3550 329
rect 3584 316 3598 350
rect 3464 313 3598 316
rect 3034 208 3100 249
rect 3034 174 3050 208
rect 3084 174 3100 208
rect 3034 158 3100 174
rect 3134 269 3312 279
rect 3134 235 3206 269
rect 3240 235 3312 269
rect 3134 201 3312 235
rect 3134 167 3206 201
rect 3240 167 3312 201
rect 2856 85 2894 119
rect 2928 85 2966 119
rect 3134 119 3312 167
rect 3346 249 3362 283
rect 3396 249 3412 283
rect 3658 283 3724 451
rect 3758 735 3936 751
rect 3758 729 3830 735
rect 3864 729 3936 735
rect 3792 695 3830 729
rect 3864 695 3902 729
rect 3758 656 3936 695
rect 3758 622 3830 656
rect 3864 622 3936 656
rect 3758 576 3936 622
rect 3758 542 3830 576
rect 3864 542 3936 576
rect 3758 485 3936 542
rect 3758 451 3830 485
rect 3864 451 3936 485
rect 3758 435 3936 451
rect 3970 735 4052 751
rect 3970 701 3986 735
rect 4020 701 4052 735
rect 3970 656 4052 701
rect 3970 622 3986 656
rect 4020 622 4052 656
rect 3970 576 4052 622
rect 3970 542 3986 576
rect 4020 542 4052 576
rect 3970 498 4052 542
rect 3970 451 3986 498
rect 4020 451 4052 498
rect 3776 363 3910 379
rect 3776 350 3792 363
rect 3776 316 3790 350
rect 3826 329 3860 363
rect 3894 350 3910 363
rect 3824 316 3862 329
rect 3896 316 3910 350
rect 3776 313 3910 316
rect 3346 208 3412 249
rect 3346 174 3362 208
rect 3396 174 3412 208
rect 3346 158 3412 174
rect 3446 269 3624 279
rect 3446 235 3518 269
rect 3552 235 3624 269
rect 3446 201 3624 235
rect 3446 167 3518 201
rect 3552 167 3624 201
rect 3168 85 3206 119
rect 3240 85 3278 119
rect 3446 119 3624 167
rect 3658 249 3674 283
rect 3708 249 3724 283
rect 3970 283 4052 451
rect 4086 731 4192 751
rect 4086 729 4142 731
rect 4176 729 4192 731
rect 4120 697 4142 729
rect 4120 695 4158 697
rect 4086 656 4192 695
rect 4086 622 4142 656
rect 4176 622 4192 656
rect 4086 576 4192 622
rect 4086 542 4142 576
rect 4176 542 4192 576
rect 4086 489 4192 542
rect 4086 455 4142 489
rect 4176 455 4192 489
rect 4086 435 4192 455
rect 4282 735 4348 751
rect 4282 701 4298 735
rect 4332 701 4348 735
rect 4282 656 4348 701
rect 4282 622 4298 656
rect 4332 622 4348 656
rect 4282 576 4348 622
rect 4282 542 4298 576
rect 4332 542 4348 576
rect 4282 498 4348 542
rect 4282 451 4298 498
rect 4332 451 4348 498
rect 4086 363 4220 379
rect 4086 350 4102 363
rect 4086 316 4100 350
rect 4136 329 4170 363
rect 4204 350 4220 363
rect 4134 316 4172 329
rect 4206 316 4220 350
rect 4086 313 4220 316
rect 3658 208 3724 249
rect 3658 174 3674 208
rect 3708 174 3724 208
rect 3658 158 3724 174
rect 3758 269 3936 279
rect 3758 235 3830 269
rect 3864 235 3936 269
rect 3758 201 3936 235
rect 3758 167 3830 201
rect 3864 167 3936 201
rect 3480 85 3518 119
rect 3552 85 3590 119
rect 3758 119 3936 167
rect 3970 249 3986 283
rect 4020 249 4052 283
rect 4282 283 4348 451
rect 4382 735 4560 751
rect 4382 729 4454 735
rect 4488 729 4560 735
rect 4416 695 4454 729
rect 4488 695 4526 729
rect 4382 656 4560 695
rect 4382 622 4454 656
rect 4488 622 4560 656
rect 4382 576 4560 622
rect 4382 542 4454 576
rect 4488 542 4560 576
rect 4382 485 4560 542
rect 4382 451 4454 485
rect 4488 451 4560 485
rect 4382 435 4560 451
rect 4594 735 4660 751
rect 4594 701 4610 735
rect 4644 701 4660 735
rect 4594 656 4660 701
rect 4594 622 4610 656
rect 4644 622 4660 656
rect 4594 576 4660 622
rect 4594 542 4610 576
rect 4644 542 4660 576
rect 4594 498 4660 542
rect 4594 451 4610 498
rect 4644 451 4660 498
rect 4400 363 4534 379
rect 4400 350 4416 363
rect 4400 316 4414 350
rect 4450 329 4484 363
rect 4518 350 4534 363
rect 4448 316 4486 329
rect 4520 316 4534 350
rect 4400 313 4534 316
rect 3970 208 4052 249
rect 3970 174 3986 208
rect 4020 174 4052 208
rect 3970 158 4052 174
rect 4086 269 4192 279
rect 4086 235 4142 269
rect 4176 235 4192 269
rect 4086 198 4192 235
rect 4086 164 4142 198
rect 4176 164 4192 198
rect 3792 85 3830 119
rect 3864 85 3902 119
rect 4086 119 4192 164
rect 4282 249 4298 283
rect 4332 249 4348 283
rect 4594 283 4660 451
rect 4694 735 4872 751
rect 4694 729 4766 735
rect 4800 729 4872 735
rect 4728 695 4766 729
rect 4800 695 4838 729
rect 4694 656 4872 695
rect 4694 622 4766 656
rect 4800 622 4872 656
rect 4694 576 4872 622
rect 4694 542 4766 576
rect 4800 542 4872 576
rect 4694 485 4872 542
rect 4694 451 4766 485
rect 4800 451 4872 485
rect 4694 435 4872 451
rect 4906 735 4972 751
rect 4906 701 4922 735
rect 4956 701 4972 735
rect 4906 656 4972 701
rect 4906 622 4922 656
rect 4956 622 4972 656
rect 4906 576 4972 622
rect 4906 542 4922 576
rect 4956 542 4972 576
rect 4906 498 4972 542
rect 4906 451 4922 498
rect 4956 451 4972 498
rect 4712 363 4846 379
rect 4712 350 4728 363
rect 4712 316 4726 350
rect 4762 329 4796 363
rect 4830 350 4846 363
rect 4760 316 4798 329
rect 4832 316 4846 350
rect 4712 313 4846 316
rect 4282 208 4348 249
rect 4282 174 4298 208
rect 4332 174 4348 208
rect 4282 158 4348 174
rect 4382 269 4560 279
rect 4382 235 4454 269
rect 4488 235 4560 269
rect 4382 201 4560 235
rect 4382 167 4454 201
rect 4488 167 4560 201
rect 4120 85 4158 119
rect 4382 119 4560 167
rect 4594 249 4610 283
rect 4644 249 4660 283
rect 4906 283 4972 451
rect 5006 735 5184 751
rect 5006 729 5078 735
rect 5112 729 5184 735
rect 5040 695 5078 729
rect 5112 695 5150 729
rect 5006 656 5184 695
rect 5006 622 5078 656
rect 5112 622 5184 656
rect 5006 576 5184 622
rect 5006 542 5078 576
rect 5112 542 5184 576
rect 5006 485 5184 542
rect 5006 451 5078 485
rect 5112 451 5184 485
rect 5006 435 5184 451
rect 5218 735 5284 751
rect 5218 701 5234 735
rect 5268 701 5284 735
rect 5218 656 5284 701
rect 5218 622 5234 656
rect 5268 622 5284 656
rect 5218 576 5284 622
rect 5218 542 5234 576
rect 5268 542 5284 576
rect 5218 498 5284 542
rect 5218 451 5234 498
rect 5268 451 5284 498
rect 5024 363 5158 379
rect 5024 350 5040 363
rect 5024 316 5038 350
rect 5074 329 5108 363
rect 5142 350 5158 363
rect 5072 316 5110 329
rect 5144 316 5158 350
rect 5024 313 5158 316
rect 4594 208 4660 249
rect 4594 174 4610 208
rect 4644 174 4660 208
rect 4594 158 4660 174
rect 4694 269 4872 279
rect 4694 235 4766 269
rect 4800 235 4872 269
rect 4694 201 4872 235
rect 4694 167 4766 201
rect 4800 167 4872 201
rect 4416 85 4454 119
rect 4488 85 4526 119
rect 4694 119 4872 167
rect 4906 249 4922 283
rect 4956 249 4972 283
rect 5218 283 5284 451
rect 5318 735 5496 751
rect 5318 729 5390 735
rect 5424 729 5496 735
rect 5352 695 5390 729
rect 5424 695 5462 729
rect 5318 656 5496 695
rect 5318 622 5390 656
rect 5424 622 5496 656
rect 5318 576 5496 622
rect 5318 542 5390 576
rect 5424 542 5496 576
rect 5318 485 5496 542
rect 5318 451 5390 485
rect 5424 451 5496 485
rect 5318 435 5496 451
rect 5530 735 5596 751
rect 5530 701 5546 735
rect 5580 701 5596 735
rect 5530 656 5596 701
rect 5530 622 5546 656
rect 5580 622 5596 656
rect 5530 576 5596 622
rect 5530 542 5546 576
rect 5580 542 5596 576
rect 5530 498 5596 542
rect 5530 451 5546 498
rect 5580 451 5596 498
rect 5336 363 5470 379
rect 5336 350 5352 363
rect 5336 316 5350 350
rect 5386 329 5420 363
rect 5454 350 5470 363
rect 5384 316 5422 329
rect 5456 316 5470 350
rect 5336 313 5470 316
rect 4906 208 4972 249
rect 4906 174 4922 208
rect 4956 174 4972 208
rect 4906 158 4972 174
rect 5006 269 5184 279
rect 5006 235 5078 269
rect 5112 235 5184 269
rect 5006 201 5184 235
rect 5006 167 5078 201
rect 5112 167 5184 201
rect 4728 85 4766 119
rect 4800 85 4838 119
rect 5006 119 5184 167
rect 5218 249 5234 283
rect 5268 249 5284 283
rect 5530 283 5596 451
rect 5630 735 5808 751
rect 5630 729 5702 735
rect 5736 729 5808 735
rect 5664 695 5702 729
rect 5736 695 5774 729
rect 5630 656 5808 695
rect 5630 622 5702 656
rect 5736 622 5808 656
rect 5630 576 5808 622
rect 5630 542 5702 576
rect 5736 542 5808 576
rect 5630 485 5808 542
rect 5630 451 5702 485
rect 5736 451 5808 485
rect 5630 435 5808 451
rect 5842 735 5908 751
rect 5842 701 5858 735
rect 5892 701 5908 735
rect 5842 656 5908 701
rect 5842 622 5858 656
rect 5892 622 5908 656
rect 5842 576 5908 622
rect 5842 542 5858 576
rect 5892 542 5908 576
rect 5842 498 5908 542
rect 5842 451 5858 498
rect 5892 451 5908 498
rect 5648 363 5782 379
rect 5648 350 5664 363
rect 5648 316 5662 350
rect 5698 329 5732 363
rect 5766 350 5782 363
rect 5696 316 5734 329
rect 5768 316 5782 350
rect 5648 313 5782 316
rect 5218 208 5284 249
rect 5218 174 5234 208
rect 5268 174 5284 208
rect 5218 158 5284 174
rect 5318 269 5496 279
rect 5318 235 5390 269
rect 5424 235 5496 269
rect 5318 201 5496 235
rect 5318 167 5390 201
rect 5424 167 5496 201
rect 5040 85 5078 119
rect 5112 85 5150 119
rect 5318 119 5496 167
rect 5530 249 5546 283
rect 5580 249 5596 283
rect 5842 283 5908 451
rect 5942 735 6120 751
rect 5942 729 6014 735
rect 6048 729 6120 735
rect 5976 695 6014 729
rect 6048 695 6086 729
rect 5942 656 6120 695
rect 5942 622 6014 656
rect 6048 622 6120 656
rect 5942 576 6120 622
rect 5942 542 6014 576
rect 6048 542 6120 576
rect 5942 485 6120 542
rect 5942 451 6014 485
rect 6048 451 6120 485
rect 5942 435 6120 451
rect 6154 735 6220 751
rect 6154 701 6170 735
rect 6204 701 6220 735
rect 6154 656 6220 701
rect 6154 622 6170 656
rect 6204 622 6220 656
rect 6154 576 6220 622
rect 6154 542 6170 576
rect 6204 542 6220 576
rect 6154 498 6220 542
rect 6154 451 6170 498
rect 6204 451 6220 498
rect 5960 363 6094 379
rect 5960 350 5976 363
rect 5960 316 5974 350
rect 6010 329 6044 363
rect 6078 350 6094 363
rect 6008 316 6046 329
rect 6080 316 6094 350
rect 5960 313 6094 316
rect 5530 208 5596 249
rect 5530 174 5546 208
rect 5580 174 5596 208
rect 5530 158 5596 174
rect 5630 269 5808 279
rect 5630 235 5702 269
rect 5736 235 5808 269
rect 5630 201 5808 235
rect 5630 167 5702 201
rect 5736 167 5808 201
rect 5352 85 5390 119
rect 5424 85 5462 119
rect 5630 119 5808 167
rect 5842 249 5858 283
rect 5892 249 5908 283
rect 6154 283 6220 451
rect 6254 735 6432 751
rect 6254 729 6326 735
rect 6360 729 6432 735
rect 6288 695 6326 729
rect 6360 695 6398 729
rect 6254 656 6432 695
rect 6254 622 6326 656
rect 6360 622 6432 656
rect 6254 576 6432 622
rect 6254 542 6326 576
rect 6360 542 6432 576
rect 6254 485 6432 542
rect 6254 451 6326 485
rect 6360 451 6432 485
rect 6254 435 6432 451
rect 6466 735 6548 751
rect 6466 701 6482 735
rect 6516 701 6548 735
rect 6466 656 6548 701
rect 6466 622 6482 656
rect 6516 622 6548 656
rect 6466 576 6548 622
rect 6466 542 6482 576
rect 6516 542 6548 576
rect 6466 498 6548 542
rect 6466 451 6482 498
rect 6516 451 6548 498
rect 6272 363 6406 379
rect 6272 350 6288 363
rect 6272 316 6286 350
rect 6322 329 6356 363
rect 6390 350 6406 363
rect 6320 316 6358 329
rect 6392 316 6406 350
rect 6272 313 6406 316
rect 5842 208 5908 249
rect 5842 174 5858 208
rect 5892 174 5908 208
rect 5842 158 5908 174
rect 5942 269 6120 279
rect 5942 235 6014 269
rect 6048 235 6120 269
rect 5942 201 6120 235
rect 5942 167 6014 201
rect 6048 167 6120 201
rect 5664 85 5702 119
rect 5736 85 5774 119
rect 5942 119 6120 167
rect 6154 249 6170 283
rect 6204 249 6220 283
rect 6466 283 6548 451
rect 6582 731 6688 751
rect 6582 729 6638 731
rect 6672 729 6688 731
rect 6616 697 6638 729
rect 6616 695 6654 697
rect 6582 656 6688 695
rect 6582 622 6638 656
rect 6672 622 6688 656
rect 6582 576 6688 622
rect 6582 542 6638 576
rect 6672 542 6688 576
rect 6582 489 6688 542
rect 6582 455 6638 489
rect 6672 455 6688 489
rect 6582 435 6688 455
rect 6154 208 6220 249
rect 6154 174 6170 208
rect 6204 174 6220 208
rect 6154 158 6220 174
rect 6254 269 6432 279
rect 6254 235 6326 269
rect 6360 235 6432 269
rect 6254 201 6432 235
rect 6254 167 6326 201
rect 6360 167 6432 201
rect 5976 85 6014 119
rect 6048 85 6086 119
rect 6254 119 6432 167
rect 6466 249 6482 283
rect 6516 249 6548 283
rect 6466 208 6548 249
rect 6466 174 6482 208
rect 6516 174 6548 208
rect 6466 158 6548 174
rect 6582 279 6688 299
rect 6582 245 6638 279
rect 6672 245 6688 279
rect 6582 208 6688 245
rect 6582 174 6638 208
rect 6672 174 6688 208
rect 6288 85 6326 119
rect 6360 85 6398 119
rect 6582 119 6688 174
rect 6616 85 6654 119
rect 268 83 446 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 5023 17
rect 5057 -17 5119 17
rect 5153 -17 5215 17
rect 5249 -17 5311 17
rect 5345 -17 5407 17
rect 5441 -17 5503 17
rect 5537 -17 5599 17
rect 5633 -17 5695 17
rect 5729 -17 5791 17
rect 5825 -17 5887 17
rect 5921 -17 5983 17
rect 6017 -17 6079 17
rect 6113 -17 6175 17
rect 6209 -17 6271 17
rect 6305 -17 6367 17
rect 6401 -17 6463 17
rect 6497 -17 6559 17
rect 6593 -17 6655 17
rect 6689 -17 6720 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
rect 4063 797 4097 831
rect 4159 797 4193 831
rect 4255 797 4289 831
rect 4351 797 4385 831
rect 4447 797 4481 831
rect 4543 797 4577 831
rect 4639 797 4673 831
rect 4735 797 4769 831
rect 4831 797 4865 831
rect 4927 797 4961 831
rect 5023 797 5057 831
rect 5119 797 5153 831
rect 5215 797 5249 831
rect 5311 797 5345 831
rect 5407 797 5441 831
rect 5503 797 5537 831
rect 5599 797 5633 831
rect 5695 797 5729 831
rect 5791 797 5825 831
rect 5887 797 5921 831
rect 5983 797 6017 831
rect 6079 797 6113 831
rect 6175 797 6209 831
rect 6271 797 6305 831
rect 6367 797 6401 831
rect 6463 797 6497 831
rect 6559 797 6593 831
rect 6655 797 6689 831
rect 30 697 38 729
rect 38 697 64 729
rect 30 695 64 697
rect 102 695 136 729
rect 268 695 302 729
rect 340 697 350 729
rect 350 697 374 729
rect 340 695 374 697
rect 412 695 446 729
rect 576 695 610 729
rect 648 697 662 729
rect 662 697 682 729
rect 648 695 682 697
rect 720 695 754 729
rect 892 695 926 729
rect 964 697 974 729
rect 974 697 998 729
rect 964 695 998 697
rect 1036 695 1070 729
rect 1200 695 1234 729
rect 1272 697 1286 729
rect 1286 697 1306 729
rect 1272 695 1306 697
rect 1344 695 1378 729
rect 1516 695 1550 729
rect 1588 697 1598 729
rect 1598 697 1622 729
rect 1588 695 1622 697
rect 1660 695 1694 729
rect 1802 485 1836 498
rect 1802 464 1836 485
rect 1004 316 1038 350
rect 1076 316 1110 350
rect 1148 316 1182 350
rect 1220 316 1254 350
rect 1292 316 1326 350
rect 1364 316 1398 350
rect 1436 316 1470 350
rect 1886 695 1920 729
rect 1958 701 1992 729
rect 1958 695 1992 701
rect 2030 695 2064 729
rect 2114 485 2148 498
rect 2114 464 2148 485
rect 1918 329 1920 350
rect 1920 329 1952 350
rect 1990 329 2022 350
rect 2022 329 2024 350
rect 1918 316 1952 329
rect 1990 316 2024 329
rect 23 85 57 119
rect 95 85 129 119
rect 268 85 302 119
rect 340 85 374 119
rect 412 85 446 119
rect 592 85 626 119
rect 664 85 698 119
rect 736 85 770 119
rect 888 85 922 119
rect 960 85 994 119
rect 1032 85 1066 119
rect 1216 85 1250 119
rect 1288 85 1322 119
rect 1360 85 1394 119
rect 2198 695 2232 729
rect 2270 701 2304 729
rect 2270 695 2304 701
rect 2342 695 2376 729
rect 2426 485 2460 498
rect 2426 464 2460 485
rect 2230 329 2232 350
rect 2232 329 2264 350
rect 2302 329 2334 350
rect 2334 329 2336 350
rect 2230 316 2264 329
rect 2302 316 2336 329
rect 1512 85 1546 119
rect 1584 85 1618 119
rect 1656 85 1690 119
rect 2510 695 2544 729
rect 2582 701 2616 729
rect 2582 695 2616 701
rect 2654 695 2688 729
rect 2738 485 2772 498
rect 2738 464 2772 485
rect 2542 329 2544 350
rect 2544 329 2576 350
rect 2614 329 2646 350
rect 2646 329 2648 350
rect 2542 316 2576 329
rect 2614 316 2648 329
rect 1886 85 1920 119
rect 1958 85 1992 119
rect 2030 85 2064 119
rect 2822 695 2856 729
rect 2894 701 2928 729
rect 2894 695 2928 701
rect 2966 695 3000 729
rect 3050 485 3084 498
rect 3050 464 3084 485
rect 2854 329 2856 350
rect 2856 329 2888 350
rect 2926 329 2958 350
rect 2958 329 2960 350
rect 2854 316 2888 329
rect 2926 316 2960 329
rect 2198 85 2232 119
rect 2270 85 2304 119
rect 2342 85 2376 119
rect 3134 695 3168 729
rect 3206 701 3240 729
rect 3206 695 3240 701
rect 3278 695 3312 729
rect 3362 485 3396 498
rect 3362 464 3396 485
rect 3166 329 3168 350
rect 3168 329 3200 350
rect 3238 329 3270 350
rect 3270 329 3272 350
rect 3166 316 3200 329
rect 3238 316 3272 329
rect 2510 85 2544 119
rect 2582 85 2616 119
rect 2654 85 2688 119
rect 3446 695 3480 729
rect 3518 701 3552 729
rect 3518 695 3552 701
rect 3590 695 3624 729
rect 3674 485 3708 498
rect 3674 464 3708 485
rect 3478 329 3480 350
rect 3480 329 3512 350
rect 3550 329 3582 350
rect 3582 329 3584 350
rect 3478 316 3512 329
rect 3550 316 3584 329
rect 2822 85 2856 119
rect 2894 85 2928 119
rect 2966 85 3000 119
rect 3758 695 3792 729
rect 3830 701 3864 729
rect 3830 695 3864 701
rect 3902 695 3936 729
rect 3986 485 4020 498
rect 3986 464 4020 485
rect 3790 329 3792 350
rect 3792 329 3824 350
rect 3862 329 3894 350
rect 3894 329 3896 350
rect 3790 316 3824 329
rect 3862 316 3896 329
rect 3134 85 3168 119
rect 3206 85 3240 119
rect 3278 85 3312 119
rect 4086 695 4120 729
rect 4158 697 4176 729
rect 4176 697 4192 729
rect 4158 695 4192 697
rect 4298 485 4332 498
rect 4298 464 4332 485
rect 4100 329 4102 350
rect 4102 329 4134 350
rect 4172 329 4204 350
rect 4204 329 4206 350
rect 4100 316 4134 329
rect 4172 316 4206 329
rect 3446 85 3480 119
rect 3518 85 3552 119
rect 3590 85 3624 119
rect 4382 695 4416 729
rect 4454 701 4488 729
rect 4454 695 4488 701
rect 4526 695 4560 729
rect 4610 485 4644 498
rect 4610 464 4644 485
rect 4414 329 4416 350
rect 4416 329 4448 350
rect 4486 329 4518 350
rect 4518 329 4520 350
rect 4414 316 4448 329
rect 4486 316 4520 329
rect 3758 85 3792 119
rect 3830 85 3864 119
rect 3902 85 3936 119
rect 4694 695 4728 729
rect 4766 701 4800 729
rect 4766 695 4800 701
rect 4838 695 4872 729
rect 4922 485 4956 498
rect 4922 464 4956 485
rect 4726 329 4728 350
rect 4728 329 4760 350
rect 4798 329 4830 350
rect 4830 329 4832 350
rect 4726 316 4760 329
rect 4798 316 4832 329
rect 4086 85 4120 119
rect 4158 85 4192 119
rect 5006 695 5040 729
rect 5078 701 5112 729
rect 5078 695 5112 701
rect 5150 695 5184 729
rect 5234 485 5268 498
rect 5234 464 5268 485
rect 5038 329 5040 350
rect 5040 329 5072 350
rect 5110 329 5142 350
rect 5142 329 5144 350
rect 5038 316 5072 329
rect 5110 316 5144 329
rect 4382 85 4416 119
rect 4454 85 4488 119
rect 4526 85 4560 119
rect 5318 695 5352 729
rect 5390 701 5424 729
rect 5390 695 5424 701
rect 5462 695 5496 729
rect 5546 485 5580 498
rect 5546 464 5580 485
rect 5350 329 5352 350
rect 5352 329 5384 350
rect 5422 329 5454 350
rect 5454 329 5456 350
rect 5350 316 5384 329
rect 5422 316 5456 329
rect 4694 85 4728 119
rect 4766 85 4800 119
rect 4838 85 4872 119
rect 5630 695 5664 729
rect 5702 701 5736 729
rect 5702 695 5736 701
rect 5774 695 5808 729
rect 5858 485 5892 498
rect 5858 464 5892 485
rect 5662 329 5664 350
rect 5664 329 5696 350
rect 5734 329 5766 350
rect 5766 329 5768 350
rect 5662 316 5696 329
rect 5734 316 5768 329
rect 5006 85 5040 119
rect 5078 85 5112 119
rect 5150 85 5184 119
rect 5942 695 5976 729
rect 6014 701 6048 729
rect 6014 695 6048 701
rect 6086 695 6120 729
rect 6170 485 6204 498
rect 6170 464 6204 485
rect 5974 329 5976 350
rect 5976 329 6008 350
rect 6046 329 6078 350
rect 6078 329 6080 350
rect 5974 316 6008 329
rect 6046 316 6080 329
rect 5318 85 5352 119
rect 5390 85 5424 119
rect 5462 85 5496 119
rect 6254 695 6288 729
rect 6326 701 6360 729
rect 6326 695 6360 701
rect 6398 695 6432 729
rect 6482 485 6516 498
rect 6482 464 6516 485
rect 6286 329 6288 350
rect 6288 329 6320 350
rect 6358 329 6390 350
rect 6390 329 6392 350
rect 6286 316 6320 329
rect 6358 316 6392 329
rect 5630 85 5664 119
rect 5702 85 5736 119
rect 5774 85 5808 119
rect 6582 695 6616 729
rect 6654 697 6672 729
rect 6672 697 6688 729
rect 6654 695 6688 697
rect 5942 85 5976 119
rect 6014 85 6048 119
rect 6086 85 6120 119
rect 6254 85 6288 119
rect 6326 85 6360 119
rect 6398 85 6432 119
rect 6582 85 6616 119
rect 6654 85 6688 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect 4927 -17 4961 17
rect 5023 -17 5057 17
rect 5119 -17 5153 17
rect 5215 -17 5249 17
rect 5311 -17 5345 17
rect 5407 -17 5441 17
rect 5503 -17 5537 17
rect 5599 -17 5633 17
rect 5695 -17 5729 17
rect 5791 -17 5825 17
rect 5887 -17 5921 17
rect 5983 -17 6017 17
rect 6079 -17 6113 17
rect 6175 -17 6209 17
rect 6271 -17 6305 17
rect 6367 -17 6401 17
rect 6463 -17 6497 17
rect 6559 -17 6593 17
rect 6655 -17 6689 17
<< metal1 >>
rect 0 831 6720 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4063 831
rect 4097 797 4159 831
rect 4193 797 4255 831
rect 4289 797 4351 831
rect 4385 797 4447 831
rect 4481 797 4543 831
rect 4577 797 4639 831
rect 4673 797 4735 831
rect 4769 797 4831 831
rect 4865 797 4927 831
rect 4961 797 5023 831
rect 5057 797 5119 831
rect 5153 797 5215 831
rect 5249 797 5311 831
rect 5345 797 5407 831
rect 5441 797 5503 831
rect 5537 797 5599 831
rect 5633 797 5695 831
rect 5729 797 5791 831
rect 5825 797 5887 831
rect 5921 797 5983 831
rect 6017 797 6079 831
rect 6113 797 6175 831
rect 6209 797 6271 831
rect 6305 797 6367 831
rect 6401 797 6463 831
rect 6497 797 6559 831
rect 6593 797 6655 831
rect 6689 797 6720 831
rect 0 791 6720 797
rect 0 729 6720 763
rect 0 695 30 729
rect 64 695 102 729
rect 136 695 268 729
rect 302 695 340 729
rect 374 695 412 729
rect 446 695 576 729
rect 610 695 648 729
rect 682 695 720 729
rect 754 695 892 729
rect 926 695 964 729
rect 998 695 1036 729
rect 1070 695 1200 729
rect 1234 695 1272 729
rect 1306 695 1344 729
rect 1378 695 1516 729
rect 1550 695 1588 729
rect 1622 695 1660 729
rect 1694 695 1886 729
rect 1920 695 1958 729
rect 1992 695 2030 729
rect 2064 695 2198 729
rect 2232 695 2270 729
rect 2304 695 2342 729
rect 2376 695 2510 729
rect 2544 695 2582 729
rect 2616 695 2654 729
rect 2688 695 2822 729
rect 2856 695 2894 729
rect 2928 695 2966 729
rect 3000 695 3134 729
rect 3168 695 3206 729
rect 3240 695 3278 729
rect 3312 695 3446 729
rect 3480 695 3518 729
rect 3552 695 3590 729
rect 3624 695 3758 729
rect 3792 695 3830 729
rect 3864 695 3902 729
rect 3936 695 4086 729
rect 4120 695 4158 729
rect 4192 695 4382 729
rect 4416 695 4454 729
rect 4488 695 4526 729
rect 4560 695 4694 729
rect 4728 695 4766 729
rect 4800 695 4838 729
rect 4872 695 5006 729
rect 5040 695 5078 729
rect 5112 695 5150 729
rect 5184 695 5318 729
rect 5352 695 5390 729
rect 5424 695 5462 729
rect 5496 695 5630 729
rect 5664 695 5702 729
rect 5736 695 5774 729
rect 5808 695 5942 729
rect 5976 695 6014 729
rect 6048 695 6086 729
rect 6120 695 6254 729
rect 6288 695 6326 729
rect 6360 695 6398 729
rect 6432 695 6582 729
rect 6616 695 6654 729
rect 6688 695 6720 729
rect 0 689 6720 695
rect 1790 498 6528 504
rect 1790 464 1802 498
rect 1836 464 2114 498
rect 2148 464 2426 498
rect 2460 464 2738 498
rect 2772 464 3050 498
rect 3084 464 3362 498
rect 3396 464 3674 498
rect 3708 464 3986 498
rect 4020 464 4298 498
rect 4332 464 4610 498
rect 4644 464 4922 498
rect 4956 464 5234 498
rect 5268 464 5546 498
rect 5580 464 5858 498
rect 5892 464 6170 498
rect 6204 464 6482 498
rect 6516 464 6528 498
rect 1790 458 6528 464
rect 992 350 6418 356
rect 992 316 1004 350
rect 1038 316 1076 350
rect 1110 316 1148 350
rect 1182 316 1220 350
rect 1254 316 1292 350
rect 1326 316 1364 350
rect 1398 316 1436 350
rect 1470 316 1918 350
rect 1952 316 1990 350
rect 2024 316 2230 350
rect 2264 316 2302 350
rect 2336 316 2542 350
rect 2576 316 2614 350
rect 2648 316 2854 350
rect 2888 316 2926 350
rect 2960 316 3166 350
rect 3200 316 3238 350
rect 3272 316 3478 350
rect 3512 316 3550 350
rect 3584 316 3790 350
rect 3824 316 3862 350
rect 3896 316 4100 350
rect 4134 316 4172 350
rect 4206 316 4414 350
rect 4448 316 4486 350
rect 4520 316 4726 350
rect 4760 316 4798 350
rect 4832 316 5038 350
rect 5072 316 5110 350
rect 5144 316 5350 350
rect 5384 316 5422 350
rect 5456 316 5662 350
rect 5696 316 5734 350
rect 5768 316 5974 350
rect 6008 316 6046 350
rect 6080 316 6286 350
rect 6320 316 6358 350
rect 6392 316 6418 350
rect 992 310 6418 316
rect 0 119 6720 125
rect 0 85 23 119
rect 57 85 95 119
rect 129 85 268 119
rect 302 85 340 119
rect 374 85 412 119
rect 446 85 592 119
rect 626 85 664 119
rect 698 85 736 119
rect 770 85 888 119
rect 922 85 960 119
rect 994 85 1032 119
rect 1066 85 1216 119
rect 1250 85 1288 119
rect 1322 85 1360 119
rect 1394 85 1512 119
rect 1546 85 1584 119
rect 1618 85 1656 119
rect 1690 85 1886 119
rect 1920 85 1958 119
rect 1992 85 2030 119
rect 2064 85 2198 119
rect 2232 85 2270 119
rect 2304 85 2342 119
rect 2376 85 2510 119
rect 2544 85 2582 119
rect 2616 85 2654 119
rect 2688 85 2822 119
rect 2856 85 2894 119
rect 2928 85 2966 119
rect 3000 85 3134 119
rect 3168 85 3206 119
rect 3240 85 3278 119
rect 3312 85 3446 119
rect 3480 85 3518 119
rect 3552 85 3590 119
rect 3624 85 3758 119
rect 3792 85 3830 119
rect 3864 85 3902 119
rect 3936 85 4086 119
rect 4120 85 4158 119
rect 4192 85 4382 119
rect 4416 85 4454 119
rect 4488 85 4526 119
rect 4560 85 4694 119
rect 4728 85 4766 119
rect 4800 85 4838 119
rect 4872 85 5006 119
rect 5040 85 5078 119
rect 5112 85 5150 119
rect 5184 85 5318 119
rect 5352 85 5390 119
rect 5424 85 5462 119
rect 5496 85 5630 119
rect 5664 85 5702 119
rect 5736 85 5774 119
rect 5808 85 5942 119
rect 5976 85 6014 119
rect 6048 85 6086 119
rect 6120 85 6254 119
rect 6288 85 6326 119
rect 6360 85 6398 119
rect 6432 85 6582 119
rect 6616 85 6654 119
rect 6688 85 6720 119
rect 0 51 6720 85
rect 0 17 6720 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 5023 17
rect 5057 -17 5119 17
rect 5153 -17 5215 17
rect 5249 -17 5311 17
rect 5345 -17 5407 17
rect 5441 -17 5503 17
rect 5537 -17 5599 17
rect 5633 -17 5695 17
rect 5729 -17 5791 17
rect 5825 -17 5887 17
rect 5921 -17 5983 17
rect 6017 -17 6079 17
rect 6113 -17 6175 17
rect 6209 -17 6271 17
rect 6305 -17 6367 17
rect 6401 -17 6463 17
rect 6497 -17 6559 17
rect 6593 -17 6655 17
rect 6689 -17 6720 17
rect 0 -23 6720 -17
<< labels >>
rlabel comment s 0 0 0 0 4 buf_16
flabel metal1 s 0 51 6720 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 6720 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 1790 458 6528 504 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel metal1 s 5049 11 5049 11 0 FreeSans 340 0 0 0 VNB
port 3 nsew
flabel metal1 s 0 689 6720 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 6720 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 5049 802 5049 802 0 FreeSans 340 0 0 0 VPB
port 4 nsew
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 6720 814
string GDS_END 1091352
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1031596
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
