magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 20955 0 21038 732
<< locali >>
rect -5487 429 -5449 463
rect -5571 291 -5537 329
rect -5385 291 -5351 329
<< viali >>
rect -5521 429 -5487 463
rect -5449 429 -5415 463
rect -5571 329 -5537 363
rect -5571 257 -5537 291
rect -5385 329 -5351 363
rect -5385 257 -5351 291
<< metal1 >>
rect -194 2003 147 2009
rect -142 1951 -130 2003
rect -78 1951 147 2003
rect -194 1935 147 1951
rect -142 1883 -130 1935
rect -78 1883 147 1935
rect -194 1866 147 1883
rect -142 1814 -130 1866
rect -78 1814 147 1866
rect 202 1826 501 2002
rect -194 1808 147 1814
rect 692 1808 808 2009
rect 3646 2003 3762 2009
rect 3698 1951 3710 2003
rect 3646 1935 3762 1951
rect 3698 1883 3710 1935
rect 3646 1866 3762 1883
rect 3698 1814 3710 1866
rect 3646 1808 3762 1814
rect 3948 2003 4064 2009
rect 4000 1951 4012 2003
rect 3948 1935 4064 1951
rect 4000 1883 4012 1935
rect 3948 1866 4064 1883
rect 4000 1814 4012 1866
rect 3948 1808 4064 1814
rect 8093 2003 8209 2009
rect 8145 1951 8157 2003
rect 8093 1935 8209 1951
rect 8145 1883 8157 1935
rect 8093 1866 8209 1883
rect 8145 1814 8157 1866
rect 8093 1808 8209 1814
rect 8984 2003 9100 2009
rect 9036 1951 9048 2003
rect 8984 1935 9100 1951
rect 9036 1883 9048 1935
rect 8984 1866 9100 1883
rect 9036 1814 9048 1866
rect 8984 1808 9100 1814
rect 11938 2003 12054 2009
rect 11990 1951 12002 2003
rect 11938 1935 12054 1951
rect 11990 1883 12002 1935
rect 11938 1866 12054 1883
rect 11990 1814 12002 1866
rect 11938 1808 12054 1814
rect 13130 2003 13246 2009
rect 13182 1951 13194 2003
rect 13130 1935 13246 1951
rect 13182 1883 13194 1935
rect 13130 1866 13246 1883
rect 13182 1814 13194 1866
rect 13130 1808 13246 1814
rect 14639 2003 14691 2009
rect 14639 1935 14691 1951
rect 14639 1866 14691 1883
rect 14639 1808 14691 1814
rect 16084 2003 16200 2009
rect 16136 1951 16148 2003
rect 16084 1935 16200 1951
rect 16136 1883 16148 1935
rect 16084 1866 16200 1883
rect 16136 1814 16148 1866
rect 16084 1808 16200 1814
rect 17276 2003 17392 2009
rect 17328 1951 17340 2003
rect 17276 1935 17392 1951
rect 17328 1883 17340 1935
rect 17276 1866 17392 1883
rect 17328 1814 17340 1866
rect 17276 1808 17392 1814
rect 18785 2003 18837 2009
rect 18785 1935 18837 1951
rect 18785 1866 18837 1883
rect 18785 1808 18837 1814
rect 20230 2003 20346 2009
rect 20282 1951 20294 2003
rect 20230 1935 20346 1951
rect 20282 1883 20294 1935
rect 20230 1866 20346 1883
rect 20282 1814 20294 1866
rect 20230 1808 20346 1814
rect 1339 1727 1345 1779
rect 1397 1727 1409 1779
rect 1461 1727 1921 1779
tri 1841 1693 1875 1727 ne
rect 1875 1632 1921 1727
rect 1876 1630 1920 1631
rect 2069 1765 2121 1771
rect 2069 1701 2121 1713
rect 2069 1632 2121 1649
rect 2070 1630 2120 1631
rect 2333 1765 2385 1771
rect 2333 1701 2385 1713
rect 2333 1632 2385 1649
rect 2334 1630 2384 1631
rect 2533 1727 2993 1779
rect 3045 1727 3057 1779
rect 3109 1727 3115 1779
rect 5485 1727 5491 1779
rect 5543 1727 5555 1779
rect 5607 1727 6067 1779
rect 2533 1632 2579 1727
tri 2579 1693 2613 1727 nw
tri 5987 1693 6021 1727 ne
rect 2534 1630 2578 1631
rect 1875 1594 1921 1630
rect 2533 1594 2579 1630
rect 1876 1593 1920 1594
rect 1875 1540 1921 1592
rect 2070 1593 2120 1594
rect 2069 1540 2121 1592
rect 2334 1593 2384 1594
rect 2333 1540 2385 1592
rect 2534 1593 2578 1594
rect 2533 1540 2579 1592
rect 6021 1632 6067 1727
rect 6022 1630 6066 1631
rect 6215 1765 6267 1771
rect 6215 1701 6267 1713
rect 6215 1632 6267 1649
rect 6216 1630 6266 1631
rect 6479 1765 6531 1771
rect 6479 1701 6531 1713
rect 6479 1632 6531 1649
rect 6480 1630 6530 1631
rect 6679 1727 7139 1779
rect 7191 1727 7203 1779
rect 7255 1727 7261 1779
rect 9631 1727 9637 1779
rect 9689 1727 9701 1779
rect 9753 1727 10213 1779
rect 6679 1632 6725 1727
tri 6725 1693 6759 1727 nw
tri 10133 1693 10167 1727 ne
rect 6680 1630 6724 1631
rect 6021 1594 6067 1630
rect 6679 1594 6725 1630
rect 6022 1593 6066 1594
rect 6021 1540 6067 1592
rect 6216 1593 6266 1594
rect 6215 1540 6267 1592
rect 6480 1593 6530 1594
rect 6479 1540 6531 1592
rect 6680 1593 6724 1594
rect 6679 1540 6725 1592
rect 10167 1632 10213 1727
rect 10168 1630 10212 1631
rect 10361 1765 10413 1771
rect 10361 1701 10413 1713
rect 10361 1632 10413 1649
rect 10362 1630 10412 1631
rect 10625 1765 10677 1771
rect 10625 1701 10677 1713
rect 10625 1632 10677 1649
rect 10626 1630 10676 1631
rect 10825 1727 11285 1779
rect 11337 1727 11349 1779
rect 11401 1727 11407 1779
rect 13777 1727 13783 1779
rect 13835 1727 13847 1779
rect 13899 1727 14359 1779
rect 10825 1632 10871 1727
tri 10871 1693 10905 1727 nw
tri 14264 1693 14298 1727 ne
rect 14298 1693 14359 1727
tri 14298 1684 14307 1693 ne
rect 10826 1630 10870 1631
rect 14307 1632 14359 1693
rect 14308 1630 14358 1631
rect 14507 1765 14559 1771
rect 14507 1701 14559 1713
rect 14507 1643 14559 1649
rect 14507 1632 14553 1643
tri 14553 1637 14559 1643 nw
rect 14771 1765 14823 1771
rect 14771 1701 14823 1713
rect 14508 1630 14552 1631
rect 14771 1632 14823 1649
rect 14772 1630 14822 1631
rect 14971 1727 15431 1779
rect 15483 1727 15495 1779
rect 15547 1727 15553 1779
rect 17923 1727 17929 1779
rect 17981 1727 17993 1779
rect 18045 1727 18505 1779
rect 14971 1632 15017 1727
tri 15017 1693 15051 1727 nw
tri 18425 1693 18459 1727 ne
rect 14972 1630 15016 1631
rect 10167 1594 10213 1630
rect 10825 1594 10871 1630
rect 14507 1594 14553 1630
rect 14971 1594 15017 1630
rect 10168 1593 10212 1594
rect 10167 1540 10213 1592
rect 10362 1593 10412 1594
rect 10361 1540 10413 1592
rect 10626 1593 10676 1594
rect 10625 1540 10677 1592
rect 10826 1593 10870 1594
rect 10825 1540 10871 1592
rect 14308 1593 14358 1594
rect 14307 1540 14359 1592
rect 14508 1593 14552 1594
rect 14507 1540 14553 1592
rect 14772 1593 14822 1594
tri 14553 1540 14559 1546 sw
rect 14771 1540 14823 1592
rect 14972 1593 15016 1594
rect 14971 1540 15017 1592
rect 18459 1632 18505 1727
rect 18460 1630 18504 1631
rect 18653 1765 18705 1771
rect 18653 1701 18705 1713
rect 18653 1632 18705 1649
rect 18654 1630 18704 1631
rect 18917 1765 18969 1771
rect 18917 1701 18969 1713
rect 18917 1632 18969 1649
rect 18918 1630 18968 1631
rect 19117 1727 19577 1779
rect 19629 1727 19641 1779
rect 19693 1727 19699 1779
rect 19117 1632 19163 1727
tri 19163 1693 19197 1727 nw
rect 19118 1630 19162 1631
rect 18459 1594 18505 1630
rect 19117 1594 19163 1630
rect 18460 1593 18504 1594
rect 18459 1540 18505 1592
rect 18654 1593 18704 1594
rect 18653 1540 18705 1592
rect 18918 1593 18968 1594
rect 18917 1540 18969 1592
rect 19118 1593 19162 1594
rect 19117 1540 19163 1592
tri 14307 1534 14313 1540 ne
rect 1875 1396 1921 1448
rect 1876 1394 1920 1395
rect 2069 1396 2121 1448
rect 2070 1394 2120 1395
rect 2069 1358 2121 1394
rect 1876 1357 1920 1358
tri 1841 1311 1875 1345 se
rect 1875 1304 1921 1356
rect 2070 1357 2120 1358
tri 1921 1311 1955 1345 sw
tri 2035 1311 2069 1345 se
rect 2069 1304 2121 1356
rect 2333 1396 2385 1448
rect 2334 1394 2384 1395
rect 2533 1396 2579 1448
rect 2534 1394 2578 1395
rect 6021 1396 6067 1448
rect 6022 1394 6066 1395
rect 6215 1396 6267 1448
rect 6216 1394 6266 1395
rect 2333 1358 2385 1394
rect 6215 1358 6267 1394
rect 2334 1357 2384 1358
tri 2327 1339 2333 1345 se
rect 2333 1339 2385 1356
rect 2534 1357 2578 1358
tri 2121 1311 2149 1339 sw
tri 2299 1311 2327 1339 se
rect 2327 1311 2385 1339
tri 2385 1311 2419 1345 sw
tri 2499 1311 2533 1345 se
rect 2333 1304 2385 1311
rect 2533 1304 2579 1356
rect 6022 1357 6066 1358
tri 2579 1311 2613 1345 sw
tri 5987 1311 6021 1345 se
rect 6021 1304 6067 1356
rect 6216 1357 6266 1358
tri 6067 1311 6101 1345 sw
tri 6181 1311 6215 1345 se
rect 6215 1304 6267 1356
rect 6479 1396 6531 1448
rect 6480 1394 6530 1395
rect 6679 1396 6725 1448
rect 6680 1394 6724 1395
rect 10167 1396 10213 1448
rect 10168 1394 10212 1395
rect 10361 1396 10413 1448
rect 10362 1394 10412 1395
rect 6479 1358 6531 1394
rect 10361 1358 10413 1394
rect 6480 1357 6530 1358
tri 6267 1311 6295 1339 sw
tri 6451 1311 6479 1339 se
rect 6479 1304 6531 1356
rect 6680 1357 6724 1358
tri 6531 1311 6565 1345 sw
tri 6645 1311 6679 1345 se
rect 6679 1304 6725 1356
rect 10168 1357 10212 1358
tri 6725 1311 6759 1345 sw
tri 10133 1311 10167 1345 se
rect 10167 1304 10213 1356
rect 10362 1357 10412 1358
tri 10213 1311 10247 1345 sw
tri 10327 1311 10361 1345 se
rect 10361 1304 10413 1356
rect 10625 1396 10677 1448
rect 10626 1394 10676 1395
rect 10825 1396 10871 1448
rect 10826 1394 10870 1395
rect 10625 1358 10677 1394
rect 10626 1357 10676 1358
tri 10413 1311 10441 1339 sw
tri 10597 1311 10625 1339 se
rect 10625 1304 10677 1356
rect 10826 1357 10870 1358
tri 10677 1311 10711 1345 sw
tri 10791 1311 10825 1345 se
rect 10825 1304 10871 1356
tri 10871 1311 10905 1345 sw
rect 14771 1298 14823 1304
rect 208 1127 499 1290
rect 14771 1234 14823 1246
rect 14771 1170 14823 1182
rect 14771 1112 14823 1118
rect 14965 1298 15017 1304
rect 14965 1234 15017 1246
rect 14965 1170 15017 1182
rect 14965 1112 15017 1118
rect 18459 1298 18511 1304
rect 18459 1234 18511 1246
rect 18459 1170 18511 1182
rect 18459 1112 18511 1118
rect 18653 1298 18705 1304
rect 18653 1234 18705 1246
rect 18653 1170 18705 1182
rect 18653 1112 18705 1118
rect 1526 722 1578 734
rect 583 670 635 676
tri 549 596 583 630 ne
rect 583 606 635 618
rect 2876 722 2928 734
rect 1526 658 1578 670
rect 2118 709 2170 715
tri 2084 629 2118 663 ne
rect 2118 645 2170 657
rect 1526 600 1578 606
rect 2118 587 2170 593
rect 2284 709 2336 715
rect 5672 722 5724 734
rect 2284 645 2336 657
tri 2336 629 2370 663 nw
rect 2876 658 2928 670
rect 2876 600 2928 606
rect 3819 670 3871 676
rect 4729 670 4781 676
rect 3819 606 3871 618
rect 2284 587 2336 593
rect 583 548 635 554
tri 3871 596 3905 630 nw
tri 4695 596 4729 630 ne
rect 4729 606 4781 618
rect 3819 548 3871 554
rect 7022 722 7074 734
rect 5672 658 5724 670
rect 6264 709 6316 715
tri 6230 629 6264 663 ne
rect 6264 645 6316 657
rect 5672 600 5724 606
rect 6264 587 6316 593
rect 6430 709 6482 715
rect 9818 722 9870 734
rect 6430 645 6482 657
tri 6482 629 6516 663 nw
rect 7022 658 7074 670
rect 7022 600 7074 606
rect 7965 670 8017 676
rect 8875 670 8927 676
rect 7965 606 8017 618
rect 6430 587 6482 593
rect 4729 548 4781 554
tri 8017 596 8051 630 nw
tri 8841 596 8875 630 ne
rect 8875 606 8927 618
rect 7965 548 8017 554
rect 11168 722 11220 734
rect 9818 658 9870 670
rect 10410 709 10462 715
tri 10376 629 10410 663 ne
rect 10410 645 10462 657
rect 9818 600 9870 606
rect 10410 587 10462 593
rect 10576 709 10628 715
rect 13964 722 14016 734
rect 10576 645 10628 657
tri 10628 629 10662 663 nw
rect 11168 658 11220 670
rect 11168 600 11220 606
rect 12111 670 12163 676
rect 13021 670 13073 676
rect 12111 606 12163 618
rect 10576 587 10628 593
rect 8875 548 8927 554
tri 12163 596 12197 630 nw
tri 12987 596 13021 630 ne
rect 13021 606 13073 618
rect 12111 548 12163 554
rect 15314 722 15366 734
rect 13964 658 14016 670
rect 14556 709 14608 715
tri 14522 629 14556 663 ne
rect 14556 645 14608 657
rect 13964 600 14016 606
rect 14556 587 14608 593
rect 14722 709 14774 715
rect 18110 722 18162 734
rect 14722 645 14774 657
tri 14774 629 14808 663 nw
rect 15314 658 15366 670
rect 15314 600 15366 606
rect 16257 670 16309 676
rect 17167 670 17219 676
rect 16257 606 16309 618
rect 14722 587 14774 593
rect 13021 548 13073 554
tri 16309 596 16343 630 nw
tri 17133 596 17167 630 ne
rect 17167 606 17219 618
rect 16257 548 16309 554
rect 19460 722 19512 734
rect 18110 658 18162 670
rect 18702 709 18754 715
tri 18668 629 18702 663 ne
rect 18702 645 18754 657
rect 18110 600 18162 606
rect 18702 587 18754 593
rect 18868 709 18920 715
rect 18868 645 18920 657
tri 18920 629 18954 663 nw
rect 19460 658 19512 670
rect 19460 600 19512 606
rect 20403 670 20455 676
rect 20403 606 20455 618
rect 18868 587 18920 593
rect 17167 548 17219 554
tri 20455 596 20489 630 nw
rect 20403 548 20455 554
rect -5619 526 -5567 532
tri 1812 504 1816 508 se
tri 2041 504 2045 508 sw
tri 2409 504 2413 508 se
tri 2638 504 2642 508 sw
tri 5958 504 5962 508 se
tri 6187 504 6191 508 sw
tri 6555 504 6559 508 se
tri 6784 504 6788 508 sw
tri 10104 504 10108 508 se
tri 10333 504 10337 508 sw
tri 10701 504 10705 508 se
tri 10930 504 10934 508 sw
tri 14250 504 14254 508 se
tri 14479 504 14483 508 sw
tri 14847 504 14851 508 se
tri 15076 504 15080 508 sw
tri 18396 504 18400 508 se
tri 18625 504 18629 508 sw
tri 18993 504 18997 508 se
tri 19222 504 19226 508 sw
tri 1782 474 1812 504 se
rect 1812 474 2045 504
tri 2045 474 2075 504 sw
tri 2379 474 2409 504 se
rect 2409 474 2642 504
tri 2642 474 2672 504 sw
tri 5928 474 5958 504 se
rect 5958 474 6191 504
tri 6191 474 6221 504 sw
tri 6525 474 6555 504 se
rect 6555 474 6788 504
tri 6788 474 6818 504 sw
tri 10074 474 10104 504 se
rect 10104 474 10337 504
tri 10337 474 10367 504 sw
tri 10671 474 10701 504 se
rect 10701 474 10934 504
tri 10934 474 10964 504 sw
tri 14220 474 14250 504 se
rect 14250 474 14483 504
tri 14483 474 14513 504 sw
tri 14817 474 14847 504 se
rect 14847 474 15080 504
tri 15080 474 15110 504 sw
tri 18366 474 18396 504 se
rect 18396 474 18629 504
tri 18629 474 18659 504 sw
tri 18963 474 18993 504 se
rect 18993 474 19226 504
tri 19226 474 19256 504 sw
rect -5619 469 -5567 474
rect -5619 463 -5403 469
rect -5619 462 -5521 463
rect -5567 429 -5521 462
rect -5487 429 -5449 463
rect -5415 429 -5403 463
rect -5567 423 -5403 429
rect -194 468 154 474
rect -5619 404 -5567 410
rect -142 416 -130 468
rect -78 416 154 468
rect -194 402 154 416
rect -5577 363 -5345 375
rect -5577 329 -5571 363
rect -5537 329 -5385 363
rect -5351 329 -5345 363
rect -142 350 -130 402
rect -78 350 154 402
rect -194 344 154 350
rect 692 344 808 474
rect 3646 468 3762 474
rect 3698 416 3710 468
rect 3646 402 3762 416
rect 3698 350 3710 402
rect 3646 344 3762 350
rect 3948 468 4064 474
rect 4000 416 4012 468
rect 3948 402 4064 416
rect 4000 350 4012 402
rect 3948 344 4064 350
rect 8093 468 8209 474
rect 8145 416 8157 468
rect 8093 402 8209 416
rect 8145 350 8157 402
rect 8093 344 8209 350
rect 8984 468 9100 474
rect 9036 416 9048 468
rect 8984 402 9100 416
rect 9036 350 9048 402
rect 8984 344 9100 350
rect 11938 468 12054 474
rect 11990 416 12002 468
rect 11938 402 12054 416
rect 11990 350 12002 402
rect 11938 344 12054 350
rect 13130 468 13246 474
rect 13182 416 13194 468
rect 13130 402 13246 416
rect 13182 350 13194 402
rect 13130 344 13246 350
rect 14639 468 14691 474
rect 14639 402 14691 416
rect 14639 344 14691 350
rect 16084 468 16200 474
rect 16136 416 16148 468
rect 16084 402 16200 416
rect 16136 350 16148 402
rect 16084 344 16200 350
rect 17276 468 17392 474
rect 17328 416 17340 468
rect 17276 402 17392 416
rect 17328 350 17340 402
rect 17276 344 17392 350
rect 18785 468 18837 474
rect 18785 402 18837 416
rect 18785 344 18837 350
rect 20230 468 20346 474
rect 20282 416 20294 468
rect 20230 402 20346 416
rect 20282 350 20294 402
rect 20230 344 20346 350
rect -5577 291 -5345 329
rect -5577 257 -5571 291
rect -5537 257 -5385 291
rect -5351 257 -5345 291
rect -5577 245 -5345 257
rect 212 132 569 298
rect 13509 -47 13515 5
rect 13567 -47 13579 5
rect 13631 -47 14853 5
rect 14905 -47 14917 5
rect 14969 -47 15507 5
rect 15559 -47 15571 5
rect 15623 -47 17853 5
rect 17905 -47 17917 5
rect 17969 -47 18486 5
rect 18538 -47 18550 5
rect 18602 -47 18608 5
rect 0 -127 1532 -75
rect 1584 -127 1596 -75
rect 1648 -127 2806 -75
rect 2858 -127 2870 -75
rect 2922 -127 5678 -75
rect 5730 -127 5742 -75
rect 5794 -127 6952 -75
rect 7004 -127 7016 -75
rect 7068 -127 9824 -75
rect 9876 -127 9888 -75
rect 9940 -127 11098 -75
rect 11150 -127 11162 -75
rect 11214 -127 13970 -75
rect 14022 -127 14034 -75
rect 14086 -127 15244 -75
rect 15296 -127 15308 -75
rect 15360 -127 18257 -75
rect 18309 -127 18321 -75
rect 18373 -127 19390 -75
rect 19442 -127 19454 -75
rect 19506 -127 20871 -75
tri -1955 -168 -1942 -155 se
rect -1942 -168 1269 -155
rect -6326 -220 -5689 -168
rect -5637 -220 -5625 -168
rect -5573 -207 1269 -168
rect 1321 -207 1333 -155
rect 1385 -207 1923 -155
rect 1975 -207 1987 -155
rect 2039 -207 2415 -155
rect 2467 -207 2479 -155
rect 2531 -207 3069 -155
rect 3121 -207 3133 -155
rect 3185 -207 5415 -155
rect 5467 -207 5479 -155
rect 5531 -207 6069 -155
rect 6121 -207 6133 -155
rect 6185 -207 6561 -155
rect 6613 -207 6625 -155
rect 6677 -207 7215 -155
rect 7267 -207 7279 -155
rect 7331 -207 9561 -155
rect 9613 -207 9625 -155
rect 9677 -207 10215 -155
rect 10267 -207 10279 -155
rect 10331 -207 10707 -155
rect 10759 -207 10771 -155
rect 10823 -207 11361 -155
rect 11413 -207 11425 -155
rect 11477 -207 13515 -155
rect 13567 -207 13579 -155
rect 13631 -207 13637 -155
rect 13701 -207 13707 -155
rect 13759 -207 13771 -155
rect 13823 -207 14361 -155
rect 14413 -207 14425 -155
rect 14477 -207 18507 -155
rect 18559 -207 18571 -155
rect 18623 -207 18999 -155
rect 19051 -207 19063 -155
rect 19115 -207 19653 -155
rect 19705 -207 19717 -155
rect 19769 -207 20871 -155
rect -5573 -220 -1933 -207
tri -1933 -220 -1920 -207 nw
rect 14245 -479 14251 -427
rect 14303 -479 14315 -427
rect 14367 -479 14373 -427
rect 14465 -479 14471 -427
rect 14523 -479 14535 -427
rect 14587 -479 14593 -427
<< rmetal1 >>
rect 1875 1631 1921 1632
rect 1875 1630 1876 1631
rect 1920 1630 1921 1631
rect 2069 1631 2121 1632
rect 2069 1630 2070 1631
rect 2120 1630 2121 1631
rect 2333 1631 2385 1632
rect 2333 1630 2334 1631
rect 2384 1630 2385 1631
rect 2533 1631 2579 1632
rect 2533 1630 2534 1631
rect 2578 1630 2579 1631
rect 1875 1593 1876 1594
rect 1920 1593 1921 1594
rect 1875 1592 1921 1593
rect 2069 1593 2070 1594
rect 2120 1593 2121 1594
rect 2069 1592 2121 1593
rect 2333 1593 2334 1594
rect 2384 1593 2385 1594
rect 2333 1592 2385 1593
rect 2533 1593 2534 1594
rect 2578 1593 2579 1594
rect 2533 1592 2579 1593
rect 6021 1631 6067 1632
rect 6021 1630 6022 1631
rect 6066 1630 6067 1631
rect 6215 1631 6267 1632
rect 6215 1630 6216 1631
rect 6266 1630 6267 1631
rect 6479 1631 6531 1632
rect 6479 1630 6480 1631
rect 6530 1630 6531 1631
rect 6679 1631 6725 1632
rect 6679 1630 6680 1631
rect 6724 1630 6725 1631
rect 6021 1593 6022 1594
rect 6066 1593 6067 1594
rect 6021 1592 6067 1593
rect 6215 1593 6216 1594
rect 6266 1593 6267 1594
rect 6215 1592 6267 1593
rect 6479 1593 6480 1594
rect 6530 1593 6531 1594
rect 6479 1592 6531 1593
rect 6679 1593 6680 1594
rect 6724 1593 6725 1594
rect 6679 1592 6725 1593
rect 10167 1631 10213 1632
rect 10167 1630 10168 1631
rect 10212 1630 10213 1631
rect 10361 1631 10413 1632
rect 10361 1630 10362 1631
rect 10412 1630 10413 1631
rect 10625 1631 10677 1632
rect 10625 1630 10626 1631
rect 10676 1630 10677 1631
rect 10825 1631 10871 1632
rect 10825 1630 10826 1631
rect 10870 1630 10871 1631
rect 14307 1631 14359 1632
rect 14307 1630 14308 1631
rect 14358 1630 14359 1631
rect 14507 1631 14553 1632
rect 14507 1630 14508 1631
rect 14552 1630 14553 1631
rect 14771 1631 14823 1632
rect 14771 1630 14772 1631
rect 14822 1630 14823 1631
rect 14971 1631 15017 1632
rect 14971 1630 14972 1631
rect 15016 1630 15017 1631
rect 10167 1593 10168 1594
rect 10212 1593 10213 1594
rect 10167 1592 10213 1593
rect 10361 1593 10362 1594
rect 10412 1593 10413 1594
rect 10361 1592 10413 1593
rect 10625 1593 10626 1594
rect 10676 1593 10677 1594
rect 10625 1592 10677 1593
rect 10825 1593 10826 1594
rect 10870 1593 10871 1594
rect 10825 1592 10871 1593
rect 14307 1593 14308 1594
rect 14358 1593 14359 1594
rect 14307 1592 14359 1593
rect 14507 1593 14508 1594
rect 14552 1593 14553 1594
rect 14507 1592 14553 1593
rect 14771 1593 14772 1594
rect 14822 1593 14823 1594
rect 14771 1592 14823 1593
rect 14971 1593 14972 1594
rect 15016 1593 15017 1594
rect 14971 1592 15017 1593
rect 18459 1631 18505 1632
rect 18459 1630 18460 1631
rect 18504 1630 18505 1631
rect 18653 1631 18705 1632
rect 18653 1630 18654 1631
rect 18704 1630 18705 1631
rect 18917 1631 18969 1632
rect 18917 1630 18918 1631
rect 18968 1630 18969 1631
rect 19117 1631 19163 1632
rect 19117 1630 19118 1631
rect 19162 1630 19163 1631
rect 18459 1593 18460 1594
rect 18504 1593 18505 1594
rect 18459 1592 18505 1593
rect 18653 1593 18654 1594
rect 18704 1593 18705 1594
rect 18653 1592 18705 1593
rect 18917 1593 18918 1594
rect 18968 1593 18969 1594
rect 18917 1592 18969 1593
rect 19117 1593 19118 1594
rect 19162 1593 19163 1594
rect 19117 1592 19163 1593
rect 1875 1395 1921 1396
rect 1875 1394 1876 1395
rect 1920 1394 1921 1395
rect 2069 1395 2121 1396
rect 2069 1394 2070 1395
rect 2120 1394 2121 1395
rect 1875 1357 1876 1358
rect 1920 1357 1921 1358
rect 1875 1356 1921 1357
rect 2069 1357 2070 1358
rect 2120 1357 2121 1358
rect 2069 1356 2121 1357
rect 2333 1395 2385 1396
rect 2333 1394 2334 1395
rect 2384 1394 2385 1395
rect 2533 1395 2579 1396
rect 2533 1394 2534 1395
rect 2578 1394 2579 1395
rect 6021 1395 6067 1396
rect 6021 1394 6022 1395
rect 6066 1394 6067 1395
rect 6215 1395 6267 1396
rect 6215 1394 6216 1395
rect 6266 1394 6267 1395
rect 2333 1357 2334 1358
rect 2384 1357 2385 1358
rect 2333 1356 2385 1357
rect 2533 1357 2534 1358
rect 2578 1357 2579 1358
rect 2533 1356 2579 1357
rect 6021 1357 6022 1358
rect 6066 1357 6067 1358
rect 6021 1356 6067 1357
rect 6215 1357 6216 1358
rect 6266 1357 6267 1358
rect 6215 1356 6267 1357
rect 6479 1395 6531 1396
rect 6479 1394 6480 1395
rect 6530 1394 6531 1395
rect 6679 1395 6725 1396
rect 6679 1394 6680 1395
rect 6724 1394 6725 1395
rect 10167 1395 10213 1396
rect 10167 1394 10168 1395
rect 10212 1394 10213 1395
rect 10361 1395 10413 1396
rect 10361 1394 10362 1395
rect 10412 1394 10413 1395
rect 6479 1357 6480 1358
rect 6530 1357 6531 1358
rect 6479 1356 6531 1357
rect 6679 1357 6680 1358
rect 6724 1357 6725 1358
rect 6679 1356 6725 1357
rect 10167 1357 10168 1358
rect 10212 1357 10213 1358
rect 10167 1356 10213 1357
rect 10361 1357 10362 1358
rect 10412 1357 10413 1358
rect 10361 1356 10413 1357
rect 10625 1395 10677 1396
rect 10625 1394 10626 1395
rect 10676 1394 10677 1395
rect 10825 1395 10871 1396
rect 10825 1394 10826 1395
rect 10870 1394 10871 1395
rect 10625 1357 10626 1358
rect 10676 1357 10677 1358
rect 10625 1356 10677 1357
rect 10825 1357 10826 1358
rect 10870 1357 10871 1358
rect 10825 1356 10871 1357
<< via1 >>
rect -194 1951 -142 2003
rect -130 1951 -78 2003
rect -194 1883 -142 1935
rect -130 1883 -78 1935
rect -194 1814 -142 1866
rect -130 1814 -78 1866
rect 3646 1951 3698 2003
rect 3710 1951 3762 2003
rect 3646 1883 3698 1935
rect 3710 1883 3762 1935
rect 3646 1814 3698 1866
rect 3710 1814 3762 1866
rect 3948 1951 4000 2003
rect 4012 1951 4064 2003
rect 3948 1883 4000 1935
rect 4012 1883 4064 1935
rect 3948 1814 4000 1866
rect 4012 1814 4064 1866
rect 8093 1951 8145 2003
rect 8157 1951 8209 2003
rect 8093 1883 8145 1935
rect 8157 1883 8209 1935
rect 8093 1814 8145 1866
rect 8157 1814 8209 1866
rect 8984 1951 9036 2003
rect 9048 1951 9100 2003
rect 8984 1883 9036 1935
rect 9048 1883 9100 1935
rect 8984 1814 9036 1866
rect 9048 1814 9100 1866
rect 11938 1951 11990 2003
rect 12002 1951 12054 2003
rect 11938 1883 11990 1935
rect 12002 1883 12054 1935
rect 11938 1814 11990 1866
rect 12002 1814 12054 1866
rect 13130 1951 13182 2003
rect 13194 1951 13246 2003
rect 13130 1883 13182 1935
rect 13194 1883 13246 1935
rect 13130 1814 13182 1866
rect 13194 1814 13246 1866
rect 14639 1951 14691 2003
rect 14639 1883 14691 1935
rect 14639 1814 14691 1866
rect 16084 1951 16136 2003
rect 16148 1951 16200 2003
rect 16084 1883 16136 1935
rect 16148 1883 16200 1935
rect 16084 1814 16136 1866
rect 16148 1814 16200 1866
rect 17276 1951 17328 2003
rect 17340 1951 17392 2003
rect 17276 1883 17328 1935
rect 17340 1883 17392 1935
rect 17276 1814 17328 1866
rect 17340 1814 17392 1866
rect 18785 1951 18837 2003
rect 18785 1883 18837 1935
rect 18785 1814 18837 1866
rect 20230 1951 20282 2003
rect 20294 1951 20346 2003
rect 20230 1883 20282 1935
rect 20294 1883 20346 1935
rect 20230 1814 20282 1866
rect 20294 1814 20346 1866
rect 1345 1727 1397 1779
rect 1409 1727 1461 1779
rect 2069 1713 2121 1765
rect 2069 1649 2121 1701
rect 2333 1713 2385 1765
rect 2333 1649 2385 1701
rect 2993 1727 3045 1779
rect 3057 1727 3109 1779
rect 5491 1727 5543 1779
rect 5555 1727 5607 1779
rect 6215 1713 6267 1765
rect 6215 1649 6267 1701
rect 6479 1713 6531 1765
rect 6479 1649 6531 1701
rect 7139 1727 7191 1779
rect 7203 1727 7255 1779
rect 9637 1727 9689 1779
rect 9701 1727 9753 1779
rect 10361 1713 10413 1765
rect 10361 1649 10413 1701
rect 10625 1713 10677 1765
rect 10625 1649 10677 1701
rect 11285 1727 11337 1779
rect 11349 1727 11401 1779
rect 13783 1727 13835 1779
rect 13847 1727 13899 1779
rect 14507 1713 14559 1765
rect 14507 1649 14559 1701
rect 14771 1713 14823 1765
rect 14771 1649 14823 1701
rect 15431 1727 15483 1779
rect 15495 1727 15547 1779
rect 17929 1727 17981 1779
rect 17993 1727 18045 1779
rect 18653 1713 18705 1765
rect 18653 1649 18705 1701
rect 18917 1713 18969 1765
rect 18917 1649 18969 1701
rect 19577 1727 19629 1779
rect 19641 1727 19693 1779
rect 14771 1246 14823 1298
rect 14771 1182 14823 1234
rect 14771 1118 14823 1170
rect 14965 1246 15017 1298
rect 14965 1182 15017 1234
rect 14965 1118 15017 1170
rect 18459 1246 18511 1298
rect 18459 1182 18511 1234
rect 18459 1118 18511 1170
rect 18653 1246 18705 1298
rect 18653 1182 18705 1234
rect 18653 1118 18705 1170
rect 583 618 635 670
rect 583 554 635 606
rect 1526 670 1578 722
rect 1526 606 1578 658
rect 2118 657 2170 709
rect 2118 593 2170 645
rect 2284 657 2336 709
rect 2876 670 2928 722
rect 2284 593 2336 645
rect 2876 606 2928 658
rect 3819 618 3871 670
rect 3819 554 3871 606
rect 4729 618 4781 670
rect 4729 554 4781 606
rect 5672 670 5724 722
rect 5672 606 5724 658
rect 6264 657 6316 709
rect 6264 593 6316 645
rect 6430 657 6482 709
rect 7022 670 7074 722
rect 6430 593 6482 645
rect 7022 606 7074 658
rect 7965 618 8017 670
rect 7965 554 8017 606
rect 8875 618 8927 670
rect 8875 554 8927 606
rect 9818 670 9870 722
rect 9818 606 9870 658
rect 10410 657 10462 709
rect 10410 593 10462 645
rect 10576 657 10628 709
rect 11168 670 11220 722
rect 10576 593 10628 645
rect 11168 606 11220 658
rect 12111 618 12163 670
rect 12111 554 12163 606
rect 13021 618 13073 670
rect 13021 554 13073 606
rect 13964 670 14016 722
rect 13964 606 14016 658
rect 14556 657 14608 709
rect 14556 593 14608 645
rect 14722 657 14774 709
rect 15314 670 15366 722
rect 14722 593 14774 645
rect 15314 606 15366 658
rect 16257 618 16309 670
rect 16257 554 16309 606
rect 17167 618 17219 670
rect 17167 554 17219 606
rect 18110 670 18162 722
rect 18110 606 18162 658
rect 18702 657 18754 709
rect 18702 593 18754 645
rect 18868 657 18920 709
rect 19460 670 19512 722
rect 18868 593 18920 645
rect 19460 606 19512 658
rect 20403 618 20455 670
rect 20403 554 20455 606
rect -5619 474 -5567 526
rect -5619 410 -5567 462
rect -194 416 -142 468
rect -130 416 -78 468
rect -194 350 -142 402
rect -130 350 -78 402
rect 3646 416 3698 468
rect 3710 416 3762 468
rect 3646 350 3698 402
rect 3710 350 3762 402
rect 3948 416 4000 468
rect 4012 416 4064 468
rect 3948 350 4000 402
rect 4012 350 4064 402
rect 8093 416 8145 468
rect 8157 416 8209 468
rect 8093 350 8145 402
rect 8157 350 8209 402
rect 8984 416 9036 468
rect 9048 416 9100 468
rect 8984 350 9036 402
rect 9048 350 9100 402
rect 11938 416 11990 468
rect 12002 416 12054 468
rect 11938 350 11990 402
rect 12002 350 12054 402
rect 13130 416 13182 468
rect 13194 416 13246 468
rect 13130 350 13182 402
rect 13194 350 13246 402
rect 14639 416 14691 468
rect 14639 350 14691 402
rect 16084 416 16136 468
rect 16148 416 16200 468
rect 16084 350 16136 402
rect 16148 350 16200 402
rect 17276 416 17328 468
rect 17340 416 17392 468
rect 17276 350 17328 402
rect 17340 350 17392 402
rect 18785 416 18837 468
rect 18785 350 18837 402
rect 20230 416 20282 468
rect 20294 416 20346 468
rect 20230 350 20282 402
rect 20294 350 20346 402
rect 13515 -47 13567 5
rect 13579 -47 13631 5
rect 14853 -47 14905 5
rect 14917 -47 14969 5
rect 15507 -47 15559 5
rect 15571 -47 15623 5
rect 17853 -47 17905 5
rect 17917 -47 17969 5
rect 18486 -47 18538 5
rect 18550 -47 18602 5
rect 1532 -127 1584 -75
rect 1596 -127 1648 -75
rect 2806 -127 2858 -75
rect 2870 -127 2922 -75
rect 5678 -127 5730 -75
rect 5742 -127 5794 -75
rect 6952 -127 7004 -75
rect 7016 -127 7068 -75
rect 9824 -127 9876 -75
rect 9888 -127 9940 -75
rect 11098 -127 11150 -75
rect 11162 -127 11214 -75
rect 13970 -127 14022 -75
rect 14034 -127 14086 -75
rect 15244 -127 15296 -75
rect 15308 -127 15360 -75
rect 18257 -127 18309 -75
rect 18321 -127 18373 -75
rect 19390 -127 19442 -75
rect 19454 -127 19506 -75
rect -5689 -220 -5637 -168
rect -5625 -220 -5573 -168
rect 1269 -207 1321 -155
rect 1333 -207 1385 -155
rect 1923 -207 1975 -155
rect 1987 -207 2039 -155
rect 2415 -207 2467 -155
rect 2479 -207 2531 -155
rect 3069 -207 3121 -155
rect 3133 -207 3185 -155
rect 5415 -207 5467 -155
rect 5479 -207 5531 -155
rect 6069 -207 6121 -155
rect 6133 -207 6185 -155
rect 6561 -207 6613 -155
rect 6625 -207 6677 -155
rect 7215 -207 7267 -155
rect 7279 -207 7331 -155
rect 9561 -207 9613 -155
rect 9625 -207 9677 -155
rect 10215 -207 10267 -155
rect 10279 -207 10331 -155
rect 10707 -207 10759 -155
rect 10771 -207 10823 -155
rect 11361 -207 11413 -155
rect 11425 -207 11477 -155
rect 13515 -207 13567 -155
rect 13579 -207 13631 -155
rect 13707 -207 13759 -155
rect 13771 -207 13823 -155
rect 14361 -207 14413 -155
rect 14425 -207 14477 -155
rect 18507 -207 18559 -155
rect 18571 -207 18623 -155
rect 18999 -207 19051 -155
rect 19063 -207 19115 -155
rect 19653 -207 19705 -155
rect 19717 -207 19769 -155
rect 14251 -479 14303 -427
rect 14315 -479 14367 -427
rect 14471 -479 14523 -427
rect 14535 -479 14587 -427
<< metal2 >>
rect -194 2003 -78 2009
rect -142 1951 -130 2003
rect -194 1935 -78 1951
rect -142 1883 -130 1935
rect -194 1866 -78 1883
rect -142 1814 -130 1866
rect -5619 526 -5567 532
rect -5619 462 -5567 474
rect -5619 -168 -5567 410
rect -194 468 -78 1814
rect 3646 2003 3762 2009
rect 3698 1951 3710 2003
rect 3646 1935 3762 1951
rect 3698 1883 3710 1935
rect 3646 1866 3762 1883
rect 3698 1814 3710 1866
rect 1339 1727 1345 1779
rect 1397 1727 1409 1779
rect 1461 1727 1467 1779
rect 1993 1765 2121 1771
rect 1339 1713 1411 1727
tri 1411 1713 1425 1727 nw
rect 1993 1713 2069 1765
rect 1339 1701 1399 1713
tri 1399 1701 1411 1713 nw
rect 1993 1701 2121 1713
rect -142 416 -130 468
rect -194 402 -78 416
rect -142 350 -130 402
rect -194 344 -78 350
rect 583 670 635 676
rect 583 606 635 618
rect 583 0 635 554
rect 879 0 931 547
tri 1333 -127 1339 -121 se
rect 1339 -127 1391 1701
tri 1391 1693 1399 1701 nw
rect 1993 1649 2069 1701
rect 1993 1643 2121 1649
rect 2333 1765 2461 1771
rect 2385 1713 2461 1765
rect 2987 1727 2993 1779
rect 3045 1727 3057 1779
rect 3109 1727 3115 1779
tri 3029 1713 3043 1727 ne
rect 3043 1713 3115 1727
rect 2333 1701 2461 1713
tri 3043 1701 3055 1713 ne
rect 3055 1701 3115 1713
rect 2385 1649 2461 1701
tri 3055 1693 3063 1701 ne
rect 2333 1643 2461 1649
rect 1526 722 1578 728
rect 1526 658 1578 670
rect 1526 -47 1578 606
tri 1578 -47 1584 -41 sw
rect 1526 -75 1584 -47
tri 1584 -75 1612 -47 sw
rect 1526 -127 1532 -75
rect 1584 -127 1596 -75
rect 1648 -127 1654 -75
tri 1987 -127 1993 -121 se
rect 1993 -127 2045 1643
tri 2045 1609 2079 1643 nw
tri 2375 1609 2409 1643 ne
rect 2118 709 2170 715
rect 2118 645 2170 657
rect 2118 0 2170 593
rect 2284 709 2336 715
rect 2284 645 2336 657
rect 2284 0 2336 593
tri 1305 -155 1333 -127 se
rect 1333 -155 1391 -127
tri 1959 -155 1987 -127 se
rect 1987 -155 2045 -127
rect -5695 -220 -5689 -168
rect -5637 -220 -5625 -168
rect -5573 -220 -5567 -168
rect 1263 -207 1269 -155
rect 1321 -207 1333 -155
rect 1385 -207 1391 -155
rect 1917 -207 1923 -155
rect 1975 -207 1987 -155
rect 2039 -207 2045 -155
rect 2409 -127 2461 1643
rect 2876 722 2928 728
rect 2876 658 2928 670
tri 2870 -47 2876 -41 se
rect 2876 -47 2928 606
tri 2842 -75 2870 -47 se
rect 2870 -75 2928 -47
tri 2461 -127 2467 -121 sw
rect 2800 -127 2806 -75
rect 2858 -127 2870 -75
rect 2922 -127 2928 -75
rect 3063 -127 3115 1701
rect 3523 0 3575 547
rect 3646 468 3762 1814
rect 3948 2003 4064 2009
rect 4000 1951 4012 2003
rect 3948 1935 4064 1951
rect 4000 1883 4012 1935
rect 3948 1866 4064 1883
rect 4000 1814 4012 1866
rect 3698 416 3710 468
rect 3646 402 3762 416
rect 3698 350 3710 402
rect 3646 344 3762 350
rect 3819 670 3871 676
rect 3819 606 3871 618
rect 3819 0 3871 554
rect 3948 468 4064 1814
rect 8093 2003 8209 2009
rect 8145 1951 8157 2003
rect 8093 1935 8209 1951
rect 8145 1883 8157 1935
rect 8093 1866 8209 1883
rect 8145 1814 8157 1866
rect 5485 1727 5491 1779
rect 5543 1727 5555 1779
rect 5607 1727 5613 1779
rect 6139 1765 6267 1771
rect 5485 1713 5557 1727
tri 5557 1713 5571 1727 nw
rect 6139 1713 6215 1765
rect 5485 1701 5545 1713
tri 5545 1701 5557 1713 nw
rect 6139 1701 6267 1713
rect 4000 416 4012 468
rect 3948 402 4064 416
rect 4000 350 4012 402
rect 3948 344 4064 350
rect 4729 670 4781 676
rect 4729 606 4781 618
rect 4729 0 4781 554
rect 5025 0 5077 547
tri 3115 -127 3121 -121 sw
tri 5479 -127 5485 -121 se
rect 5485 -127 5537 1701
tri 5537 1693 5545 1701 nw
rect 6139 1649 6215 1701
rect 6139 1643 6267 1649
rect 6479 1765 6607 1771
rect 6531 1713 6607 1765
rect 7133 1727 7139 1779
rect 7191 1727 7203 1779
rect 7255 1727 7261 1779
tri 7175 1713 7189 1727 ne
rect 7189 1713 7261 1727
rect 6479 1701 6607 1713
tri 7189 1701 7201 1713 ne
rect 7201 1701 7261 1713
rect 6531 1649 6607 1701
tri 7201 1693 7209 1701 ne
rect 6479 1643 6607 1649
rect 5672 722 5724 728
rect 5672 658 5724 670
rect 5672 -47 5724 606
tri 5724 -47 5730 -41 sw
rect 5672 -75 5730 -47
tri 5730 -75 5758 -47 sw
rect 5672 -127 5678 -75
rect 5730 -127 5742 -75
rect 5794 -127 5800 -75
tri 6133 -127 6139 -121 se
rect 6139 -127 6191 1643
tri 6191 1609 6225 1643 nw
tri 6521 1609 6555 1643 ne
rect 6264 709 6316 715
rect 6264 645 6316 657
rect 6264 0 6316 593
rect 6430 709 6482 715
rect 6430 645 6482 657
rect 6430 0 6482 593
rect 2409 -155 2467 -127
tri 2467 -155 2495 -127 sw
rect 3063 -155 3121 -127
tri 3121 -155 3149 -127 sw
tri 5451 -155 5479 -127 se
rect 5479 -155 5537 -127
tri 6105 -155 6133 -127 se
rect 6133 -155 6191 -127
rect 2409 -207 2415 -155
rect 2467 -207 2479 -155
rect 2531 -207 2537 -155
rect 3063 -207 3069 -155
rect 3121 -207 3133 -155
rect 3185 -207 3191 -155
rect 5409 -207 5415 -155
rect 5467 -207 5479 -155
rect 5531 -207 5537 -155
rect 6063 -207 6069 -155
rect 6121 -207 6133 -155
rect 6185 -207 6191 -155
rect 6555 -127 6607 1643
rect 7022 722 7074 728
rect 7022 658 7074 670
tri 7016 -47 7022 -41 se
rect 7022 -47 7074 606
tri 6988 -75 7016 -47 se
rect 7016 -75 7074 -47
tri 6607 -127 6613 -121 sw
rect 6946 -127 6952 -75
rect 7004 -127 7016 -75
rect 7068 -127 7074 -75
rect 7209 -127 7261 1701
rect 7965 670 8017 676
rect 7965 606 8017 618
rect 7669 0 7721 547
rect 7965 0 8017 554
rect 8093 468 8209 1814
rect 8984 2003 9100 2009
rect 9036 1951 9048 2003
rect 8984 1935 9100 1951
rect 9036 1883 9048 1935
rect 8984 1866 9100 1883
rect 9036 1814 9048 1866
rect 8145 416 8157 468
rect 8093 402 8209 416
rect 8145 350 8157 402
rect 8093 344 8209 350
rect 8875 670 8927 676
rect 8875 606 8927 618
rect 8875 0 8927 554
rect 8984 468 9100 1814
rect 11938 2003 12054 2009
rect 11990 1951 12002 2003
rect 11938 1935 12054 1951
rect 11990 1883 12002 1935
rect 11938 1866 12054 1883
rect 11990 1814 12002 1866
rect 9631 1727 9637 1779
rect 9689 1727 9701 1779
rect 9753 1727 9759 1779
rect 10285 1765 10413 1771
rect 9631 1713 9703 1727
tri 9703 1713 9717 1727 nw
rect 10285 1713 10361 1765
rect 9631 1701 9691 1713
tri 9691 1701 9703 1713 nw
rect 10285 1701 10413 1713
rect 9036 416 9048 468
rect 8984 402 9100 416
rect 9036 350 9048 402
rect 8984 344 9100 350
rect 9171 0 9223 547
tri 7261 -127 7267 -121 sw
tri 9625 -127 9631 -121 se
rect 9631 -127 9683 1701
tri 9683 1693 9691 1701 nw
rect 10285 1649 10361 1701
rect 10285 1643 10413 1649
rect 10625 1765 10753 1771
rect 10677 1713 10753 1765
rect 11279 1727 11285 1779
rect 11337 1727 11349 1779
rect 11401 1727 11407 1779
tri 11321 1713 11335 1727 ne
rect 11335 1713 11407 1727
rect 10625 1701 10753 1713
tri 11335 1701 11347 1713 ne
rect 11347 1701 11407 1713
rect 10677 1649 10753 1701
tri 11347 1693 11355 1701 ne
rect 10625 1643 10753 1649
rect 9818 722 9870 728
rect 9818 658 9870 670
rect 9818 -47 9870 606
tri 9870 -47 9876 -41 sw
rect 9818 -75 9876 -47
tri 9876 -75 9904 -47 sw
rect 9818 -127 9824 -75
rect 9876 -127 9888 -75
rect 9940 -127 9946 -75
tri 10279 -127 10285 -121 se
rect 10285 -127 10337 1643
tri 10337 1609 10371 1643 nw
tri 10667 1609 10701 1643 ne
rect 10410 709 10462 715
rect 10410 645 10462 657
rect 10410 0 10462 593
rect 10576 709 10628 715
rect 10576 645 10628 657
rect 10576 0 10628 593
rect 6555 -155 6613 -127
tri 6613 -155 6641 -127 sw
rect 7209 -155 7267 -127
tri 7267 -155 7295 -127 sw
tri 9597 -155 9625 -127 se
rect 9625 -155 9683 -127
tri 10251 -155 10279 -127 se
rect 10279 -155 10337 -127
rect 6555 -207 6561 -155
rect 6613 -207 6625 -155
rect 6677 -207 6683 -155
rect 7209 -207 7215 -155
rect 7267 -207 7279 -155
rect 7331 -207 7337 -155
rect 9555 -207 9561 -155
rect 9613 -207 9625 -155
rect 9677 -207 9683 -155
rect 10209 -207 10215 -155
rect 10267 -207 10279 -155
rect 10331 -207 10337 -155
rect 10701 -127 10753 1643
rect 11168 722 11220 728
rect 11168 658 11220 670
tri 11162 -47 11168 -41 se
rect 11168 -47 11220 606
tri 11134 -75 11162 -47 se
rect 11162 -75 11220 -47
tri 10753 -127 10759 -121 sw
rect 11092 -127 11098 -75
rect 11150 -127 11162 -75
rect 11214 -127 11220 -75
rect 11355 -127 11407 1701
rect 11815 0 11867 547
rect 11938 468 12054 1814
rect 13130 2003 13246 2009
rect 13182 1951 13194 2003
rect 13130 1935 13246 1951
rect 13182 1883 13194 1935
rect 13130 1866 13246 1883
rect 13182 1814 13194 1866
rect 11990 416 12002 468
rect 11938 402 12054 416
rect 11990 350 12002 402
rect 11938 344 12054 350
rect 12111 670 12163 676
rect 12111 606 12163 618
rect 12111 0 12163 554
rect 13021 670 13073 676
rect 13021 606 13073 618
rect 13021 0 13073 554
rect 13130 468 13246 1814
rect 14639 2003 14691 2009
rect 14639 1935 14691 1951
rect 14639 1866 14691 1883
rect 13777 1727 13783 1779
rect 13835 1727 13847 1779
rect 13899 1727 13905 1779
rect 14422 1765 14559 1771
rect 13777 1713 13849 1727
tri 13849 1713 13863 1727 nw
rect 14422 1713 14507 1765
rect 13777 1701 13837 1713
tri 13837 1701 13849 1713 nw
rect 14422 1701 14559 1713
rect 13182 416 13194 468
rect 13130 402 13246 416
rect 13182 350 13194 402
rect 13130 344 13246 350
rect 13317 0 13369 547
rect 13509 -47 13515 5
rect 13567 -47 13579 5
rect 13631 -47 13637 5
tri 11407 -127 11413 -121 sw
rect 10701 -155 10759 -127
tri 10759 -155 10787 -127 sw
rect 11355 -133 11413 -127
tri 11413 -133 11419 -127 sw
rect 11355 -155 11419 -133
tri 11419 -155 11441 -133 sw
rect 13509 -155 13637 -47
tri 13771 -127 13777 -121 se
rect 13777 -127 13829 1701
tri 13829 1693 13837 1701 nw
rect 14422 1649 14507 1701
rect 14422 1643 14559 1649
rect 14313 1396 14365 1448
rect 14314 1394 14364 1395
rect 14313 1358 14365 1394
rect 14314 1357 14364 1358
rect 14313 1304 14365 1356
tri 14365 1304 14382 1321 sw
tri 14313 1298 14319 1304 ne
rect 14319 1298 14382 1304
tri 14382 1298 14388 1304 sw
tri 14319 1274 14343 1298 ne
rect 13964 722 14016 728
rect 13964 658 14016 670
rect 13964 -47 14016 606
tri 14339 5 14343 9 se
rect 14343 5 14388 1298
tri 14293 -41 14339 5 se
rect 14339 -13 14388 5
rect 14339 -41 14354 -13
tri 14016 -47 14022 -41 sw
tri 14287 -47 14293 -41 se
rect 14293 -47 14354 -41
tri 14354 -47 14388 -13 nw
rect 13964 -75 14022 -47
tri 14022 -75 14050 -47 sw
tri 14282 -52 14287 -47 se
rect 14287 -52 14349 -47
tri 14349 -52 14354 -47 nw
rect 13964 -127 13970 -75
rect 14022 -127 14034 -75
rect 14086 -127 14092 -75
tri 13765 -133 13771 -127 se
rect 13771 -133 13829 -127
tri 13743 -155 13765 -133 se
rect 13765 -155 13829 -133
rect 10701 -207 10707 -155
rect 10759 -207 10771 -155
rect 10823 -207 10829 -155
rect 11355 -207 11361 -155
rect 11413 -207 11425 -155
rect 11477 -207 11483 -155
rect 13509 -207 13515 -155
rect 13567 -207 13579 -155
rect 13631 -207 13637 -155
rect 13701 -207 13707 -155
rect 13759 -207 13771 -155
rect 13823 -207 13829 -155
rect 14282 -427 14326 -52
tri 14326 -75 14349 -52 nw
tri 14416 -127 14422 -121 se
rect 14422 -127 14463 1643
tri 14463 1598 14508 1643 nw
rect 14507 1396 14559 1448
rect 14508 1394 14558 1395
rect 14508 1357 14558 1358
tri 14501 1298 14507 1304 se
rect 14507 1298 14559 1356
tri 14492 1289 14501 1298 se
rect 14501 1289 14559 1298
rect 14492 1287 14559 1289
rect 14492 -75 14526 1287
tri 14526 1254 14559 1287 nw
rect 14556 709 14608 715
rect 14556 645 14608 657
rect 14556 0 14608 593
rect 14639 468 14691 1814
rect 16084 2003 16200 2009
rect 16136 1951 16148 2003
rect 16084 1935 16200 1951
rect 16136 1883 16148 1935
rect 16084 1866 16200 1883
rect 16136 1814 16148 1866
rect 14771 1765 14912 1771
rect 14823 1713 14912 1765
rect 15425 1727 15431 1779
rect 15483 1727 15495 1779
rect 15547 1727 15553 1779
tri 15467 1713 15481 1727 ne
rect 15481 1713 15553 1727
rect 14771 1701 14912 1713
tri 15481 1701 15493 1713 ne
rect 15493 1701 15553 1713
rect 14823 1649 14912 1701
tri 15493 1693 15501 1701 ne
rect 14771 1643 14912 1649
tri 14826 1600 14869 1643 ne
rect 14771 1396 14823 1448
rect 14772 1394 14822 1395
rect 14771 1358 14823 1394
rect 14772 1357 14822 1358
rect 14771 1298 14823 1356
rect 14771 1234 14823 1246
rect 14771 1170 14823 1182
rect 14771 1112 14823 1118
rect 14639 402 14691 416
rect 14639 344 14691 350
rect 14722 709 14774 715
rect 14722 645 14774 657
rect 14722 0 14774 593
tri 14847 5 14869 27 se
rect 14869 5 14912 1643
rect 14965 1396 15017 1448
rect 14966 1394 15016 1395
rect 14966 1357 15016 1358
rect 14965 1298 15017 1356
rect 14965 1234 15017 1246
rect 14965 1170 15017 1182
rect 14965 1112 15017 1118
rect 15314 722 15366 728
rect 15314 658 15366 670
tri 14912 5 14946 39 sw
rect 14847 -47 14853 5
rect 14905 -47 14917 5
rect 14969 -47 14975 5
tri 15308 -47 15314 -41 se
rect 15314 -47 15366 606
rect 15501 5 15553 1701
tri 15553 5 15587 39 sw
rect 15501 -47 15507 5
rect 15559 -47 15571 5
rect 15623 -47 15629 5
rect 15961 0 16013 547
rect 16084 468 16200 1814
rect 17276 2003 17392 2009
rect 17328 1951 17340 2003
rect 17276 1935 17392 1951
rect 17328 1883 17340 1935
rect 17276 1866 17392 1883
rect 17328 1814 17340 1866
rect 16136 416 16148 468
rect 16084 402 16200 416
rect 16136 350 16148 402
rect 16084 344 16200 350
rect 16257 670 16309 676
rect 16257 606 16309 618
rect 16257 0 16309 554
rect 17167 670 17219 676
rect 17167 606 17219 618
rect 17167 0 17219 554
rect 17276 468 17392 1814
rect 18785 2003 18837 2009
rect 18785 1935 18837 1951
rect 18785 1866 18837 1883
rect 17923 1727 17929 1779
rect 17981 1727 17993 1779
rect 18045 1727 18051 1779
rect 18565 1765 18705 1771
rect 17923 1713 17995 1727
tri 17995 1713 18009 1727 nw
rect 18565 1713 18653 1765
rect 17923 1701 17983 1713
tri 17983 1701 17995 1713 nw
rect 18565 1701 18705 1713
rect 17328 416 17340 468
rect 17276 402 17392 416
rect 17328 350 17340 402
rect 17276 344 17392 350
rect 17463 0 17515 547
tri 17889 5 17923 39 se
rect 17923 5 17975 1701
tri 17975 1693 17983 1701 nw
rect 18565 1649 18653 1701
rect 18565 1643 18705 1649
rect 18459 1396 18511 1448
rect 18460 1394 18510 1395
rect 18460 1357 18510 1358
rect 18459 1298 18511 1356
rect 18459 1234 18511 1246
rect 18459 1170 18511 1182
rect 18459 1112 18511 1118
rect 18110 722 18162 728
rect 18110 658 18162 670
rect 18110 468 18162 606
tri 18162 468 18179 485 sw
rect 18110 465 18179 468
tri 18179 465 18182 468 sw
rect 18110 453 18356 465
tri 18110 442 18121 453 ne
rect 18121 442 18356 453
tri 18356 442 18379 465 sw
tri 18121 416 18147 442 ne
rect 18147 416 18379 442
tri 18147 415 18148 416 ne
rect 18148 415 18379 416
tri 18298 402 18311 415 ne
rect 18311 402 18379 415
tri 18311 390 18323 402 ne
rect 17847 -47 17853 5
rect 17905 -47 17917 5
rect 17969 -47 17975 5
tri 18317 -47 18323 -41 se
rect 18323 -47 18379 402
tri 18531 5 18565 39 se
rect 18565 5 18608 1643
tri 18608 1600 18651 1643 nw
rect 18653 1396 18705 1448
rect 18654 1394 18704 1395
rect 18653 1358 18705 1394
rect 18654 1357 18704 1358
rect 18653 1298 18705 1356
rect 18653 1234 18705 1246
rect 18653 1170 18705 1182
rect 18653 1112 18705 1118
rect 18479 -47 18486 5
rect 18538 -47 18550 5
rect 18602 -47 18608 5
rect 18702 709 18754 715
rect 18702 645 18754 657
rect 18702 0 18754 593
rect 18785 468 18837 1814
rect 20230 2003 20346 2009
rect 20282 1951 20294 2003
rect 20230 1935 20346 1951
rect 20282 1883 20294 1935
rect 20230 1866 20346 1883
rect 20282 1814 20294 1866
rect 18917 1765 19058 1771
rect 18969 1713 19058 1765
rect 19571 1727 19577 1779
rect 19629 1727 19641 1779
rect 19693 1727 19699 1779
rect 18917 1701 19058 1713
rect 18969 1649 19058 1701
tri 19613 1693 19647 1727 ne
rect 18917 1643 19058 1649
tri 18981 1609 19015 1643 ne
rect 18917 1396 18969 1448
rect 18918 1394 18968 1395
rect 18917 1358 18969 1394
rect 18918 1357 18968 1358
rect 18917 1289 18969 1356
tri 18969 1289 18984 1304 sw
rect 18917 1287 18984 1289
tri 18917 1254 18950 1287 ne
rect 18785 402 18837 416
rect 18785 344 18837 350
rect 18868 709 18920 715
rect 18868 645 18920 657
rect 18868 0 18920 593
tri 15301 -54 15308 -47 se
rect 15308 -54 15366 -47
tri 14526 -75 14547 -54 sw
tri 15280 -75 15301 -54 se
rect 15301 -75 15366 -54
tri 18289 -75 18317 -47 se
rect 18317 -75 18379 -47
tri 18947 -75 18950 -72 se
rect 18950 -75 18984 1287
rect 14492 -79 14547 -75
tri 14547 -79 14551 -75 sw
tri 14492 -108 14521 -79 ne
rect 14521 -84 14551 -79
tri 14551 -84 14556 -79 sw
tri 14410 -133 14416 -127 se
rect 14416 -133 14463 -127
tri 14388 -155 14410 -133 se
rect 14410 -155 14463 -133
tri 14463 -155 14483 -135 sw
rect 14355 -207 14361 -155
rect 14413 -207 14425 -155
rect 14477 -207 14483 -155
rect 14521 -427 14556 -84
rect 15238 -127 15244 -75
rect 15296 -127 15308 -75
rect 15360 -127 15366 -75
rect 18251 -127 18257 -75
rect 18309 -127 18321 -75
rect 18373 -127 18379 -75
tri 18928 -94 18947 -75 se
rect 18947 -94 18984 -75
rect 18928 -97 18984 -94
rect 18501 -207 18507 -155
rect 18559 -207 18571 -155
rect 18623 -207 18629 -155
rect 14245 -479 14251 -427
rect 14303 -479 14315 -427
rect 14367 -479 14373 -427
rect 14465 -479 14471 -427
rect 14523 -479 14535 -427
rect 14587 -479 14593 -427
rect 18928 -935 18963 -97
tri 18963 -118 18984 -97 nw
rect 19015 -127 19058 1643
rect 19111 1396 19163 1448
rect 19112 1394 19162 1395
rect 19112 1357 19162 1358
tri 19094 1304 19111 1321 se
rect 19111 1304 19163 1356
tri 19088 1298 19094 1304 se
rect 19094 1298 19133 1304
rect 19088 -13 19133 1298
tri 19133 1274 19163 1304 nw
rect 19460 722 19512 728
rect 19460 658 19512 670
tri 19088 -52 19127 -13 ne
rect 19127 -41 19133 -13
tri 19133 -41 19183 9 sw
rect 19127 -47 19183 -41
tri 19183 -47 19189 -41 sw
tri 19454 -47 19460 -41 se
rect 19460 -47 19512 606
rect 19127 -52 19189 -47
tri 19189 -52 19194 -47 sw
tri 19127 -58 19133 -52 ne
rect 19133 -58 19194 -52
tri 19133 -75 19150 -58 ne
tri 19058 -127 19073 -112 sw
tri 18993 -155 19015 -133 se
rect 19015 -155 19073 -127
tri 19073 -155 19101 -127 sw
rect 18993 -207 18999 -155
rect 19051 -207 19063 -155
rect 19115 -207 19121 -155
tri 19089 -300 19150 -239 se
rect 19150 -264 19194 -58
tri 19426 -75 19454 -47 se
rect 19454 -75 19512 -47
rect 19384 -127 19390 -75
rect 19442 -127 19454 -75
rect 19506 -127 19512 -75
rect 19647 -127 19699 1727
rect 20107 0 20159 547
rect 20230 468 20346 1814
rect 20282 416 20294 468
rect 20230 402 20346 416
rect 20282 350 20294 402
rect 20230 344 20346 350
rect 20403 670 20455 676
rect 20403 606 20455 618
rect 20403 0 20455 554
tri 19699 -127 19705 -121 sw
rect 19647 -155 19705 -127
tri 19705 -155 19733 -127 sw
rect 19647 -207 19653 -155
rect 19705 -207 19717 -155
rect 19769 -207 19775 -155
rect 19150 -300 19158 -264
tri 19158 -300 19194 -264 nw
rect 19089 -939 19124 -300
tri 19124 -334 19158 -300 nw
<< rmetal2 >>
rect 14313 1395 14365 1396
rect 14313 1394 14314 1395
rect 14364 1394 14365 1395
rect 14313 1357 14314 1358
rect 14364 1357 14365 1358
rect 14313 1356 14365 1357
rect 14507 1395 14559 1396
rect 14507 1394 14508 1395
rect 14558 1394 14559 1395
rect 14507 1357 14508 1358
rect 14558 1357 14559 1358
rect 14507 1356 14559 1357
rect 14771 1395 14823 1396
rect 14771 1394 14772 1395
rect 14822 1394 14823 1395
rect 14771 1357 14772 1358
rect 14822 1357 14823 1358
rect 14771 1356 14823 1357
rect 14965 1395 15017 1396
rect 14965 1394 14966 1395
rect 15016 1394 15017 1395
rect 14965 1357 14966 1358
rect 15016 1357 15017 1358
rect 14965 1356 15017 1357
rect 18459 1395 18511 1396
rect 18459 1394 18460 1395
rect 18510 1394 18511 1395
rect 18459 1357 18460 1358
rect 18510 1357 18511 1358
rect 18459 1356 18511 1357
rect 18653 1395 18705 1396
rect 18653 1394 18654 1395
rect 18704 1394 18705 1395
rect 18653 1357 18654 1358
rect 18704 1357 18705 1358
rect 18653 1356 18705 1357
rect 18917 1395 18969 1396
rect 18917 1394 18918 1395
rect 18968 1394 18969 1395
rect 18917 1357 18918 1358
rect 18968 1357 18969 1358
rect 18917 1356 18969 1357
rect 19111 1395 19163 1396
rect 19111 1394 19112 1395
rect 19162 1394 19163 1395
rect 19111 1357 19112 1358
rect 19162 1357 19163 1358
rect 19111 1356 19163 1357
use sky130_fd_io__com_ctl_ls_ovt  sky130_fd_io__com_ctl_ls_ovt_0
timestamp 1648127584
transform -1 0 12592 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovt  sky130_fd_io__com_ctl_ls_ovt_1
timestamp 1648127584
transform 1 0 8446 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovt  sky130_fd_io__com_ctl_ls_ovt_2
timestamp 1648127584
transform -1 0 8446 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovt  sky130_fd_io__com_ctl_ls_ovt_3
timestamp 1648127584
transform 1 0 4300 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovt  sky130_fd_io__com_ctl_ls_ovt_4
timestamp 1648127584
transform 1 0 154 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovt  sky130_fd_io__com_ctl_ls_ovt_5
timestamp 1648127584
transform -1 0 4300 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovtv2  sky130_fd_io__com_ctl_ls_ovtv2_0
timestamp 1648127584
transform 1 0 16738 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovtv2  sky130_fd_io__com_ctl_ls_ovtv2_1
timestamp 1648127584
transform -1 0 20884 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovtv2  sky130_fd_io__com_ctl_ls_ovtv2_2
timestamp 1648127584
transform 1 0 12592 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls_ovtv2  sky130_fd_io__com_ctl_ls_ovtv2_3
timestamp 1648127584
transform -1 0 16738 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x2  sky130_fd_io__hvsbt_inv_x2_0
timestamp 1648127584
transform -1 0 -5199 0 1 -74
box 0 24 534 1116
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_0
timestamp 1648127584
transform 0 1 10825 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_1
timestamp 1648127584
transform 0 -1 10213 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_2
timestamp 1648127584
transform 0 1 6679 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_3
timestamp 1648127584
transform 0 -1 6067 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_4
timestamp 1648127584
transform 0 1 2533 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_5
timestamp 1648127584
transform 0 -1 1921 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1648127584
transform 0 1 18917 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1648127584
transform 0 -1 18705 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_2
timestamp 1648127584
transform 0 1 14771 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_3
timestamp 1648127584
transform 0 1 14307 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_4
timestamp 1648127584
transform 0 1 10625 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_5
timestamp 1648127584
transform 0 -1 10413 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_6
timestamp 1648127584
transform 0 1 6479 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_7
timestamp 1648127584
transform 0 -1 6267 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_8
timestamp 1648127584
transform 0 1 2333 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_9
timestamp 1648127584
transform 0 -1 2121 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_0
timestamp 1648127584
transform 0 1 19117 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_1
timestamp 1648127584
transform 0 -1 18505 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_2
timestamp 1648127584
transform 0 1 14971 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_3
timestamp 1648127584
transform 0 1 14507 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_4
timestamp 1648127584
transform 0 1 10825 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_5
timestamp 1648127584
transform 0 -1 10213 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_6
timestamp 1648127584
transform 0 1 6679 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_7
timestamp 1648127584
transform 0 -1 6067 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_8
timestamp 1648127584
transform 0 1 2533 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_9
timestamp 1648127584
transform 0 -1 1921 -1 0 1684
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1648127584
transform 0 1 10625 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1648127584
transform 0 -1 10413 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_2
timestamp 1648127584
transform 0 1 6479 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_3
timestamp 1648127584
transform 0 -1 6267 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_4
timestamp 1648127584
transform 0 1 2333 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_5
timestamp 1648127584
transform 0 -1 2121 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2o_cdns_55959141808439  sky130_fd_io__tk_em2o_cdns_55959141808439_0
timestamp 1648127584
transform 0 1 19111 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2o_cdns_55959141808439  sky130_fd_io__tk_em2o_cdns_55959141808439_1
timestamp 1648127584
transform 0 -1 18511 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2o_cdns_55959141808439  sky130_fd_io__tk_em2o_cdns_55959141808439_2
timestamp 1648127584
transform 0 1 14965 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2o_cdns_55959141808439  sky130_fd_io__tk_em2o_cdns_55959141808439_3
timestamp 1648127584
transform 0 1 14507 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2s_cdns_55959141808438  sky130_fd_io__tk_em2s_cdns_55959141808438_0
timestamp 1648127584
transform 0 1 18917 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2s_cdns_55959141808438  sky130_fd_io__tk_em2s_cdns_55959141808438_1
timestamp 1648127584
transform 0 -1 18705 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2s_cdns_55959141808438  sky130_fd_io__tk_em2s_cdns_55959141808438_2
timestamp 1648127584
transform 0 1 14771 -1 0 1448
box 0 24 144 28
use sky130_fd_io__tk_em2s_cdns_55959141808438  sky130_fd_io__tk_em2s_cdns_55959141808438_3
timestamp 1648127584
transform 0 1 14313 -1 0 1448
box 0 24 144 28
<< labels >>
flabel metal2 s 14727 13 14768 105 3 FreeSans 200 0 0 0 DM[2]
port 1 nsew
flabel metal2 s 18707 16 18742 139 3 FreeSans 200 0 0 0 DM[1]
port 2 nsew
flabel metal2 s 18876 20 18913 127 3 FreeSans 200 0 0 0 DM[0]
port 3 nsew
flabel metal2 s 14560 9 14600 89 3 FreeSans 200 0 0 0 INP_DIS
port 4 nsew
flabel metal2 s 10581 8 10620 93 3 FreeSans 200 0 0 0 VTRIP_SEL
port 5 nsew
flabel metal2 s 10415 11 10452 103 3 FreeSans 200 180 0 0 IB_MODE_SEL[0]
port 6 nsew
flabel metal2 s 6437 14 6475 108 3 FreeSans 200 0 0 0 IB_MODE_SEL[1]
port 7 nsew
flabel metal2 s 6276 22 6307 93 3 FreeSans 200 0 0 0 SLEW_CTL[0]
port 8 nsew
flabel metal2 s 2292 20 2327 113 3 FreeSans 200 0 0 0 SLEW_CTL[1]
port 9 nsew
flabel metal2 s 2121 14 2166 106 3 FreeSans 200 0 0 0 HYST_TRIM
port 10 nsew
flabel metal2 s 20115 24 20152 142 3 FreeSans 200 0 0 0 DM_H_N[0]
port 11 nsew
flabel metal2 s 17475 24 17505 152 3 FreeSans 200 0 0 0 DM_H_N[1]
port 12 nsew
flabel metal2 s 15972 18 16005 141 3 FreeSans 200 0 0 0 DM_H_N[2]
port 13 nsew
flabel metal2 s 20409 23 20447 109 3 FreeSans 200 0 0 0 DM_H[0]
port 14 nsew
flabel metal2 s 17172 19 17206 110 3 FreeSans 200 0 0 0 DM_H[1]
port 15 nsew
flabel metal2 s 16260 30 16303 124 3 FreeSans 200 0 0 0 DM_H[2]
port 16 nsew
flabel metal2 s 13026 8 13066 95 3 FreeSans 200 0 0 0 INP_DIS_H
port 17 nsew
flabel metal2 s 13324 13 13363 103 3 FreeSans 200 0 0 0 INP_DIS_H_N
port 18 nsew
flabel metal2 s 12113 12 12155 104 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 19 nsew
flabel metal2 s 11818 20 11862 104 3 FreeSans 200 0 0 0 VTRIP_SEL_H_N
port 20 nsew
flabel metal2 s 8880 12 8918 97 3 FreeSans 200 0 0 0 IB_MODE_SEL_H[0]
port 21 nsew
flabel metal2 s 7971 16 8009 126 3 FreeSans 200 0 0 0 IB_MODE_SEL_H[1]
port 22 nsew
flabel metal2 s 9179 19 9217 115 3 FreeSans 200 0 0 0 IB_MODE_SEL_H_N[0]
port 23 nsew
flabel metal2 s 7675 19 7711 146 3 FreeSans 200 0 0 0 IB_MODE_SEL_H_N[1]
port 24 nsew
flabel metal2 s 4733 10 4771 120 3 FreeSans 200 0 0 0 SLEW_CTL_H[0]
port 25 nsew
flabel metal2 s 3825 16 3863 125 3 FreeSans 200 0 0 0 SLEW_CTL_H[1]
port 26 nsew
flabel metal2 s 5031 17 5067 147 3 FreeSans 200 0 0 0 SLEW_CTL_H_N[0]
port 27 nsew
flabel metal2 s 3530 18 3569 155 3 FreeSans 200 0 0 0 SLEW_CTL_H_N[1]
port 28 nsew
flabel metal2 s 587 7 629 121 3 FreeSans 200 0 0 0 HYST_TRIM_H
port 29 nsew
flabel metal2 s 882 6 927 124 3 FreeSans 200 0 0 0 HYST_TRIM_H_N
port 30 nsew
flabel metal2 s 19090 -476 19122 -444 3 FreeSans 520 90 0 0 STARTUP_ST_H
port 31 nsew
flabel metal2 s 18930 -476 18962 -444 3 FreeSans 520 90 0 0 STARTUP_ST_H
port 31 nsew
flabel metal2 s 14284 -476 14316 -444 3 FreeSans 520 90 0 0 STARTUP_ST_H
port 31 nsew
flabel metal2 s 14526 -468 14558 -436 3 FreeSans 520 0 0 0 STARTUP_ST_H
port 31 nsew
flabel metal2 s 14403 -193 14453 -164 3 FreeSans 520 90 0 0 STARTUP_RST_H
port 32 nsew
flabel metal1 s 208 1127 499 1290 3 FreeSans 400 0 0 0 VGND
port 33 nsew
flabel metal1 s 212 132 569 298 3 FreeSans 400 0 0 0 VCC_IO
port 34 nsew
flabel metal1 s 202 1826 501 2002 3 FreeSans 400 0 0 0 VPWR
port 35 nsew
flabel metal1 s 6 -119 117 -85 3 FreeSans 400 0 0 0 HLD_I_H_N
port 36 nsew
flabel metal1 s -5502 884 -5502 884 0 FreeSans 440 0 0 0 VCC_IO
port 34 nsew
flabel metal1 s -5485 87 -5485 87 0 FreeSans 440 0 0 0 VGND
port 33 nsew
flabel metal1 s -5570 298 -5544 336 3 FreeSans 520 0 0 0 OD_I_H_N
port 37 nsew
<< properties >>
string GDS_END 35906586
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35846530
<< end >>
