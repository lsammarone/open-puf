magic
tech sky130A
magscale 1 2
timestamp 1654402208
<< metal3 >>
rect -3150 12522 3149 12550
rect -3150 12458 3065 12522
rect 3129 12458 3149 12522
rect -3150 12442 3149 12458
rect -3150 12378 3065 12442
rect 3129 12378 3149 12442
rect -3150 12362 3149 12378
rect -3150 12298 3065 12362
rect 3129 12298 3149 12362
rect -3150 12282 3149 12298
rect -3150 12218 3065 12282
rect 3129 12218 3149 12282
rect -3150 12202 3149 12218
rect -3150 12138 3065 12202
rect 3129 12138 3149 12202
rect -3150 12122 3149 12138
rect -3150 12058 3065 12122
rect 3129 12058 3149 12122
rect -3150 12042 3149 12058
rect -3150 11978 3065 12042
rect 3129 11978 3149 12042
rect -3150 11962 3149 11978
rect -3150 11898 3065 11962
rect 3129 11898 3149 11962
rect -3150 11882 3149 11898
rect -3150 11818 3065 11882
rect 3129 11818 3149 11882
rect -3150 11802 3149 11818
rect -3150 11738 3065 11802
rect 3129 11738 3149 11802
rect -3150 11722 3149 11738
rect -3150 11658 3065 11722
rect 3129 11658 3149 11722
rect -3150 11642 3149 11658
rect -3150 11578 3065 11642
rect 3129 11578 3149 11642
rect -3150 11562 3149 11578
rect -3150 11498 3065 11562
rect 3129 11498 3149 11562
rect -3150 11482 3149 11498
rect -3150 11418 3065 11482
rect 3129 11418 3149 11482
rect -3150 11402 3149 11418
rect -3150 11338 3065 11402
rect 3129 11338 3149 11402
rect -3150 11322 3149 11338
rect -3150 11258 3065 11322
rect 3129 11258 3149 11322
rect -3150 11242 3149 11258
rect -3150 11178 3065 11242
rect 3129 11178 3149 11242
rect -3150 11162 3149 11178
rect -3150 11098 3065 11162
rect 3129 11098 3149 11162
rect -3150 11082 3149 11098
rect -3150 11018 3065 11082
rect 3129 11018 3149 11082
rect -3150 11002 3149 11018
rect -3150 10938 3065 11002
rect 3129 10938 3149 11002
rect -3150 10922 3149 10938
rect -3150 10858 3065 10922
rect 3129 10858 3149 10922
rect -3150 10842 3149 10858
rect -3150 10778 3065 10842
rect 3129 10778 3149 10842
rect -3150 10762 3149 10778
rect -3150 10698 3065 10762
rect 3129 10698 3149 10762
rect -3150 10682 3149 10698
rect -3150 10618 3065 10682
rect 3129 10618 3149 10682
rect -3150 10602 3149 10618
rect -3150 10538 3065 10602
rect 3129 10538 3149 10602
rect -3150 10522 3149 10538
rect -3150 10458 3065 10522
rect 3129 10458 3149 10522
rect -3150 10442 3149 10458
rect -3150 10378 3065 10442
rect 3129 10378 3149 10442
rect -3150 10362 3149 10378
rect -3150 10298 3065 10362
rect 3129 10298 3149 10362
rect -3150 10282 3149 10298
rect -3150 10218 3065 10282
rect 3129 10218 3149 10282
rect -3150 10202 3149 10218
rect -3150 10138 3065 10202
rect 3129 10138 3149 10202
rect -3150 10122 3149 10138
rect -3150 10058 3065 10122
rect 3129 10058 3149 10122
rect -3150 10042 3149 10058
rect -3150 9978 3065 10042
rect 3129 9978 3149 10042
rect -3150 9962 3149 9978
rect -3150 9898 3065 9962
rect 3129 9898 3149 9962
rect -3150 9882 3149 9898
rect -3150 9818 3065 9882
rect 3129 9818 3149 9882
rect -3150 9802 3149 9818
rect -3150 9738 3065 9802
rect 3129 9738 3149 9802
rect -3150 9722 3149 9738
rect -3150 9658 3065 9722
rect 3129 9658 3149 9722
rect -3150 9642 3149 9658
rect -3150 9578 3065 9642
rect 3129 9578 3149 9642
rect -3150 9562 3149 9578
rect -3150 9498 3065 9562
rect 3129 9498 3149 9562
rect -3150 9482 3149 9498
rect -3150 9418 3065 9482
rect 3129 9418 3149 9482
rect -3150 9402 3149 9418
rect -3150 9338 3065 9402
rect 3129 9338 3149 9402
rect -3150 9322 3149 9338
rect -3150 9258 3065 9322
rect 3129 9258 3149 9322
rect -3150 9242 3149 9258
rect -3150 9178 3065 9242
rect 3129 9178 3149 9242
rect -3150 9162 3149 9178
rect -3150 9098 3065 9162
rect 3129 9098 3149 9162
rect -3150 9082 3149 9098
rect -3150 9018 3065 9082
rect 3129 9018 3149 9082
rect -3150 9002 3149 9018
rect -3150 8938 3065 9002
rect 3129 8938 3149 9002
rect -3150 8922 3149 8938
rect -3150 8858 3065 8922
rect 3129 8858 3149 8922
rect -3150 8842 3149 8858
rect -3150 8778 3065 8842
rect 3129 8778 3149 8842
rect -3150 8762 3149 8778
rect -3150 8698 3065 8762
rect 3129 8698 3149 8762
rect -3150 8682 3149 8698
rect -3150 8618 3065 8682
rect 3129 8618 3149 8682
rect -3150 8602 3149 8618
rect -3150 8538 3065 8602
rect 3129 8538 3149 8602
rect -3150 8522 3149 8538
rect -3150 8458 3065 8522
rect 3129 8458 3149 8522
rect -3150 8442 3149 8458
rect -3150 8378 3065 8442
rect 3129 8378 3149 8442
rect -3150 8362 3149 8378
rect -3150 8298 3065 8362
rect 3129 8298 3149 8362
rect -3150 8282 3149 8298
rect -3150 8218 3065 8282
rect 3129 8218 3149 8282
rect -3150 8202 3149 8218
rect -3150 8138 3065 8202
rect 3129 8138 3149 8202
rect -3150 8122 3149 8138
rect -3150 8058 3065 8122
rect 3129 8058 3149 8122
rect -3150 8042 3149 8058
rect -3150 7978 3065 8042
rect 3129 7978 3149 8042
rect -3150 7962 3149 7978
rect -3150 7898 3065 7962
rect 3129 7898 3149 7962
rect -3150 7882 3149 7898
rect -3150 7818 3065 7882
rect 3129 7818 3149 7882
rect -3150 7802 3149 7818
rect -3150 7738 3065 7802
rect 3129 7738 3149 7802
rect -3150 7722 3149 7738
rect -3150 7658 3065 7722
rect 3129 7658 3149 7722
rect -3150 7642 3149 7658
rect -3150 7578 3065 7642
rect 3129 7578 3149 7642
rect -3150 7562 3149 7578
rect -3150 7498 3065 7562
rect 3129 7498 3149 7562
rect -3150 7482 3149 7498
rect -3150 7418 3065 7482
rect 3129 7418 3149 7482
rect -3150 7402 3149 7418
rect -3150 7338 3065 7402
rect 3129 7338 3149 7402
rect -3150 7322 3149 7338
rect -3150 7258 3065 7322
rect 3129 7258 3149 7322
rect -3150 7242 3149 7258
rect -3150 7178 3065 7242
rect 3129 7178 3149 7242
rect -3150 7162 3149 7178
rect -3150 7098 3065 7162
rect 3129 7098 3149 7162
rect -3150 7082 3149 7098
rect -3150 7018 3065 7082
rect 3129 7018 3149 7082
rect -3150 7002 3149 7018
rect -3150 6938 3065 7002
rect 3129 6938 3149 7002
rect -3150 6922 3149 6938
rect -3150 6858 3065 6922
rect 3129 6858 3149 6922
rect -3150 6842 3149 6858
rect -3150 6778 3065 6842
rect 3129 6778 3149 6842
rect -3150 6762 3149 6778
rect -3150 6698 3065 6762
rect 3129 6698 3149 6762
rect -3150 6682 3149 6698
rect -3150 6618 3065 6682
rect 3129 6618 3149 6682
rect -3150 6602 3149 6618
rect -3150 6538 3065 6602
rect 3129 6538 3149 6602
rect -3150 6522 3149 6538
rect -3150 6458 3065 6522
rect 3129 6458 3149 6522
rect -3150 6442 3149 6458
rect -3150 6378 3065 6442
rect 3129 6378 3149 6442
rect -3150 6350 3149 6378
rect -3150 6222 3149 6250
rect -3150 6158 3065 6222
rect 3129 6158 3149 6222
rect -3150 6142 3149 6158
rect -3150 6078 3065 6142
rect 3129 6078 3149 6142
rect -3150 6062 3149 6078
rect -3150 5998 3065 6062
rect 3129 5998 3149 6062
rect -3150 5982 3149 5998
rect -3150 5918 3065 5982
rect 3129 5918 3149 5982
rect -3150 5902 3149 5918
rect -3150 5838 3065 5902
rect 3129 5838 3149 5902
rect -3150 5822 3149 5838
rect -3150 5758 3065 5822
rect 3129 5758 3149 5822
rect -3150 5742 3149 5758
rect -3150 5678 3065 5742
rect 3129 5678 3149 5742
rect -3150 5662 3149 5678
rect -3150 5598 3065 5662
rect 3129 5598 3149 5662
rect -3150 5582 3149 5598
rect -3150 5518 3065 5582
rect 3129 5518 3149 5582
rect -3150 5502 3149 5518
rect -3150 5438 3065 5502
rect 3129 5438 3149 5502
rect -3150 5422 3149 5438
rect -3150 5358 3065 5422
rect 3129 5358 3149 5422
rect -3150 5342 3149 5358
rect -3150 5278 3065 5342
rect 3129 5278 3149 5342
rect -3150 5262 3149 5278
rect -3150 5198 3065 5262
rect 3129 5198 3149 5262
rect -3150 5182 3149 5198
rect -3150 5118 3065 5182
rect 3129 5118 3149 5182
rect -3150 5102 3149 5118
rect -3150 5038 3065 5102
rect 3129 5038 3149 5102
rect -3150 5022 3149 5038
rect -3150 4958 3065 5022
rect 3129 4958 3149 5022
rect -3150 4942 3149 4958
rect -3150 4878 3065 4942
rect 3129 4878 3149 4942
rect -3150 4862 3149 4878
rect -3150 4798 3065 4862
rect 3129 4798 3149 4862
rect -3150 4782 3149 4798
rect -3150 4718 3065 4782
rect 3129 4718 3149 4782
rect -3150 4702 3149 4718
rect -3150 4638 3065 4702
rect 3129 4638 3149 4702
rect -3150 4622 3149 4638
rect -3150 4558 3065 4622
rect 3129 4558 3149 4622
rect -3150 4542 3149 4558
rect -3150 4478 3065 4542
rect 3129 4478 3149 4542
rect -3150 4462 3149 4478
rect -3150 4398 3065 4462
rect 3129 4398 3149 4462
rect -3150 4382 3149 4398
rect -3150 4318 3065 4382
rect 3129 4318 3149 4382
rect -3150 4302 3149 4318
rect -3150 4238 3065 4302
rect 3129 4238 3149 4302
rect -3150 4222 3149 4238
rect -3150 4158 3065 4222
rect 3129 4158 3149 4222
rect -3150 4142 3149 4158
rect -3150 4078 3065 4142
rect 3129 4078 3149 4142
rect -3150 4062 3149 4078
rect -3150 3998 3065 4062
rect 3129 3998 3149 4062
rect -3150 3982 3149 3998
rect -3150 3918 3065 3982
rect 3129 3918 3149 3982
rect -3150 3902 3149 3918
rect -3150 3838 3065 3902
rect 3129 3838 3149 3902
rect -3150 3822 3149 3838
rect -3150 3758 3065 3822
rect 3129 3758 3149 3822
rect -3150 3742 3149 3758
rect -3150 3678 3065 3742
rect 3129 3678 3149 3742
rect -3150 3662 3149 3678
rect -3150 3598 3065 3662
rect 3129 3598 3149 3662
rect -3150 3582 3149 3598
rect -3150 3518 3065 3582
rect 3129 3518 3149 3582
rect -3150 3502 3149 3518
rect -3150 3438 3065 3502
rect 3129 3438 3149 3502
rect -3150 3422 3149 3438
rect -3150 3358 3065 3422
rect 3129 3358 3149 3422
rect -3150 3342 3149 3358
rect -3150 3278 3065 3342
rect 3129 3278 3149 3342
rect -3150 3262 3149 3278
rect -3150 3198 3065 3262
rect 3129 3198 3149 3262
rect -3150 3182 3149 3198
rect -3150 3118 3065 3182
rect 3129 3118 3149 3182
rect -3150 3102 3149 3118
rect -3150 3038 3065 3102
rect 3129 3038 3149 3102
rect -3150 3022 3149 3038
rect -3150 2958 3065 3022
rect 3129 2958 3149 3022
rect -3150 2942 3149 2958
rect -3150 2878 3065 2942
rect 3129 2878 3149 2942
rect -3150 2862 3149 2878
rect -3150 2798 3065 2862
rect 3129 2798 3149 2862
rect -3150 2782 3149 2798
rect -3150 2718 3065 2782
rect 3129 2718 3149 2782
rect -3150 2702 3149 2718
rect -3150 2638 3065 2702
rect 3129 2638 3149 2702
rect -3150 2622 3149 2638
rect -3150 2558 3065 2622
rect 3129 2558 3149 2622
rect -3150 2542 3149 2558
rect -3150 2478 3065 2542
rect 3129 2478 3149 2542
rect -3150 2462 3149 2478
rect -3150 2398 3065 2462
rect 3129 2398 3149 2462
rect -3150 2382 3149 2398
rect -3150 2318 3065 2382
rect 3129 2318 3149 2382
rect -3150 2302 3149 2318
rect -3150 2238 3065 2302
rect 3129 2238 3149 2302
rect -3150 2222 3149 2238
rect -3150 2158 3065 2222
rect 3129 2158 3149 2222
rect -3150 2142 3149 2158
rect -3150 2078 3065 2142
rect 3129 2078 3149 2142
rect -3150 2062 3149 2078
rect -3150 1998 3065 2062
rect 3129 1998 3149 2062
rect -3150 1982 3149 1998
rect -3150 1918 3065 1982
rect 3129 1918 3149 1982
rect -3150 1902 3149 1918
rect -3150 1838 3065 1902
rect 3129 1838 3149 1902
rect -3150 1822 3149 1838
rect -3150 1758 3065 1822
rect 3129 1758 3149 1822
rect -3150 1742 3149 1758
rect -3150 1678 3065 1742
rect 3129 1678 3149 1742
rect -3150 1662 3149 1678
rect -3150 1598 3065 1662
rect 3129 1598 3149 1662
rect -3150 1582 3149 1598
rect -3150 1518 3065 1582
rect 3129 1518 3149 1582
rect -3150 1502 3149 1518
rect -3150 1438 3065 1502
rect 3129 1438 3149 1502
rect -3150 1422 3149 1438
rect -3150 1358 3065 1422
rect 3129 1358 3149 1422
rect -3150 1342 3149 1358
rect -3150 1278 3065 1342
rect 3129 1278 3149 1342
rect -3150 1262 3149 1278
rect -3150 1198 3065 1262
rect 3129 1198 3149 1262
rect -3150 1182 3149 1198
rect -3150 1118 3065 1182
rect 3129 1118 3149 1182
rect -3150 1102 3149 1118
rect -3150 1038 3065 1102
rect 3129 1038 3149 1102
rect -3150 1022 3149 1038
rect -3150 958 3065 1022
rect 3129 958 3149 1022
rect -3150 942 3149 958
rect -3150 878 3065 942
rect 3129 878 3149 942
rect -3150 862 3149 878
rect -3150 798 3065 862
rect 3129 798 3149 862
rect -3150 782 3149 798
rect -3150 718 3065 782
rect 3129 718 3149 782
rect -3150 702 3149 718
rect -3150 638 3065 702
rect 3129 638 3149 702
rect -3150 622 3149 638
rect -3150 558 3065 622
rect 3129 558 3149 622
rect -3150 542 3149 558
rect -3150 478 3065 542
rect 3129 478 3149 542
rect -3150 462 3149 478
rect -3150 398 3065 462
rect 3129 398 3149 462
rect -3150 382 3149 398
rect -3150 318 3065 382
rect 3129 318 3149 382
rect -3150 302 3149 318
rect -3150 238 3065 302
rect 3129 238 3149 302
rect -3150 222 3149 238
rect -3150 158 3065 222
rect 3129 158 3149 222
rect -3150 142 3149 158
rect -3150 78 3065 142
rect 3129 78 3149 142
rect -3150 50 3149 78
rect -3150 -78 3149 -50
rect -3150 -142 3065 -78
rect 3129 -142 3149 -78
rect -3150 -158 3149 -142
rect -3150 -222 3065 -158
rect 3129 -222 3149 -158
rect -3150 -238 3149 -222
rect -3150 -302 3065 -238
rect 3129 -302 3149 -238
rect -3150 -318 3149 -302
rect -3150 -382 3065 -318
rect 3129 -382 3149 -318
rect -3150 -398 3149 -382
rect -3150 -462 3065 -398
rect 3129 -462 3149 -398
rect -3150 -478 3149 -462
rect -3150 -542 3065 -478
rect 3129 -542 3149 -478
rect -3150 -558 3149 -542
rect -3150 -622 3065 -558
rect 3129 -622 3149 -558
rect -3150 -638 3149 -622
rect -3150 -702 3065 -638
rect 3129 -702 3149 -638
rect -3150 -718 3149 -702
rect -3150 -782 3065 -718
rect 3129 -782 3149 -718
rect -3150 -798 3149 -782
rect -3150 -862 3065 -798
rect 3129 -862 3149 -798
rect -3150 -878 3149 -862
rect -3150 -942 3065 -878
rect 3129 -942 3149 -878
rect -3150 -958 3149 -942
rect -3150 -1022 3065 -958
rect 3129 -1022 3149 -958
rect -3150 -1038 3149 -1022
rect -3150 -1102 3065 -1038
rect 3129 -1102 3149 -1038
rect -3150 -1118 3149 -1102
rect -3150 -1182 3065 -1118
rect 3129 -1182 3149 -1118
rect -3150 -1198 3149 -1182
rect -3150 -1262 3065 -1198
rect 3129 -1262 3149 -1198
rect -3150 -1278 3149 -1262
rect -3150 -1342 3065 -1278
rect 3129 -1342 3149 -1278
rect -3150 -1358 3149 -1342
rect -3150 -1422 3065 -1358
rect 3129 -1422 3149 -1358
rect -3150 -1438 3149 -1422
rect -3150 -1502 3065 -1438
rect 3129 -1502 3149 -1438
rect -3150 -1518 3149 -1502
rect -3150 -1582 3065 -1518
rect 3129 -1582 3149 -1518
rect -3150 -1598 3149 -1582
rect -3150 -1662 3065 -1598
rect 3129 -1662 3149 -1598
rect -3150 -1678 3149 -1662
rect -3150 -1742 3065 -1678
rect 3129 -1742 3149 -1678
rect -3150 -1758 3149 -1742
rect -3150 -1822 3065 -1758
rect 3129 -1822 3149 -1758
rect -3150 -1838 3149 -1822
rect -3150 -1902 3065 -1838
rect 3129 -1902 3149 -1838
rect -3150 -1918 3149 -1902
rect -3150 -1982 3065 -1918
rect 3129 -1982 3149 -1918
rect -3150 -1998 3149 -1982
rect -3150 -2062 3065 -1998
rect 3129 -2062 3149 -1998
rect -3150 -2078 3149 -2062
rect -3150 -2142 3065 -2078
rect 3129 -2142 3149 -2078
rect -3150 -2158 3149 -2142
rect -3150 -2222 3065 -2158
rect 3129 -2222 3149 -2158
rect -3150 -2238 3149 -2222
rect -3150 -2302 3065 -2238
rect 3129 -2302 3149 -2238
rect -3150 -2318 3149 -2302
rect -3150 -2382 3065 -2318
rect 3129 -2382 3149 -2318
rect -3150 -2398 3149 -2382
rect -3150 -2462 3065 -2398
rect 3129 -2462 3149 -2398
rect -3150 -2478 3149 -2462
rect -3150 -2542 3065 -2478
rect 3129 -2542 3149 -2478
rect -3150 -2558 3149 -2542
rect -3150 -2622 3065 -2558
rect 3129 -2622 3149 -2558
rect -3150 -2638 3149 -2622
rect -3150 -2702 3065 -2638
rect 3129 -2702 3149 -2638
rect -3150 -2718 3149 -2702
rect -3150 -2782 3065 -2718
rect 3129 -2782 3149 -2718
rect -3150 -2798 3149 -2782
rect -3150 -2862 3065 -2798
rect 3129 -2862 3149 -2798
rect -3150 -2878 3149 -2862
rect -3150 -2942 3065 -2878
rect 3129 -2942 3149 -2878
rect -3150 -2958 3149 -2942
rect -3150 -3022 3065 -2958
rect 3129 -3022 3149 -2958
rect -3150 -3038 3149 -3022
rect -3150 -3102 3065 -3038
rect 3129 -3102 3149 -3038
rect -3150 -3118 3149 -3102
rect -3150 -3182 3065 -3118
rect 3129 -3182 3149 -3118
rect -3150 -3198 3149 -3182
rect -3150 -3262 3065 -3198
rect 3129 -3262 3149 -3198
rect -3150 -3278 3149 -3262
rect -3150 -3342 3065 -3278
rect 3129 -3342 3149 -3278
rect -3150 -3358 3149 -3342
rect -3150 -3422 3065 -3358
rect 3129 -3422 3149 -3358
rect -3150 -3438 3149 -3422
rect -3150 -3502 3065 -3438
rect 3129 -3502 3149 -3438
rect -3150 -3518 3149 -3502
rect -3150 -3582 3065 -3518
rect 3129 -3582 3149 -3518
rect -3150 -3598 3149 -3582
rect -3150 -3662 3065 -3598
rect 3129 -3662 3149 -3598
rect -3150 -3678 3149 -3662
rect -3150 -3742 3065 -3678
rect 3129 -3742 3149 -3678
rect -3150 -3758 3149 -3742
rect -3150 -3822 3065 -3758
rect 3129 -3822 3149 -3758
rect -3150 -3838 3149 -3822
rect -3150 -3902 3065 -3838
rect 3129 -3902 3149 -3838
rect -3150 -3918 3149 -3902
rect -3150 -3982 3065 -3918
rect 3129 -3982 3149 -3918
rect -3150 -3998 3149 -3982
rect -3150 -4062 3065 -3998
rect 3129 -4062 3149 -3998
rect -3150 -4078 3149 -4062
rect -3150 -4142 3065 -4078
rect 3129 -4142 3149 -4078
rect -3150 -4158 3149 -4142
rect -3150 -4222 3065 -4158
rect 3129 -4222 3149 -4158
rect -3150 -4238 3149 -4222
rect -3150 -4302 3065 -4238
rect 3129 -4302 3149 -4238
rect -3150 -4318 3149 -4302
rect -3150 -4382 3065 -4318
rect 3129 -4382 3149 -4318
rect -3150 -4398 3149 -4382
rect -3150 -4462 3065 -4398
rect 3129 -4462 3149 -4398
rect -3150 -4478 3149 -4462
rect -3150 -4542 3065 -4478
rect 3129 -4542 3149 -4478
rect -3150 -4558 3149 -4542
rect -3150 -4622 3065 -4558
rect 3129 -4622 3149 -4558
rect -3150 -4638 3149 -4622
rect -3150 -4702 3065 -4638
rect 3129 -4702 3149 -4638
rect -3150 -4718 3149 -4702
rect -3150 -4782 3065 -4718
rect 3129 -4782 3149 -4718
rect -3150 -4798 3149 -4782
rect -3150 -4862 3065 -4798
rect 3129 -4862 3149 -4798
rect -3150 -4878 3149 -4862
rect -3150 -4942 3065 -4878
rect 3129 -4942 3149 -4878
rect -3150 -4958 3149 -4942
rect -3150 -5022 3065 -4958
rect 3129 -5022 3149 -4958
rect -3150 -5038 3149 -5022
rect -3150 -5102 3065 -5038
rect 3129 -5102 3149 -5038
rect -3150 -5118 3149 -5102
rect -3150 -5182 3065 -5118
rect 3129 -5182 3149 -5118
rect -3150 -5198 3149 -5182
rect -3150 -5262 3065 -5198
rect 3129 -5262 3149 -5198
rect -3150 -5278 3149 -5262
rect -3150 -5342 3065 -5278
rect 3129 -5342 3149 -5278
rect -3150 -5358 3149 -5342
rect -3150 -5422 3065 -5358
rect 3129 -5422 3149 -5358
rect -3150 -5438 3149 -5422
rect -3150 -5502 3065 -5438
rect 3129 -5502 3149 -5438
rect -3150 -5518 3149 -5502
rect -3150 -5582 3065 -5518
rect 3129 -5582 3149 -5518
rect -3150 -5598 3149 -5582
rect -3150 -5662 3065 -5598
rect 3129 -5662 3149 -5598
rect -3150 -5678 3149 -5662
rect -3150 -5742 3065 -5678
rect 3129 -5742 3149 -5678
rect -3150 -5758 3149 -5742
rect -3150 -5822 3065 -5758
rect 3129 -5822 3149 -5758
rect -3150 -5838 3149 -5822
rect -3150 -5902 3065 -5838
rect 3129 -5902 3149 -5838
rect -3150 -5918 3149 -5902
rect -3150 -5982 3065 -5918
rect 3129 -5982 3149 -5918
rect -3150 -5998 3149 -5982
rect -3150 -6062 3065 -5998
rect 3129 -6062 3149 -5998
rect -3150 -6078 3149 -6062
rect -3150 -6142 3065 -6078
rect 3129 -6142 3149 -6078
rect -3150 -6158 3149 -6142
rect -3150 -6222 3065 -6158
rect 3129 -6222 3149 -6158
rect -3150 -6250 3149 -6222
rect -3150 -6378 3149 -6350
rect -3150 -6442 3065 -6378
rect 3129 -6442 3149 -6378
rect -3150 -6458 3149 -6442
rect -3150 -6522 3065 -6458
rect 3129 -6522 3149 -6458
rect -3150 -6538 3149 -6522
rect -3150 -6602 3065 -6538
rect 3129 -6602 3149 -6538
rect -3150 -6618 3149 -6602
rect -3150 -6682 3065 -6618
rect 3129 -6682 3149 -6618
rect -3150 -6698 3149 -6682
rect -3150 -6762 3065 -6698
rect 3129 -6762 3149 -6698
rect -3150 -6778 3149 -6762
rect -3150 -6842 3065 -6778
rect 3129 -6842 3149 -6778
rect -3150 -6858 3149 -6842
rect -3150 -6922 3065 -6858
rect 3129 -6922 3149 -6858
rect -3150 -6938 3149 -6922
rect -3150 -7002 3065 -6938
rect 3129 -7002 3149 -6938
rect -3150 -7018 3149 -7002
rect -3150 -7082 3065 -7018
rect 3129 -7082 3149 -7018
rect -3150 -7098 3149 -7082
rect -3150 -7162 3065 -7098
rect 3129 -7162 3149 -7098
rect -3150 -7178 3149 -7162
rect -3150 -7242 3065 -7178
rect 3129 -7242 3149 -7178
rect -3150 -7258 3149 -7242
rect -3150 -7322 3065 -7258
rect 3129 -7322 3149 -7258
rect -3150 -7338 3149 -7322
rect -3150 -7402 3065 -7338
rect 3129 -7402 3149 -7338
rect -3150 -7418 3149 -7402
rect -3150 -7482 3065 -7418
rect 3129 -7482 3149 -7418
rect -3150 -7498 3149 -7482
rect -3150 -7562 3065 -7498
rect 3129 -7562 3149 -7498
rect -3150 -7578 3149 -7562
rect -3150 -7642 3065 -7578
rect 3129 -7642 3149 -7578
rect -3150 -7658 3149 -7642
rect -3150 -7722 3065 -7658
rect 3129 -7722 3149 -7658
rect -3150 -7738 3149 -7722
rect -3150 -7802 3065 -7738
rect 3129 -7802 3149 -7738
rect -3150 -7818 3149 -7802
rect -3150 -7882 3065 -7818
rect 3129 -7882 3149 -7818
rect -3150 -7898 3149 -7882
rect -3150 -7962 3065 -7898
rect 3129 -7962 3149 -7898
rect -3150 -7978 3149 -7962
rect -3150 -8042 3065 -7978
rect 3129 -8042 3149 -7978
rect -3150 -8058 3149 -8042
rect -3150 -8122 3065 -8058
rect 3129 -8122 3149 -8058
rect -3150 -8138 3149 -8122
rect -3150 -8202 3065 -8138
rect 3129 -8202 3149 -8138
rect -3150 -8218 3149 -8202
rect -3150 -8282 3065 -8218
rect 3129 -8282 3149 -8218
rect -3150 -8298 3149 -8282
rect -3150 -8362 3065 -8298
rect 3129 -8362 3149 -8298
rect -3150 -8378 3149 -8362
rect -3150 -8442 3065 -8378
rect 3129 -8442 3149 -8378
rect -3150 -8458 3149 -8442
rect -3150 -8522 3065 -8458
rect 3129 -8522 3149 -8458
rect -3150 -8538 3149 -8522
rect -3150 -8602 3065 -8538
rect 3129 -8602 3149 -8538
rect -3150 -8618 3149 -8602
rect -3150 -8682 3065 -8618
rect 3129 -8682 3149 -8618
rect -3150 -8698 3149 -8682
rect -3150 -8762 3065 -8698
rect 3129 -8762 3149 -8698
rect -3150 -8778 3149 -8762
rect -3150 -8842 3065 -8778
rect 3129 -8842 3149 -8778
rect -3150 -8858 3149 -8842
rect -3150 -8922 3065 -8858
rect 3129 -8922 3149 -8858
rect -3150 -8938 3149 -8922
rect -3150 -9002 3065 -8938
rect 3129 -9002 3149 -8938
rect -3150 -9018 3149 -9002
rect -3150 -9082 3065 -9018
rect 3129 -9082 3149 -9018
rect -3150 -9098 3149 -9082
rect -3150 -9162 3065 -9098
rect 3129 -9162 3149 -9098
rect -3150 -9178 3149 -9162
rect -3150 -9242 3065 -9178
rect 3129 -9242 3149 -9178
rect -3150 -9258 3149 -9242
rect -3150 -9322 3065 -9258
rect 3129 -9322 3149 -9258
rect -3150 -9338 3149 -9322
rect -3150 -9402 3065 -9338
rect 3129 -9402 3149 -9338
rect -3150 -9418 3149 -9402
rect -3150 -9482 3065 -9418
rect 3129 -9482 3149 -9418
rect -3150 -9498 3149 -9482
rect -3150 -9562 3065 -9498
rect 3129 -9562 3149 -9498
rect -3150 -9578 3149 -9562
rect -3150 -9642 3065 -9578
rect 3129 -9642 3149 -9578
rect -3150 -9658 3149 -9642
rect -3150 -9722 3065 -9658
rect 3129 -9722 3149 -9658
rect -3150 -9738 3149 -9722
rect -3150 -9802 3065 -9738
rect 3129 -9802 3149 -9738
rect -3150 -9818 3149 -9802
rect -3150 -9882 3065 -9818
rect 3129 -9882 3149 -9818
rect -3150 -9898 3149 -9882
rect -3150 -9962 3065 -9898
rect 3129 -9962 3149 -9898
rect -3150 -9978 3149 -9962
rect -3150 -10042 3065 -9978
rect 3129 -10042 3149 -9978
rect -3150 -10058 3149 -10042
rect -3150 -10122 3065 -10058
rect 3129 -10122 3149 -10058
rect -3150 -10138 3149 -10122
rect -3150 -10202 3065 -10138
rect 3129 -10202 3149 -10138
rect -3150 -10218 3149 -10202
rect -3150 -10282 3065 -10218
rect 3129 -10282 3149 -10218
rect -3150 -10298 3149 -10282
rect -3150 -10362 3065 -10298
rect 3129 -10362 3149 -10298
rect -3150 -10378 3149 -10362
rect -3150 -10442 3065 -10378
rect 3129 -10442 3149 -10378
rect -3150 -10458 3149 -10442
rect -3150 -10522 3065 -10458
rect 3129 -10522 3149 -10458
rect -3150 -10538 3149 -10522
rect -3150 -10602 3065 -10538
rect 3129 -10602 3149 -10538
rect -3150 -10618 3149 -10602
rect -3150 -10682 3065 -10618
rect 3129 -10682 3149 -10618
rect -3150 -10698 3149 -10682
rect -3150 -10762 3065 -10698
rect 3129 -10762 3149 -10698
rect -3150 -10778 3149 -10762
rect -3150 -10842 3065 -10778
rect 3129 -10842 3149 -10778
rect -3150 -10858 3149 -10842
rect -3150 -10922 3065 -10858
rect 3129 -10922 3149 -10858
rect -3150 -10938 3149 -10922
rect -3150 -11002 3065 -10938
rect 3129 -11002 3149 -10938
rect -3150 -11018 3149 -11002
rect -3150 -11082 3065 -11018
rect 3129 -11082 3149 -11018
rect -3150 -11098 3149 -11082
rect -3150 -11162 3065 -11098
rect 3129 -11162 3149 -11098
rect -3150 -11178 3149 -11162
rect -3150 -11242 3065 -11178
rect 3129 -11242 3149 -11178
rect -3150 -11258 3149 -11242
rect -3150 -11322 3065 -11258
rect 3129 -11322 3149 -11258
rect -3150 -11338 3149 -11322
rect -3150 -11402 3065 -11338
rect 3129 -11402 3149 -11338
rect -3150 -11418 3149 -11402
rect -3150 -11482 3065 -11418
rect 3129 -11482 3149 -11418
rect -3150 -11498 3149 -11482
rect -3150 -11562 3065 -11498
rect 3129 -11562 3149 -11498
rect -3150 -11578 3149 -11562
rect -3150 -11642 3065 -11578
rect 3129 -11642 3149 -11578
rect -3150 -11658 3149 -11642
rect -3150 -11722 3065 -11658
rect 3129 -11722 3149 -11658
rect -3150 -11738 3149 -11722
rect -3150 -11802 3065 -11738
rect 3129 -11802 3149 -11738
rect -3150 -11818 3149 -11802
rect -3150 -11882 3065 -11818
rect 3129 -11882 3149 -11818
rect -3150 -11898 3149 -11882
rect -3150 -11962 3065 -11898
rect 3129 -11962 3149 -11898
rect -3150 -11978 3149 -11962
rect -3150 -12042 3065 -11978
rect 3129 -12042 3149 -11978
rect -3150 -12058 3149 -12042
rect -3150 -12122 3065 -12058
rect 3129 -12122 3149 -12058
rect -3150 -12138 3149 -12122
rect -3150 -12202 3065 -12138
rect 3129 -12202 3149 -12138
rect -3150 -12218 3149 -12202
rect -3150 -12282 3065 -12218
rect 3129 -12282 3149 -12218
rect -3150 -12298 3149 -12282
rect -3150 -12362 3065 -12298
rect 3129 -12362 3149 -12298
rect -3150 -12378 3149 -12362
rect -3150 -12442 3065 -12378
rect 3129 -12442 3149 -12378
rect -3150 -12458 3149 -12442
rect -3150 -12522 3065 -12458
rect 3129 -12522 3149 -12458
rect -3150 -12550 3149 -12522
<< via3 >>
rect 3065 12458 3129 12522
rect 3065 12378 3129 12442
rect 3065 12298 3129 12362
rect 3065 12218 3129 12282
rect 3065 12138 3129 12202
rect 3065 12058 3129 12122
rect 3065 11978 3129 12042
rect 3065 11898 3129 11962
rect 3065 11818 3129 11882
rect 3065 11738 3129 11802
rect 3065 11658 3129 11722
rect 3065 11578 3129 11642
rect 3065 11498 3129 11562
rect 3065 11418 3129 11482
rect 3065 11338 3129 11402
rect 3065 11258 3129 11322
rect 3065 11178 3129 11242
rect 3065 11098 3129 11162
rect 3065 11018 3129 11082
rect 3065 10938 3129 11002
rect 3065 10858 3129 10922
rect 3065 10778 3129 10842
rect 3065 10698 3129 10762
rect 3065 10618 3129 10682
rect 3065 10538 3129 10602
rect 3065 10458 3129 10522
rect 3065 10378 3129 10442
rect 3065 10298 3129 10362
rect 3065 10218 3129 10282
rect 3065 10138 3129 10202
rect 3065 10058 3129 10122
rect 3065 9978 3129 10042
rect 3065 9898 3129 9962
rect 3065 9818 3129 9882
rect 3065 9738 3129 9802
rect 3065 9658 3129 9722
rect 3065 9578 3129 9642
rect 3065 9498 3129 9562
rect 3065 9418 3129 9482
rect 3065 9338 3129 9402
rect 3065 9258 3129 9322
rect 3065 9178 3129 9242
rect 3065 9098 3129 9162
rect 3065 9018 3129 9082
rect 3065 8938 3129 9002
rect 3065 8858 3129 8922
rect 3065 8778 3129 8842
rect 3065 8698 3129 8762
rect 3065 8618 3129 8682
rect 3065 8538 3129 8602
rect 3065 8458 3129 8522
rect 3065 8378 3129 8442
rect 3065 8298 3129 8362
rect 3065 8218 3129 8282
rect 3065 8138 3129 8202
rect 3065 8058 3129 8122
rect 3065 7978 3129 8042
rect 3065 7898 3129 7962
rect 3065 7818 3129 7882
rect 3065 7738 3129 7802
rect 3065 7658 3129 7722
rect 3065 7578 3129 7642
rect 3065 7498 3129 7562
rect 3065 7418 3129 7482
rect 3065 7338 3129 7402
rect 3065 7258 3129 7322
rect 3065 7178 3129 7242
rect 3065 7098 3129 7162
rect 3065 7018 3129 7082
rect 3065 6938 3129 7002
rect 3065 6858 3129 6922
rect 3065 6778 3129 6842
rect 3065 6698 3129 6762
rect 3065 6618 3129 6682
rect 3065 6538 3129 6602
rect 3065 6458 3129 6522
rect 3065 6378 3129 6442
rect 3065 6158 3129 6222
rect 3065 6078 3129 6142
rect 3065 5998 3129 6062
rect 3065 5918 3129 5982
rect 3065 5838 3129 5902
rect 3065 5758 3129 5822
rect 3065 5678 3129 5742
rect 3065 5598 3129 5662
rect 3065 5518 3129 5582
rect 3065 5438 3129 5502
rect 3065 5358 3129 5422
rect 3065 5278 3129 5342
rect 3065 5198 3129 5262
rect 3065 5118 3129 5182
rect 3065 5038 3129 5102
rect 3065 4958 3129 5022
rect 3065 4878 3129 4942
rect 3065 4798 3129 4862
rect 3065 4718 3129 4782
rect 3065 4638 3129 4702
rect 3065 4558 3129 4622
rect 3065 4478 3129 4542
rect 3065 4398 3129 4462
rect 3065 4318 3129 4382
rect 3065 4238 3129 4302
rect 3065 4158 3129 4222
rect 3065 4078 3129 4142
rect 3065 3998 3129 4062
rect 3065 3918 3129 3982
rect 3065 3838 3129 3902
rect 3065 3758 3129 3822
rect 3065 3678 3129 3742
rect 3065 3598 3129 3662
rect 3065 3518 3129 3582
rect 3065 3438 3129 3502
rect 3065 3358 3129 3422
rect 3065 3278 3129 3342
rect 3065 3198 3129 3262
rect 3065 3118 3129 3182
rect 3065 3038 3129 3102
rect 3065 2958 3129 3022
rect 3065 2878 3129 2942
rect 3065 2798 3129 2862
rect 3065 2718 3129 2782
rect 3065 2638 3129 2702
rect 3065 2558 3129 2622
rect 3065 2478 3129 2542
rect 3065 2398 3129 2462
rect 3065 2318 3129 2382
rect 3065 2238 3129 2302
rect 3065 2158 3129 2222
rect 3065 2078 3129 2142
rect 3065 1998 3129 2062
rect 3065 1918 3129 1982
rect 3065 1838 3129 1902
rect 3065 1758 3129 1822
rect 3065 1678 3129 1742
rect 3065 1598 3129 1662
rect 3065 1518 3129 1582
rect 3065 1438 3129 1502
rect 3065 1358 3129 1422
rect 3065 1278 3129 1342
rect 3065 1198 3129 1262
rect 3065 1118 3129 1182
rect 3065 1038 3129 1102
rect 3065 958 3129 1022
rect 3065 878 3129 942
rect 3065 798 3129 862
rect 3065 718 3129 782
rect 3065 638 3129 702
rect 3065 558 3129 622
rect 3065 478 3129 542
rect 3065 398 3129 462
rect 3065 318 3129 382
rect 3065 238 3129 302
rect 3065 158 3129 222
rect 3065 78 3129 142
rect 3065 -142 3129 -78
rect 3065 -222 3129 -158
rect 3065 -302 3129 -238
rect 3065 -382 3129 -318
rect 3065 -462 3129 -398
rect 3065 -542 3129 -478
rect 3065 -622 3129 -558
rect 3065 -702 3129 -638
rect 3065 -782 3129 -718
rect 3065 -862 3129 -798
rect 3065 -942 3129 -878
rect 3065 -1022 3129 -958
rect 3065 -1102 3129 -1038
rect 3065 -1182 3129 -1118
rect 3065 -1262 3129 -1198
rect 3065 -1342 3129 -1278
rect 3065 -1422 3129 -1358
rect 3065 -1502 3129 -1438
rect 3065 -1582 3129 -1518
rect 3065 -1662 3129 -1598
rect 3065 -1742 3129 -1678
rect 3065 -1822 3129 -1758
rect 3065 -1902 3129 -1838
rect 3065 -1982 3129 -1918
rect 3065 -2062 3129 -1998
rect 3065 -2142 3129 -2078
rect 3065 -2222 3129 -2158
rect 3065 -2302 3129 -2238
rect 3065 -2382 3129 -2318
rect 3065 -2462 3129 -2398
rect 3065 -2542 3129 -2478
rect 3065 -2622 3129 -2558
rect 3065 -2702 3129 -2638
rect 3065 -2782 3129 -2718
rect 3065 -2862 3129 -2798
rect 3065 -2942 3129 -2878
rect 3065 -3022 3129 -2958
rect 3065 -3102 3129 -3038
rect 3065 -3182 3129 -3118
rect 3065 -3262 3129 -3198
rect 3065 -3342 3129 -3278
rect 3065 -3422 3129 -3358
rect 3065 -3502 3129 -3438
rect 3065 -3582 3129 -3518
rect 3065 -3662 3129 -3598
rect 3065 -3742 3129 -3678
rect 3065 -3822 3129 -3758
rect 3065 -3902 3129 -3838
rect 3065 -3982 3129 -3918
rect 3065 -4062 3129 -3998
rect 3065 -4142 3129 -4078
rect 3065 -4222 3129 -4158
rect 3065 -4302 3129 -4238
rect 3065 -4382 3129 -4318
rect 3065 -4462 3129 -4398
rect 3065 -4542 3129 -4478
rect 3065 -4622 3129 -4558
rect 3065 -4702 3129 -4638
rect 3065 -4782 3129 -4718
rect 3065 -4862 3129 -4798
rect 3065 -4942 3129 -4878
rect 3065 -5022 3129 -4958
rect 3065 -5102 3129 -5038
rect 3065 -5182 3129 -5118
rect 3065 -5262 3129 -5198
rect 3065 -5342 3129 -5278
rect 3065 -5422 3129 -5358
rect 3065 -5502 3129 -5438
rect 3065 -5582 3129 -5518
rect 3065 -5662 3129 -5598
rect 3065 -5742 3129 -5678
rect 3065 -5822 3129 -5758
rect 3065 -5902 3129 -5838
rect 3065 -5982 3129 -5918
rect 3065 -6062 3129 -5998
rect 3065 -6142 3129 -6078
rect 3065 -6222 3129 -6158
rect 3065 -6442 3129 -6378
rect 3065 -6522 3129 -6458
rect 3065 -6602 3129 -6538
rect 3065 -6682 3129 -6618
rect 3065 -6762 3129 -6698
rect 3065 -6842 3129 -6778
rect 3065 -6922 3129 -6858
rect 3065 -7002 3129 -6938
rect 3065 -7082 3129 -7018
rect 3065 -7162 3129 -7098
rect 3065 -7242 3129 -7178
rect 3065 -7322 3129 -7258
rect 3065 -7402 3129 -7338
rect 3065 -7482 3129 -7418
rect 3065 -7562 3129 -7498
rect 3065 -7642 3129 -7578
rect 3065 -7722 3129 -7658
rect 3065 -7802 3129 -7738
rect 3065 -7882 3129 -7818
rect 3065 -7962 3129 -7898
rect 3065 -8042 3129 -7978
rect 3065 -8122 3129 -8058
rect 3065 -8202 3129 -8138
rect 3065 -8282 3129 -8218
rect 3065 -8362 3129 -8298
rect 3065 -8442 3129 -8378
rect 3065 -8522 3129 -8458
rect 3065 -8602 3129 -8538
rect 3065 -8682 3129 -8618
rect 3065 -8762 3129 -8698
rect 3065 -8842 3129 -8778
rect 3065 -8922 3129 -8858
rect 3065 -9002 3129 -8938
rect 3065 -9082 3129 -9018
rect 3065 -9162 3129 -9098
rect 3065 -9242 3129 -9178
rect 3065 -9322 3129 -9258
rect 3065 -9402 3129 -9338
rect 3065 -9482 3129 -9418
rect 3065 -9562 3129 -9498
rect 3065 -9642 3129 -9578
rect 3065 -9722 3129 -9658
rect 3065 -9802 3129 -9738
rect 3065 -9882 3129 -9818
rect 3065 -9962 3129 -9898
rect 3065 -10042 3129 -9978
rect 3065 -10122 3129 -10058
rect 3065 -10202 3129 -10138
rect 3065 -10282 3129 -10218
rect 3065 -10362 3129 -10298
rect 3065 -10442 3129 -10378
rect 3065 -10522 3129 -10458
rect 3065 -10602 3129 -10538
rect 3065 -10682 3129 -10618
rect 3065 -10762 3129 -10698
rect 3065 -10842 3129 -10778
rect 3065 -10922 3129 -10858
rect 3065 -11002 3129 -10938
rect 3065 -11082 3129 -11018
rect 3065 -11162 3129 -11098
rect 3065 -11242 3129 -11178
rect 3065 -11322 3129 -11258
rect 3065 -11402 3129 -11338
rect 3065 -11482 3129 -11418
rect 3065 -11562 3129 -11498
rect 3065 -11642 3129 -11578
rect 3065 -11722 3129 -11658
rect 3065 -11802 3129 -11738
rect 3065 -11882 3129 -11818
rect 3065 -11962 3129 -11898
rect 3065 -12042 3129 -11978
rect 3065 -12122 3129 -12058
rect 3065 -12202 3129 -12138
rect 3065 -12282 3129 -12218
rect 3065 -12362 3129 -12298
rect 3065 -12442 3129 -12378
rect 3065 -12522 3129 -12458
<< mimcap >>
rect -3050 12402 2950 12450
rect -3050 6498 -3002 12402
rect 2902 6498 2950 12402
rect -3050 6450 2950 6498
rect -3050 6102 2950 6150
rect -3050 198 -3002 6102
rect 2902 198 2950 6102
rect -3050 150 2950 198
rect -3050 -198 2950 -150
rect -3050 -6102 -3002 -198
rect 2902 -6102 2950 -198
rect -3050 -6150 2950 -6102
rect -3050 -6498 2950 -6450
rect -3050 -12402 -3002 -6498
rect 2902 -12402 2950 -6498
rect -3050 -12450 2950 -12402
<< mimcapcontact >>
rect -3002 6498 2902 12402
rect -3002 198 2902 6102
rect -3002 -6102 2902 -198
rect -3002 -12402 2902 -6498
<< metal4 >>
rect -102 12411 2 12600
rect 3018 12538 3122 12600
rect 3018 12522 3145 12538
rect 3018 12458 3065 12522
rect 3129 12458 3145 12522
rect 3018 12442 3145 12458
rect -3011 12402 2911 12411
rect -3011 6498 -3002 12402
rect 2902 6498 2911 12402
rect -3011 6489 2911 6498
rect 3018 12378 3065 12442
rect 3129 12378 3145 12442
rect 3018 12362 3145 12378
rect 3018 12298 3065 12362
rect 3129 12298 3145 12362
rect 3018 12282 3145 12298
rect 3018 12218 3065 12282
rect 3129 12218 3145 12282
rect 3018 12202 3145 12218
rect 3018 12138 3065 12202
rect 3129 12138 3145 12202
rect 3018 12122 3145 12138
rect 3018 12058 3065 12122
rect 3129 12058 3145 12122
rect 3018 12042 3145 12058
rect 3018 11978 3065 12042
rect 3129 11978 3145 12042
rect 3018 11962 3145 11978
rect 3018 11898 3065 11962
rect 3129 11898 3145 11962
rect 3018 11882 3145 11898
rect 3018 11818 3065 11882
rect 3129 11818 3145 11882
rect 3018 11802 3145 11818
rect 3018 11738 3065 11802
rect 3129 11738 3145 11802
rect 3018 11722 3145 11738
rect 3018 11658 3065 11722
rect 3129 11658 3145 11722
rect 3018 11642 3145 11658
rect 3018 11578 3065 11642
rect 3129 11578 3145 11642
rect 3018 11562 3145 11578
rect 3018 11498 3065 11562
rect 3129 11498 3145 11562
rect 3018 11482 3145 11498
rect 3018 11418 3065 11482
rect 3129 11418 3145 11482
rect 3018 11402 3145 11418
rect 3018 11338 3065 11402
rect 3129 11338 3145 11402
rect 3018 11322 3145 11338
rect 3018 11258 3065 11322
rect 3129 11258 3145 11322
rect 3018 11242 3145 11258
rect 3018 11178 3065 11242
rect 3129 11178 3145 11242
rect 3018 11162 3145 11178
rect 3018 11098 3065 11162
rect 3129 11098 3145 11162
rect 3018 11082 3145 11098
rect 3018 11018 3065 11082
rect 3129 11018 3145 11082
rect 3018 11002 3145 11018
rect 3018 10938 3065 11002
rect 3129 10938 3145 11002
rect 3018 10922 3145 10938
rect 3018 10858 3065 10922
rect 3129 10858 3145 10922
rect 3018 10842 3145 10858
rect 3018 10778 3065 10842
rect 3129 10778 3145 10842
rect 3018 10762 3145 10778
rect 3018 10698 3065 10762
rect 3129 10698 3145 10762
rect 3018 10682 3145 10698
rect 3018 10618 3065 10682
rect 3129 10618 3145 10682
rect 3018 10602 3145 10618
rect 3018 10538 3065 10602
rect 3129 10538 3145 10602
rect 3018 10522 3145 10538
rect 3018 10458 3065 10522
rect 3129 10458 3145 10522
rect 3018 10442 3145 10458
rect 3018 10378 3065 10442
rect 3129 10378 3145 10442
rect 3018 10362 3145 10378
rect 3018 10298 3065 10362
rect 3129 10298 3145 10362
rect 3018 10282 3145 10298
rect 3018 10218 3065 10282
rect 3129 10218 3145 10282
rect 3018 10202 3145 10218
rect 3018 10138 3065 10202
rect 3129 10138 3145 10202
rect 3018 10122 3145 10138
rect 3018 10058 3065 10122
rect 3129 10058 3145 10122
rect 3018 10042 3145 10058
rect 3018 9978 3065 10042
rect 3129 9978 3145 10042
rect 3018 9962 3145 9978
rect 3018 9898 3065 9962
rect 3129 9898 3145 9962
rect 3018 9882 3145 9898
rect 3018 9818 3065 9882
rect 3129 9818 3145 9882
rect 3018 9802 3145 9818
rect 3018 9738 3065 9802
rect 3129 9738 3145 9802
rect 3018 9722 3145 9738
rect 3018 9658 3065 9722
rect 3129 9658 3145 9722
rect 3018 9642 3145 9658
rect 3018 9578 3065 9642
rect 3129 9578 3145 9642
rect 3018 9562 3145 9578
rect 3018 9498 3065 9562
rect 3129 9498 3145 9562
rect 3018 9482 3145 9498
rect 3018 9418 3065 9482
rect 3129 9418 3145 9482
rect 3018 9402 3145 9418
rect 3018 9338 3065 9402
rect 3129 9338 3145 9402
rect 3018 9322 3145 9338
rect 3018 9258 3065 9322
rect 3129 9258 3145 9322
rect 3018 9242 3145 9258
rect 3018 9178 3065 9242
rect 3129 9178 3145 9242
rect 3018 9162 3145 9178
rect 3018 9098 3065 9162
rect 3129 9098 3145 9162
rect 3018 9082 3145 9098
rect 3018 9018 3065 9082
rect 3129 9018 3145 9082
rect 3018 9002 3145 9018
rect 3018 8938 3065 9002
rect 3129 8938 3145 9002
rect 3018 8922 3145 8938
rect 3018 8858 3065 8922
rect 3129 8858 3145 8922
rect 3018 8842 3145 8858
rect 3018 8778 3065 8842
rect 3129 8778 3145 8842
rect 3018 8762 3145 8778
rect 3018 8698 3065 8762
rect 3129 8698 3145 8762
rect 3018 8682 3145 8698
rect 3018 8618 3065 8682
rect 3129 8618 3145 8682
rect 3018 8602 3145 8618
rect 3018 8538 3065 8602
rect 3129 8538 3145 8602
rect 3018 8522 3145 8538
rect 3018 8458 3065 8522
rect 3129 8458 3145 8522
rect 3018 8442 3145 8458
rect 3018 8378 3065 8442
rect 3129 8378 3145 8442
rect 3018 8362 3145 8378
rect 3018 8298 3065 8362
rect 3129 8298 3145 8362
rect 3018 8282 3145 8298
rect 3018 8218 3065 8282
rect 3129 8218 3145 8282
rect 3018 8202 3145 8218
rect 3018 8138 3065 8202
rect 3129 8138 3145 8202
rect 3018 8122 3145 8138
rect 3018 8058 3065 8122
rect 3129 8058 3145 8122
rect 3018 8042 3145 8058
rect 3018 7978 3065 8042
rect 3129 7978 3145 8042
rect 3018 7962 3145 7978
rect 3018 7898 3065 7962
rect 3129 7898 3145 7962
rect 3018 7882 3145 7898
rect 3018 7818 3065 7882
rect 3129 7818 3145 7882
rect 3018 7802 3145 7818
rect 3018 7738 3065 7802
rect 3129 7738 3145 7802
rect 3018 7722 3145 7738
rect 3018 7658 3065 7722
rect 3129 7658 3145 7722
rect 3018 7642 3145 7658
rect 3018 7578 3065 7642
rect 3129 7578 3145 7642
rect 3018 7562 3145 7578
rect 3018 7498 3065 7562
rect 3129 7498 3145 7562
rect 3018 7482 3145 7498
rect 3018 7418 3065 7482
rect 3129 7418 3145 7482
rect 3018 7402 3145 7418
rect 3018 7338 3065 7402
rect 3129 7338 3145 7402
rect 3018 7322 3145 7338
rect 3018 7258 3065 7322
rect 3129 7258 3145 7322
rect 3018 7242 3145 7258
rect 3018 7178 3065 7242
rect 3129 7178 3145 7242
rect 3018 7162 3145 7178
rect 3018 7098 3065 7162
rect 3129 7098 3145 7162
rect 3018 7082 3145 7098
rect 3018 7018 3065 7082
rect 3129 7018 3145 7082
rect 3018 7002 3145 7018
rect 3018 6938 3065 7002
rect 3129 6938 3145 7002
rect 3018 6922 3145 6938
rect 3018 6858 3065 6922
rect 3129 6858 3145 6922
rect 3018 6842 3145 6858
rect 3018 6778 3065 6842
rect 3129 6778 3145 6842
rect 3018 6762 3145 6778
rect 3018 6698 3065 6762
rect 3129 6698 3145 6762
rect 3018 6682 3145 6698
rect 3018 6618 3065 6682
rect 3129 6618 3145 6682
rect 3018 6602 3145 6618
rect 3018 6538 3065 6602
rect 3129 6538 3145 6602
rect 3018 6522 3145 6538
rect -102 6111 2 6489
rect 3018 6458 3065 6522
rect 3129 6458 3145 6522
rect 3018 6442 3145 6458
rect 3018 6378 3065 6442
rect 3129 6378 3145 6442
rect 3018 6362 3145 6378
rect 3018 6238 3122 6362
rect 3018 6222 3145 6238
rect 3018 6158 3065 6222
rect 3129 6158 3145 6222
rect 3018 6142 3145 6158
rect -3011 6102 2911 6111
rect -3011 198 -3002 6102
rect 2902 198 2911 6102
rect -3011 189 2911 198
rect 3018 6078 3065 6142
rect 3129 6078 3145 6142
rect 3018 6062 3145 6078
rect 3018 5998 3065 6062
rect 3129 5998 3145 6062
rect 3018 5982 3145 5998
rect 3018 5918 3065 5982
rect 3129 5918 3145 5982
rect 3018 5902 3145 5918
rect 3018 5838 3065 5902
rect 3129 5838 3145 5902
rect 3018 5822 3145 5838
rect 3018 5758 3065 5822
rect 3129 5758 3145 5822
rect 3018 5742 3145 5758
rect 3018 5678 3065 5742
rect 3129 5678 3145 5742
rect 3018 5662 3145 5678
rect 3018 5598 3065 5662
rect 3129 5598 3145 5662
rect 3018 5582 3145 5598
rect 3018 5518 3065 5582
rect 3129 5518 3145 5582
rect 3018 5502 3145 5518
rect 3018 5438 3065 5502
rect 3129 5438 3145 5502
rect 3018 5422 3145 5438
rect 3018 5358 3065 5422
rect 3129 5358 3145 5422
rect 3018 5342 3145 5358
rect 3018 5278 3065 5342
rect 3129 5278 3145 5342
rect 3018 5262 3145 5278
rect 3018 5198 3065 5262
rect 3129 5198 3145 5262
rect 3018 5182 3145 5198
rect 3018 5118 3065 5182
rect 3129 5118 3145 5182
rect 3018 5102 3145 5118
rect 3018 5038 3065 5102
rect 3129 5038 3145 5102
rect 3018 5022 3145 5038
rect 3018 4958 3065 5022
rect 3129 4958 3145 5022
rect 3018 4942 3145 4958
rect 3018 4878 3065 4942
rect 3129 4878 3145 4942
rect 3018 4862 3145 4878
rect 3018 4798 3065 4862
rect 3129 4798 3145 4862
rect 3018 4782 3145 4798
rect 3018 4718 3065 4782
rect 3129 4718 3145 4782
rect 3018 4702 3145 4718
rect 3018 4638 3065 4702
rect 3129 4638 3145 4702
rect 3018 4622 3145 4638
rect 3018 4558 3065 4622
rect 3129 4558 3145 4622
rect 3018 4542 3145 4558
rect 3018 4478 3065 4542
rect 3129 4478 3145 4542
rect 3018 4462 3145 4478
rect 3018 4398 3065 4462
rect 3129 4398 3145 4462
rect 3018 4382 3145 4398
rect 3018 4318 3065 4382
rect 3129 4318 3145 4382
rect 3018 4302 3145 4318
rect 3018 4238 3065 4302
rect 3129 4238 3145 4302
rect 3018 4222 3145 4238
rect 3018 4158 3065 4222
rect 3129 4158 3145 4222
rect 3018 4142 3145 4158
rect 3018 4078 3065 4142
rect 3129 4078 3145 4142
rect 3018 4062 3145 4078
rect 3018 3998 3065 4062
rect 3129 3998 3145 4062
rect 3018 3982 3145 3998
rect 3018 3918 3065 3982
rect 3129 3918 3145 3982
rect 3018 3902 3145 3918
rect 3018 3838 3065 3902
rect 3129 3838 3145 3902
rect 3018 3822 3145 3838
rect 3018 3758 3065 3822
rect 3129 3758 3145 3822
rect 3018 3742 3145 3758
rect 3018 3678 3065 3742
rect 3129 3678 3145 3742
rect 3018 3662 3145 3678
rect 3018 3598 3065 3662
rect 3129 3598 3145 3662
rect 3018 3582 3145 3598
rect 3018 3518 3065 3582
rect 3129 3518 3145 3582
rect 3018 3502 3145 3518
rect 3018 3438 3065 3502
rect 3129 3438 3145 3502
rect 3018 3422 3145 3438
rect 3018 3358 3065 3422
rect 3129 3358 3145 3422
rect 3018 3342 3145 3358
rect 3018 3278 3065 3342
rect 3129 3278 3145 3342
rect 3018 3262 3145 3278
rect 3018 3198 3065 3262
rect 3129 3198 3145 3262
rect 3018 3182 3145 3198
rect 3018 3118 3065 3182
rect 3129 3118 3145 3182
rect 3018 3102 3145 3118
rect 3018 3038 3065 3102
rect 3129 3038 3145 3102
rect 3018 3022 3145 3038
rect 3018 2958 3065 3022
rect 3129 2958 3145 3022
rect 3018 2942 3145 2958
rect 3018 2878 3065 2942
rect 3129 2878 3145 2942
rect 3018 2862 3145 2878
rect 3018 2798 3065 2862
rect 3129 2798 3145 2862
rect 3018 2782 3145 2798
rect 3018 2718 3065 2782
rect 3129 2718 3145 2782
rect 3018 2702 3145 2718
rect 3018 2638 3065 2702
rect 3129 2638 3145 2702
rect 3018 2622 3145 2638
rect 3018 2558 3065 2622
rect 3129 2558 3145 2622
rect 3018 2542 3145 2558
rect 3018 2478 3065 2542
rect 3129 2478 3145 2542
rect 3018 2462 3145 2478
rect 3018 2398 3065 2462
rect 3129 2398 3145 2462
rect 3018 2382 3145 2398
rect 3018 2318 3065 2382
rect 3129 2318 3145 2382
rect 3018 2302 3145 2318
rect 3018 2238 3065 2302
rect 3129 2238 3145 2302
rect 3018 2222 3145 2238
rect 3018 2158 3065 2222
rect 3129 2158 3145 2222
rect 3018 2142 3145 2158
rect 3018 2078 3065 2142
rect 3129 2078 3145 2142
rect 3018 2062 3145 2078
rect 3018 1998 3065 2062
rect 3129 1998 3145 2062
rect 3018 1982 3145 1998
rect 3018 1918 3065 1982
rect 3129 1918 3145 1982
rect 3018 1902 3145 1918
rect 3018 1838 3065 1902
rect 3129 1838 3145 1902
rect 3018 1822 3145 1838
rect 3018 1758 3065 1822
rect 3129 1758 3145 1822
rect 3018 1742 3145 1758
rect 3018 1678 3065 1742
rect 3129 1678 3145 1742
rect 3018 1662 3145 1678
rect 3018 1598 3065 1662
rect 3129 1598 3145 1662
rect 3018 1582 3145 1598
rect 3018 1518 3065 1582
rect 3129 1518 3145 1582
rect 3018 1502 3145 1518
rect 3018 1438 3065 1502
rect 3129 1438 3145 1502
rect 3018 1422 3145 1438
rect 3018 1358 3065 1422
rect 3129 1358 3145 1422
rect 3018 1342 3145 1358
rect 3018 1278 3065 1342
rect 3129 1278 3145 1342
rect 3018 1262 3145 1278
rect 3018 1198 3065 1262
rect 3129 1198 3145 1262
rect 3018 1182 3145 1198
rect 3018 1118 3065 1182
rect 3129 1118 3145 1182
rect 3018 1102 3145 1118
rect 3018 1038 3065 1102
rect 3129 1038 3145 1102
rect 3018 1022 3145 1038
rect 3018 958 3065 1022
rect 3129 958 3145 1022
rect 3018 942 3145 958
rect 3018 878 3065 942
rect 3129 878 3145 942
rect 3018 862 3145 878
rect 3018 798 3065 862
rect 3129 798 3145 862
rect 3018 782 3145 798
rect 3018 718 3065 782
rect 3129 718 3145 782
rect 3018 702 3145 718
rect 3018 638 3065 702
rect 3129 638 3145 702
rect 3018 622 3145 638
rect 3018 558 3065 622
rect 3129 558 3145 622
rect 3018 542 3145 558
rect 3018 478 3065 542
rect 3129 478 3145 542
rect 3018 462 3145 478
rect 3018 398 3065 462
rect 3129 398 3145 462
rect 3018 382 3145 398
rect 3018 318 3065 382
rect 3129 318 3145 382
rect 3018 302 3145 318
rect 3018 238 3065 302
rect 3129 238 3145 302
rect 3018 222 3145 238
rect -102 -189 2 189
rect 3018 158 3065 222
rect 3129 158 3145 222
rect 3018 142 3145 158
rect 3018 78 3065 142
rect 3129 78 3145 142
rect 3018 62 3145 78
rect 3018 -62 3122 62
rect 3018 -78 3145 -62
rect 3018 -142 3065 -78
rect 3129 -142 3145 -78
rect 3018 -158 3145 -142
rect -3011 -198 2911 -189
rect -3011 -6102 -3002 -198
rect 2902 -6102 2911 -198
rect -3011 -6111 2911 -6102
rect 3018 -222 3065 -158
rect 3129 -222 3145 -158
rect 3018 -238 3145 -222
rect 3018 -302 3065 -238
rect 3129 -302 3145 -238
rect 3018 -318 3145 -302
rect 3018 -382 3065 -318
rect 3129 -382 3145 -318
rect 3018 -398 3145 -382
rect 3018 -462 3065 -398
rect 3129 -462 3145 -398
rect 3018 -478 3145 -462
rect 3018 -542 3065 -478
rect 3129 -542 3145 -478
rect 3018 -558 3145 -542
rect 3018 -622 3065 -558
rect 3129 -622 3145 -558
rect 3018 -638 3145 -622
rect 3018 -702 3065 -638
rect 3129 -702 3145 -638
rect 3018 -718 3145 -702
rect 3018 -782 3065 -718
rect 3129 -782 3145 -718
rect 3018 -798 3145 -782
rect 3018 -862 3065 -798
rect 3129 -862 3145 -798
rect 3018 -878 3145 -862
rect 3018 -942 3065 -878
rect 3129 -942 3145 -878
rect 3018 -958 3145 -942
rect 3018 -1022 3065 -958
rect 3129 -1022 3145 -958
rect 3018 -1038 3145 -1022
rect 3018 -1102 3065 -1038
rect 3129 -1102 3145 -1038
rect 3018 -1118 3145 -1102
rect 3018 -1182 3065 -1118
rect 3129 -1182 3145 -1118
rect 3018 -1198 3145 -1182
rect 3018 -1262 3065 -1198
rect 3129 -1262 3145 -1198
rect 3018 -1278 3145 -1262
rect 3018 -1342 3065 -1278
rect 3129 -1342 3145 -1278
rect 3018 -1358 3145 -1342
rect 3018 -1422 3065 -1358
rect 3129 -1422 3145 -1358
rect 3018 -1438 3145 -1422
rect 3018 -1502 3065 -1438
rect 3129 -1502 3145 -1438
rect 3018 -1518 3145 -1502
rect 3018 -1582 3065 -1518
rect 3129 -1582 3145 -1518
rect 3018 -1598 3145 -1582
rect 3018 -1662 3065 -1598
rect 3129 -1662 3145 -1598
rect 3018 -1678 3145 -1662
rect 3018 -1742 3065 -1678
rect 3129 -1742 3145 -1678
rect 3018 -1758 3145 -1742
rect 3018 -1822 3065 -1758
rect 3129 -1822 3145 -1758
rect 3018 -1838 3145 -1822
rect 3018 -1902 3065 -1838
rect 3129 -1902 3145 -1838
rect 3018 -1918 3145 -1902
rect 3018 -1982 3065 -1918
rect 3129 -1982 3145 -1918
rect 3018 -1998 3145 -1982
rect 3018 -2062 3065 -1998
rect 3129 -2062 3145 -1998
rect 3018 -2078 3145 -2062
rect 3018 -2142 3065 -2078
rect 3129 -2142 3145 -2078
rect 3018 -2158 3145 -2142
rect 3018 -2222 3065 -2158
rect 3129 -2222 3145 -2158
rect 3018 -2238 3145 -2222
rect 3018 -2302 3065 -2238
rect 3129 -2302 3145 -2238
rect 3018 -2318 3145 -2302
rect 3018 -2382 3065 -2318
rect 3129 -2382 3145 -2318
rect 3018 -2398 3145 -2382
rect 3018 -2462 3065 -2398
rect 3129 -2462 3145 -2398
rect 3018 -2478 3145 -2462
rect 3018 -2542 3065 -2478
rect 3129 -2542 3145 -2478
rect 3018 -2558 3145 -2542
rect 3018 -2622 3065 -2558
rect 3129 -2622 3145 -2558
rect 3018 -2638 3145 -2622
rect 3018 -2702 3065 -2638
rect 3129 -2702 3145 -2638
rect 3018 -2718 3145 -2702
rect 3018 -2782 3065 -2718
rect 3129 -2782 3145 -2718
rect 3018 -2798 3145 -2782
rect 3018 -2862 3065 -2798
rect 3129 -2862 3145 -2798
rect 3018 -2878 3145 -2862
rect 3018 -2942 3065 -2878
rect 3129 -2942 3145 -2878
rect 3018 -2958 3145 -2942
rect 3018 -3022 3065 -2958
rect 3129 -3022 3145 -2958
rect 3018 -3038 3145 -3022
rect 3018 -3102 3065 -3038
rect 3129 -3102 3145 -3038
rect 3018 -3118 3145 -3102
rect 3018 -3182 3065 -3118
rect 3129 -3182 3145 -3118
rect 3018 -3198 3145 -3182
rect 3018 -3262 3065 -3198
rect 3129 -3262 3145 -3198
rect 3018 -3278 3145 -3262
rect 3018 -3342 3065 -3278
rect 3129 -3342 3145 -3278
rect 3018 -3358 3145 -3342
rect 3018 -3422 3065 -3358
rect 3129 -3422 3145 -3358
rect 3018 -3438 3145 -3422
rect 3018 -3502 3065 -3438
rect 3129 -3502 3145 -3438
rect 3018 -3518 3145 -3502
rect 3018 -3582 3065 -3518
rect 3129 -3582 3145 -3518
rect 3018 -3598 3145 -3582
rect 3018 -3662 3065 -3598
rect 3129 -3662 3145 -3598
rect 3018 -3678 3145 -3662
rect 3018 -3742 3065 -3678
rect 3129 -3742 3145 -3678
rect 3018 -3758 3145 -3742
rect 3018 -3822 3065 -3758
rect 3129 -3822 3145 -3758
rect 3018 -3838 3145 -3822
rect 3018 -3902 3065 -3838
rect 3129 -3902 3145 -3838
rect 3018 -3918 3145 -3902
rect 3018 -3982 3065 -3918
rect 3129 -3982 3145 -3918
rect 3018 -3998 3145 -3982
rect 3018 -4062 3065 -3998
rect 3129 -4062 3145 -3998
rect 3018 -4078 3145 -4062
rect 3018 -4142 3065 -4078
rect 3129 -4142 3145 -4078
rect 3018 -4158 3145 -4142
rect 3018 -4222 3065 -4158
rect 3129 -4222 3145 -4158
rect 3018 -4238 3145 -4222
rect 3018 -4302 3065 -4238
rect 3129 -4302 3145 -4238
rect 3018 -4318 3145 -4302
rect 3018 -4382 3065 -4318
rect 3129 -4382 3145 -4318
rect 3018 -4398 3145 -4382
rect 3018 -4462 3065 -4398
rect 3129 -4462 3145 -4398
rect 3018 -4478 3145 -4462
rect 3018 -4542 3065 -4478
rect 3129 -4542 3145 -4478
rect 3018 -4558 3145 -4542
rect 3018 -4622 3065 -4558
rect 3129 -4622 3145 -4558
rect 3018 -4638 3145 -4622
rect 3018 -4702 3065 -4638
rect 3129 -4702 3145 -4638
rect 3018 -4718 3145 -4702
rect 3018 -4782 3065 -4718
rect 3129 -4782 3145 -4718
rect 3018 -4798 3145 -4782
rect 3018 -4862 3065 -4798
rect 3129 -4862 3145 -4798
rect 3018 -4878 3145 -4862
rect 3018 -4942 3065 -4878
rect 3129 -4942 3145 -4878
rect 3018 -4958 3145 -4942
rect 3018 -5022 3065 -4958
rect 3129 -5022 3145 -4958
rect 3018 -5038 3145 -5022
rect 3018 -5102 3065 -5038
rect 3129 -5102 3145 -5038
rect 3018 -5118 3145 -5102
rect 3018 -5182 3065 -5118
rect 3129 -5182 3145 -5118
rect 3018 -5198 3145 -5182
rect 3018 -5262 3065 -5198
rect 3129 -5262 3145 -5198
rect 3018 -5278 3145 -5262
rect 3018 -5342 3065 -5278
rect 3129 -5342 3145 -5278
rect 3018 -5358 3145 -5342
rect 3018 -5422 3065 -5358
rect 3129 -5422 3145 -5358
rect 3018 -5438 3145 -5422
rect 3018 -5502 3065 -5438
rect 3129 -5502 3145 -5438
rect 3018 -5518 3145 -5502
rect 3018 -5582 3065 -5518
rect 3129 -5582 3145 -5518
rect 3018 -5598 3145 -5582
rect 3018 -5662 3065 -5598
rect 3129 -5662 3145 -5598
rect 3018 -5678 3145 -5662
rect 3018 -5742 3065 -5678
rect 3129 -5742 3145 -5678
rect 3018 -5758 3145 -5742
rect 3018 -5822 3065 -5758
rect 3129 -5822 3145 -5758
rect 3018 -5838 3145 -5822
rect 3018 -5902 3065 -5838
rect 3129 -5902 3145 -5838
rect 3018 -5918 3145 -5902
rect 3018 -5982 3065 -5918
rect 3129 -5982 3145 -5918
rect 3018 -5998 3145 -5982
rect 3018 -6062 3065 -5998
rect 3129 -6062 3145 -5998
rect 3018 -6078 3145 -6062
rect -102 -6489 2 -6111
rect 3018 -6142 3065 -6078
rect 3129 -6142 3145 -6078
rect 3018 -6158 3145 -6142
rect 3018 -6222 3065 -6158
rect 3129 -6222 3145 -6158
rect 3018 -6238 3145 -6222
rect 3018 -6362 3122 -6238
rect 3018 -6378 3145 -6362
rect 3018 -6442 3065 -6378
rect 3129 -6442 3145 -6378
rect 3018 -6458 3145 -6442
rect -3011 -6498 2911 -6489
rect -3011 -12402 -3002 -6498
rect 2902 -12402 2911 -6498
rect -3011 -12411 2911 -12402
rect 3018 -6522 3065 -6458
rect 3129 -6522 3145 -6458
rect 3018 -6538 3145 -6522
rect 3018 -6602 3065 -6538
rect 3129 -6602 3145 -6538
rect 3018 -6618 3145 -6602
rect 3018 -6682 3065 -6618
rect 3129 -6682 3145 -6618
rect 3018 -6698 3145 -6682
rect 3018 -6762 3065 -6698
rect 3129 -6762 3145 -6698
rect 3018 -6778 3145 -6762
rect 3018 -6842 3065 -6778
rect 3129 -6842 3145 -6778
rect 3018 -6858 3145 -6842
rect 3018 -6922 3065 -6858
rect 3129 -6922 3145 -6858
rect 3018 -6938 3145 -6922
rect 3018 -7002 3065 -6938
rect 3129 -7002 3145 -6938
rect 3018 -7018 3145 -7002
rect 3018 -7082 3065 -7018
rect 3129 -7082 3145 -7018
rect 3018 -7098 3145 -7082
rect 3018 -7162 3065 -7098
rect 3129 -7162 3145 -7098
rect 3018 -7178 3145 -7162
rect 3018 -7242 3065 -7178
rect 3129 -7242 3145 -7178
rect 3018 -7258 3145 -7242
rect 3018 -7322 3065 -7258
rect 3129 -7322 3145 -7258
rect 3018 -7338 3145 -7322
rect 3018 -7402 3065 -7338
rect 3129 -7402 3145 -7338
rect 3018 -7418 3145 -7402
rect 3018 -7482 3065 -7418
rect 3129 -7482 3145 -7418
rect 3018 -7498 3145 -7482
rect 3018 -7562 3065 -7498
rect 3129 -7562 3145 -7498
rect 3018 -7578 3145 -7562
rect 3018 -7642 3065 -7578
rect 3129 -7642 3145 -7578
rect 3018 -7658 3145 -7642
rect 3018 -7722 3065 -7658
rect 3129 -7722 3145 -7658
rect 3018 -7738 3145 -7722
rect 3018 -7802 3065 -7738
rect 3129 -7802 3145 -7738
rect 3018 -7818 3145 -7802
rect 3018 -7882 3065 -7818
rect 3129 -7882 3145 -7818
rect 3018 -7898 3145 -7882
rect 3018 -7962 3065 -7898
rect 3129 -7962 3145 -7898
rect 3018 -7978 3145 -7962
rect 3018 -8042 3065 -7978
rect 3129 -8042 3145 -7978
rect 3018 -8058 3145 -8042
rect 3018 -8122 3065 -8058
rect 3129 -8122 3145 -8058
rect 3018 -8138 3145 -8122
rect 3018 -8202 3065 -8138
rect 3129 -8202 3145 -8138
rect 3018 -8218 3145 -8202
rect 3018 -8282 3065 -8218
rect 3129 -8282 3145 -8218
rect 3018 -8298 3145 -8282
rect 3018 -8362 3065 -8298
rect 3129 -8362 3145 -8298
rect 3018 -8378 3145 -8362
rect 3018 -8442 3065 -8378
rect 3129 -8442 3145 -8378
rect 3018 -8458 3145 -8442
rect 3018 -8522 3065 -8458
rect 3129 -8522 3145 -8458
rect 3018 -8538 3145 -8522
rect 3018 -8602 3065 -8538
rect 3129 -8602 3145 -8538
rect 3018 -8618 3145 -8602
rect 3018 -8682 3065 -8618
rect 3129 -8682 3145 -8618
rect 3018 -8698 3145 -8682
rect 3018 -8762 3065 -8698
rect 3129 -8762 3145 -8698
rect 3018 -8778 3145 -8762
rect 3018 -8842 3065 -8778
rect 3129 -8842 3145 -8778
rect 3018 -8858 3145 -8842
rect 3018 -8922 3065 -8858
rect 3129 -8922 3145 -8858
rect 3018 -8938 3145 -8922
rect 3018 -9002 3065 -8938
rect 3129 -9002 3145 -8938
rect 3018 -9018 3145 -9002
rect 3018 -9082 3065 -9018
rect 3129 -9082 3145 -9018
rect 3018 -9098 3145 -9082
rect 3018 -9162 3065 -9098
rect 3129 -9162 3145 -9098
rect 3018 -9178 3145 -9162
rect 3018 -9242 3065 -9178
rect 3129 -9242 3145 -9178
rect 3018 -9258 3145 -9242
rect 3018 -9322 3065 -9258
rect 3129 -9322 3145 -9258
rect 3018 -9338 3145 -9322
rect 3018 -9402 3065 -9338
rect 3129 -9402 3145 -9338
rect 3018 -9418 3145 -9402
rect 3018 -9482 3065 -9418
rect 3129 -9482 3145 -9418
rect 3018 -9498 3145 -9482
rect 3018 -9562 3065 -9498
rect 3129 -9562 3145 -9498
rect 3018 -9578 3145 -9562
rect 3018 -9642 3065 -9578
rect 3129 -9642 3145 -9578
rect 3018 -9658 3145 -9642
rect 3018 -9722 3065 -9658
rect 3129 -9722 3145 -9658
rect 3018 -9738 3145 -9722
rect 3018 -9802 3065 -9738
rect 3129 -9802 3145 -9738
rect 3018 -9818 3145 -9802
rect 3018 -9882 3065 -9818
rect 3129 -9882 3145 -9818
rect 3018 -9898 3145 -9882
rect 3018 -9962 3065 -9898
rect 3129 -9962 3145 -9898
rect 3018 -9978 3145 -9962
rect 3018 -10042 3065 -9978
rect 3129 -10042 3145 -9978
rect 3018 -10058 3145 -10042
rect 3018 -10122 3065 -10058
rect 3129 -10122 3145 -10058
rect 3018 -10138 3145 -10122
rect 3018 -10202 3065 -10138
rect 3129 -10202 3145 -10138
rect 3018 -10218 3145 -10202
rect 3018 -10282 3065 -10218
rect 3129 -10282 3145 -10218
rect 3018 -10298 3145 -10282
rect 3018 -10362 3065 -10298
rect 3129 -10362 3145 -10298
rect 3018 -10378 3145 -10362
rect 3018 -10442 3065 -10378
rect 3129 -10442 3145 -10378
rect 3018 -10458 3145 -10442
rect 3018 -10522 3065 -10458
rect 3129 -10522 3145 -10458
rect 3018 -10538 3145 -10522
rect 3018 -10602 3065 -10538
rect 3129 -10602 3145 -10538
rect 3018 -10618 3145 -10602
rect 3018 -10682 3065 -10618
rect 3129 -10682 3145 -10618
rect 3018 -10698 3145 -10682
rect 3018 -10762 3065 -10698
rect 3129 -10762 3145 -10698
rect 3018 -10778 3145 -10762
rect 3018 -10842 3065 -10778
rect 3129 -10842 3145 -10778
rect 3018 -10858 3145 -10842
rect 3018 -10922 3065 -10858
rect 3129 -10922 3145 -10858
rect 3018 -10938 3145 -10922
rect 3018 -11002 3065 -10938
rect 3129 -11002 3145 -10938
rect 3018 -11018 3145 -11002
rect 3018 -11082 3065 -11018
rect 3129 -11082 3145 -11018
rect 3018 -11098 3145 -11082
rect 3018 -11162 3065 -11098
rect 3129 -11162 3145 -11098
rect 3018 -11178 3145 -11162
rect 3018 -11242 3065 -11178
rect 3129 -11242 3145 -11178
rect 3018 -11258 3145 -11242
rect 3018 -11322 3065 -11258
rect 3129 -11322 3145 -11258
rect 3018 -11338 3145 -11322
rect 3018 -11402 3065 -11338
rect 3129 -11402 3145 -11338
rect 3018 -11418 3145 -11402
rect 3018 -11482 3065 -11418
rect 3129 -11482 3145 -11418
rect 3018 -11498 3145 -11482
rect 3018 -11562 3065 -11498
rect 3129 -11562 3145 -11498
rect 3018 -11578 3145 -11562
rect 3018 -11642 3065 -11578
rect 3129 -11642 3145 -11578
rect 3018 -11658 3145 -11642
rect 3018 -11722 3065 -11658
rect 3129 -11722 3145 -11658
rect 3018 -11738 3145 -11722
rect 3018 -11802 3065 -11738
rect 3129 -11802 3145 -11738
rect 3018 -11818 3145 -11802
rect 3018 -11882 3065 -11818
rect 3129 -11882 3145 -11818
rect 3018 -11898 3145 -11882
rect 3018 -11962 3065 -11898
rect 3129 -11962 3145 -11898
rect 3018 -11978 3145 -11962
rect 3018 -12042 3065 -11978
rect 3129 -12042 3145 -11978
rect 3018 -12058 3145 -12042
rect 3018 -12122 3065 -12058
rect 3129 -12122 3145 -12058
rect 3018 -12138 3145 -12122
rect 3018 -12202 3065 -12138
rect 3129 -12202 3145 -12138
rect 3018 -12218 3145 -12202
rect 3018 -12282 3065 -12218
rect 3129 -12282 3145 -12218
rect 3018 -12298 3145 -12282
rect 3018 -12362 3065 -12298
rect 3129 -12362 3145 -12298
rect 3018 -12378 3145 -12362
rect -102 -12600 2 -12411
rect 3018 -12442 3065 -12378
rect 3129 -12442 3145 -12378
rect 3018 -12458 3145 -12442
rect 3018 -12522 3065 -12458
rect 3129 -12522 3145 -12458
rect 3018 -12538 3145 -12522
rect 3018 -12600 3122 -12538
<< properties >>
string FIXED_BBOX -3150 6350 3050 12550
<< end >>
