magic
tech sky130A
magscale 1 2
timestamp 1654206378
<< nwell >>
rect 30736 4124 31114 5272
rect 14749 3456 15131 3777
rect 44891 3616 45273 3937
<< nsubdiff >>
rect 45016 3789 45150 3808
rect 45016 3755 45088 3789
rect 45122 3755 45150 3789
rect 45016 3738 45150 3755
rect 14874 3629 15008 3648
rect 14874 3595 14946 3629
rect 14980 3595 15008 3629
rect 14874 3578 15008 3595
<< nsubdiffcont >>
rect 45088 3755 45122 3789
rect 14946 3595 14980 3629
<< locali >>
rect 29711 3830 30067 3836
rect 29711 3796 29758 3830
rect 29792 3796 29846 3830
rect 29880 3796 30067 3830
rect 29711 3786 30067 3796
rect 44813 3789 45356 3809
rect 44813 3755 45088 3789
rect 45122 3755 45356 3789
rect 44813 3737 45356 3755
rect 14671 3629 15214 3649
rect 14671 3595 14946 3629
rect 14980 3595 15214 3629
rect 14671 3577 15214 3595
<< viali >>
rect 29758 3796 29792 3830
rect 29846 3796 29880 3830
rect 30423 3828 30457 3862
rect 30606 3792 30640 3826
rect 30694 3792 30728 3826
rect 30782 3792 30816 3826
rect 30870 3792 30904 3826
rect 30958 3792 30992 3826
rect 31046 3792 31080 3826
rect 31134 3792 31168 3826
rect 31222 3792 31256 3826
rect 31310 3792 31344 3826
rect 30423 3748 30457 3782
rect 31029 3690 31063 3724
rect 31195 3686 31229 3720
rect 31363 3692 31397 3726
rect 31530 3690 31564 3724
rect 31700 3691 31734 3725
rect 31864 3692 31898 3726
rect 43514 3669 43548 3714
rect 43682 3676 43716 3721
rect 43850 3666 43884 3711
rect 44018 3678 44052 3723
rect 44184 3676 44218 3721
rect 44350 3678 44384 3723
rect 44518 3678 44552 3723
rect 44692 3676 44726 3721
rect 45448 3670 45482 3715
rect 45610 3674 45644 3719
rect 45780 3678 45814 3723
rect 45944 3674 45978 3719
rect 46114 3674 46148 3719
rect 46282 3670 46316 3715
rect 46450 3674 46484 3719
rect 46624 3670 46658 3715
rect 43714 3578 43748 3612
rect 43814 3578 43848 3612
rect 43914 3578 43948 3612
rect 44014 3578 44048 3612
rect 44114 3578 44148 3612
rect 44214 3578 44248 3612
rect 44314 3578 44348 3612
rect 44414 3578 44448 3612
rect 45374 3578 45408 3612
rect 45474 3578 45508 3612
rect 45574 3578 45608 3612
rect 45674 3578 45708 3612
rect 45774 3578 45808 3612
rect 45874 3578 45908 3612
rect 45974 3578 46008 3612
rect 46074 3578 46108 3612
rect 13372 3509 13406 3554
rect 13540 3516 13574 3561
rect 13708 3506 13742 3551
rect 13876 3518 13910 3563
rect 14042 3516 14076 3561
rect 14208 3518 14242 3563
rect 14376 3518 14410 3563
rect 14550 3516 14584 3561
rect 15306 3510 15340 3555
rect 15468 3514 15502 3559
rect 15638 3518 15672 3563
rect 15802 3514 15836 3559
rect 15972 3514 16006 3559
rect 16140 3510 16174 3555
rect 16308 3514 16342 3559
rect 16482 3510 16516 3555
rect 13572 3418 13606 3452
rect 13672 3418 13706 3452
rect 13772 3418 13806 3452
rect 13872 3418 13906 3452
rect 13972 3418 14006 3452
rect 14072 3418 14106 3452
rect 14172 3418 14206 3452
rect 14272 3418 14306 3452
rect 15232 3418 15266 3452
rect 15332 3418 15366 3452
rect 15432 3418 15466 3452
rect 15532 3418 15566 3452
rect 15632 3418 15666 3452
rect 15732 3418 15766 3452
rect 15832 3418 15866 3452
rect 15932 3418 15966 3452
<< metal1 >>
rect 14423 4747 14678 5103
rect 30359 4770 30693 5094
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14678 4747
rect 7079 4606 7615 4690
rect 14423 4665 14678 4695
rect 30359 4718 30402 4770
rect 30454 4718 30515 4770
rect 30567 4718 30616 4770
rect 30668 4718 30693 4770
rect 30359 4674 30693 4718
rect 44563 4747 44790 5115
rect 44563 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 52529 4785 52735 4812
rect 52529 4733 52575 4785
rect 52627 4733 52670 4785
rect 52722 4733 52735 4785
rect 52529 4723 52735 4733
rect 22113 4615 22721 4673
rect 37217 4623 37841 4681
rect 44563 4661 44790 4695
rect 52223 4629 52956 4687
rect 30487 4150 30555 4163
rect 30487 4098 30517 4150
rect 30487 4067 30555 4098
rect 32027 4067 32062 4163
rect -907 3931 17093 3997
rect 17027 3845 17093 3931
rect 44732 3923 45399 3932
rect 30408 3862 30487 3890
rect 44742 3874 45399 3923
rect 17027 3830 29974 3845
rect 17027 3796 29758 3830
rect 29792 3796 29846 3830
rect 29880 3796 29974 3830
rect 17027 3779 29974 3796
rect 30408 3828 30423 3862
rect 30457 3834 30487 3862
rect 30457 3828 31406 3834
rect 30408 3826 31406 3828
rect 30408 3792 30606 3826
rect 30640 3792 30694 3826
rect 30728 3792 30782 3826
rect 30816 3792 30870 3826
rect 30904 3792 30958 3826
rect 30992 3792 31046 3826
rect 31080 3792 31134 3826
rect 31168 3792 31222 3826
rect 31256 3792 31310 3826
rect 31344 3792 31406 3826
rect 30408 3786 31406 3792
rect 30408 3782 30490 3786
rect 14642 3718 15291 3768
rect 30408 3748 30423 3782
rect 30457 3748 30490 3782
rect 30408 3730 30490 3748
rect 30979 3741 31924 3754
rect 14590 3710 15291 3718
rect 30979 3724 31195 3741
rect 30979 3690 31029 3724
rect 31063 3690 31195 3724
rect 30979 3686 31195 3690
rect 31247 3689 31355 3741
rect 31407 3689 31488 3741
rect 31540 3724 31601 3741
rect 31564 3690 31601 3724
rect 31540 3689 31601 3690
rect 31653 3726 31924 3741
rect 31653 3725 31864 3726
rect 31653 3691 31700 3725
rect 31734 3692 31864 3725
rect 31898 3692 31924 3726
rect 31734 3691 31924 3692
rect 31653 3689 31924 3691
rect 31229 3686 31924 3689
rect 30979 3671 31924 3686
rect 37381 3723 52816 3733
rect 37381 3721 44018 3723
rect 37381 3714 43682 3721
rect 37381 3713 37563 3714
rect 37381 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3669 43514 3714
rect 43548 3676 43682 3714
rect 43716 3711 44018 3721
rect 43716 3676 43850 3711
rect 43548 3669 43850 3676
rect 37615 3666 43850 3669
rect 43884 3678 44018 3711
rect 44052 3721 44350 3723
rect 44052 3678 44184 3721
rect 43884 3676 44184 3678
rect 44218 3678 44350 3721
rect 44384 3678 44518 3723
rect 44552 3721 45780 3723
rect 44552 3678 44692 3721
rect 44218 3676 44692 3678
rect 44726 3719 45780 3721
rect 44726 3715 45610 3719
rect 44726 3676 45448 3715
rect 43884 3670 45448 3676
rect 45482 3674 45610 3715
rect 45644 3678 45780 3719
rect 45814 3719 52816 3723
rect 45814 3678 45944 3719
rect 45644 3674 45944 3678
rect 45978 3674 46114 3719
rect 46148 3715 46450 3719
rect 46148 3674 46282 3715
rect 45482 3670 46282 3674
rect 46316 3674 46450 3715
rect 46484 3715 52816 3719
rect 46484 3674 46624 3715
rect 46316 3670 46624 3674
rect 46658 3714 52816 3715
rect 46658 3709 52664 3714
rect 46658 3670 52573 3709
rect 43884 3666 52573 3670
rect 37615 3662 52573 3666
rect 37512 3661 52573 3662
rect 37381 3657 52573 3661
rect 52625 3662 52664 3709
rect 52716 3662 52816 3714
rect 52625 3657 52816 3662
rect 37381 3652 52816 3657
rect 30487 3597 30555 3619
rect 7224 3563 22590 3573
rect 7224 3561 13876 3563
rect 7224 3558 13540 3561
rect 7224 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3554 13540 3558
rect 7413 3509 13372 3554
rect 13406 3516 13540 3554
rect 13574 3551 13876 3561
rect 13574 3516 13708 3551
rect 13406 3509 13708 3516
rect 7413 3506 13708 3509
rect 13742 3518 13876 3551
rect 13910 3561 14208 3563
rect 13910 3518 14042 3561
rect 13742 3516 14042 3518
rect 14076 3518 14208 3561
rect 14242 3518 14376 3563
rect 14410 3561 15638 3563
rect 14410 3518 14550 3561
rect 14076 3516 14550 3518
rect 14584 3559 15638 3561
rect 14584 3555 15468 3559
rect 14584 3516 15306 3555
rect 13742 3510 15306 3516
rect 15340 3514 15468 3555
rect 15502 3518 15638 3559
rect 15672 3559 22590 3563
rect 15672 3518 15802 3559
rect 15502 3514 15802 3518
rect 15836 3514 15972 3559
rect 16006 3555 16308 3559
rect 16006 3514 16140 3555
rect 15340 3510 16140 3514
rect 16174 3514 16308 3555
rect 16342 3556 22590 3559
rect 16342 3555 22475 3556
rect 16342 3514 16482 3555
rect 16174 3510 16482 3514
rect 16516 3549 22475 3555
rect 16516 3510 22376 3549
rect 13742 3506 22376 3510
rect 7224 3497 22376 3506
rect 22428 3504 22475 3549
rect 22527 3504 22590 3556
rect 30518 3545 30555 3597
rect 30487 3523 30555 3545
rect 32027 3523 32062 3619
rect 43682 3612 46285 3618
rect 43682 3578 43714 3612
rect 43748 3578 43814 3612
rect 43848 3578 43914 3612
rect 43948 3578 44014 3612
rect 44048 3578 44114 3612
rect 44148 3578 44214 3612
rect 44248 3578 44314 3612
rect 44348 3578 44414 3612
rect 44448 3578 45374 3612
rect 45408 3578 45474 3612
rect 45508 3578 45574 3612
rect 45608 3578 45674 3612
rect 45708 3578 45774 3612
rect 45808 3578 45874 3612
rect 45908 3578 45974 3612
rect 46008 3578 46074 3612
rect 46108 3578 46285 3612
rect 43682 3573 46285 3578
rect 43682 3570 45128 3573
rect 44978 3569 45128 3570
rect 22428 3497 22590 3504
rect 7224 3492 22590 3497
rect 44978 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3570 46285 3573
rect 45180 3521 45206 3570
rect 45075 3517 45206 3521
rect 44978 3478 45206 3517
rect 13540 3452 16143 3458
rect 13540 3418 13572 3452
rect 13606 3418 13672 3452
rect 13706 3418 13772 3452
rect 13806 3418 13872 3452
rect 13906 3418 13972 3452
rect 14006 3418 14072 3452
rect 14106 3418 14172 3452
rect 14206 3418 14272 3452
rect 14306 3418 15232 3452
rect 15266 3418 15332 3452
rect 15366 3418 15432 3452
rect 15466 3418 15532 3452
rect 15566 3418 15632 3452
rect 15666 3418 15732 3452
rect 15766 3418 15832 3452
rect 15866 3418 15932 3452
rect 15966 3418 16143 3452
rect 13540 3413 16143 3418
rect 13540 3410 14986 3413
rect 14836 3409 14986 3410
rect 14836 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3410 16143 3413
rect 15038 3361 15064 3410
rect 14933 3357 15064 3361
rect 14836 3318 15064 3357
rect 44732 3326 45484 3384
rect 13202 3148 13253 3244
rect 14590 3172 15271 3230
rect 19721 3175 45232 3219
rect 19721 3173 45120 3175
rect 13202 3147 13252 3148
rect 19721 3121 31184 3173
rect 31236 3121 31328 3173
rect 31380 3121 31472 3173
rect 31524 3172 45120 3173
rect 31524 3121 45031 3172
rect 19721 3120 45031 3121
rect 45083 3123 45120 3172
rect 45172 3123 45232 3175
rect 45083 3120 45232 3123
rect 19721 3096 45232 3120
rect 19721 3089 45031 3096
rect 19721 3037 31183 3089
rect 31235 3037 31327 3089
rect 31379 3037 31471 3089
rect 31523 3044 45031 3089
rect 45083 3044 45124 3096
rect 45176 3044 45232 3096
rect 31523 3037 45232 3044
rect 14848 3013 45232 3037
rect 14848 2992 19927 3013
rect 14848 2940 14885 2992
rect 14937 2987 19927 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 19927 2987
rect 14848 2914 19927 2935
rect 14848 2912 14979 2914
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 19927 2914
rect 14937 2860 19927 2862
rect 14848 2831 19927 2860
rect 7015 2762 7678 2820
rect 22113 2774 22741 2832
rect 37125 2774 37888 2832
rect 52315 2765 52966 2823
rect 52547 2665 52745 2669
rect 52547 2613 52576 2665
rect 52628 2613 52659 2665
rect 52711 2613 52745 2665
rect 52547 2576 52745 2613
rect 60382 780 60604 858
<< via1 >>
rect 7264 4761 7316 4813
rect 7345 4760 7397 4812
rect 22380 4758 22432 4810
rect 22475 4758 22527 4810
rect 14443 4695 14495 4747
rect 14521 4695 14573 4747
rect 14614 4695 14666 4747
rect 6272 4615 6324 4667
rect 6379 4617 6431 4669
rect 6481 4617 6533 4669
rect 6581 4618 6633 4670
rect 30402 4718 30454 4770
rect 30515 4718 30567 4770
rect 30616 4718 30668 4770
rect 37457 4760 37509 4812
rect 37559 4760 37611 4812
rect 44594 4695 44646 4747
rect 44677 4695 44729 4747
rect 52575 4733 52627 4785
rect 52670 4733 52722 4785
rect 21302 4621 21354 4673
rect 21405 4621 21457 4673
rect 21488 4621 21540 4673
rect 21589 4621 21641 4673
rect 21676 4621 21728 4673
rect 36434 4617 36486 4669
rect 36522 4617 36574 4669
rect 36607 4622 36659 4674
rect 53350 4614 53402 4666
rect 53444 4614 53496 4666
rect 53521 4614 53573 4666
rect 53601 4613 53653 4665
rect 53675 4614 53727 4666
rect 30414 4095 30466 4147
rect 30517 4098 30569 4150
rect 30618 4098 30670 4150
rect 44600 3870 44652 3922
rect 44690 3871 44742 3923
rect 14467 3718 14519 3770
rect 14590 3718 14642 3770
rect 31195 3720 31247 3741
rect 31195 3689 31229 3720
rect 31229 3689 31247 3720
rect 31355 3726 31407 3741
rect 31355 3692 31363 3726
rect 31363 3692 31397 3726
rect 31397 3692 31407 3726
rect 31355 3689 31407 3692
rect 31488 3724 31540 3741
rect 31488 3690 31530 3724
rect 31530 3690 31540 3724
rect 31488 3689 31540 3690
rect 31601 3689 31653 3741
rect 37460 3661 37512 3713
rect 37563 3662 37615 3714
rect 52573 3657 52625 3709
rect 52664 3662 52716 3714
rect 7265 3506 7317 3558
rect 7361 3506 7413 3558
rect 22376 3497 22428 3549
rect 22475 3504 22527 3556
rect 30370 3543 30422 3595
rect 30466 3545 30518 3597
rect 30577 3548 30629 3600
rect 30669 3545 30721 3597
rect 45023 3517 45075 3569
rect 45128 3521 45180 3573
rect 14881 3357 14933 3409
rect 14986 3361 15038 3413
rect 46035 3330 46087 3382
rect 46127 3331 46179 3383
rect 46217 3330 46269 3382
rect 46305 3329 46357 3381
rect 13680 3169 13732 3221
rect 13764 3169 13816 3221
rect 13857 3170 13909 3222
rect 31184 3121 31236 3173
rect 31328 3121 31380 3173
rect 31472 3121 31524 3173
rect 45031 3120 45083 3172
rect 45120 3123 45172 3175
rect 31183 3037 31235 3089
rect 31327 3037 31379 3089
rect 31471 3037 31523 3089
rect 45031 3044 45083 3096
rect 45124 3044 45176 3096
rect 14885 2940 14937 2992
rect 14979 2935 15031 2987
rect 14885 2860 14937 2912
rect 14979 2862 15031 2914
rect 6266 2765 6318 2817
rect 6364 2765 6416 2817
rect 6459 2765 6511 2817
rect 6564 2765 6616 2817
rect 21316 2770 21368 2822
rect 21416 2770 21468 2822
rect 21515 2770 21567 2822
rect 21618 2770 21670 2822
rect 36424 2764 36476 2816
rect 36512 2764 36564 2816
rect 36610 2760 36662 2812
rect 53346 2761 53398 2813
rect 53434 2761 53486 2813
rect 53517 2761 53569 2813
rect 53604 2761 53656 2813
rect 7265 2623 7317 2675
rect 7345 2621 7397 2673
rect 22381 2638 22433 2690
rect 22464 2638 22516 2690
rect 37459 2628 37511 2680
rect 37550 2628 37602 2680
rect 52576 2613 52628 2665
rect 52659 2613 52711 2665
<< metal2 >>
rect 1390 6648 1434 7270
rect 3278 6648 3322 7270
rect 5166 6648 5210 7270
rect 7054 6648 7098 7270
rect 8942 6648 8986 7270
rect 10830 6648 10874 7270
rect 12718 6648 12762 7270
rect 14606 6648 14650 7270
rect 16494 6648 16538 7270
rect 18382 6648 18426 7270
rect 20270 6648 20314 7270
rect 22158 6648 22202 7270
rect 24046 6648 24090 7270
rect 25934 6648 25978 7270
rect 27822 6648 27866 7270
rect 29710 6648 29754 7270
rect 31598 6648 31642 7270
rect 33486 6648 33530 7270
rect 35374 6648 35418 7270
rect 37262 6648 37306 7270
rect 39150 6648 39194 7270
rect 41038 6648 41082 7270
rect 42926 6648 42970 7270
rect 44814 6648 44858 7270
rect 46702 6648 46746 7270
rect 48590 6648 48634 7270
rect 50478 6648 50522 7270
rect 52366 6648 52410 7270
rect 54254 6648 54298 7270
rect 56142 6648 56186 7270
rect 58030 6648 58074 7270
rect 59918 6648 59962 7270
rect 60491 5966 60605 6013
rect -636 5930 -394 5966
rect 59938 5930 60605 5966
rect -636 5876 -520 5930
rect -629 1510 -539 5876
rect 7240 4813 7429 4843
rect 7240 4761 7264 4813
rect 7316 4812 7429 4813
rect 7316 4761 7345 4812
rect 7240 4760 7345 4761
rect 7397 4760 7429 4812
rect 6208 4670 6692 4719
rect 6208 4669 6581 4670
rect 6208 4667 6379 4669
rect 6208 4615 6272 4667
rect 6324 4617 6379 4667
rect 6431 4617 6481 4669
rect 6533 4618 6581 4669
rect 6633 4618 6692 4670
rect 6533 4617 6692 4618
rect 6324 4615 6692 4617
rect 6208 3372 6692 4615
rect 6208 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6692 3372
rect 6208 3257 6692 3316
rect 6208 3201 6275 3257
rect 6331 3201 6389 3257
rect 6445 3201 6503 3257
rect 6559 3201 6692 3257
rect 6208 3142 6692 3201
rect 6208 3086 6275 3142
rect 6331 3086 6389 3142
rect 6445 3086 6503 3142
rect 6559 3086 6692 3142
rect 6208 2817 6692 3086
rect 6208 2765 6266 2817
rect 6318 2765 6364 2817
rect 6416 2765 6459 2817
rect 6511 2765 6564 2817
rect 6616 2765 6692 2817
rect 6208 2729 6692 2765
rect 7240 3558 7429 4760
rect 14423 4747 14683 4818
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14683 4747
rect 22351 4810 22540 4833
rect 22351 4758 22380 4810
rect 22432 4758 22475 4810
rect 22527 4758 22540 4810
rect 14423 3770 14683 4695
rect 14423 3718 14467 3770
rect 14519 3718 14590 3770
rect 14642 3718 14683 3770
rect 14423 3674 14683 3718
rect 21264 4673 21731 4697
rect 21264 4621 21302 4673
rect 21354 4621 21405 4673
rect 21457 4621 21488 4673
rect 21540 4621 21589 4673
rect 21641 4621 21676 4673
rect 21728 4621 21731 4673
rect 7240 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3506 7429 3558
rect 7240 2675 7429 3506
rect 14848 3413 15054 3458
rect 14848 3409 14986 3413
rect 14848 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3361 15054 3413
rect 14933 3357 15054 3361
rect 7240 2623 7265 2675
rect 7317 2673 7429 2675
rect 7317 2623 7345 2673
rect 7240 2621 7345 2623
rect 7397 2621 7429 2673
rect 13629 3222 13982 3268
rect 13629 3221 13857 3222
rect 13629 3169 13680 3221
rect 13732 3169 13764 3221
rect 13816 3170 13857 3221
rect 13909 3170 13982 3222
rect 13816 3169 13982 3170
rect 13629 2811 13982 3169
rect 14848 2992 15054 3357
rect 14848 2940 14885 2992
rect 14937 2987 15054 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 15054 2987
rect 14848 2914 15054 2935
rect 14848 2912 14979 2914
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 15054 2914
rect 14937 2860 15054 2862
rect 14848 2831 15054 2860
rect 21264 3282 21731 4621
rect 21264 3226 21314 3282
rect 21370 3226 21418 3282
rect 21474 3226 21522 3282
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21264 3166 21731 3226
rect 21264 3110 21314 3166
rect 21370 3110 21418 3166
rect 21474 3110 21522 3166
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3050 21731 3110
rect 21264 2994 21314 3050
rect 21370 2994 21418 3050
rect 21474 2994 21522 3050
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 13629 2755 13669 2811
rect 13725 2755 13777 2811
rect 13833 2755 13885 2811
rect 13941 2755 13982 2811
rect 13629 2717 13982 2755
rect 21264 2822 21731 2994
rect 21264 2770 21316 2822
rect 21368 2770 21416 2822
rect 21468 2770 21515 2822
rect 21567 2770 21618 2822
rect 21670 2770 21731 2822
rect 21264 2746 21731 2770
rect 22351 3556 22540 4758
rect 30356 4770 30691 4813
rect 30356 4718 30402 4770
rect 30454 4718 30515 4770
rect 30567 4718 30616 4770
rect 30668 4718 30691 4770
rect 30356 4150 30691 4718
rect 37442 4812 37629 4831
rect 37442 4760 37457 4812
rect 37509 4760 37559 4812
rect 37611 4760 37629 4812
rect 30356 4147 30517 4150
rect 30356 4095 30414 4147
rect 30466 4098 30517 4147
rect 30569 4098 30618 4150
rect 30670 4098 30691 4150
rect 30466 4095 30691 4098
rect 30356 4063 30691 4095
rect 36380 4674 36680 4695
rect 36380 4669 36607 4674
rect 36380 4617 36434 4669
rect 36486 4617 36522 4669
rect 36574 4622 36607 4669
rect 36659 4622 36680 4674
rect 36574 4617 36680 4622
rect 31127 3741 31666 3764
rect 31127 3689 31195 3741
rect 31247 3689 31355 3741
rect 31407 3689 31488 3741
rect 31540 3689 31601 3741
rect 31653 3689 31666 3741
rect 22351 3549 22475 3556
rect 22351 3497 22376 3549
rect 22428 3504 22475 3549
rect 22527 3504 22540 3556
rect 22428 3497 22540 3504
rect 13629 2661 13669 2717
rect 13725 2661 13777 2717
rect 13833 2661 13885 2717
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 22351 2690 22540 3497
rect 30318 3600 30743 3618
rect 30318 3597 30577 3600
rect 30318 3595 30466 3597
rect 30318 3543 30370 3595
rect 30422 3545 30466 3595
rect 30518 3548 30577 3597
rect 30629 3597 30743 3600
rect 30629 3548 30669 3597
rect 30518 3545 30669 3548
rect 30721 3545 30743 3597
rect 30422 3543 30743 3545
rect 30318 2931 30743 3543
rect 31127 3173 31666 3689
rect 31127 3121 31184 3173
rect 31236 3121 31328 3173
rect 31380 3121 31472 3173
rect 31524 3121 31666 3173
rect 31127 3089 31666 3121
rect 31127 3037 31183 3089
rect 31235 3037 31327 3089
rect 31379 3037 31471 3089
rect 31523 3037 31666 3089
rect 31127 2963 31666 3037
rect 36380 3631 36680 4617
rect 36380 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36680 3631
rect 36380 3543 36680 3575
rect 36380 3487 36401 3543
rect 36457 3487 36495 3543
rect 36551 3487 36589 3543
rect 36645 3487 36680 3543
rect 36380 3455 36680 3487
rect 36380 3399 36401 3455
rect 36457 3399 36495 3455
rect 36551 3399 36589 3455
rect 36645 3399 36680 3455
rect 30318 2875 30364 2931
rect 30420 2875 30489 2931
rect 30545 2875 30614 2931
rect 30670 2875 30743 2931
rect 30318 2835 30743 2875
rect 30318 2779 30364 2835
rect 30420 2779 30489 2835
rect 30545 2779 30614 2835
rect 30670 2779 30743 2835
rect 30318 2747 30743 2779
rect 36380 2816 36680 3399
rect 36380 2764 36424 2816
rect 36476 2764 36512 2816
rect 36564 2812 36680 2816
rect 36564 2764 36610 2812
rect 36380 2760 36610 2764
rect 36662 2760 36680 2812
rect 36380 2743 36680 2760
rect 37442 3714 37629 4760
rect 44571 4747 44790 4800
rect 44571 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 44571 3923 44790 4695
rect 44571 3922 44690 3923
rect 44571 3870 44600 3922
rect 44652 3871 44690 3922
rect 44742 3871 44790 3923
rect 44652 3870 44790 3871
rect 44571 3835 44790 3870
rect 52546 4785 52735 4808
rect 52546 4733 52575 4785
rect 52627 4733 52670 4785
rect 52722 4733 52735 4785
rect 37442 3713 37563 3714
rect 37442 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3662 37629 3714
rect 37512 3661 37629 3662
rect 22351 2638 22381 2690
rect 22433 2638 22464 2690
rect 22516 2638 22540 2690
rect 22351 2625 22540 2638
rect 37442 2680 37629 3661
rect 52546 3714 52735 4733
rect 52546 3709 52664 3714
rect 52546 3657 52573 3709
rect 52625 3662 52664 3709
rect 52716 3662 52735 3714
rect 52625 3657 52735 3662
rect 44990 3573 45196 3618
rect 44990 3569 45128 3573
rect 44990 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3521 45196 3573
rect 45075 3517 45196 3521
rect 44990 3175 45196 3517
rect 44990 3172 45120 3175
rect 44990 3120 45031 3172
rect 45083 3123 45120 3172
rect 45172 3123 45196 3175
rect 45083 3120 45196 3123
rect 44990 3096 45196 3120
rect 44990 3044 45031 3096
rect 45083 3044 45124 3096
rect 45176 3044 45196 3096
rect 44990 3001 45196 3044
rect 45998 3383 46412 3405
rect 45998 3382 46127 3383
rect 45998 3330 46035 3382
rect 46087 3331 46127 3382
rect 46179 3382 46412 3383
rect 46179 3331 46217 3382
rect 46087 3330 46217 3331
rect 46269 3381 46412 3382
rect 46269 3330 46305 3381
rect 45998 3329 46305 3330
rect 46357 3329 46412 3381
rect 37442 2628 37459 2680
rect 37511 2628 37550 2680
rect 37602 2628 37629 2680
rect 7240 2603 7429 2621
rect 37442 2620 37629 2628
rect 45998 2784 46412 3329
rect 45998 2728 46035 2784
rect 46091 2728 46128 2784
rect 46184 2728 46221 2784
rect 46277 2728 46314 2784
rect 46370 2728 46412 2784
rect 45998 2702 46412 2728
rect 45998 2646 46035 2702
rect 46091 2646 46128 2702
rect 46184 2646 46221 2702
rect 46277 2646 46314 2702
rect 46370 2646 46412 2702
rect 45998 2609 46412 2646
rect 52546 2665 52735 3657
rect 53311 4666 53732 4695
rect 53311 4614 53350 4666
rect 53402 4614 53444 4666
rect 53496 4614 53521 4666
rect 53573 4665 53675 4666
rect 53573 4614 53601 4665
rect 53311 4613 53601 4614
rect 53653 4614 53675 4665
rect 53727 4614 53732 4666
rect 53653 4613 53732 4614
rect 53311 3176 53732 4613
rect 53311 3120 53348 3176
rect 53404 3120 53452 3176
rect 53508 3120 53556 3176
rect 53612 3120 53660 3176
rect 53716 3120 53732 3176
rect 53311 3086 53732 3120
rect 53311 3030 53348 3086
rect 53404 3030 53452 3086
rect 53508 3030 53556 3086
rect 53612 3030 53660 3086
rect 53716 3030 53732 3086
rect 53311 2813 53732 3030
rect 53311 2761 53346 2813
rect 53398 2761 53434 2813
rect 53486 2761 53517 2813
rect 53569 2761 53604 2813
rect 53656 2761 53732 2813
rect 53311 2745 53732 2761
rect 52546 2613 52576 2665
rect 52628 2613 52659 2665
rect 52711 2613 52735 2665
rect 52546 2600 52735 2613
rect 60491 1588 60605 5930
rect 60448 1510 60642 1588
rect -634 1474 51 1510
rect 60376 1474 60642 1510
rect -629 1391 -539 1474
rect 20 170 64 792
rect 1908 170 1952 792
rect 3796 170 3840 792
rect 5684 170 5728 792
rect 7572 170 7616 792
rect 9460 170 9504 792
rect 11348 170 11392 792
rect 13236 170 13280 792
rect 15124 170 15168 792
rect 17012 170 17056 792
rect 18900 170 18944 792
rect 20788 170 20832 792
rect 22676 170 22720 792
rect 24564 170 24608 792
rect 26452 170 26496 792
rect 28340 170 28384 792
rect 30228 170 30272 792
rect 32116 170 32160 792
rect 34004 170 34048 792
rect 35892 170 35936 792
rect 37780 170 37824 792
rect 39668 170 39712 792
rect 41556 170 41600 792
rect 43444 170 43488 792
rect 45332 170 45376 792
rect 47220 170 47264 792
rect 49108 170 49152 792
rect 50996 170 51040 792
rect 52884 170 52928 792
rect 54772 170 54816 792
rect 56660 170 56704 792
rect 58548 170 58592 792
<< via2 >>
rect 6275 3316 6331 3372
rect 6389 3316 6445 3372
rect 6503 3316 6559 3372
rect 6275 3201 6331 3257
rect 6389 3201 6445 3257
rect 6503 3201 6559 3257
rect 6275 3086 6331 3142
rect 6389 3086 6445 3142
rect 6503 3086 6559 3142
rect 21314 3226 21370 3282
rect 21418 3226 21474 3282
rect 21522 3226 21578 3282
rect 21626 3226 21682 3282
rect 21314 3110 21370 3166
rect 21418 3110 21474 3166
rect 21522 3110 21578 3166
rect 21626 3110 21682 3166
rect 21314 2994 21370 3050
rect 21418 2994 21474 3050
rect 21522 2994 21578 3050
rect 21626 2994 21682 3050
rect 13669 2755 13725 2811
rect 13777 2755 13833 2811
rect 13885 2755 13941 2811
rect 13669 2661 13725 2717
rect 13777 2661 13833 2717
rect 13885 2661 13941 2717
rect 36401 3575 36457 3631
rect 36495 3575 36551 3631
rect 36589 3575 36645 3631
rect 36401 3487 36457 3543
rect 36495 3487 36551 3543
rect 36589 3487 36645 3543
rect 36401 3399 36457 3455
rect 36495 3399 36551 3455
rect 36589 3399 36645 3455
rect 30364 2875 30420 2931
rect 30489 2875 30545 2931
rect 30614 2875 30670 2931
rect 30364 2779 30420 2835
rect 30489 2779 30545 2835
rect 30614 2779 30670 2835
rect 46035 2728 46091 2784
rect 46128 2728 46184 2784
rect 46221 2728 46277 2784
rect 46314 2728 46370 2784
rect 46035 2646 46091 2702
rect 46128 2646 46184 2702
rect 46221 2646 46277 2702
rect 46314 2646 46370 2702
rect 53348 3120 53404 3176
rect 53452 3120 53508 3176
rect 53556 3120 53612 3176
rect 53660 3120 53716 3176
rect 53348 3030 53404 3086
rect 53452 3030 53508 3086
rect 53556 3030 53612 3086
rect 53660 3030 53716 3086
<< metal3 >>
rect 36378 3631 36682 3645
rect 36378 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36682 3631
rect 36378 3543 36682 3575
rect 36378 3487 36401 3543
rect 36457 3532 36495 3543
rect 36551 3533 36589 3543
rect 36645 3533 36682 3543
rect 36551 3487 36568 3533
rect 36378 3455 36414 3487
rect 36501 3455 36568 3487
rect 6274 3398 6616 3431
rect 36378 3399 36401 3455
rect 36551 3421 36568 3455
rect 36655 3421 36682 3533
rect 36457 3399 36495 3420
rect 36551 3399 36589 3421
rect 36645 3399 36682 3421
rect 6206 3372 6695 3398
rect 36378 3379 36682 3399
rect 6206 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6695 3372
rect 6206 3257 6695 3316
rect 6206 3229 6275 3257
rect 6331 3229 6389 3257
rect 6445 3235 6503 3257
rect 6559 3235 6695 3257
rect 6206 3138 6272 3229
rect 6358 3201 6389 3229
rect 6559 3201 6568 3235
rect 6358 3144 6423 3201
rect 6509 3144 6568 3201
rect 6654 3144 6695 3235
rect 6358 3142 6695 3144
rect 6358 3138 6389 3142
rect 6206 3086 6275 3138
rect 6331 3086 6389 3138
rect 6445 3086 6503 3142
rect 6559 3086 6695 3142
rect 6206 3031 6695 3086
rect 21264 3282 21731 3336
rect 21264 3239 21314 3282
rect 21370 3239 21418 3282
rect 21264 3155 21312 3239
rect 21405 3226 21418 3239
rect 21474 3239 21522 3282
rect 21474 3226 21479 3239
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21405 3166 21479 3226
rect 21572 3166 21731 3226
rect 21405 3155 21418 3166
rect 21264 3110 21314 3155
rect 21370 3110 21418 3155
rect 21474 3155 21479 3166
rect 21474 3110 21522 3155
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3078 21731 3110
rect 21264 2994 21312 3078
rect 21405 3050 21479 3078
rect 21572 3050 21731 3078
rect 21405 2994 21418 3050
rect 21474 2994 21479 3050
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 53311 3183 53733 3204
rect 53311 3176 53355 3183
rect 53439 3176 53476 3183
rect 53560 3176 53614 3183
rect 53698 3176 53733 3183
rect 53311 3120 53348 3176
rect 53439 3120 53452 3176
rect 53612 3120 53614 3176
rect 53716 3120 53733 3176
rect 53311 3086 53355 3120
rect 53439 3086 53476 3120
rect 53560 3086 53614 3120
rect 53698 3086 53733 3120
rect 53311 3030 53348 3086
rect 53439 3030 53452 3086
rect 53612 3030 53614 3086
rect 53716 3030 53733 3086
rect 53311 3025 53355 3030
rect 53439 3025 53476 3030
rect 53560 3025 53614 3030
rect 53698 3025 53733 3030
rect 53311 2996 53733 3025
rect 21264 2950 21731 2994
rect 30316 2931 30741 2969
rect 30316 2892 30364 2931
rect 30420 2892 30489 2931
rect 30545 2892 30614 2931
rect 30670 2892 30741 2931
rect 13629 2811 13982 2834
rect 13629 2763 13669 2811
rect 13725 2763 13777 2811
rect 13833 2763 13885 2811
rect 13629 2694 13653 2763
rect 13730 2694 13756 2763
rect 13833 2694 13859 2763
rect 13941 2755 13982 2811
rect 13936 2717 13982 2755
rect 30316 2780 30362 2892
rect 30449 2780 30481 2892
rect 30568 2780 30600 2892
rect 30687 2780 30741 2892
rect 30316 2779 30364 2780
rect 30420 2779 30489 2780
rect 30545 2779 30614 2780
rect 30670 2779 30741 2780
rect 30316 2742 30741 2779
rect 45998 2808 46413 2851
rect 45998 2807 46176 2808
rect 45998 2784 46036 2807
rect 46120 2784 46176 2807
rect 46260 2784 46304 2808
rect 13629 2661 13669 2694
rect 13725 2661 13777 2694
rect 13833 2661 13885 2694
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 45998 2728 46035 2784
rect 46120 2728 46128 2784
rect 46277 2728 46304 2784
rect 45998 2702 46036 2728
rect 46120 2702 46176 2728
rect 46260 2702 46304 2728
rect 45998 2646 46035 2702
rect 46120 2649 46128 2702
rect 46277 2650 46304 2702
rect 46388 2650 46413 2808
rect 46091 2646 46128 2649
rect 46184 2646 46221 2650
rect 46277 2646 46314 2650
rect 46370 2646 46413 2650
rect 45998 2610 46413 2646
<< via3 >>
rect 2518 7211 2624 7389
rect 2727 7210 2833 7388
rect 2893 7210 2999 7388
rect 3073 7212 3179 7390
rect 1284 5093 1390 5271
rect 1456 5094 1562 5272
rect 1630 5093 1736 5271
rect 36414 3487 36457 3532
rect 36457 3487 36495 3532
rect 36495 3487 36501 3532
rect 36568 3487 36589 3533
rect 36589 3487 36645 3533
rect 36645 3487 36655 3533
rect 36414 3455 36501 3487
rect 36568 3455 36655 3487
rect 36414 3420 36457 3455
rect 36457 3420 36495 3455
rect 36495 3420 36501 3455
rect 36568 3421 36589 3455
rect 36589 3421 36645 3455
rect 36645 3421 36655 3455
rect 6272 3201 6275 3229
rect 6275 3201 6331 3229
rect 6331 3201 6358 3229
rect 6423 3201 6445 3235
rect 6445 3201 6503 3235
rect 6503 3201 6509 3235
rect 6272 3142 6358 3201
rect 6423 3144 6509 3201
rect 6568 3144 6654 3235
rect 6272 3138 6275 3142
rect 6275 3138 6331 3142
rect 6331 3138 6358 3142
rect 21312 3226 21314 3239
rect 21314 3226 21370 3239
rect 21370 3226 21405 3239
rect 21479 3226 21522 3239
rect 21522 3226 21572 3239
rect 21312 3166 21405 3226
rect 21479 3166 21572 3226
rect 21312 3155 21314 3166
rect 21314 3155 21370 3166
rect 21370 3155 21405 3166
rect 21479 3155 21522 3166
rect 21522 3155 21572 3166
rect 21312 3050 21405 3078
rect 21479 3050 21572 3078
rect 21312 2994 21314 3050
rect 21314 2994 21370 3050
rect 21370 2994 21405 3050
rect 21479 2994 21522 3050
rect 21522 2994 21572 3050
rect 53355 3176 53439 3183
rect 53476 3176 53560 3183
rect 53614 3176 53698 3183
rect 53355 3120 53404 3176
rect 53404 3120 53439 3176
rect 53476 3120 53508 3176
rect 53508 3120 53556 3176
rect 53556 3120 53560 3176
rect 53614 3120 53660 3176
rect 53660 3120 53698 3176
rect 53355 3086 53439 3120
rect 53476 3086 53560 3120
rect 53614 3086 53698 3120
rect 53355 3030 53404 3086
rect 53404 3030 53439 3086
rect 53476 3030 53508 3086
rect 53508 3030 53556 3086
rect 53556 3030 53560 3086
rect 53614 3030 53660 3086
rect 53660 3030 53698 3086
rect 53355 3025 53439 3030
rect 53476 3025 53560 3030
rect 53614 3025 53698 3030
rect 13653 2755 13669 2763
rect 13669 2755 13725 2763
rect 13725 2755 13730 2763
rect 13653 2717 13730 2755
rect 13653 2694 13669 2717
rect 13669 2694 13725 2717
rect 13725 2694 13730 2717
rect 13756 2755 13777 2763
rect 13777 2755 13833 2763
rect 13756 2717 13833 2755
rect 13756 2694 13777 2717
rect 13777 2694 13833 2717
rect 13859 2755 13885 2763
rect 13885 2755 13936 2763
rect 13859 2717 13936 2755
rect 30362 2875 30364 2892
rect 30364 2875 30420 2892
rect 30420 2875 30449 2892
rect 30362 2835 30449 2875
rect 30362 2780 30364 2835
rect 30364 2780 30420 2835
rect 30420 2780 30449 2835
rect 30481 2875 30489 2892
rect 30489 2875 30545 2892
rect 30545 2875 30568 2892
rect 30481 2835 30568 2875
rect 30481 2780 30489 2835
rect 30489 2780 30545 2835
rect 30545 2780 30568 2835
rect 30600 2875 30614 2892
rect 30614 2875 30670 2892
rect 30670 2875 30687 2892
rect 30600 2835 30687 2875
rect 30600 2780 30614 2835
rect 30614 2780 30670 2835
rect 30670 2780 30687 2835
rect 46036 2784 46120 2807
rect 46176 2784 46260 2808
rect 46304 2784 46388 2808
rect 13859 2694 13885 2717
rect 13885 2694 13936 2717
rect 46036 2728 46091 2784
rect 46091 2728 46120 2784
rect 46176 2728 46184 2784
rect 46184 2728 46221 2784
rect 46221 2728 46260 2784
rect 46304 2728 46314 2784
rect 46314 2728 46370 2784
rect 46370 2728 46388 2784
rect 46036 2702 46120 2728
rect 46176 2702 46260 2728
rect 46304 2702 46388 2728
rect 46036 2649 46091 2702
rect 46091 2649 46120 2702
rect 46176 2650 46184 2702
rect 46184 2650 46221 2702
rect 46221 2650 46260 2702
rect 46304 2650 46314 2702
rect 46314 2650 46370 2702
rect 46370 2650 46388 2702
rect 1286 2145 1392 2323
rect 1491 2147 1597 2325
rect 1690 2147 1796 2325
rect 2532 34 2638 212
rect 2753 34 2859 212
rect 2962 34 3068 212
rect 3136 34 3242 212
rect 6260 66 6346 157
rect 6408 66 6494 157
rect 6556 66 6642 157
rect 13779 140 13856 209
rect 13802 21 13879 90
rect 21317 61 21413 169
rect 21450 61 21546 169
rect 21583 61 21679 169
rect 30383 48 30470 160
rect 30506 48 30593 160
rect 30638 48 30725 160
rect 36412 45 36499 157
rect 36581 45 36668 157
rect 46038 32 46122 190
rect 46151 32 46235 190
rect 46266 32 46350 190
rect 53361 42 53445 200
rect 53480 42 53564 200
rect 53609 42 53693 200
<< metal4 >>
rect 2467 7390 3251 7443
rect 2467 7389 3073 7390
rect 2467 7211 2518 7389
rect 2624 7388 3073 7389
rect 2624 7211 2727 7388
rect 2467 7210 2727 7211
rect 2833 7210 2893 7388
rect 2999 7212 3073 7388
rect 3179 7212 3251 7390
rect 2999 7210 3251 7212
rect 1234 5272 1852 5401
rect 1234 5271 1456 5272
rect 1234 5093 1284 5271
rect 1390 5094 1456 5271
rect 1562 5271 1852 5272
rect 1562 5094 1630 5271
rect 1390 5093 1630 5094
rect 1736 5093 1852 5271
rect 1234 2325 1852 5093
rect 1234 2323 1491 2325
rect 1234 2145 1286 2323
rect 1392 2147 1491 2323
rect 1597 2147 1690 2325
rect 1796 2147 1852 2325
rect 1392 2145 1852 2147
rect 1234 2095 1852 2145
rect 2467 212 3251 7210
rect 36378 3533 36683 3690
rect 36378 3532 36568 3533
rect 36378 3420 36414 3532
rect 36501 3421 36568 3532
rect 36655 3421 36683 3533
rect 36501 3420 36683 3421
rect 2467 34 2532 212
rect 2638 34 2753 212
rect 2859 34 2962 212
rect 3068 34 3136 212
rect 3242 34 3251 212
rect 2467 -55 3251 34
rect 6214 3235 6683 3350
rect 6214 3229 6423 3235
rect 6214 3138 6272 3229
rect 6358 3144 6423 3229
rect 6509 3144 6568 3235
rect 6654 3144 6683 3235
rect 6358 3138 6683 3144
rect 6214 157 6683 3138
rect 21264 3239 21731 3364
rect 21264 3155 21312 3239
rect 21405 3155 21479 3239
rect 21572 3155 21731 3239
rect 21264 3078 21731 3155
rect 21264 2994 21312 3078
rect 21405 2994 21479 3078
rect 21572 2994 21731 3078
rect 13629 2763 13983 2835
rect 13629 2694 13653 2763
rect 13730 2694 13756 2763
rect 13833 2694 13859 2763
rect 13936 2694 13983 2763
rect 13629 2634 13983 2694
rect 6214 66 6260 157
rect 6346 66 6408 157
rect 6494 66 6556 157
rect 6642 66 6683 157
rect 6214 -33 6683 66
rect 13705 209 13906 2634
rect 13705 140 13779 209
rect 13856 140 13906 209
rect 13705 90 13906 140
rect 13705 21 13802 90
rect 13879 21 13906 90
rect 13705 -58 13906 21
rect 21264 169 21731 2994
rect 21264 61 21317 169
rect 21413 61 21450 169
rect 21546 61 21583 169
rect 21679 61 21731 169
rect 21264 -8 21731 61
rect 30316 2892 30741 2971
rect 30316 2780 30362 2892
rect 30449 2780 30481 2892
rect 30568 2780 30600 2892
rect 30687 2780 30741 2892
rect 30316 160 30741 2780
rect 30316 48 30383 160
rect 30470 48 30506 160
rect 30593 48 30638 160
rect 30725 48 30741 160
rect 30316 6 30741 48
rect 36378 157 36683 3420
rect 53311 3183 53736 3206
rect 53311 3025 53355 3183
rect 53439 3025 53476 3183
rect 53560 3025 53614 3183
rect 53698 3025 53736 3183
rect 36378 45 36412 157
rect 36499 45 36581 157
rect 36668 45 36683 157
rect 36378 -3 36683 45
rect 45998 2808 46412 2897
rect 45998 2807 46176 2808
rect 45998 2649 46036 2807
rect 46120 2650 46176 2807
rect 46260 2650 46304 2808
rect 46388 2650 46412 2808
rect 46120 2649 46412 2650
rect 45998 190 46412 2649
rect 45998 32 46038 190
rect 46122 32 46151 190
rect 46235 32 46266 190
rect 46350 32 46412 190
rect 45998 -56 46412 32
rect 53311 200 53736 3025
rect 53311 42 53361 200
rect 53445 42 53480 200
rect 53564 42 53609 200
rect 53693 42 53736 200
rect 53311 -44 53736 42
use brbufhalf  brbufhalf_0
timestamp 1654123708
transform 1 0 3552 0 1 -2528
box -3552 2527 26658 5370
use brbufhalf  brbufhalf_1
timestamp 1654123708
transform 1 0 33754 0 1 -2528
box -3552 2527 26658 5370
use brbufhalf  brbufhalf_2
timestamp 1654123708
transform -1 0 56430 0 -1 9968
box -3552 2527 26658 5370
use brbufhalf  brbufhalf_3
timestamp 1654123708
transform -1 0 26228 0 -1 9968
box -3552 2527 26658 5370
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1653697408
transform 1 0 30027 0 1 3571
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654066915
transform 1 0 15169 0 1 3195
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654066915
transform 1 0 13239 0 1 3195
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1654066915
transform 1 0 30555 0 1 3571
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1654066915
transform 1 0 45311 0 1 3355
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1654066915
transform 1 0 43381 0 1 3355
box -38 -48 1510 592
<< labels >>
flabel metal4 1234 2325 1852 5093 1 FreeSans 1600 0 0 0 VDD
port 1 n
flabel metal4 2467 212 3251 7210 1 FreeSans 1600 0 0 0 VSS
port 2 n
flabel metal1 60382 780 60604 858 1 FreeSans 1600 0 0 0 OUT
port 3 n
flabel metal2 59918 6648 59962 7270 1 FreeSans 800 0 0 0 C[0]
port 67 n
flabel metal2 58030 6648 58074 7270 1 FreeSans 800 0 0 0 C[1]
port 66 n
flabel metal2 56142 6648 56186 7270 1 FreeSans 800 0 0 0 C[2]
port 65 n
flabel metal2 54254 6648 54298 7270 1 FreeSans 800 0 0 0 C[3]
port 64 n
flabel metal2 52366 6648 52410 7270 1 FreeSans 800 0 0 0 C[4]
port 63 n
flabel metal2 50478 6648 50522 7270 1 FreeSans 800 0 0 0 C[5]
port 62 n
flabel metal2 48590 6648 48634 7270 1 FreeSans 800 0 0 0 C[6]
port 61 n
flabel metal2 46702 6648 46746 7270 1 FreeSans 800 0 0 0 C[7]
port 60 n
flabel metal2 44814 6648 44858 7270 1 FreeSans 800 0 0 0 C[8]
port 59 n
flabel metal2 42926 6648 42970 7270 1 FreeSans 800 0 0 0 C[9]
port 58 n
flabel metal2 41038 6648 41082 7270 1 FreeSans 800 0 0 0 C[10]
port 57 n
flabel metal2 39150 6648 39194 7270 1 FreeSans 800 0 0 0 C[11]
port 56 n
flabel metal2 37262 6648 37306 7270 1 FreeSans 800 0 0 0 C[12]
port 55 n
flabel metal2 35374 6648 35418 7270 1 FreeSans 800 0 0 0 C[13]
port 54 n
flabel metal2 33486 6648 33530 7270 1 FreeSans 800 0 0 0 C[14]
port 53 n
flabel metal2 31598 6648 31642 7270 1 FreeSans 800 0 0 0 C[15]
port 52 n
flabel metal2 29710 6648 29754 7270 1 FreeSans 800 0 0 0 C[16]
port 51 n
flabel metal2 27822 6648 27866 7270 1 FreeSans 800 0 0 0 C[17]
port 50 n
flabel metal2 25934 6648 25978 7270 1 FreeSans 800 0 0 0 C[18]
port 49 n
flabel metal2 24046 6648 24090 7270 1 FreeSans 800 0 0 0 C[19]
port 48 n
flabel metal2 22158 6648 22202 7270 1 FreeSans 800 0 0 0 C[20]
port 47 n
flabel metal2 20270 6648 20314 7270 1 FreeSans 800 0 0 0 C[21]
port 46 n
flabel metal2 18382 6648 18426 7270 1 FreeSans 800 0 0 0 C[22]
port 45 n
flabel metal2 16494 6648 16538 7270 1 FreeSans 800 0 0 0 C[23]
port 44 n
flabel metal2 14606 6648 14650 7270 1 FreeSans 800 0 0 0 C[24]
port 43 n
flabel metal2 12718 6648 12762 7270 1 FreeSans 800 0 0 0 C[25]
port 42 n
flabel metal2 10830 6648 10874 7270 1 FreeSans 800 0 0 0 C[26]
port 41 n
flabel metal2 8942 6648 8986 7270 1 FreeSans 800 0 0 0 C[27]
port 40 n
flabel metal2 7054 6648 7098 7270 1 FreeSans 800 0 0 0 C[28]
port 39 n
flabel metal2 5166 6648 5210 7270 1 FreeSans 800 0 0 0 C[29]
port 38 n
flabel metal2 3278 6648 3322 7270 1 FreeSans 800 0 0 0 C[30]
port 37 n
flabel metal2 1390 6648 1434 7270 1 FreeSans 800 0 0 0 C[31]
port 36 n
flabel metal2 20 170 64 792 1 FreeSans 800 0 0 0 C[32]
port 35 n
flabel metal2 1908 170 1952 792 1 FreeSans 800 0 0 0 C[33]
port 34 n
flabel metal2 3796 170 3840 792 1 FreeSans 800 0 0 0 C[34]
port 33 n
flabel metal2 5684 170 5728 792 1 FreeSans 800 0 0 0 C[35]
port 32 n
flabel metal2 7572 170 7616 792 1 FreeSans 800 0 0 0 C[36]
port 31 n
flabel metal2 9460 170 9504 792 1 FreeSans 800 0 0 0 C[37]
port 30 n
flabel metal2 11348 170 11392 792 1 FreeSans 800 0 0 0 C[38]
port 29 n
flabel metal2 13236 170 13280 792 1 FreeSans 800 0 0 0 C[39]
port 28 n
flabel metal2 15124 170 15168 792 1 FreeSans 800 0 0 0 C[40]
port 27 n
flabel metal2 17012 170 17056 792 1 FreeSans 800 0 0 0 C[41]
port 26 n
flabel metal2 18900 170 18944 792 1 FreeSans 800 0 0 0 C[42]
port 25 n
flabel metal2 20788 170 20832 792 1 FreeSans 800 0 0 0 C[43]
port 24 n
flabel metal2 22676 170 22720 792 1 FreeSans 800 0 0 0 C[44]
port 23 n
flabel metal2 24564 170 24608 792 1 FreeSans 800 0 0 0 C[45]
port 22 n
flabel metal2 26452 170 26496 792 1 FreeSans 800 0 0 0 C[46]
port 21 n
flabel metal2 28340 170 28384 792 1 FreeSans 800 0 0 0 C[47]
port 20 n
flabel metal2 30228 170 30272 792 1 FreeSans 800 0 0 0 C[48]
port 19 n
flabel metal2 32116 170 32160 792 1 FreeSans 800 0 0 0 C[49]
port 18 n
flabel metal2 34004 170 34048 792 1 FreeSans 800 0 0 0 C[50]
port 17 n
flabel metal2 35892 170 35936 792 1 FreeSans 800 0 0 0 C[51]
port 16 n
flabel metal2 37780 170 37824 792 1 FreeSans 800 0 0 0 C[52]
port 15 n
flabel metal2 39668 170 39712 792 1 FreeSans 800 0 0 0 C[53]
port 14 n
flabel metal2 41556 170 41600 792 1 FreeSans 800 0 0 0 C[54]
port 13 n
flabel metal2 43444 170 43488 792 1 FreeSans 800 0 0 0 C[55]
port 12 n
flabel metal2 45332 170 45376 792 1 FreeSans 800 0 0 0 C[56]
port 11 n
flabel metal2 47220 170 47264 792 1 FreeSans 800 0 0 0 C[57]
port 10 n
flabel metal2 49108 170 49152 792 1 FreeSans 800 0 0 0 C[58]
port 9 n
flabel metal2 50996 170 51040 792 1 FreeSans 800 0 0 0 C[59]
port 8 n
flabel metal2 52884 170 52928 792 1 FreeSans 800 0 0 0 C[60]
port 7 n
flabel metal2 54772 170 54816 792 1 FreeSans 800 0 0 0 C[61]
port 6 n
flabel metal2 56660 170 56704 792 1 FreeSans 800 0 0 0 C[62]
port 5 n
flabel metal2 58548 170 58592 792 1 FreeSans 800 0 0 0 C[63]
port 4 n
flabel metal1 -907 3931 -653 3997 1 FreeSans 1600 0 0 0 RESET
port 68 n
<< end >>
