magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 549 157 735 203
rect 1 21 735 157
rect 29 -17 63 21
<< locali >>
rect 17 199 90 335
rect 304 84 360 339
rect 405 84 459 339
rect 497 133 565 339
rect 667 299 719 493
rect 685 161 719 299
rect 651 68 719 161
rect 651 59 718 68
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 34 403 69 493
rect 103 439 169 527
rect 230 409 264 493
rect 311 445 445 527
rect 488 409 522 493
rect 562 445 628 527
rect 34 369 160 403
rect 126 265 160 369
rect 230 375 633 409
rect 126 199 196 265
rect 126 165 160 199
rect 34 131 160 165
rect 34 51 69 131
rect 230 117 264 375
rect 103 17 169 93
rect 218 51 264 117
rect 599 265 633 375
rect 599 199 651 265
rect 551 17 617 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 17 199 90 335 6 A_N
port 1 nsew signal input
rlabel locali s 304 84 360 339 6 B
port 2 nsew signal input
rlabel locali s 405 84 459 339 6 C
port 3 nsew signal input
rlabel locali s 497 133 565 339 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 735 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 549 157 735 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 651 59 718 68 6 X
port 9 nsew signal output
rlabel locali s 651 68 719 161 6 X
port 9 nsew signal output
rlabel locali s 685 161 719 299 6 X
port 9 nsew signal output
rlabel locali s 667 299 719 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3042500
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3034946
<< end >>
