magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 11772 -270 23593 34
<< pwell >>
rect 10099 -220 11657 4351
<< obsli1 >>
rect 9522 0 23971 39532
rect 9522 -194 11631 0
rect 11807 -23 12009 0
rect 23346 -23 23536 0
rect 11807 -213 23536 -23
<< obsm1 >>
rect 9437 0 23983 39538
rect 10125 -181 11171 0
rect 11807 -23 12070 0
tri 12070 -23 12093 0 sw
tri 23285 -23 23308 0 se
rect 23308 -23 23536 0
rect 11807 -213 23536 -23
<< metal2 >>
rect 9499 -407 14279 4
rect 19478 -407 24258 4725
<< obsm2 >>
rect 9453 4781 24258 38608
rect 9453 60 19422 4781
rect 14335 0 19422 60
rect 14579 -407 14979 -23
<< metal3 >>
rect 0 -407 14279 2730
rect 14579 -407 16779 138
rect 16978 -407 19178 1859
rect 19478 -407 33800 2730
<< obsm3 >>
rect 0 2810 33800 39593
rect 14359 1939 19398 2810
rect 14359 218 16898 1939
rect 14359 138 14499 218
rect 16859 138 16898 218
rect 19258 138 19398 1939
<< metal4 >>
rect 0 34750 9641 39593
rect 25649 34750 33800 39593
rect 0 13600 9543 18593
rect 25177 13600 33800 18593
rect 0 12410 9543 13300
rect 25177 12410 33800 13300
rect 0 11240 9543 12130
rect 25177 11240 33800 12130
rect 0 10874 33800 10940
rect 0 10218 33800 10814
rect 0 9922 9448 10158
rect 25177 9922 33800 10158
rect 0 9266 33800 9862
rect 0 9140 33800 9206
rect 0 7910 9450 8840
rect 25177 7910 33800 8840
rect 0 6940 9543 7630
rect 25177 6940 33800 7630
rect 0 5970 9543 6660
rect 25177 5970 33800 6660
rect 0 4760 9543 5690
rect 25177 4760 33800 5690
rect 0 3550 9543 4480
rect 24241 3550 33800 4480
rect 0 2580 9543 3270
rect 24241 2580 33800 3270
rect 0 1370 9543 2300
rect 25177 1370 33800 2300
rect 0 0 9543 1090
rect 25177 0 33800 1090
<< obsm4 >>
rect 9721 34670 25569 39593
rect 9448 18673 25649 34670
rect 9623 13520 25097 18673
rect 9448 13380 25649 13520
rect 9623 12330 25097 13380
rect 9448 12210 25649 12330
rect 9623 11160 25097 12210
rect 9448 11020 25649 11160
rect 9528 9942 25097 10138
rect 9448 8920 25649 9060
rect 9530 7830 25097 8920
rect 9448 7710 25649 7830
rect 9623 6860 25097 7710
rect 9448 6740 25649 6860
rect 9623 5890 25097 6740
rect 9448 5770 25649 5890
rect 9623 4680 25097 5770
rect 9448 4560 25649 4680
rect 9623 3470 24161 4560
rect 9448 3350 25649 3470
rect 9623 2500 24161 3350
rect 9448 2380 25649 2500
rect 9623 1290 25097 2380
rect 9448 1170 25649 1290
rect 9623 0 25097 1170
<< metal5 >>
rect 10810 20617 22978 32782
rect 0 13600 9543 18590
rect 0 12430 9543 13280
rect 0 11260 9543 12110
rect 25177 13600 33800 18590
rect 25177 12430 33800 13280
rect 25177 11260 33800 12110
rect 0 9140 9448 10940
rect 25177 9140 33800 10940
rect 0 7930 9543 8820
rect 0 6960 9543 7610
rect 0 5990 9543 6640
rect 0 4780 9543 5670
rect 0 3570 9543 4460
rect 25177 7930 33800 8820
rect 25177 6960 33800 7610
rect 25177 5990 33800 6640
rect 25177 4780 33800 5670
rect 25177 3570 33800 4460
rect 0 2600 9543 3250
rect 24241 2600 33800 3250
rect 0 1390 9543 2280
rect 0 20 9543 1070
rect 25177 1390 33800 2280
rect 25177 20 33800 1070
<< obsm5 >>
rect 0 33102 33800 39593
rect 0 20297 10490 33102
rect 23298 20297 33800 33102
rect 0 18910 33800 20297
rect 9863 10940 24857 18910
rect 9768 9140 24857 10940
rect 9863 3570 24857 9140
rect 9863 2280 23921 3570
rect 9863 20 24857 2280
<< labels >>
rlabel metal4 s 0 10218 33800 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 10218 254 10814 6 AMUXBUS_A
port 1 nsew signal bidirectional
rlabel metal4 s 0 9266 33800 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal4 s 0 9266 254 9862 6 AMUXBUS_B
port 2 nsew signal bidirectional
rlabel metal2 s 19478 -407 24258 4725 6 DRN_HVC
port 3 nsew power bidirectional
rlabel metal3 s 16978 -407 19178 1859 6 DRN_HVC
port 3 nsew power bidirectional
rlabel metal3 s 0 -407 14279 2730 6 P_CORE
port 4 nsew power bidirectional
rlabel metal3 s 19478 -407 33800 2730 6 P_CORE
port 4 nsew power bidirectional
rlabel metal5 s 10810 20617 22978 32782 6 P_PAD
port 5 nsew power bidirectional
rlabel metal2 s 9499 -407 14279 4 8 SRC_BDY_HVC
port 6 nsew ground bidirectional
rlabel metal3 s 14579 -407 16779 138 8 SRC_BDY_HVC
port 6 nsew ground bidirectional
rlabel metal5 s 25177 9140 33800 10940 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 25177 6960 33800 7610 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 25177 9922 33800 10158 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 10874 33800 10940 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 9140 33800 9206 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 25177 6940 33800 7630 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 9140 9448 10940 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 0 6960 9543 7610 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 9140 254 9206 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 9922 9448 10158 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 10874 254 10940 6 VSSA
port 7 nsew ground bidirectional
rlabel metal4 s 0 6940 9543 7630 6 VSSA
port 7 nsew ground bidirectional
rlabel metal5 s 24241 2600 33800 3250 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 24241 2580 33800 3270 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 2600 9543 3250 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 2580 9543 3270 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 25177 5990 33800 6640 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal4 s 25177 5970 33800 6660 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal5 s 0 5990 9543 6640 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal4 s 0 5970 9543 6660 6 VSWITCH
port 9 nsew power bidirectional
rlabel metal5 s 25177 12430 33800 13280 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 25177 12410 33800 13300 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 0 12430 9543 13280 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal4 s 0 12410 9543 13300 6 VDDIO_Q
port 10 nsew power bidirectional
rlabel metal5 s 25177 20 33800 1070 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 25177 0 33800 1090 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal5 s 0 20 9543 1070 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal4 s 0 0 9543 1090 6 VCCHIB
port 11 nsew power bidirectional
rlabel metal5 s 25177 13600 33800 18590 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 25177 3570 33800 4460 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 24241 3550 33800 4480 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 25177 13600 33800 18593 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 0 13600 9543 18590 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 0 3570 9543 4460 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 0 3550 9543 4480 6 VDDIO
port 12 nsew power bidirectional
rlabel metal4 s 0 13600 9543 18593 6 VDDIO
port 12 nsew power bidirectional
rlabel metal5 s 25177 1390 33800 2280 6 VCCD
port 13 nsew power bidirectional
rlabel metal4 s 25177 1370 33800 2300 6 VCCD
port 13 nsew power bidirectional
rlabel metal5 s 0 1390 9543 2280 6 VCCD
port 13 nsew power bidirectional
rlabel metal4 s 0 1370 9543 2300 6 VCCD
port 13 nsew power bidirectional
rlabel metal4 s 25649 34750 33800 39593 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 33672 37913 33674 37915 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal5 s 25177 4780 33800 5670 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 25177 4760 33800 5690 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 33546 34750 33800 39593 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 0 34750 9641 39593 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 126 37913 128 37915 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal5 s 0 4780 9543 5670 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 0 34750 254 39593 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal4 s 0 4760 9543 5690 6 VSSIO
port 14 nsew ground bidirectional
rlabel metal5 s 25177 7930 33800 8820 6 VSSD
port 15 nsew ground bidirectional
rlabel metal4 s 25177 7910 33800 8840 6 VSSD
port 15 nsew ground bidirectional
rlabel metal5 s 0 7930 9543 8820 6 VSSD
port 15 nsew ground bidirectional
rlabel metal4 s 0 7910 9450 8840 6 VSSD
port 15 nsew ground bidirectional
rlabel metal5 s 25177 11260 33800 12110 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal4 s 25177 11240 33800 12130 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal5 s 0 11260 9543 12110 6 VSSIO_Q
port 16 nsew ground bidirectional
rlabel metal4 s 0 11240 9543 12130 6 VSSIO_Q
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 33800 39593
string LEFclass PAD POWER
string LEFview TRUE
string GDS_END 2340684
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 2324050
<< end >>
