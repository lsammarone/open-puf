magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 98 157 800 203
rect 1 21 800 157
rect 30 -17 64 21
<< locali >>
rect 17 215 85 328
rect 187 283 444 340
rect 480 283 544 340
rect 187 181 221 283
rect 187 147 405 181
rect 200 57 266 147
rect 371 117 405 147
rect 507 199 544 283
rect 578 199 640 340
rect 371 51 418 117
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 408 69 444
rect 110 442 182 527
rect 284 442 350 527
rect 451 442 519 527
rect 704 442 811 485
rect 17 374 724 408
rect 17 362 153 374
rect 119 181 153 362
rect 17 147 153 181
rect 255 215 473 249
rect 17 58 69 147
rect 124 17 158 113
rect 439 178 473 215
rect 678 265 724 374
rect 678 199 736 265
rect 439 165 480 178
rect 770 165 811 442
rect 439 144 811 165
rect 450 131 811 144
rect 300 17 334 113
rect 452 17 518 97
rect 552 61 586 131
rect 732 121 811 131
rect 620 17 698 97
rect 732 61 783 121
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 507 199 544 283 6 A
port 1 nsew signal input
rlabel locali s 480 283 544 340 6 A
port 1 nsew signal input
rlabel locali s 578 199 640 340 6 B
port 2 nsew signal input
rlabel locali s 17 215 85 328 6 C_N
port 3 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 800 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 98 157 800 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 371 51 418 117 6 X
port 8 nsew signal output
rlabel locali s 371 117 405 147 6 X
port 8 nsew signal output
rlabel locali s 200 57 266 147 6 X
port 8 nsew signal output
rlabel locali s 187 147 405 181 6 X
port 8 nsew signal output
rlabel locali s 187 181 221 283 6 X
port 8 nsew signal output
rlabel locali s 187 283 444 340 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1045250
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1038816
<< end >>
