magic
tech sky130A
timestamp 1652772933
<< locali >>
rect 1258 2746 1380 2767
<< viali >>
rect 1488 3089 1505 3106
rect 1537 2749 1555 2768
rect 1488 2686 1507 2704
rect 1481 2468 1498 2486
<< metal1 >>
rect 1481 3114 1513 3116
rect 1481 3111 1484 3114
rect 1480 3088 1484 3111
rect 1510 3088 1513 3114
rect 1480 3085 1513 3088
rect 1481 3084 1513 3085
rect 1529 2768 1563 2775
rect 1529 2749 1537 2768
rect 1555 2749 1563 2768
rect 1529 2742 1563 2749
rect 1482 2709 1515 2712
rect 1482 2683 1486 2709
rect 1512 2683 1515 2709
rect 1482 2680 1515 2683
rect 1471 2490 1505 2494
rect 1471 2464 1475 2490
rect 1502 2464 1507 2490
rect 1471 2461 1505 2464
<< via1 >>
rect 1484 3106 1510 3114
rect 1484 3089 1488 3106
rect 1488 3089 1505 3106
rect 1505 3089 1510 3106
rect 1484 3088 1510 3089
rect 1486 2704 1512 2709
rect 1486 2686 1488 2704
rect 1488 2686 1507 2704
rect 1507 2686 1512 2704
rect 1486 2683 1512 2686
rect 1475 2486 1502 2490
rect 1475 2468 1481 2486
rect 1481 2468 1498 2486
rect 1498 2468 1502 2486
rect 1475 2464 1502 2468
<< metal2 >>
rect 1481 3114 1513 3116
rect 1481 3088 1484 3114
rect 1510 3088 1513 3114
rect 1481 3084 1513 3088
rect 1481 2712 1496 3084
rect 1481 2709 1515 2712
rect 1481 2694 1486 2709
rect 1482 2683 1486 2694
rect 1512 2683 1515 2709
rect 1482 2680 1515 2683
rect 1482 2494 1496 2680
rect 1471 2490 1505 2494
rect 1471 2464 1475 2490
rect 1502 2464 1505 2490
rect 1471 2461 1505 2464
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 1176 0 1 2638
box -19 -24 157 296
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 1342 0 1 2637
box -19 -24 249 296
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 1172 0 -1 3218
box -19 -24 433 296
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_1
timestamp 1650294714
transform 1 0 1170 0 -1 2597
box -19 -24 433 296
<< end >>
