/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/r+c/res_high__cap_high__lin.spice