magic
tech sky130A
magscale 1 2
timestamp 1654197755
<< nwell >>
rect 684 6800 910 6838
rect 588 6678 910 6800
rect 262 6607 1126 6678
rect 2572 6800 2798 6838
rect 2476 6678 2798 6800
rect 2150 6607 3014 6678
rect 4460 6800 4686 6838
rect 4364 6678 4686 6800
rect 4038 6607 4902 6678
rect 6348 6800 6574 6838
rect 6252 6678 6574 6800
rect 5926 6607 6790 6678
rect 8236 6800 8462 6838
rect 8140 6678 8462 6800
rect 7814 6607 8678 6678
rect 10124 6800 10350 6838
rect 10028 6678 10350 6800
rect 9702 6607 10566 6678
rect 12012 6800 12238 6838
rect 11916 6678 12238 6800
rect 11590 6607 12454 6678
rect 13900 6800 14126 6838
rect 13804 6678 14126 6800
rect 13478 6607 14342 6678
rect 15782 6800 16008 6838
rect 15686 6678 16008 6800
rect 15360 6607 16224 6678
rect 17670 6800 17896 6838
rect 17574 6678 17896 6800
rect 17248 6607 18112 6678
rect 19558 6800 19784 6838
rect 19462 6678 19784 6800
rect 19136 6607 20000 6678
rect 21446 6800 21672 6838
rect 21350 6678 21672 6800
rect 21024 6607 21888 6678
rect 23334 6800 23560 6838
rect 23238 6678 23560 6800
rect 22912 6607 23776 6678
rect 25222 6800 25448 6838
rect 25126 6678 25448 6800
rect 24800 6607 25664 6678
rect 27110 6800 27336 6838
rect 27014 6678 27336 6800
rect 26688 6607 27552 6678
rect 28998 6800 29224 6838
rect 28902 6678 29224 6800
rect 28576 6607 29440 6678
rect 30886 6800 31112 6838
rect 30790 6678 31112 6800
rect 30464 6607 31328 6678
rect 32774 6800 33000 6838
rect 32678 6678 33000 6800
rect 32352 6607 33216 6678
rect 34662 6800 34888 6838
rect 34566 6678 34888 6800
rect 34240 6607 35104 6678
rect 36550 6800 36776 6838
rect 36454 6678 36776 6800
rect 36128 6607 36992 6678
rect 38438 6800 38664 6838
rect 38342 6678 38664 6800
rect 38016 6607 38880 6678
rect 40326 6800 40552 6838
rect 40230 6678 40552 6800
rect 39904 6607 40768 6678
rect 42214 6800 42440 6838
rect 42118 6678 42440 6800
rect 41792 6607 42656 6678
rect 44102 6800 44328 6838
rect 44006 6678 44328 6800
rect 43680 6607 44544 6678
rect 45984 6800 46210 6838
rect 45888 6678 46210 6800
rect 45562 6607 46426 6678
rect 47872 6800 48098 6838
rect 47776 6678 48098 6800
rect 47450 6607 48314 6678
rect 49760 6800 49986 6838
rect 49664 6678 49986 6800
rect 49338 6607 50202 6678
rect 51648 6800 51874 6838
rect 51552 6678 51874 6800
rect 51226 6607 52090 6678
rect 53536 6800 53762 6838
rect 53440 6678 53762 6800
rect 53114 6607 53978 6678
rect 55424 6800 55650 6838
rect 55328 6678 55650 6800
rect 55002 6607 55866 6678
rect 57312 6800 57538 6838
rect 57216 6678 57538 6800
rect 56890 6607 57754 6678
rect 59200 6800 59426 6838
rect 59104 6678 59426 6800
rect 58778 6607 59642 6678
rect 262 6601 1464 6607
rect 2150 6601 3352 6607
rect 4038 6601 5240 6607
rect 5926 6601 7128 6607
rect 7814 6601 9016 6607
rect 9702 6601 10904 6607
rect 11590 6601 12792 6607
rect 13478 6601 14680 6607
rect 15360 6601 16562 6607
rect 17248 6601 18450 6607
rect 19136 6601 20338 6607
rect 21024 6601 22226 6607
rect 22912 6601 24114 6607
rect 24800 6601 26002 6607
rect 26688 6601 27890 6607
rect 28576 6601 29778 6607
rect 30464 6601 31666 6607
rect 32352 6601 33554 6607
rect 34240 6601 35442 6607
rect 36128 6601 37330 6607
rect 38016 6601 39218 6607
rect 39904 6601 41106 6607
rect 41792 6601 42994 6607
rect 43680 6601 44882 6607
rect 45562 6601 46764 6607
rect 47450 6601 48652 6607
rect 49338 6601 50540 6607
rect 51226 6601 52428 6607
rect 53114 6601 54316 6607
rect 55002 6601 56204 6607
rect 56890 6601 58092 6607
rect -430 6599 -78 6601
rect 262 6599 1810 6601
rect 2150 6599 3698 6601
rect 4038 6599 5586 6601
rect 5926 6599 7474 6601
rect 7814 6599 9362 6601
rect 9702 6599 11250 6601
rect 11590 6599 13138 6601
rect 13478 6599 15020 6601
rect 15360 6599 16908 6601
rect 17248 6599 18796 6601
rect 19136 6599 20684 6601
rect 21024 6599 22572 6601
rect 22912 6599 24460 6601
rect 24800 6599 26348 6601
rect 26688 6599 28236 6601
rect 28576 6599 30124 6601
rect 30464 6599 32012 6601
rect 32352 6599 33900 6601
rect 34240 6599 35788 6601
rect 36128 6599 37676 6601
rect 38016 6599 39564 6601
rect 39904 6599 41452 6601
rect 41792 6599 43340 6601
rect 43680 6599 45222 6601
rect 45562 6599 47110 6601
rect 47450 6599 48998 6601
rect 49338 6599 50886 6601
rect 51226 6599 52774 6601
rect 53114 6599 54662 6601
rect 55002 6599 56550 6601
rect 56890 6599 58438 6601
rect 58778 6599 59980 6607
rect -430 6286 59980 6599
rect -430 6280 1126 6286
rect 1458 6280 3014 6286
rect 3346 6280 4902 6286
rect 5234 6280 6790 6286
rect 7122 6280 8678 6286
rect 9010 6280 10566 6286
rect 10898 6280 12454 6286
rect 12786 6280 14342 6286
rect 14668 6280 16224 6286
rect 16556 6280 18112 6286
rect 18444 6280 20000 6286
rect 20332 6280 21888 6286
rect 22220 6280 23776 6286
rect 24108 6280 25664 6286
rect 25996 6280 27552 6286
rect 27884 6280 29440 6286
rect 29772 6280 31328 6286
rect 31660 6280 33216 6286
rect 33548 6280 35104 6286
rect 35436 6280 36992 6286
rect 37324 6280 38880 6286
rect 39212 6280 40768 6286
rect 41100 6280 42656 6286
rect 42988 6280 44544 6286
rect 44870 6280 46426 6286
rect 46758 6280 48314 6286
rect 48646 6280 50202 6286
rect 50534 6280 52090 6286
rect 52422 6280 53978 6286
rect 54310 6280 55866 6286
rect 56198 6280 57754 6286
rect 58086 6280 59642 6286
rect -84 6278 1126 6280
rect 1804 6278 3014 6280
rect 3692 6278 4902 6280
rect 5580 6278 6790 6280
rect 7468 6278 8678 6280
rect 9356 6278 10566 6280
rect 11244 6278 12454 6280
rect 13132 6278 14342 6280
rect 15014 6278 16224 6280
rect 16902 6278 18112 6280
rect 18790 6278 20000 6280
rect 20678 6278 21888 6280
rect 22566 6278 23776 6280
rect 24454 6278 25664 6280
rect 26342 6278 27552 6280
rect 28230 6278 29440 6280
rect 30118 6278 31328 6280
rect 32006 6278 33216 6280
rect 33894 6278 35104 6280
rect 35782 6278 36992 6280
rect 37670 6278 38880 6280
rect 39558 6278 40768 6280
rect 41446 6278 42656 6280
rect 43334 6278 44544 6280
rect 45216 6278 46426 6280
rect 47104 6278 48314 6280
rect 48992 6278 50202 6280
rect 50880 6278 52090 6280
rect 52768 6278 53978 6280
rect 54656 6278 55866 6280
rect 56544 6278 57754 6280
rect 58432 6278 59642 6280
rect 682 5744 908 5782
rect 586 5556 908 5744
rect 2570 5744 2796 5782
rect 2474 5556 2796 5744
rect 4458 5744 4684 5782
rect 4362 5556 4684 5744
rect 6346 5744 6572 5782
rect 6250 5556 6572 5744
rect 8234 5744 8460 5782
rect 8138 5556 8460 5744
rect 10122 5744 10348 5782
rect 10026 5556 10348 5744
rect 12010 5744 12236 5782
rect 11914 5556 12236 5744
rect 13898 5744 14124 5782
rect 13802 5556 14124 5744
rect 15780 5744 16006 5782
rect 15684 5556 16006 5744
rect 17668 5744 17894 5782
rect 17572 5556 17894 5744
rect 19556 5744 19782 5782
rect 19460 5556 19782 5744
rect 21444 5744 21670 5782
rect 21348 5556 21670 5744
rect 23332 5744 23558 5782
rect 23236 5556 23558 5744
rect 25220 5744 25446 5782
rect 25124 5556 25446 5744
rect 27108 5744 27334 5782
rect 27012 5556 27334 5744
rect 28996 5744 29222 5782
rect 28900 5556 29222 5744
rect 30884 5744 31110 5782
rect 30788 5556 31110 5744
rect 32772 5744 32998 5782
rect 32676 5556 32998 5744
rect 34660 5744 34886 5782
rect 34564 5556 34886 5744
rect 36548 5744 36774 5782
rect 36452 5556 36774 5744
rect 38436 5744 38662 5782
rect 38340 5556 38662 5744
rect 40324 5744 40550 5782
rect 40228 5556 40550 5744
rect 42212 5744 42438 5782
rect 42116 5556 42438 5744
rect 44100 5744 44326 5782
rect 44004 5556 44326 5744
rect 45982 5744 46208 5782
rect 45886 5556 46208 5744
rect 47870 5744 48096 5782
rect 47774 5556 48096 5744
rect 49758 5744 49984 5782
rect 49662 5556 49984 5744
rect 51646 5744 51872 5782
rect 51550 5556 51872 5744
rect 53534 5744 53760 5782
rect 53438 5556 53760 5744
rect 55422 5744 55648 5782
rect 55326 5556 55648 5744
rect 57310 5744 57536 5782
rect 57214 5556 57536 5744
rect 59198 5744 59424 5782
rect 59102 5556 59424 5744
rect 120 5222 1288 5556
rect 2008 5222 3176 5556
rect 3896 5222 5064 5556
rect 5784 5230 6952 5556
rect 5626 4909 7174 5230
rect 7672 5228 8840 5556
rect 7508 4907 9056 5228
rect 9560 5222 10728 5556
rect 11448 5222 12616 5556
rect 13336 5222 14504 5556
rect 15218 5222 16386 5556
rect 17106 5222 18274 5556
rect 18994 5222 20162 5556
rect 20882 5230 22050 5556
rect 15460 3777 15956 5222
rect 20724 4909 22272 5230
rect 22770 5228 23938 5556
rect 22606 4907 24154 5228
rect 24658 5222 25826 5556
rect 26546 5222 27714 5556
rect 28434 5222 29602 5556
rect 30322 5222 31490 5556
rect 32210 5222 33378 5556
rect 34098 5222 35266 5556
rect 35986 5230 37154 5556
rect 30782 4153 31162 5222
rect 35828 4909 37376 5230
rect 37874 5228 39042 5556
rect 37710 4907 39258 5228
rect 39762 5222 40930 5556
rect 41650 5222 42818 5556
rect 43538 5222 44706 5556
rect 45420 5222 46588 5556
rect 47308 5222 48476 5556
rect 49196 5222 50364 5556
rect 51084 5230 52252 5556
rect 29989 4152 32065 4153
rect 29989 3832 32102 4152
rect 45704 3937 46200 5222
rect 50926 4909 52474 5230
rect 52972 5228 54140 5556
rect 52808 4907 54356 5228
rect 54860 5222 56028 5556
rect 56748 5222 57916 5556
rect 58636 5222 59804 5556
rect 13201 3456 16679 3777
rect 43343 3616 46821 3937
rect 178 1884 1346 2218
rect 2066 1884 3234 2218
rect 3954 1884 5122 2218
rect 5626 2212 7174 2533
rect 5842 1884 7010 2212
rect 7508 2210 9056 2531
rect 7730 1884 8898 2210
rect 9618 1884 10786 2218
rect 11506 1884 12674 2218
rect 13394 1884 14562 2218
rect 15276 1884 16444 2218
rect 17164 1884 18332 2218
rect 19052 1884 20220 2218
rect 20724 2212 22272 2533
rect 20940 1884 22108 2212
rect 22606 2210 24154 2531
rect 22828 1884 23996 2210
rect 24716 1884 25884 2218
rect 26604 1884 27772 2218
rect 28492 1884 29660 2218
rect 30380 1884 31548 2218
rect 32268 1884 33436 2218
rect 34156 1884 35324 2218
rect 35828 2212 37376 2533
rect 36044 1884 37212 2212
rect 37710 2210 39258 2531
rect 37932 1884 39100 2210
rect 39820 1884 40988 2218
rect 41708 1884 42876 2218
rect 43596 1884 44764 2218
rect 45478 1884 46646 2218
rect 47366 1884 48534 2218
rect 49254 1884 50422 2218
rect 50926 2212 52474 2533
rect 51142 1884 52310 2212
rect 52808 2210 54356 2531
rect 53030 1884 54198 2210
rect 54918 1884 56086 2218
rect 56806 1884 57974 2218
rect 58694 1884 59862 2218
rect 558 1696 880 1884
rect 558 1658 784 1696
rect 2446 1696 2768 1884
rect 2446 1658 2672 1696
rect 4334 1696 4656 1884
rect 4334 1658 4560 1696
rect 6222 1696 6544 1884
rect 6222 1658 6448 1696
rect 8110 1696 8432 1884
rect 8110 1658 8336 1696
rect 9998 1696 10320 1884
rect 9998 1658 10224 1696
rect 11886 1696 12208 1884
rect 11886 1658 12112 1696
rect 13774 1696 14096 1884
rect 13774 1658 14000 1696
rect 15656 1696 15978 1884
rect 15656 1658 15882 1696
rect 17544 1696 17866 1884
rect 17544 1658 17770 1696
rect 19432 1696 19754 1884
rect 19432 1658 19658 1696
rect 21320 1696 21642 1884
rect 21320 1658 21546 1696
rect 23208 1696 23530 1884
rect 23208 1658 23434 1696
rect 25096 1696 25418 1884
rect 25096 1658 25322 1696
rect 26984 1696 27306 1884
rect 26984 1658 27210 1696
rect 28872 1696 29194 1884
rect 28872 1658 29098 1696
rect 30760 1696 31082 1884
rect 30760 1658 30986 1696
rect 32648 1696 32970 1884
rect 32648 1658 32874 1696
rect 34536 1696 34858 1884
rect 34536 1658 34762 1696
rect 36424 1696 36746 1884
rect 36424 1658 36650 1696
rect 38312 1696 38634 1884
rect 38312 1658 38538 1696
rect 40200 1696 40522 1884
rect 40200 1658 40426 1696
rect 42088 1696 42410 1884
rect 42088 1658 42314 1696
rect 43976 1696 44298 1884
rect 43976 1658 44202 1696
rect 45858 1696 46180 1884
rect 45858 1658 46084 1696
rect 47746 1696 48068 1884
rect 47746 1658 47972 1696
rect 49634 1696 49956 1884
rect 49634 1658 49860 1696
rect 51522 1696 51844 1884
rect 51522 1658 51748 1696
rect 53410 1696 53732 1884
rect 53410 1658 53636 1696
rect 55298 1696 55620 1884
rect 55298 1658 55524 1696
rect 57186 1696 57508 1884
rect 57186 1658 57412 1696
rect 59074 1696 59396 1884
rect 59074 1658 59300 1696
rect 340 1160 1550 1162
rect 2228 1160 3438 1162
rect 4116 1160 5326 1162
rect 6004 1160 7214 1162
rect 7892 1160 9102 1162
rect 9780 1160 10990 1162
rect 11668 1160 12878 1162
rect 13556 1160 14766 1162
rect 15438 1160 16648 1162
rect 17326 1160 18536 1162
rect 19214 1160 20424 1162
rect 21102 1160 22312 1162
rect 22990 1160 24200 1162
rect 24878 1160 26088 1162
rect 26766 1160 27976 1162
rect 28654 1160 29864 1162
rect 30542 1160 31752 1162
rect 32430 1160 33640 1162
rect 34318 1160 35528 1162
rect 36206 1160 37416 1162
rect 38094 1160 39304 1162
rect 39982 1160 41192 1162
rect 41870 1160 43080 1162
rect 43758 1160 44968 1162
rect 45640 1160 46850 1162
rect 47528 1160 48738 1162
rect 49416 1160 50626 1162
rect 51304 1160 52514 1162
rect 53192 1160 54402 1162
rect 55080 1160 56290 1162
rect 56968 1160 58178 1162
rect 58856 1160 60066 1162
rect 340 1154 1896 1160
rect 2228 1154 3784 1160
rect 4116 1154 5672 1160
rect 6004 1154 7560 1160
rect 7892 1154 9448 1160
rect 9780 1154 11336 1160
rect 11668 1154 13224 1160
rect 13556 1154 15112 1160
rect 15438 1154 16994 1160
rect 17326 1154 18882 1160
rect 19214 1154 20770 1160
rect 21102 1154 22658 1160
rect 22990 1154 24546 1160
rect 24878 1154 26434 1160
rect 26766 1154 28322 1160
rect 28654 1154 30210 1160
rect 30542 1154 32098 1160
rect 32430 1154 33986 1160
rect 34318 1154 35874 1160
rect 36206 1154 37762 1160
rect 38094 1154 39650 1160
rect 39982 1154 41538 1160
rect 41870 1154 43426 1160
rect 43758 1154 45314 1160
rect 45640 1154 47196 1160
rect 47528 1154 49084 1160
rect 49416 1154 50972 1160
rect 51304 1154 52860 1160
rect 53192 1154 54748 1160
rect 55080 1154 56636 1160
rect 56968 1154 58524 1160
rect 58856 1154 60412 1160
rect 2 841 60412 1154
rect 2 833 1204 841
rect 1544 839 3092 841
rect 3432 839 4980 841
rect 5320 839 6868 841
rect 7208 839 8756 841
rect 9096 839 10644 841
rect 10984 839 12532 841
rect 12872 839 14420 841
rect 14760 839 16302 841
rect 16642 839 18190 841
rect 18530 839 20078 841
rect 20418 839 21966 841
rect 22306 839 23854 841
rect 24194 839 25742 841
rect 26082 839 27630 841
rect 27970 839 29518 841
rect 29858 839 31406 841
rect 31746 839 33294 841
rect 33634 839 35182 841
rect 35522 839 37070 841
rect 37410 839 38958 841
rect 39298 839 40846 841
rect 41186 839 42734 841
rect 43074 839 44622 841
rect 44962 839 46504 841
rect 46844 839 48392 841
rect 48732 839 50280 841
rect 50620 839 52168 841
rect 52508 839 54056 841
rect 54396 839 55944 841
rect 56284 839 57832 841
rect 58172 839 59720 841
rect 60060 839 60412 841
rect 1890 833 3092 839
rect 3778 833 4980 839
rect 5666 833 6868 839
rect 7554 833 8756 839
rect 9442 833 10644 839
rect 11330 833 12532 839
rect 13218 833 14420 839
rect 15100 833 16302 839
rect 16988 833 18190 839
rect 18876 833 20078 839
rect 20764 833 21966 839
rect 22652 833 23854 839
rect 24540 833 25742 839
rect 26428 833 27630 839
rect 28316 833 29518 839
rect 30204 833 31406 839
rect 32092 833 33294 839
rect 33980 833 35182 839
rect 35868 833 37070 839
rect 37756 833 38958 839
rect 39644 833 40846 839
rect 41532 833 42734 839
rect 43420 833 44622 839
rect 45302 833 46504 839
rect 47190 833 48392 839
rect 49078 833 50280 839
rect 50966 833 52168 839
rect 52854 833 54056 839
rect 54742 833 55944 839
rect 56630 833 57832 839
rect 58518 833 59720 839
rect 340 762 1204 833
rect 556 640 878 762
rect 556 602 782 640
rect 2228 762 3092 833
rect 2444 640 2766 762
rect 2444 602 2670 640
rect 4116 762 4980 833
rect 4332 640 4654 762
rect 4332 602 4558 640
rect 6004 762 6868 833
rect 6220 640 6542 762
rect 6220 602 6446 640
rect 7892 762 8756 833
rect 8108 640 8430 762
rect 8108 602 8334 640
rect 9780 762 10644 833
rect 9996 640 10318 762
rect 9996 602 10222 640
rect 11668 762 12532 833
rect 11884 640 12206 762
rect 11884 602 12110 640
rect 13556 762 14420 833
rect 13772 640 14094 762
rect 13772 602 13998 640
rect 15438 762 16302 833
rect 15654 640 15976 762
rect 15654 602 15880 640
rect 17326 762 18190 833
rect 17542 640 17864 762
rect 17542 602 17768 640
rect 19214 762 20078 833
rect 19430 640 19752 762
rect 19430 602 19656 640
rect 21102 762 21966 833
rect 21318 640 21640 762
rect 21318 602 21544 640
rect 22990 762 23854 833
rect 23206 640 23528 762
rect 23206 602 23432 640
rect 24878 762 25742 833
rect 25094 640 25416 762
rect 25094 602 25320 640
rect 26766 762 27630 833
rect 26982 640 27304 762
rect 26982 602 27208 640
rect 28654 762 29518 833
rect 28870 640 29192 762
rect 28870 602 29096 640
rect 30542 762 31406 833
rect 30758 640 31080 762
rect 30758 602 30984 640
rect 32430 762 33294 833
rect 32646 640 32968 762
rect 32646 602 32872 640
rect 34318 762 35182 833
rect 34534 640 34856 762
rect 34534 602 34760 640
rect 36206 762 37070 833
rect 36422 640 36744 762
rect 36422 602 36648 640
rect 38094 762 38958 833
rect 38310 640 38632 762
rect 38310 602 38536 640
rect 39982 762 40846 833
rect 40198 640 40520 762
rect 40198 602 40424 640
rect 41870 762 42734 833
rect 42086 640 42408 762
rect 42086 602 42312 640
rect 43758 762 44622 833
rect 43974 640 44296 762
rect 43974 602 44200 640
rect 45640 762 46504 833
rect 45856 640 46178 762
rect 45856 602 46082 640
rect 47528 762 48392 833
rect 47744 640 48066 762
rect 47744 602 47970 640
rect 49416 762 50280 833
rect 49632 640 49954 762
rect 49632 602 49858 640
rect 51304 762 52168 833
rect 51520 640 51842 762
rect 51520 602 51746 640
rect 53192 762 54056 833
rect 53408 640 53730 762
rect 53408 602 53634 640
rect 55080 762 55944 833
rect 55296 640 55618 762
rect 55296 602 55522 640
rect 56968 762 57832 833
rect 57184 640 57506 762
rect 57184 602 57410 640
rect 58856 762 59720 833
rect 59072 640 59394 762
rect 59072 602 59298 640
<< pwell >>
rect 628 7178 840 7278
rect 2516 7178 2728 7278
rect 4404 7178 4616 7278
rect 6292 7178 6504 7278
rect 8180 7178 8392 7278
rect 10068 7178 10280 7278
rect 11956 7178 12168 7278
rect 13844 7178 14056 7278
rect 15726 7178 15938 7278
rect 17614 7178 17826 7278
rect 19502 7178 19714 7278
rect 21390 7178 21602 7278
rect 23278 7178 23490 7278
rect 25166 7178 25378 7278
rect 27054 7178 27266 7278
rect 28942 7178 29154 7278
rect 30830 7178 31042 7278
rect 32718 7178 32930 7278
rect 34606 7178 34818 7278
rect 36494 7178 36706 7278
rect 38382 7178 38594 7278
rect 40270 7178 40482 7278
rect 42158 7178 42370 7278
rect 44046 7178 44258 7278
rect 45928 7178 46140 7278
rect 47816 7178 48028 7278
rect 49704 7178 49916 7278
rect 51592 7178 51804 7278
rect 53480 7178 53692 7278
rect 55368 7178 55580 7278
rect 57256 7178 57468 7278
rect 59144 7178 59356 7278
rect 582 6912 884 7094
rect 2470 6912 2772 7094
rect 4358 6912 4660 7094
rect 6246 6912 6548 7094
rect 8134 6912 8436 7094
rect 10022 6912 10324 7094
rect 11910 6912 12212 7094
rect 13798 6912 14100 7094
rect 15680 6912 15982 7094
rect 17568 6912 17870 7094
rect 19456 6912 19758 7094
rect 21344 6912 21646 7094
rect 23232 6912 23534 7094
rect 25120 6912 25422 7094
rect 27008 6912 27310 7094
rect 28896 6912 29198 7094
rect 30784 6912 31086 7094
rect 32672 6912 32974 7094
rect 34560 6912 34862 7094
rect 36448 6912 36750 7094
rect 38336 6912 38638 7094
rect 40224 6912 40526 7094
rect 42112 6912 42414 7094
rect 44000 6912 44302 7094
rect 45882 6912 46184 7094
rect 47770 6912 48072 7094
rect 49658 6912 49960 7094
rect 51546 6912 51848 7094
rect 53434 6912 53736 7094
rect 55322 6912 55624 7094
rect 57210 6912 57512 7094
rect 59098 6912 59400 7094
rect -391 6685 -117 6841
rect 2 6657 188 6839
rect 1198 6665 1384 6847
rect 1497 6685 1771 6841
rect 1890 6657 2076 6839
rect 3086 6665 3272 6847
rect 3385 6685 3659 6841
rect 3778 6657 3964 6839
rect 4974 6665 5160 6847
rect 5273 6685 5547 6841
rect 5666 6657 5852 6839
rect 6862 6665 7048 6847
rect 7161 6685 7435 6841
rect 7554 6657 7740 6839
rect 8750 6665 8936 6847
rect 9049 6685 9323 6841
rect 9442 6657 9628 6839
rect 10638 6665 10824 6847
rect 10937 6685 11211 6841
rect 11330 6657 11516 6839
rect 12526 6665 12712 6847
rect 12825 6685 13099 6841
rect 13218 6657 13404 6839
rect 14414 6665 14600 6847
rect 14707 6685 14981 6841
rect 15100 6657 15286 6839
rect 16296 6665 16482 6847
rect 16595 6685 16869 6841
rect 16988 6657 17174 6839
rect 18184 6665 18370 6847
rect 18483 6685 18757 6841
rect 18876 6657 19062 6839
rect 20072 6665 20258 6847
rect 20371 6685 20645 6841
rect 20764 6657 20950 6839
rect 21960 6665 22146 6847
rect 22259 6685 22533 6841
rect 22652 6657 22838 6839
rect 23848 6665 24034 6847
rect 24147 6685 24421 6841
rect 24540 6657 24726 6839
rect 25736 6665 25922 6847
rect 26035 6685 26309 6841
rect 26428 6657 26614 6839
rect 27624 6665 27810 6847
rect 27923 6685 28197 6841
rect 28316 6657 28502 6839
rect 29512 6665 29698 6847
rect 29811 6685 30085 6841
rect 30204 6657 30390 6839
rect 31400 6665 31586 6847
rect 31699 6685 31973 6841
rect 32092 6657 32278 6839
rect 33288 6665 33474 6847
rect 33587 6685 33861 6841
rect 33980 6657 34166 6839
rect 35176 6665 35362 6847
rect 35475 6685 35749 6841
rect 35868 6657 36054 6839
rect 37064 6665 37250 6847
rect 37363 6685 37637 6841
rect 37756 6657 37942 6839
rect 38952 6665 39138 6847
rect 39251 6685 39525 6841
rect 39644 6657 39830 6839
rect 40840 6665 41026 6847
rect 41139 6685 41413 6841
rect 41532 6657 41718 6839
rect 42728 6665 42914 6847
rect 43027 6685 43301 6841
rect 43420 6657 43606 6839
rect 44616 6665 44802 6847
rect 44909 6685 45183 6841
rect 45302 6657 45488 6839
rect 46498 6665 46684 6847
rect 46797 6685 47071 6841
rect 47190 6657 47376 6839
rect 48386 6665 48572 6847
rect 48685 6685 48959 6841
rect 49078 6657 49264 6839
rect 50274 6665 50460 6847
rect 50573 6685 50847 6841
rect 50966 6657 51152 6839
rect 52162 6665 52348 6847
rect 52461 6685 52735 6841
rect 52854 6657 53040 6839
rect 54050 6665 54236 6847
rect 54349 6685 54623 6841
rect 54742 6657 54928 6839
rect 55938 6665 56124 6847
rect 56237 6685 56511 6841
rect 56630 6657 56816 6839
rect 57826 6665 58012 6847
rect 58125 6685 58399 6841
rect 58518 6657 58704 6839
rect 59714 6665 59900 6847
rect 626 6122 838 6222
rect 2514 6122 2726 6222
rect 4402 6122 4614 6222
rect 6290 6122 6502 6222
rect 8178 6122 8390 6222
rect 10066 6122 10278 6222
rect 11954 6122 12166 6222
rect 13842 6122 14054 6222
rect 15724 6122 15936 6222
rect 17612 6122 17824 6222
rect 19500 6122 19712 6222
rect 21388 6122 21600 6222
rect 23276 6122 23488 6222
rect 25164 6122 25376 6222
rect 27052 6122 27264 6222
rect 28940 6122 29152 6222
rect 30828 6122 31040 6222
rect 32716 6122 32928 6222
rect 34604 6122 34816 6222
rect 36492 6122 36704 6222
rect 38380 6122 38592 6222
rect 40268 6122 40480 6222
rect 42156 6122 42368 6222
rect 44044 6122 44256 6222
rect 45926 6122 46138 6222
rect 47814 6122 48026 6222
rect 49702 6122 49914 6222
rect 51590 6122 51802 6222
rect 53478 6122 53690 6222
rect 55366 6122 55578 6222
rect 57254 6122 57466 6222
rect 59142 6122 59354 6222
rect 580 5856 882 6038
rect 2468 5856 2770 6038
rect 4356 5856 4658 6038
rect 6244 5856 6546 6038
rect 8132 5856 8434 6038
rect 10020 5856 10322 6038
rect 11908 5856 12210 6038
rect 13796 5856 14098 6038
rect 15678 5856 15980 6038
rect 17566 5856 17868 6038
rect 19454 5856 19756 6038
rect 21342 5856 21644 6038
rect 23230 5856 23532 6038
rect 25118 5856 25420 6038
rect 27006 5856 27308 6038
rect 28894 5856 29196 6038
rect 30782 5856 31084 6038
rect 32670 5856 32972 6038
rect 34558 5856 34860 6038
rect 36446 5856 36748 6038
rect 38334 5856 38636 6038
rect 40222 5856 40524 6038
rect 42110 5856 42412 6038
rect 43998 5856 44300 6038
rect 45880 5856 46182 6038
rect 47768 5856 48070 6038
rect 49656 5856 49958 6038
rect 51544 5856 51846 6038
rect 53432 5856 53734 6038
rect 55320 5856 55622 6038
rect 57208 5856 57510 6038
rect 59096 5856 59398 6038
rect 163 5611 433 5793
rect 977 5611 1247 5793
rect 2051 5611 2321 5793
rect 2865 5611 3135 5793
rect 3939 5611 4209 5793
rect 4753 5611 5023 5793
rect 5827 5611 6097 5793
rect 6641 5611 6911 5793
rect 7715 5611 7985 5793
rect 8529 5611 8799 5793
rect 9603 5611 9873 5793
rect 10417 5611 10687 5793
rect 11491 5611 11761 5793
rect 12305 5611 12575 5793
rect 13379 5611 13649 5793
rect 14193 5611 14463 5793
rect 15261 5611 15531 5793
rect 16075 5611 16345 5793
rect 17149 5611 17419 5793
rect 17963 5611 18233 5793
rect 19037 5611 19307 5793
rect 19851 5611 20121 5793
rect 20925 5611 21195 5793
rect 21739 5611 22009 5793
rect 22813 5611 23083 5793
rect 23627 5611 23897 5793
rect 24701 5611 24971 5793
rect 25515 5611 25785 5793
rect 26589 5611 26859 5793
rect 27403 5611 27673 5793
rect 28477 5611 28747 5793
rect 29291 5611 29561 5793
rect 30365 5611 30635 5793
rect 31179 5611 31449 5793
rect 32253 5611 32523 5793
rect 33067 5611 33337 5793
rect 34141 5611 34411 5793
rect 34955 5611 35225 5793
rect 36029 5611 36299 5793
rect 36843 5611 37113 5793
rect 37917 5611 38187 5793
rect 38731 5611 39001 5793
rect 39805 5611 40075 5793
rect 40619 5611 40889 5793
rect 41693 5611 41963 5793
rect 42507 5611 42777 5793
rect 43581 5611 43851 5793
rect 44395 5611 44665 5793
rect 45463 5611 45733 5793
rect 46277 5611 46547 5793
rect 47351 5611 47621 5793
rect 48165 5611 48435 5793
rect 49239 5611 49509 5793
rect 50053 5611 50323 5793
rect 51127 5611 51397 5793
rect 51941 5611 52211 5793
rect 53015 5611 53285 5793
rect 53829 5611 54099 5793
rect 54903 5611 55173 5793
rect 55717 5611 55987 5793
rect 56791 5611 57061 5793
rect 57605 5611 57875 5793
rect 58679 5611 58949 5793
rect 59493 5611 59763 5793
rect 5676 4669 7122 4851
rect 7558 4667 9004 4849
rect 20774 4669 22220 4851
rect 22656 4667 24102 4849
rect 35878 4669 37324 4851
rect 37760 4667 39206 4849
rect 50976 4669 52422 4851
rect 52858 4667 54304 4849
rect 30038 3592 30476 3774
rect 30569 3592 32015 3774
rect 30056 3554 30090 3592
rect 13253 3216 14699 3398
rect 15183 3216 16629 3398
rect 43395 3376 44841 3558
rect 45325 3376 46771 3558
rect 5678 2591 7124 2773
rect 7560 2589 9006 2771
rect 20776 2591 22222 2773
rect 22658 2589 24104 2771
rect 35880 2591 37326 2773
rect 37762 2589 39208 2771
rect 50978 2591 52424 2773
rect 52860 2589 54306 2771
rect 219 1647 489 1829
rect 1033 1647 1303 1829
rect 2107 1647 2377 1829
rect 2921 1647 3191 1829
rect 3995 1647 4265 1829
rect 4809 1647 5079 1829
rect 5883 1647 6153 1829
rect 6697 1647 6967 1829
rect 7771 1647 8041 1829
rect 8585 1647 8855 1829
rect 9659 1647 9929 1829
rect 10473 1647 10743 1829
rect 11547 1647 11817 1829
rect 12361 1647 12631 1829
rect 13435 1647 13705 1829
rect 14249 1647 14519 1829
rect 15317 1647 15587 1829
rect 16131 1647 16401 1829
rect 17205 1647 17475 1829
rect 18019 1647 18289 1829
rect 19093 1647 19363 1829
rect 19907 1647 20177 1829
rect 20981 1647 21251 1829
rect 21795 1647 22065 1829
rect 22869 1647 23139 1829
rect 23683 1647 23953 1829
rect 24757 1647 25027 1829
rect 25571 1647 25841 1829
rect 26645 1647 26915 1829
rect 27459 1647 27729 1829
rect 28533 1647 28803 1829
rect 29347 1647 29617 1829
rect 30421 1647 30691 1829
rect 31235 1647 31505 1829
rect 32309 1647 32579 1829
rect 33123 1647 33393 1829
rect 34197 1647 34467 1829
rect 35011 1647 35281 1829
rect 36085 1647 36355 1829
rect 36899 1647 37169 1829
rect 37973 1647 38243 1829
rect 38787 1647 39057 1829
rect 39861 1647 40131 1829
rect 40675 1647 40945 1829
rect 41749 1647 42019 1829
rect 42563 1647 42833 1829
rect 43637 1647 43907 1829
rect 44451 1647 44721 1829
rect 45519 1647 45789 1829
rect 46333 1647 46603 1829
rect 47407 1647 47677 1829
rect 48221 1647 48491 1829
rect 49295 1647 49565 1829
rect 50109 1647 50379 1829
rect 51183 1647 51453 1829
rect 51997 1647 52267 1829
rect 53071 1647 53341 1829
rect 53885 1647 54155 1829
rect 54959 1647 55229 1829
rect 55773 1647 56043 1829
rect 56847 1647 57117 1829
rect 57661 1647 57931 1829
rect 58735 1647 59005 1829
rect 59549 1647 59819 1829
rect 584 1402 886 1584
rect 2472 1402 2774 1584
rect 4360 1402 4662 1584
rect 6248 1402 6550 1584
rect 8136 1402 8438 1584
rect 10024 1402 10326 1584
rect 11912 1402 12214 1584
rect 13800 1402 14102 1584
rect 15682 1402 15984 1584
rect 17570 1402 17872 1584
rect 19458 1402 19760 1584
rect 21346 1402 21648 1584
rect 23234 1402 23536 1584
rect 25122 1402 25424 1584
rect 27010 1402 27312 1584
rect 28898 1402 29200 1584
rect 30786 1402 31088 1584
rect 32674 1402 32976 1584
rect 34562 1402 34864 1584
rect 36450 1402 36752 1584
rect 38338 1402 38640 1584
rect 40226 1402 40528 1584
rect 42114 1402 42416 1584
rect 44002 1402 44304 1584
rect 45884 1402 46186 1584
rect 47772 1402 48074 1584
rect 49660 1402 49962 1584
rect 51548 1402 51850 1584
rect 53436 1402 53738 1584
rect 55324 1402 55626 1584
rect 57212 1402 57514 1584
rect 59100 1402 59402 1584
rect 628 1218 840 1318
rect 2516 1218 2728 1318
rect 4404 1218 4616 1318
rect 6292 1218 6504 1318
rect 8180 1218 8392 1318
rect 10068 1218 10280 1318
rect 11956 1218 12168 1318
rect 13844 1218 14056 1318
rect 15726 1218 15938 1318
rect 17614 1218 17826 1318
rect 19502 1218 19714 1318
rect 21390 1218 21602 1318
rect 23278 1218 23490 1318
rect 25166 1218 25378 1318
rect 27054 1218 27266 1318
rect 28942 1218 29154 1318
rect 30830 1218 31042 1318
rect 32718 1218 32930 1318
rect 34606 1218 34818 1318
rect 36494 1218 36706 1318
rect 38382 1218 38594 1318
rect 40270 1218 40482 1318
rect 42158 1218 42370 1318
rect 44046 1218 44258 1318
rect 45928 1218 46140 1318
rect 47816 1218 48028 1318
rect 49704 1218 49916 1318
rect 51592 1218 51804 1318
rect 53480 1218 53692 1318
rect 55368 1218 55580 1318
rect 57256 1218 57468 1318
rect 59144 1218 59356 1318
rect 82 593 268 775
rect 1278 601 1464 783
rect 1583 599 1857 755
rect 1970 593 2156 775
rect 3166 601 3352 783
rect 3471 599 3745 755
rect 3858 593 4044 775
rect 5054 601 5240 783
rect 5359 599 5633 755
rect 5746 593 5932 775
rect 6942 601 7128 783
rect 7247 599 7521 755
rect 7634 593 7820 775
rect 8830 601 9016 783
rect 9135 599 9409 755
rect 9522 593 9708 775
rect 10718 601 10904 783
rect 11023 599 11297 755
rect 11410 593 11596 775
rect 12606 601 12792 783
rect 12911 599 13185 755
rect 13298 593 13484 775
rect 14494 601 14680 783
rect 14799 599 15073 755
rect 15180 593 15366 775
rect 16376 601 16562 783
rect 16681 599 16955 755
rect 17068 593 17254 775
rect 18264 601 18450 783
rect 18569 599 18843 755
rect 18956 593 19142 775
rect 20152 601 20338 783
rect 20457 599 20731 755
rect 20844 593 21030 775
rect 22040 601 22226 783
rect 22345 599 22619 755
rect 22732 593 22918 775
rect 23928 601 24114 783
rect 24233 599 24507 755
rect 24620 593 24806 775
rect 25816 601 26002 783
rect 26121 599 26395 755
rect 26508 593 26694 775
rect 27704 601 27890 783
rect 28009 599 28283 755
rect 28396 593 28582 775
rect 29592 601 29778 783
rect 29897 599 30171 755
rect 30284 593 30470 775
rect 31480 601 31666 783
rect 31785 599 32059 755
rect 32172 593 32358 775
rect 33368 601 33554 783
rect 33673 599 33947 755
rect 34060 593 34246 775
rect 35256 601 35442 783
rect 35561 599 35835 755
rect 35948 593 36134 775
rect 37144 601 37330 783
rect 37449 599 37723 755
rect 37836 593 38022 775
rect 39032 601 39218 783
rect 39337 599 39611 755
rect 39724 593 39910 775
rect 40920 601 41106 783
rect 41225 599 41499 755
rect 41612 593 41798 775
rect 42808 601 42994 783
rect 43113 599 43387 755
rect 43500 593 43686 775
rect 44696 601 44882 783
rect 45001 599 45275 755
rect 45382 593 45568 775
rect 46578 601 46764 783
rect 46883 599 47157 755
rect 47270 593 47456 775
rect 48466 601 48652 783
rect 48771 599 49045 755
rect 49158 593 49344 775
rect 50354 601 50540 783
rect 50659 599 50933 755
rect 51046 593 51232 775
rect 52242 601 52428 783
rect 52547 599 52821 755
rect 52934 593 53120 775
rect 54130 601 54316 783
rect 54435 599 54709 755
rect 54822 593 55008 775
rect 56018 601 56204 783
rect 56323 599 56597 755
rect 56710 593 56896 775
rect 57906 601 58092 783
rect 58211 599 58485 755
rect 58598 593 58784 775
rect 59794 601 59980 783
rect 60099 599 60373 755
rect 582 346 884 528
rect 2470 346 2772 528
rect 4358 346 4660 528
rect 6246 346 6548 528
rect 8134 346 8436 528
rect 10022 346 10324 528
rect 11910 346 12212 528
rect 13798 346 14100 528
rect 15680 346 15982 528
rect 17568 346 17870 528
rect 19456 346 19758 528
rect 21344 346 21646 528
rect 23232 346 23534 528
rect 25120 346 25422 528
rect 27008 346 27310 528
rect 28896 346 29198 528
rect 30784 346 31086 528
rect 32672 346 32974 528
rect 34560 346 34862 528
rect 36448 346 36750 528
rect 38336 346 38638 528
rect 40224 346 40526 528
rect 42112 346 42414 528
rect 44000 346 44302 528
rect 45882 346 46184 528
rect 47770 346 48072 528
rect 49658 346 49960 528
rect 51546 346 51848 528
rect 53434 346 53736 528
rect 55322 346 55624 528
rect 57210 346 57512 528
rect 59098 346 59400 528
rect 626 162 838 262
rect 2514 162 2726 262
rect 4402 162 4614 262
rect 6290 162 6502 262
rect 8178 162 8390 262
rect 10066 162 10278 262
rect 11954 162 12166 262
rect 13842 162 14054 262
rect 15724 162 15936 262
rect 17612 162 17824 262
rect 19500 162 19712 262
rect 21388 162 21600 262
rect 23276 162 23488 262
rect 25164 162 25376 262
rect 27052 162 27264 262
rect 28940 162 29152 262
rect 30828 162 31040 262
rect 32716 162 32928 262
rect 34604 162 34816 262
rect 36492 162 36704 262
rect 38380 162 38592 262
rect 40268 162 40480 262
rect 42156 162 42368 262
rect 44044 162 44256 262
rect 45926 162 46138 262
rect 47814 162 48026 262
rect 49702 162 49914 262
rect 51590 162 51802 262
rect 53478 162 53690 262
rect 55366 162 55578 262
rect 57254 162 57466 262
rect 59142 162 59354 262
<< nmos >>
rect 670 6938 700 7068
rect 766 6938 796 7068
rect 2558 6938 2588 7068
rect 2654 6938 2684 7068
rect 4446 6938 4476 7068
rect 4542 6938 4572 7068
rect 6334 6938 6364 7068
rect 6430 6938 6460 7068
rect 8222 6938 8252 7068
rect 8318 6938 8348 7068
rect 10110 6938 10140 7068
rect 10206 6938 10236 7068
rect 11998 6938 12028 7068
rect 12094 6938 12124 7068
rect 13886 6938 13916 7068
rect 13982 6938 14012 7068
rect 15768 6938 15798 7068
rect 15864 6938 15894 7068
rect 17656 6938 17686 7068
rect 17752 6938 17782 7068
rect 19544 6938 19574 7068
rect 19640 6938 19670 7068
rect 21432 6938 21462 7068
rect 21528 6938 21558 7068
rect 23320 6938 23350 7068
rect 23416 6938 23446 7068
rect 25208 6938 25238 7068
rect 25304 6938 25334 7068
rect 27096 6938 27126 7068
rect 27192 6938 27222 7068
rect 28984 6938 29014 7068
rect 29080 6938 29110 7068
rect 30872 6938 30902 7068
rect 30968 6938 30998 7068
rect 32760 6938 32790 7068
rect 32856 6938 32886 7068
rect 34648 6938 34678 7068
rect 34744 6938 34774 7068
rect 36536 6938 36566 7068
rect 36632 6938 36662 7068
rect 38424 6938 38454 7068
rect 38520 6938 38550 7068
rect 40312 6938 40342 7068
rect 40408 6938 40438 7068
rect 42200 6938 42230 7068
rect 42296 6938 42326 7068
rect 44088 6938 44118 7068
rect 44184 6938 44214 7068
rect 45970 6938 46000 7068
rect 46066 6938 46096 7068
rect 47858 6938 47888 7068
rect 47954 6938 47984 7068
rect 49746 6938 49776 7068
rect 49842 6938 49872 7068
rect 51634 6938 51664 7068
rect 51730 6938 51760 7068
rect 53522 6938 53552 7068
rect 53618 6938 53648 7068
rect 55410 6938 55440 7068
rect 55506 6938 55536 7068
rect 57298 6938 57328 7068
rect 57394 6938 57424 7068
rect 59186 6938 59216 7068
rect 59282 6938 59312 7068
rect 668 5882 698 6012
rect 764 5882 794 6012
rect 2556 5882 2586 6012
rect 2652 5882 2682 6012
rect 4444 5882 4474 6012
rect 4540 5882 4570 6012
rect 6332 5882 6362 6012
rect 6428 5882 6458 6012
rect 8220 5882 8250 6012
rect 8316 5882 8346 6012
rect 10108 5882 10138 6012
rect 10204 5882 10234 6012
rect 11996 5882 12026 6012
rect 12092 5882 12122 6012
rect 13884 5882 13914 6012
rect 13980 5882 14010 6012
rect 15766 5882 15796 6012
rect 15862 5882 15892 6012
rect 17654 5882 17684 6012
rect 17750 5882 17780 6012
rect 19542 5882 19572 6012
rect 19638 5882 19668 6012
rect 21430 5882 21460 6012
rect 21526 5882 21556 6012
rect 23318 5882 23348 6012
rect 23414 5882 23444 6012
rect 25206 5882 25236 6012
rect 25302 5882 25332 6012
rect 27094 5882 27124 6012
rect 27190 5882 27220 6012
rect 28982 5882 29012 6012
rect 29078 5882 29108 6012
rect 30870 5882 30900 6012
rect 30966 5882 30996 6012
rect 32758 5882 32788 6012
rect 32854 5882 32884 6012
rect 34646 5882 34676 6012
rect 34742 5882 34772 6012
rect 36534 5882 36564 6012
rect 36630 5882 36660 6012
rect 38422 5882 38452 6012
rect 38518 5882 38548 6012
rect 40310 5882 40340 6012
rect 40406 5882 40436 6012
rect 42198 5882 42228 6012
rect 42294 5882 42324 6012
rect 44086 5882 44116 6012
rect 44182 5882 44212 6012
rect 45968 5882 45998 6012
rect 46064 5882 46094 6012
rect 47856 5882 47886 6012
rect 47952 5882 47982 6012
rect 49744 5882 49774 6012
rect 49840 5882 49870 6012
rect 51632 5882 51662 6012
rect 51728 5882 51758 6012
rect 53520 5882 53550 6012
rect 53616 5882 53646 6012
rect 55408 5882 55438 6012
rect 55504 5882 55534 6012
rect 57296 5882 57326 6012
rect 57392 5882 57422 6012
rect 59184 5882 59214 6012
rect 59280 5882 59310 6012
rect 672 1428 702 1558
rect 768 1428 798 1558
rect 2560 1428 2590 1558
rect 2656 1428 2686 1558
rect 4448 1428 4478 1558
rect 4544 1428 4574 1558
rect 6336 1428 6366 1558
rect 6432 1428 6462 1558
rect 8224 1428 8254 1558
rect 8320 1428 8350 1558
rect 10112 1428 10142 1558
rect 10208 1428 10238 1558
rect 12000 1428 12030 1558
rect 12096 1428 12126 1558
rect 13888 1428 13918 1558
rect 13984 1428 14014 1558
rect 15770 1428 15800 1558
rect 15866 1428 15896 1558
rect 17658 1428 17688 1558
rect 17754 1428 17784 1558
rect 19546 1428 19576 1558
rect 19642 1428 19672 1558
rect 21434 1428 21464 1558
rect 21530 1428 21560 1558
rect 23322 1428 23352 1558
rect 23418 1428 23448 1558
rect 25210 1428 25240 1558
rect 25306 1428 25336 1558
rect 27098 1428 27128 1558
rect 27194 1428 27224 1558
rect 28986 1428 29016 1558
rect 29082 1428 29112 1558
rect 30874 1428 30904 1558
rect 30970 1428 31000 1558
rect 32762 1428 32792 1558
rect 32858 1428 32888 1558
rect 34650 1428 34680 1558
rect 34746 1428 34776 1558
rect 36538 1428 36568 1558
rect 36634 1428 36664 1558
rect 38426 1428 38456 1558
rect 38522 1428 38552 1558
rect 40314 1428 40344 1558
rect 40410 1428 40440 1558
rect 42202 1428 42232 1558
rect 42298 1428 42328 1558
rect 44090 1428 44120 1558
rect 44186 1428 44216 1558
rect 45972 1428 46002 1558
rect 46068 1428 46098 1558
rect 47860 1428 47890 1558
rect 47956 1428 47986 1558
rect 49748 1428 49778 1558
rect 49844 1428 49874 1558
rect 51636 1428 51666 1558
rect 51732 1428 51762 1558
rect 53524 1428 53554 1558
rect 53620 1428 53650 1558
rect 55412 1428 55442 1558
rect 55508 1428 55538 1558
rect 57300 1428 57330 1558
rect 57396 1428 57426 1558
rect 59188 1428 59218 1558
rect 59284 1428 59314 1558
rect 670 372 700 502
rect 766 372 796 502
rect 2558 372 2588 502
rect 2654 372 2684 502
rect 4446 372 4476 502
rect 4542 372 4572 502
rect 6334 372 6364 502
rect 6430 372 6460 502
rect 8222 372 8252 502
rect 8318 372 8348 502
rect 10110 372 10140 502
rect 10206 372 10236 502
rect 11998 372 12028 502
rect 12094 372 12124 502
rect 13886 372 13916 502
rect 13982 372 14012 502
rect 15768 372 15798 502
rect 15864 372 15894 502
rect 17656 372 17686 502
rect 17752 372 17782 502
rect 19544 372 19574 502
rect 19640 372 19670 502
rect 21432 372 21462 502
rect 21528 372 21558 502
rect 23320 372 23350 502
rect 23416 372 23446 502
rect 25208 372 25238 502
rect 25304 372 25334 502
rect 27096 372 27126 502
rect 27192 372 27222 502
rect 28984 372 29014 502
rect 29080 372 29110 502
rect 30872 372 30902 502
rect 30968 372 30998 502
rect 32760 372 32790 502
rect 32856 372 32886 502
rect 34648 372 34678 502
rect 34744 372 34774 502
rect 36536 372 36566 502
rect 36632 372 36662 502
rect 38424 372 38454 502
rect 38520 372 38550 502
rect 40312 372 40342 502
rect 40408 372 40438 502
rect 42200 372 42230 502
rect 42296 372 42326 502
rect 44088 372 44118 502
rect 44184 372 44214 502
rect 45970 372 46000 502
rect 46066 372 46096 502
rect 47858 372 47888 502
rect 47954 372 47984 502
rect 49746 372 49776 502
rect 49842 372 49872 502
rect 51634 372 51664 502
rect 51730 372 51760 502
rect 53522 372 53552 502
rect 53618 372 53648 502
rect 55410 372 55440 502
rect 55506 372 55536 502
rect 57298 372 57328 502
rect 57394 372 57424 502
rect 59186 372 59216 502
rect 59282 372 59312 502
<< scnmos >>
rect -313 6711 -283 6815
rect -225 6711 -195 6815
rect 80 6683 110 6813
rect 1276 6691 1306 6821
rect 1575 6711 1605 6815
rect 1663 6711 1693 6815
rect 1968 6683 1998 6813
rect 3164 6691 3194 6821
rect 3463 6711 3493 6815
rect 3551 6711 3581 6815
rect 3856 6683 3886 6813
rect 5052 6691 5082 6821
rect 5351 6711 5381 6815
rect 5439 6711 5469 6815
rect 5744 6683 5774 6813
rect 6940 6691 6970 6821
rect 7239 6711 7269 6815
rect 7327 6711 7357 6815
rect 7632 6683 7662 6813
rect 8828 6691 8858 6821
rect 9127 6711 9157 6815
rect 9215 6711 9245 6815
rect 9520 6683 9550 6813
rect 10716 6691 10746 6821
rect 11015 6711 11045 6815
rect 11103 6711 11133 6815
rect 11408 6683 11438 6813
rect 12604 6691 12634 6821
rect 12903 6711 12933 6815
rect 12991 6711 13021 6815
rect 13296 6683 13326 6813
rect 14492 6691 14522 6821
rect 14785 6711 14815 6815
rect 14873 6711 14903 6815
rect 15178 6683 15208 6813
rect 16374 6691 16404 6821
rect 16673 6711 16703 6815
rect 16761 6711 16791 6815
rect 17066 6683 17096 6813
rect 18262 6691 18292 6821
rect 18561 6711 18591 6815
rect 18649 6711 18679 6815
rect 18954 6683 18984 6813
rect 20150 6691 20180 6821
rect 20449 6711 20479 6815
rect 20537 6711 20567 6815
rect 20842 6683 20872 6813
rect 22038 6691 22068 6821
rect 22337 6711 22367 6815
rect 22425 6711 22455 6815
rect 22730 6683 22760 6813
rect 23926 6691 23956 6821
rect 24225 6711 24255 6815
rect 24313 6711 24343 6815
rect 24618 6683 24648 6813
rect 25814 6691 25844 6821
rect 26113 6711 26143 6815
rect 26201 6711 26231 6815
rect 26506 6683 26536 6813
rect 27702 6691 27732 6821
rect 28001 6711 28031 6815
rect 28089 6711 28119 6815
rect 28394 6683 28424 6813
rect 29590 6691 29620 6821
rect 29889 6711 29919 6815
rect 29977 6711 30007 6815
rect 30282 6683 30312 6813
rect 31478 6691 31508 6821
rect 31777 6711 31807 6815
rect 31865 6711 31895 6815
rect 32170 6683 32200 6813
rect 33366 6691 33396 6821
rect 33665 6711 33695 6815
rect 33753 6711 33783 6815
rect 34058 6683 34088 6813
rect 35254 6691 35284 6821
rect 35553 6711 35583 6815
rect 35641 6711 35671 6815
rect 35946 6683 35976 6813
rect 37142 6691 37172 6821
rect 37441 6711 37471 6815
rect 37529 6711 37559 6815
rect 37834 6683 37864 6813
rect 39030 6691 39060 6821
rect 39329 6711 39359 6815
rect 39417 6711 39447 6815
rect 39722 6683 39752 6813
rect 40918 6691 40948 6821
rect 41217 6711 41247 6815
rect 41305 6711 41335 6815
rect 41610 6683 41640 6813
rect 42806 6691 42836 6821
rect 43105 6711 43135 6815
rect 43193 6711 43223 6815
rect 43498 6683 43528 6813
rect 44694 6691 44724 6821
rect 44987 6711 45017 6815
rect 45075 6711 45105 6815
rect 45380 6683 45410 6813
rect 46576 6691 46606 6821
rect 46875 6711 46905 6815
rect 46963 6711 46993 6815
rect 47268 6683 47298 6813
rect 48464 6691 48494 6821
rect 48763 6711 48793 6815
rect 48851 6711 48881 6815
rect 49156 6683 49186 6813
rect 50352 6691 50382 6821
rect 50651 6711 50681 6815
rect 50739 6711 50769 6815
rect 51044 6683 51074 6813
rect 52240 6691 52270 6821
rect 52539 6711 52569 6815
rect 52627 6711 52657 6815
rect 52932 6683 52962 6813
rect 54128 6691 54158 6821
rect 54427 6711 54457 6815
rect 54515 6711 54545 6815
rect 54820 6683 54850 6813
rect 56016 6691 56046 6821
rect 56315 6711 56345 6815
rect 56403 6711 56433 6815
rect 56708 6683 56738 6813
rect 57904 6691 57934 6821
rect 58203 6711 58233 6815
rect 58291 6711 58321 6815
rect 58596 6683 58626 6813
rect 59792 6691 59822 6821
rect 241 5637 271 5767
rect 325 5637 355 5767
rect 1055 5637 1085 5767
rect 1139 5637 1169 5767
rect 2129 5637 2159 5767
rect 2213 5637 2243 5767
rect 2943 5637 2973 5767
rect 3027 5637 3057 5767
rect 4017 5637 4047 5767
rect 4101 5637 4131 5767
rect 4831 5637 4861 5767
rect 4915 5637 4945 5767
rect 5905 5637 5935 5767
rect 5989 5637 6019 5767
rect 6719 5637 6749 5767
rect 6803 5637 6833 5767
rect 7793 5637 7823 5767
rect 7877 5637 7907 5767
rect 8607 5637 8637 5767
rect 8691 5637 8721 5767
rect 9681 5637 9711 5767
rect 9765 5637 9795 5767
rect 10495 5637 10525 5767
rect 10579 5637 10609 5767
rect 11569 5637 11599 5767
rect 11653 5637 11683 5767
rect 12383 5637 12413 5767
rect 12467 5637 12497 5767
rect 13457 5637 13487 5767
rect 13541 5637 13571 5767
rect 14271 5637 14301 5767
rect 14355 5637 14385 5767
rect 15339 5637 15369 5767
rect 15423 5637 15453 5767
rect 16153 5637 16183 5767
rect 16237 5637 16267 5767
rect 17227 5637 17257 5767
rect 17311 5637 17341 5767
rect 18041 5637 18071 5767
rect 18125 5637 18155 5767
rect 19115 5637 19145 5767
rect 19199 5637 19229 5767
rect 19929 5637 19959 5767
rect 20013 5637 20043 5767
rect 21003 5637 21033 5767
rect 21087 5637 21117 5767
rect 21817 5637 21847 5767
rect 21901 5637 21931 5767
rect 22891 5637 22921 5767
rect 22975 5637 23005 5767
rect 23705 5637 23735 5767
rect 23789 5637 23819 5767
rect 24779 5637 24809 5767
rect 24863 5637 24893 5767
rect 25593 5637 25623 5767
rect 25677 5637 25707 5767
rect 26667 5637 26697 5767
rect 26751 5637 26781 5767
rect 27481 5637 27511 5767
rect 27565 5637 27595 5767
rect 28555 5637 28585 5767
rect 28639 5637 28669 5767
rect 29369 5637 29399 5767
rect 29453 5637 29483 5767
rect 30443 5637 30473 5767
rect 30527 5637 30557 5767
rect 31257 5637 31287 5767
rect 31341 5637 31371 5767
rect 32331 5637 32361 5767
rect 32415 5637 32445 5767
rect 33145 5637 33175 5767
rect 33229 5637 33259 5767
rect 34219 5637 34249 5767
rect 34303 5637 34333 5767
rect 35033 5637 35063 5767
rect 35117 5637 35147 5767
rect 36107 5637 36137 5767
rect 36191 5637 36221 5767
rect 36921 5637 36951 5767
rect 37005 5637 37035 5767
rect 37995 5637 38025 5767
rect 38079 5637 38109 5767
rect 38809 5637 38839 5767
rect 38893 5637 38923 5767
rect 39883 5637 39913 5767
rect 39967 5637 39997 5767
rect 40697 5637 40727 5767
rect 40781 5637 40811 5767
rect 41771 5637 41801 5767
rect 41855 5637 41885 5767
rect 42585 5637 42615 5767
rect 42669 5637 42699 5767
rect 43659 5637 43689 5767
rect 43743 5637 43773 5767
rect 44473 5637 44503 5767
rect 44557 5637 44587 5767
rect 45541 5637 45571 5767
rect 45625 5637 45655 5767
rect 46355 5637 46385 5767
rect 46439 5637 46469 5767
rect 47429 5637 47459 5767
rect 47513 5637 47543 5767
rect 48243 5637 48273 5767
rect 48327 5637 48357 5767
rect 49317 5637 49347 5767
rect 49401 5637 49431 5767
rect 50131 5637 50161 5767
rect 50215 5637 50245 5767
rect 51205 5637 51235 5767
rect 51289 5637 51319 5767
rect 52019 5637 52049 5767
rect 52103 5637 52133 5767
rect 53093 5637 53123 5767
rect 53177 5637 53207 5767
rect 53907 5637 53937 5767
rect 53991 5637 54021 5767
rect 54981 5637 55011 5767
rect 55065 5637 55095 5767
rect 55795 5637 55825 5767
rect 55879 5637 55909 5767
rect 56869 5637 56899 5767
rect 56953 5637 56983 5767
rect 57683 5637 57713 5767
rect 57767 5637 57797 5767
rect 58757 5637 58787 5767
rect 58841 5637 58871 5767
rect 59571 5637 59601 5767
rect 59655 5637 59685 5767
rect 5754 4695 5784 4825
rect 5838 4695 5868 4825
rect 5922 4695 5952 4825
rect 6006 4695 6036 4825
rect 6090 4695 6120 4825
rect 6174 4695 6204 4825
rect 6258 4695 6288 4825
rect 6342 4695 6372 4825
rect 6426 4695 6456 4825
rect 6510 4695 6540 4825
rect 6594 4695 6624 4825
rect 6678 4695 6708 4825
rect 6762 4695 6792 4825
rect 6846 4695 6876 4825
rect 6930 4695 6960 4825
rect 7014 4695 7044 4825
rect 7636 4693 7666 4823
rect 7720 4693 7750 4823
rect 7804 4693 7834 4823
rect 7888 4693 7918 4823
rect 7972 4693 8002 4823
rect 8056 4693 8086 4823
rect 8140 4693 8170 4823
rect 8224 4693 8254 4823
rect 8308 4693 8338 4823
rect 8392 4693 8422 4823
rect 8476 4693 8506 4823
rect 8560 4693 8590 4823
rect 8644 4693 8674 4823
rect 8728 4693 8758 4823
rect 8812 4693 8842 4823
rect 8896 4693 8926 4823
rect 20852 4695 20882 4825
rect 20936 4695 20966 4825
rect 21020 4695 21050 4825
rect 21104 4695 21134 4825
rect 21188 4695 21218 4825
rect 21272 4695 21302 4825
rect 21356 4695 21386 4825
rect 21440 4695 21470 4825
rect 21524 4695 21554 4825
rect 21608 4695 21638 4825
rect 21692 4695 21722 4825
rect 21776 4695 21806 4825
rect 21860 4695 21890 4825
rect 21944 4695 21974 4825
rect 22028 4695 22058 4825
rect 22112 4695 22142 4825
rect 22734 4693 22764 4823
rect 22818 4693 22848 4823
rect 22902 4693 22932 4823
rect 22986 4693 23016 4823
rect 23070 4693 23100 4823
rect 23154 4693 23184 4823
rect 23238 4693 23268 4823
rect 23322 4693 23352 4823
rect 23406 4693 23436 4823
rect 23490 4693 23520 4823
rect 23574 4693 23604 4823
rect 23658 4693 23688 4823
rect 23742 4693 23772 4823
rect 23826 4693 23856 4823
rect 23910 4693 23940 4823
rect 23994 4693 24024 4823
rect 35956 4695 35986 4825
rect 36040 4695 36070 4825
rect 36124 4695 36154 4825
rect 36208 4695 36238 4825
rect 36292 4695 36322 4825
rect 36376 4695 36406 4825
rect 36460 4695 36490 4825
rect 36544 4695 36574 4825
rect 36628 4695 36658 4825
rect 36712 4695 36742 4825
rect 36796 4695 36826 4825
rect 36880 4695 36910 4825
rect 36964 4695 36994 4825
rect 37048 4695 37078 4825
rect 37132 4695 37162 4825
rect 37216 4695 37246 4825
rect 37838 4693 37868 4823
rect 37922 4693 37952 4823
rect 38006 4693 38036 4823
rect 38090 4693 38120 4823
rect 38174 4693 38204 4823
rect 38258 4693 38288 4823
rect 38342 4693 38372 4823
rect 38426 4693 38456 4823
rect 38510 4693 38540 4823
rect 38594 4693 38624 4823
rect 38678 4693 38708 4823
rect 38762 4693 38792 4823
rect 38846 4693 38876 4823
rect 38930 4693 38960 4823
rect 39014 4693 39044 4823
rect 39098 4693 39128 4823
rect 51054 4695 51084 4825
rect 51138 4695 51168 4825
rect 51222 4695 51252 4825
rect 51306 4695 51336 4825
rect 51390 4695 51420 4825
rect 51474 4695 51504 4825
rect 51558 4695 51588 4825
rect 51642 4695 51672 4825
rect 51726 4695 51756 4825
rect 51810 4695 51840 4825
rect 51894 4695 51924 4825
rect 51978 4695 52008 4825
rect 52062 4695 52092 4825
rect 52146 4695 52176 4825
rect 52230 4695 52260 4825
rect 52314 4695 52344 4825
rect 52936 4693 52966 4823
rect 53020 4693 53050 4823
rect 53104 4693 53134 4823
rect 53188 4693 53218 4823
rect 53272 4693 53302 4823
rect 53356 4693 53386 4823
rect 53440 4693 53470 4823
rect 53524 4693 53554 4823
rect 53608 4693 53638 4823
rect 53692 4693 53722 4823
rect 53776 4693 53806 4823
rect 53860 4693 53890 4823
rect 53944 4693 53974 4823
rect 54028 4693 54058 4823
rect 54112 4693 54142 4823
rect 54196 4693 54226 4823
rect 30116 3618 30146 3748
rect 30200 3618 30230 3748
rect 30284 3618 30314 3748
rect 30368 3618 30398 3748
rect 30647 3618 30677 3748
rect 30731 3618 30761 3748
rect 30815 3618 30845 3748
rect 30899 3618 30929 3748
rect 30983 3618 31013 3748
rect 31067 3618 31097 3748
rect 31151 3618 31181 3748
rect 31235 3618 31265 3748
rect 31319 3618 31349 3748
rect 31403 3618 31433 3748
rect 31487 3618 31517 3748
rect 31571 3618 31601 3748
rect 31655 3618 31685 3748
rect 31739 3618 31769 3748
rect 31823 3618 31853 3748
rect 31907 3618 31937 3748
rect 43473 3402 43503 3532
rect 43557 3402 43587 3532
rect 43641 3402 43671 3532
rect 43725 3402 43755 3532
rect 43809 3402 43839 3532
rect 43893 3402 43923 3532
rect 43977 3402 44007 3532
rect 44061 3402 44091 3532
rect 44145 3402 44175 3532
rect 44229 3402 44259 3532
rect 44313 3402 44343 3532
rect 44397 3402 44427 3532
rect 44481 3402 44511 3532
rect 44565 3402 44595 3532
rect 44649 3402 44679 3532
rect 44733 3402 44763 3532
rect 45403 3402 45433 3532
rect 45487 3402 45517 3532
rect 45571 3402 45601 3532
rect 45655 3402 45685 3532
rect 45739 3402 45769 3532
rect 45823 3402 45853 3532
rect 45907 3402 45937 3532
rect 45991 3402 46021 3532
rect 46075 3402 46105 3532
rect 46159 3402 46189 3532
rect 46243 3402 46273 3532
rect 46327 3402 46357 3532
rect 46411 3402 46441 3532
rect 46495 3402 46525 3532
rect 46579 3402 46609 3532
rect 46663 3402 46693 3532
rect 13331 3242 13361 3372
rect 13415 3242 13445 3372
rect 13499 3242 13529 3372
rect 13583 3242 13613 3372
rect 13667 3242 13697 3372
rect 13751 3242 13781 3372
rect 13835 3242 13865 3372
rect 13919 3242 13949 3372
rect 14003 3242 14033 3372
rect 14087 3242 14117 3372
rect 14171 3242 14201 3372
rect 14255 3242 14285 3372
rect 14339 3242 14369 3372
rect 14423 3242 14453 3372
rect 14507 3242 14537 3372
rect 14591 3242 14621 3372
rect 15261 3242 15291 3372
rect 15345 3242 15375 3372
rect 15429 3242 15459 3372
rect 15513 3242 15543 3372
rect 15597 3242 15627 3372
rect 15681 3242 15711 3372
rect 15765 3242 15795 3372
rect 15849 3242 15879 3372
rect 15933 3242 15963 3372
rect 16017 3242 16047 3372
rect 16101 3242 16131 3372
rect 16185 3242 16215 3372
rect 16269 3242 16299 3372
rect 16353 3242 16383 3372
rect 16437 3242 16467 3372
rect 16521 3242 16551 3372
rect 5756 2617 5786 2747
rect 5840 2617 5870 2747
rect 5924 2617 5954 2747
rect 6008 2617 6038 2747
rect 6092 2617 6122 2747
rect 6176 2617 6206 2747
rect 6260 2617 6290 2747
rect 6344 2617 6374 2747
rect 6428 2617 6458 2747
rect 6512 2617 6542 2747
rect 6596 2617 6626 2747
rect 6680 2617 6710 2747
rect 6764 2617 6794 2747
rect 6848 2617 6878 2747
rect 6932 2617 6962 2747
rect 7016 2617 7046 2747
rect 7638 2615 7668 2745
rect 7722 2615 7752 2745
rect 7806 2615 7836 2745
rect 7890 2615 7920 2745
rect 7974 2615 8004 2745
rect 8058 2615 8088 2745
rect 8142 2615 8172 2745
rect 8226 2615 8256 2745
rect 8310 2615 8340 2745
rect 8394 2615 8424 2745
rect 8478 2615 8508 2745
rect 8562 2615 8592 2745
rect 8646 2615 8676 2745
rect 8730 2615 8760 2745
rect 8814 2615 8844 2745
rect 8898 2615 8928 2745
rect 20854 2617 20884 2747
rect 20938 2617 20968 2747
rect 21022 2617 21052 2747
rect 21106 2617 21136 2747
rect 21190 2617 21220 2747
rect 21274 2617 21304 2747
rect 21358 2617 21388 2747
rect 21442 2617 21472 2747
rect 21526 2617 21556 2747
rect 21610 2617 21640 2747
rect 21694 2617 21724 2747
rect 21778 2617 21808 2747
rect 21862 2617 21892 2747
rect 21946 2617 21976 2747
rect 22030 2617 22060 2747
rect 22114 2617 22144 2747
rect 22736 2615 22766 2745
rect 22820 2615 22850 2745
rect 22904 2615 22934 2745
rect 22988 2615 23018 2745
rect 23072 2615 23102 2745
rect 23156 2615 23186 2745
rect 23240 2615 23270 2745
rect 23324 2615 23354 2745
rect 23408 2615 23438 2745
rect 23492 2615 23522 2745
rect 23576 2615 23606 2745
rect 23660 2615 23690 2745
rect 23744 2615 23774 2745
rect 23828 2615 23858 2745
rect 23912 2615 23942 2745
rect 23996 2615 24026 2745
rect 35958 2617 35988 2747
rect 36042 2617 36072 2747
rect 36126 2617 36156 2747
rect 36210 2617 36240 2747
rect 36294 2617 36324 2747
rect 36378 2617 36408 2747
rect 36462 2617 36492 2747
rect 36546 2617 36576 2747
rect 36630 2617 36660 2747
rect 36714 2617 36744 2747
rect 36798 2617 36828 2747
rect 36882 2617 36912 2747
rect 36966 2617 36996 2747
rect 37050 2617 37080 2747
rect 37134 2617 37164 2747
rect 37218 2617 37248 2747
rect 37840 2615 37870 2745
rect 37924 2615 37954 2745
rect 38008 2615 38038 2745
rect 38092 2615 38122 2745
rect 38176 2615 38206 2745
rect 38260 2615 38290 2745
rect 38344 2615 38374 2745
rect 38428 2615 38458 2745
rect 38512 2615 38542 2745
rect 38596 2615 38626 2745
rect 38680 2615 38710 2745
rect 38764 2615 38794 2745
rect 38848 2615 38878 2745
rect 38932 2615 38962 2745
rect 39016 2615 39046 2745
rect 39100 2615 39130 2745
rect 51056 2617 51086 2747
rect 51140 2617 51170 2747
rect 51224 2617 51254 2747
rect 51308 2617 51338 2747
rect 51392 2617 51422 2747
rect 51476 2617 51506 2747
rect 51560 2617 51590 2747
rect 51644 2617 51674 2747
rect 51728 2617 51758 2747
rect 51812 2617 51842 2747
rect 51896 2617 51926 2747
rect 51980 2617 52010 2747
rect 52064 2617 52094 2747
rect 52148 2617 52178 2747
rect 52232 2617 52262 2747
rect 52316 2617 52346 2747
rect 52938 2615 52968 2745
rect 53022 2615 53052 2745
rect 53106 2615 53136 2745
rect 53190 2615 53220 2745
rect 53274 2615 53304 2745
rect 53358 2615 53388 2745
rect 53442 2615 53472 2745
rect 53526 2615 53556 2745
rect 53610 2615 53640 2745
rect 53694 2615 53724 2745
rect 53778 2615 53808 2745
rect 53862 2615 53892 2745
rect 53946 2615 53976 2745
rect 54030 2615 54060 2745
rect 54114 2615 54144 2745
rect 54198 2615 54228 2745
rect 297 1673 327 1803
rect 381 1673 411 1803
rect 1111 1673 1141 1803
rect 1195 1673 1225 1803
rect 2185 1673 2215 1803
rect 2269 1673 2299 1803
rect 2999 1673 3029 1803
rect 3083 1673 3113 1803
rect 4073 1673 4103 1803
rect 4157 1673 4187 1803
rect 4887 1673 4917 1803
rect 4971 1673 5001 1803
rect 5961 1673 5991 1803
rect 6045 1673 6075 1803
rect 6775 1673 6805 1803
rect 6859 1673 6889 1803
rect 7849 1673 7879 1803
rect 7933 1673 7963 1803
rect 8663 1673 8693 1803
rect 8747 1673 8777 1803
rect 9737 1673 9767 1803
rect 9821 1673 9851 1803
rect 10551 1673 10581 1803
rect 10635 1673 10665 1803
rect 11625 1673 11655 1803
rect 11709 1673 11739 1803
rect 12439 1673 12469 1803
rect 12523 1673 12553 1803
rect 13513 1673 13543 1803
rect 13597 1673 13627 1803
rect 14327 1673 14357 1803
rect 14411 1673 14441 1803
rect 15395 1673 15425 1803
rect 15479 1673 15509 1803
rect 16209 1673 16239 1803
rect 16293 1673 16323 1803
rect 17283 1673 17313 1803
rect 17367 1673 17397 1803
rect 18097 1673 18127 1803
rect 18181 1673 18211 1803
rect 19171 1673 19201 1803
rect 19255 1673 19285 1803
rect 19985 1673 20015 1803
rect 20069 1673 20099 1803
rect 21059 1673 21089 1803
rect 21143 1673 21173 1803
rect 21873 1673 21903 1803
rect 21957 1673 21987 1803
rect 22947 1673 22977 1803
rect 23031 1673 23061 1803
rect 23761 1673 23791 1803
rect 23845 1673 23875 1803
rect 24835 1673 24865 1803
rect 24919 1673 24949 1803
rect 25649 1673 25679 1803
rect 25733 1673 25763 1803
rect 26723 1673 26753 1803
rect 26807 1673 26837 1803
rect 27537 1673 27567 1803
rect 27621 1673 27651 1803
rect 28611 1673 28641 1803
rect 28695 1673 28725 1803
rect 29425 1673 29455 1803
rect 29509 1673 29539 1803
rect 30499 1673 30529 1803
rect 30583 1673 30613 1803
rect 31313 1673 31343 1803
rect 31397 1673 31427 1803
rect 32387 1673 32417 1803
rect 32471 1673 32501 1803
rect 33201 1673 33231 1803
rect 33285 1673 33315 1803
rect 34275 1673 34305 1803
rect 34359 1673 34389 1803
rect 35089 1673 35119 1803
rect 35173 1673 35203 1803
rect 36163 1673 36193 1803
rect 36247 1673 36277 1803
rect 36977 1673 37007 1803
rect 37061 1673 37091 1803
rect 38051 1673 38081 1803
rect 38135 1673 38165 1803
rect 38865 1673 38895 1803
rect 38949 1673 38979 1803
rect 39939 1673 39969 1803
rect 40023 1673 40053 1803
rect 40753 1673 40783 1803
rect 40837 1673 40867 1803
rect 41827 1673 41857 1803
rect 41911 1673 41941 1803
rect 42641 1673 42671 1803
rect 42725 1673 42755 1803
rect 43715 1673 43745 1803
rect 43799 1673 43829 1803
rect 44529 1673 44559 1803
rect 44613 1673 44643 1803
rect 45597 1673 45627 1803
rect 45681 1673 45711 1803
rect 46411 1673 46441 1803
rect 46495 1673 46525 1803
rect 47485 1673 47515 1803
rect 47569 1673 47599 1803
rect 48299 1673 48329 1803
rect 48383 1673 48413 1803
rect 49373 1673 49403 1803
rect 49457 1673 49487 1803
rect 50187 1673 50217 1803
rect 50271 1673 50301 1803
rect 51261 1673 51291 1803
rect 51345 1673 51375 1803
rect 52075 1673 52105 1803
rect 52159 1673 52189 1803
rect 53149 1673 53179 1803
rect 53233 1673 53263 1803
rect 53963 1673 53993 1803
rect 54047 1673 54077 1803
rect 55037 1673 55067 1803
rect 55121 1673 55151 1803
rect 55851 1673 55881 1803
rect 55935 1673 55965 1803
rect 56925 1673 56955 1803
rect 57009 1673 57039 1803
rect 57739 1673 57769 1803
rect 57823 1673 57853 1803
rect 58813 1673 58843 1803
rect 58897 1673 58927 1803
rect 59627 1673 59657 1803
rect 59711 1673 59741 1803
rect 160 619 190 749
rect 1356 627 1386 757
rect 1661 625 1691 729
rect 1749 625 1779 729
rect 2048 619 2078 749
rect 3244 627 3274 757
rect 3549 625 3579 729
rect 3637 625 3667 729
rect 3936 619 3966 749
rect 5132 627 5162 757
rect 5437 625 5467 729
rect 5525 625 5555 729
rect 5824 619 5854 749
rect 7020 627 7050 757
rect 7325 625 7355 729
rect 7413 625 7443 729
rect 7712 619 7742 749
rect 8908 627 8938 757
rect 9213 625 9243 729
rect 9301 625 9331 729
rect 9600 619 9630 749
rect 10796 627 10826 757
rect 11101 625 11131 729
rect 11189 625 11219 729
rect 11488 619 11518 749
rect 12684 627 12714 757
rect 12989 625 13019 729
rect 13077 625 13107 729
rect 13376 619 13406 749
rect 14572 627 14602 757
rect 14877 625 14907 729
rect 14965 625 14995 729
rect 15258 619 15288 749
rect 16454 627 16484 757
rect 16759 625 16789 729
rect 16847 625 16877 729
rect 17146 619 17176 749
rect 18342 627 18372 757
rect 18647 625 18677 729
rect 18735 625 18765 729
rect 19034 619 19064 749
rect 20230 627 20260 757
rect 20535 625 20565 729
rect 20623 625 20653 729
rect 20922 619 20952 749
rect 22118 627 22148 757
rect 22423 625 22453 729
rect 22511 625 22541 729
rect 22810 619 22840 749
rect 24006 627 24036 757
rect 24311 625 24341 729
rect 24399 625 24429 729
rect 24698 619 24728 749
rect 25894 627 25924 757
rect 26199 625 26229 729
rect 26287 625 26317 729
rect 26586 619 26616 749
rect 27782 627 27812 757
rect 28087 625 28117 729
rect 28175 625 28205 729
rect 28474 619 28504 749
rect 29670 627 29700 757
rect 29975 625 30005 729
rect 30063 625 30093 729
rect 30362 619 30392 749
rect 31558 627 31588 757
rect 31863 625 31893 729
rect 31951 625 31981 729
rect 32250 619 32280 749
rect 33446 627 33476 757
rect 33751 625 33781 729
rect 33839 625 33869 729
rect 34138 619 34168 749
rect 35334 627 35364 757
rect 35639 625 35669 729
rect 35727 625 35757 729
rect 36026 619 36056 749
rect 37222 627 37252 757
rect 37527 625 37557 729
rect 37615 625 37645 729
rect 37914 619 37944 749
rect 39110 627 39140 757
rect 39415 625 39445 729
rect 39503 625 39533 729
rect 39802 619 39832 749
rect 40998 627 41028 757
rect 41303 625 41333 729
rect 41391 625 41421 729
rect 41690 619 41720 749
rect 42886 627 42916 757
rect 43191 625 43221 729
rect 43279 625 43309 729
rect 43578 619 43608 749
rect 44774 627 44804 757
rect 45079 625 45109 729
rect 45167 625 45197 729
rect 45460 619 45490 749
rect 46656 627 46686 757
rect 46961 625 46991 729
rect 47049 625 47079 729
rect 47348 619 47378 749
rect 48544 627 48574 757
rect 48849 625 48879 729
rect 48937 625 48967 729
rect 49236 619 49266 749
rect 50432 627 50462 757
rect 50737 625 50767 729
rect 50825 625 50855 729
rect 51124 619 51154 749
rect 52320 627 52350 757
rect 52625 625 52655 729
rect 52713 625 52743 729
rect 53012 619 53042 749
rect 54208 627 54238 757
rect 54513 625 54543 729
rect 54601 625 54631 729
rect 54900 619 54930 749
rect 56096 627 56126 757
rect 56401 625 56431 729
rect 56489 625 56519 729
rect 56788 619 56818 749
rect 57984 627 58014 757
rect 58289 625 58319 729
rect 58377 625 58407 729
rect 58676 619 58706 749
rect 59872 627 59902 757
rect 60177 625 60207 729
rect 60265 625 60295 729
<< scpmoshvt >>
rect -313 6365 -283 6523
rect -225 6365 -195 6523
rect 80 6363 110 6563
rect 1276 6371 1306 6571
rect 1575 6365 1605 6523
rect 1663 6365 1693 6523
rect 1968 6363 1998 6563
rect 3164 6371 3194 6571
rect 3463 6365 3493 6523
rect 3551 6365 3581 6523
rect 3856 6363 3886 6563
rect 5052 6371 5082 6571
rect 5351 6365 5381 6523
rect 5439 6365 5469 6523
rect 5744 6363 5774 6563
rect 6940 6371 6970 6571
rect 7239 6365 7269 6523
rect 7327 6365 7357 6523
rect 7632 6363 7662 6563
rect 8828 6371 8858 6571
rect 9127 6365 9157 6523
rect 9215 6365 9245 6523
rect 9520 6363 9550 6563
rect 10716 6371 10746 6571
rect 11015 6365 11045 6523
rect 11103 6365 11133 6523
rect 11408 6363 11438 6563
rect 12604 6371 12634 6571
rect 12903 6365 12933 6523
rect 12991 6365 13021 6523
rect 13296 6363 13326 6563
rect 14492 6371 14522 6571
rect 14785 6365 14815 6523
rect 14873 6365 14903 6523
rect 15178 6363 15208 6563
rect 16374 6371 16404 6571
rect 16673 6365 16703 6523
rect 16761 6365 16791 6523
rect 17066 6363 17096 6563
rect 18262 6371 18292 6571
rect 18561 6365 18591 6523
rect 18649 6365 18679 6523
rect 18954 6363 18984 6563
rect 20150 6371 20180 6571
rect 20449 6365 20479 6523
rect 20537 6365 20567 6523
rect 20842 6363 20872 6563
rect 22038 6371 22068 6571
rect 22337 6365 22367 6523
rect 22425 6365 22455 6523
rect 22730 6363 22760 6563
rect 23926 6371 23956 6571
rect 24225 6365 24255 6523
rect 24313 6365 24343 6523
rect 24618 6363 24648 6563
rect 25814 6371 25844 6571
rect 26113 6365 26143 6523
rect 26201 6365 26231 6523
rect 26506 6363 26536 6563
rect 27702 6371 27732 6571
rect 28001 6365 28031 6523
rect 28089 6365 28119 6523
rect 28394 6363 28424 6563
rect 29590 6371 29620 6571
rect 29889 6365 29919 6523
rect 29977 6365 30007 6523
rect 30282 6363 30312 6563
rect 31478 6371 31508 6571
rect 31777 6365 31807 6523
rect 31865 6365 31895 6523
rect 32170 6363 32200 6563
rect 33366 6371 33396 6571
rect 33665 6365 33695 6523
rect 33753 6365 33783 6523
rect 34058 6363 34088 6563
rect 35254 6371 35284 6571
rect 35553 6365 35583 6523
rect 35641 6365 35671 6523
rect 35946 6363 35976 6563
rect 37142 6371 37172 6571
rect 37441 6365 37471 6523
rect 37529 6365 37559 6523
rect 37834 6363 37864 6563
rect 39030 6371 39060 6571
rect 39329 6365 39359 6523
rect 39417 6365 39447 6523
rect 39722 6363 39752 6563
rect 40918 6371 40948 6571
rect 41217 6365 41247 6523
rect 41305 6365 41335 6523
rect 41610 6363 41640 6563
rect 42806 6371 42836 6571
rect 43105 6365 43135 6523
rect 43193 6365 43223 6523
rect 43498 6363 43528 6563
rect 44694 6371 44724 6571
rect 44987 6365 45017 6523
rect 45075 6365 45105 6523
rect 45380 6363 45410 6563
rect 46576 6371 46606 6571
rect 46875 6365 46905 6523
rect 46963 6365 46993 6523
rect 47268 6363 47298 6563
rect 48464 6371 48494 6571
rect 48763 6365 48793 6523
rect 48851 6365 48881 6523
rect 49156 6363 49186 6563
rect 50352 6371 50382 6571
rect 50651 6365 50681 6523
rect 50739 6365 50769 6523
rect 51044 6363 51074 6563
rect 52240 6371 52270 6571
rect 52539 6365 52569 6523
rect 52627 6365 52657 6523
rect 52932 6363 52962 6563
rect 54128 6371 54158 6571
rect 54427 6365 54457 6523
rect 54515 6365 54545 6523
rect 54820 6363 54850 6563
rect 56016 6371 56046 6571
rect 56315 6365 56345 6523
rect 56403 6365 56433 6523
rect 56708 6363 56738 6563
rect 57904 6371 57934 6571
rect 58203 6365 58233 6523
rect 58291 6365 58321 6523
rect 58596 6363 58626 6563
rect 59792 6371 59822 6571
rect 253 5317 283 5517
rect 325 5317 355 5517
rect 1067 5317 1097 5517
rect 1139 5317 1169 5517
rect 2141 5317 2171 5517
rect 2213 5317 2243 5517
rect 2955 5317 2985 5517
rect 3027 5317 3057 5517
rect 4029 5317 4059 5517
rect 4101 5317 4131 5517
rect 4843 5317 4873 5517
rect 4915 5317 4945 5517
rect 5917 5317 5947 5517
rect 5989 5317 6019 5517
rect 6731 5317 6761 5517
rect 6803 5317 6833 5517
rect 7805 5317 7835 5517
rect 7877 5317 7907 5517
rect 8619 5317 8649 5517
rect 8691 5317 8721 5517
rect 9693 5317 9723 5517
rect 9765 5317 9795 5517
rect 10507 5317 10537 5517
rect 10579 5317 10609 5517
rect 11581 5317 11611 5517
rect 11653 5317 11683 5517
rect 12395 5317 12425 5517
rect 12467 5317 12497 5517
rect 13469 5317 13499 5517
rect 13541 5317 13571 5517
rect 14283 5317 14313 5517
rect 14355 5317 14385 5517
rect 15351 5317 15381 5517
rect 15423 5317 15453 5517
rect 16165 5317 16195 5517
rect 16237 5317 16267 5517
rect 17239 5317 17269 5517
rect 17311 5317 17341 5517
rect 18053 5317 18083 5517
rect 18125 5317 18155 5517
rect 19127 5317 19157 5517
rect 19199 5317 19229 5517
rect 19941 5317 19971 5517
rect 20013 5317 20043 5517
rect 21015 5317 21045 5517
rect 21087 5317 21117 5517
rect 21829 5317 21859 5517
rect 21901 5317 21931 5517
rect 22903 5317 22933 5517
rect 22975 5317 23005 5517
rect 23717 5317 23747 5517
rect 23789 5317 23819 5517
rect 24791 5317 24821 5517
rect 24863 5317 24893 5517
rect 25605 5317 25635 5517
rect 25677 5317 25707 5517
rect 26679 5317 26709 5517
rect 26751 5317 26781 5517
rect 27493 5317 27523 5517
rect 27565 5317 27595 5517
rect 28567 5317 28597 5517
rect 28639 5317 28669 5517
rect 29381 5317 29411 5517
rect 29453 5317 29483 5517
rect 30455 5317 30485 5517
rect 30527 5317 30557 5517
rect 31269 5317 31299 5517
rect 31341 5317 31371 5517
rect 32343 5317 32373 5517
rect 32415 5317 32445 5517
rect 33157 5317 33187 5517
rect 33229 5317 33259 5517
rect 34231 5317 34261 5517
rect 34303 5317 34333 5517
rect 35045 5317 35075 5517
rect 35117 5317 35147 5517
rect 36119 5317 36149 5517
rect 36191 5317 36221 5517
rect 36933 5317 36963 5517
rect 37005 5317 37035 5517
rect 38007 5317 38037 5517
rect 38079 5317 38109 5517
rect 38821 5317 38851 5517
rect 38893 5317 38923 5517
rect 39895 5317 39925 5517
rect 39967 5317 39997 5517
rect 40709 5317 40739 5517
rect 40781 5317 40811 5517
rect 41783 5317 41813 5517
rect 41855 5317 41885 5517
rect 42597 5317 42627 5517
rect 42669 5317 42699 5517
rect 43671 5317 43701 5517
rect 43743 5317 43773 5517
rect 44485 5317 44515 5517
rect 44557 5317 44587 5517
rect 45553 5317 45583 5517
rect 45625 5317 45655 5517
rect 46367 5317 46397 5517
rect 46439 5317 46469 5517
rect 47441 5317 47471 5517
rect 47513 5317 47543 5517
rect 48255 5317 48285 5517
rect 48327 5317 48357 5517
rect 49329 5317 49359 5517
rect 49401 5317 49431 5517
rect 50143 5317 50173 5517
rect 50215 5317 50245 5517
rect 51217 5317 51247 5517
rect 51289 5317 51319 5517
rect 52031 5317 52061 5517
rect 52103 5317 52133 5517
rect 53105 5317 53135 5517
rect 53177 5317 53207 5517
rect 53919 5317 53949 5517
rect 53991 5317 54021 5517
rect 54993 5317 55023 5517
rect 55065 5317 55095 5517
rect 55807 5317 55837 5517
rect 55879 5317 55909 5517
rect 56881 5317 56911 5517
rect 56953 5317 56983 5517
rect 57695 5317 57725 5517
rect 57767 5317 57797 5517
rect 58769 5317 58799 5517
rect 58841 5317 58871 5517
rect 59583 5317 59613 5517
rect 59655 5317 59685 5517
rect 5754 4945 5784 5145
rect 5838 4945 5868 5145
rect 5922 4945 5952 5145
rect 6006 4945 6036 5145
rect 6090 4945 6120 5145
rect 6174 4945 6204 5145
rect 6258 4945 6288 5145
rect 6342 4945 6372 5145
rect 6426 4945 6456 5145
rect 6510 4945 6540 5145
rect 6594 4945 6624 5145
rect 6678 4945 6708 5145
rect 6762 4945 6792 5145
rect 6846 4945 6876 5145
rect 6930 4945 6960 5145
rect 7014 4945 7044 5145
rect 7636 4943 7666 5143
rect 7720 4943 7750 5143
rect 7804 4943 7834 5143
rect 7888 4943 7918 5143
rect 7972 4943 8002 5143
rect 8056 4943 8086 5143
rect 8140 4943 8170 5143
rect 8224 4943 8254 5143
rect 8308 4943 8338 5143
rect 8392 4943 8422 5143
rect 8476 4943 8506 5143
rect 8560 4943 8590 5143
rect 8644 4943 8674 5143
rect 8728 4943 8758 5143
rect 8812 4943 8842 5143
rect 8896 4943 8926 5143
rect 20852 4945 20882 5145
rect 20936 4945 20966 5145
rect 21020 4945 21050 5145
rect 21104 4945 21134 5145
rect 21188 4945 21218 5145
rect 21272 4945 21302 5145
rect 21356 4945 21386 5145
rect 21440 4945 21470 5145
rect 21524 4945 21554 5145
rect 21608 4945 21638 5145
rect 21692 4945 21722 5145
rect 21776 4945 21806 5145
rect 21860 4945 21890 5145
rect 21944 4945 21974 5145
rect 22028 4945 22058 5145
rect 22112 4945 22142 5145
rect 22734 4943 22764 5143
rect 22818 4943 22848 5143
rect 22902 4943 22932 5143
rect 22986 4943 23016 5143
rect 23070 4943 23100 5143
rect 23154 4943 23184 5143
rect 23238 4943 23268 5143
rect 23322 4943 23352 5143
rect 23406 4943 23436 5143
rect 23490 4943 23520 5143
rect 23574 4943 23604 5143
rect 23658 4943 23688 5143
rect 23742 4943 23772 5143
rect 23826 4943 23856 5143
rect 23910 4943 23940 5143
rect 23994 4943 24024 5143
rect 35956 4945 35986 5145
rect 36040 4945 36070 5145
rect 36124 4945 36154 5145
rect 36208 4945 36238 5145
rect 36292 4945 36322 5145
rect 36376 4945 36406 5145
rect 36460 4945 36490 5145
rect 36544 4945 36574 5145
rect 36628 4945 36658 5145
rect 36712 4945 36742 5145
rect 36796 4945 36826 5145
rect 36880 4945 36910 5145
rect 36964 4945 36994 5145
rect 37048 4945 37078 5145
rect 37132 4945 37162 5145
rect 37216 4945 37246 5145
rect 37838 4943 37868 5143
rect 37922 4943 37952 5143
rect 38006 4943 38036 5143
rect 38090 4943 38120 5143
rect 38174 4943 38204 5143
rect 38258 4943 38288 5143
rect 38342 4943 38372 5143
rect 38426 4943 38456 5143
rect 38510 4943 38540 5143
rect 38594 4943 38624 5143
rect 38678 4943 38708 5143
rect 38762 4943 38792 5143
rect 38846 4943 38876 5143
rect 38930 4943 38960 5143
rect 39014 4943 39044 5143
rect 39098 4943 39128 5143
rect 51054 4945 51084 5145
rect 51138 4945 51168 5145
rect 51222 4945 51252 5145
rect 51306 4945 51336 5145
rect 51390 4945 51420 5145
rect 51474 4945 51504 5145
rect 51558 4945 51588 5145
rect 51642 4945 51672 5145
rect 51726 4945 51756 5145
rect 51810 4945 51840 5145
rect 51894 4945 51924 5145
rect 51978 4945 52008 5145
rect 52062 4945 52092 5145
rect 52146 4945 52176 5145
rect 52230 4945 52260 5145
rect 52314 4945 52344 5145
rect 52936 4943 52966 5143
rect 53020 4943 53050 5143
rect 53104 4943 53134 5143
rect 53188 4943 53218 5143
rect 53272 4943 53302 5143
rect 53356 4943 53386 5143
rect 53440 4943 53470 5143
rect 53524 4943 53554 5143
rect 53608 4943 53638 5143
rect 53692 4943 53722 5143
rect 53776 4943 53806 5143
rect 53860 4943 53890 5143
rect 53944 4943 53974 5143
rect 54028 4943 54058 5143
rect 54112 4943 54142 5143
rect 54196 4943 54226 5143
rect 30116 3868 30146 4068
rect 30200 3868 30230 4068
rect 30284 3868 30314 4068
rect 30368 3868 30398 4068
rect 30647 3868 30677 4068
rect 30731 3868 30761 4068
rect 30815 3868 30845 4068
rect 30899 3868 30929 4068
rect 30983 3868 31013 4068
rect 31067 3868 31097 4068
rect 31151 3868 31181 4068
rect 31235 3868 31265 4068
rect 31319 3868 31349 4068
rect 31403 3868 31433 4068
rect 31487 3868 31517 4068
rect 31571 3868 31601 4068
rect 31655 3868 31685 4068
rect 31739 3868 31769 4068
rect 31823 3868 31853 4068
rect 31907 3868 31937 4068
rect 13331 3492 13361 3692
rect 13415 3492 13445 3692
rect 13499 3492 13529 3692
rect 13583 3492 13613 3692
rect 13667 3492 13697 3692
rect 13751 3492 13781 3692
rect 13835 3492 13865 3692
rect 13919 3492 13949 3692
rect 14003 3492 14033 3692
rect 14087 3492 14117 3692
rect 14171 3492 14201 3692
rect 14255 3492 14285 3692
rect 14339 3492 14369 3692
rect 14423 3492 14453 3692
rect 14507 3492 14537 3692
rect 14591 3492 14621 3692
rect 15261 3492 15291 3692
rect 15345 3492 15375 3692
rect 15429 3492 15459 3692
rect 15513 3492 15543 3692
rect 15597 3492 15627 3692
rect 15681 3492 15711 3692
rect 15765 3492 15795 3692
rect 15849 3492 15879 3692
rect 15933 3492 15963 3692
rect 16017 3492 16047 3692
rect 16101 3492 16131 3692
rect 16185 3492 16215 3692
rect 16269 3492 16299 3692
rect 16353 3492 16383 3692
rect 16437 3492 16467 3692
rect 16521 3492 16551 3692
rect 43473 3652 43503 3852
rect 43557 3652 43587 3852
rect 43641 3652 43671 3852
rect 43725 3652 43755 3852
rect 43809 3652 43839 3852
rect 43893 3652 43923 3852
rect 43977 3652 44007 3852
rect 44061 3652 44091 3852
rect 44145 3652 44175 3852
rect 44229 3652 44259 3852
rect 44313 3652 44343 3852
rect 44397 3652 44427 3852
rect 44481 3652 44511 3852
rect 44565 3652 44595 3852
rect 44649 3652 44679 3852
rect 44733 3652 44763 3852
rect 45403 3652 45433 3852
rect 45487 3652 45517 3852
rect 45571 3652 45601 3852
rect 45655 3652 45685 3852
rect 45739 3652 45769 3852
rect 45823 3652 45853 3852
rect 45907 3652 45937 3852
rect 45991 3652 46021 3852
rect 46075 3652 46105 3852
rect 46159 3652 46189 3852
rect 46243 3652 46273 3852
rect 46327 3652 46357 3852
rect 46411 3652 46441 3852
rect 46495 3652 46525 3852
rect 46579 3652 46609 3852
rect 46663 3652 46693 3852
rect 5756 2297 5786 2497
rect 5840 2297 5870 2497
rect 5924 2297 5954 2497
rect 6008 2297 6038 2497
rect 6092 2297 6122 2497
rect 6176 2297 6206 2497
rect 6260 2297 6290 2497
rect 6344 2297 6374 2497
rect 6428 2297 6458 2497
rect 6512 2297 6542 2497
rect 6596 2297 6626 2497
rect 6680 2297 6710 2497
rect 6764 2297 6794 2497
rect 6848 2297 6878 2497
rect 6932 2297 6962 2497
rect 7016 2297 7046 2497
rect 7638 2295 7668 2495
rect 7722 2295 7752 2495
rect 7806 2295 7836 2495
rect 7890 2295 7920 2495
rect 7974 2295 8004 2495
rect 8058 2295 8088 2495
rect 8142 2295 8172 2495
rect 8226 2295 8256 2495
rect 8310 2295 8340 2495
rect 8394 2295 8424 2495
rect 8478 2295 8508 2495
rect 8562 2295 8592 2495
rect 8646 2295 8676 2495
rect 8730 2295 8760 2495
rect 8814 2295 8844 2495
rect 8898 2295 8928 2495
rect 20854 2297 20884 2497
rect 20938 2297 20968 2497
rect 21022 2297 21052 2497
rect 21106 2297 21136 2497
rect 21190 2297 21220 2497
rect 21274 2297 21304 2497
rect 21358 2297 21388 2497
rect 21442 2297 21472 2497
rect 21526 2297 21556 2497
rect 21610 2297 21640 2497
rect 21694 2297 21724 2497
rect 21778 2297 21808 2497
rect 21862 2297 21892 2497
rect 21946 2297 21976 2497
rect 22030 2297 22060 2497
rect 22114 2297 22144 2497
rect 22736 2295 22766 2495
rect 22820 2295 22850 2495
rect 22904 2295 22934 2495
rect 22988 2295 23018 2495
rect 23072 2295 23102 2495
rect 23156 2295 23186 2495
rect 23240 2295 23270 2495
rect 23324 2295 23354 2495
rect 23408 2295 23438 2495
rect 23492 2295 23522 2495
rect 23576 2295 23606 2495
rect 23660 2295 23690 2495
rect 23744 2295 23774 2495
rect 23828 2295 23858 2495
rect 23912 2295 23942 2495
rect 23996 2295 24026 2495
rect 35958 2297 35988 2497
rect 36042 2297 36072 2497
rect 36126 2297 36156 2497
rect 36210 2297 36240 2497
rect 36294 2297 36324 2497
rect 36378 2297 36408 2497
rect 36462 2297 36492 2497
rect 36546 2297 36576 2497
rect 36630 2297 36660 2497
rect 36714 2297 36744 2497
rect 36798 2297 36828 2497
rect 36882 2297 36912 2497
rect 36966 2297 36996 2497
rect 37050 2297 37080 2497
rect 37134 2297 37164 2497
rect 37218 2297 37248 2497
rect 37840 2295 37870 2495
rect 37924 2295 37954 2495
rect 38008 2295 38038 2495
rect 38092 2295 38122 2495
rect 38176 2295 38206 2495
rect 38260 2295 38290 2495
rect 38344 2295 38374 2495
rect 38428 2295 38458 2495
rect 38512 2295 38542 2495
rect 38596 2295 38626 2495
rect 38680 2295 38710 2495
rect 38764 2295 38794 2495
rect 38848 2295 38878 2495
rect 38932 2295 38962 2495
rect 39016 2295 39046 2495
rect 39100 2295 39130 2495
rect 51056 2297 51086 2497
rect 51140 2297 51170 2497
rect 51224 2297 51254 2497
rect 51308 2297 51338 2497
rect 51392 2297 51422 2497
rect 51476 2297 51506 2497
rect 51560 2297 51590 2497
rect 51644 2297 51674 2497
rect 51728 2297 51758 2497
rect 51812 2297 51842 2497
rect 51896 2297 51926 2497
rect 51980 2297 52010 2497
rect 52064 2297 52094 2497
rect 52148 2297 52178 2497
rect 52232 2297 52262 2497
rect 52316 2297 52346 2497
rect 52938 2295 52968 2495
rect 53022 2295 53052 2495
rect 53106 2295 53136 2495
rect 53190 2295 53220 2495
rect 53274 2295 53304 2495
rect 53358 2295 53388 2495
rect 53442 2295 53472 2495
rect 53526 2295 53556 2495
rect 53610 2295 53640 2495
rect 53694 2295 53724 2495
rect 53778 2295 53808 2495
rect 53862 2295 53892 2495
rect 53946 2295 53976 2495
rect 54030 2295 54060 2495
rect 54114 2295 54144 2495
rect 54198 2295 54228 2495
rect 297 1923 327 2123
rect 369 1923 399 2123
rect 1111 1923 1141 2123
rect 1183 1923 1213 2123
rect 2185 1923 2215 2123
rect 2257 1923 2287 2123
rect 2999 1923 3029 2123
rect 3071 1923 3101 2123
rect 4073 1923 4103 2123
rect 4145 1923 4175 2123
rect 4887 1923 4917 2123
rect 4959 1923 4989 2123
rect 5961 1923 5991 2123
rect 6033 1923 6063 2123
rect 6775 1923 6805 2123
rect 6847 1923 6877 2123
rect 7849 1923 7879 2123
rect 7921 1923 7951 2123
rect 8663 1923 8693 2123
rect 8735 1923 8765 2123
rect 9737 1923 9767 2123
rect 9809 1923 9839 2123
rect 10551 1923 10581 2123
rect 10623 1923 10653 2123
rect 11625 1923 11655 2123
rect 11697 1923 11727 2123
rect 12439 1923 12469 2123
rect 12511 1923 12541 2123
rect 13513 1923 13543 2123
rect 13585 1923 13615 2123
rect 14327 1923 14357 2123
rect 14399 1923 14429 2123
rect 15395 1923 15425 2123
rect 15467 1923 15497 2123
rect 16209 1923 16239 2123
rect 16281 1923 16311 2123
rect 17283 1923 17313 2123
rect 17355 1923 17385 2123
rect 18097 1923 18127 2123
rect 18169 1923 18199 2123
rect 19171 1923 19201 2123
rect 19243 1923 19273 2123
rect 19985 1923 20015 2123
rect 20057 1923 20087 2123
rect 21059 1923 21089 2123
rect 21131 1923 21161 2123
rect 21873 1923 21903 2123
rect 21945 1923 21975 2123
rect 22947 1923 22977 2123
rect 23019 1923 23049 2123
rect 23761 1923 23791 2123
rect 23833 1923 23863 2123
rect 24835 1923 24865 2123
rect 24907 1923 24937 2123
rect 25649 1923 25679 2123
rect 25721 1923 25751 2123
rect 26723 1923 26753 2123
rect 26795 1923 26825 2123
rect 27537 1923 27567 2123
rect 27609 1923 27639 2123
rect 28611 1923 28641 2123
rect 28683 1923 28713 2123
rect 29425 1923 29455 2123
rect 29497 1923 29527 2123
rect 30499 1923 30529 2123
rect 30571 1923 30601 2123
rect 31313 1923 31343 2123
rect 31385 1923 31415 2123
rect 32387 1923 32417 2123
rect 32459 1923 32489 2123
rect 33201 1923 33231 2123
rect 33273 1923 33303 2123
rect 34275 1923 34305 2123
rect 34347 1923 34377 2123
rect 35089 1923 35119 2123
rect 35161 1923 35191 2123
rect 36163 1923 36193 2123
rect 36235 1923 36265 2123
rect 36977 1923 37007 2123
rect 37049 1923 37079 2123
rect 38051 1923 38081 2123
rect 38123 1923 38153 2123
rect 38865 1923 38895 2123
rect 38937 1923 38967 2123
rect 39939 1923 39969 2123
rect 40011 1923 40041 2123
rect 40753 1923 40783 2123
rect 40825 1923 40855 2123
rect 41827 1923 41857 2123
rect 41899 1923 41929 2123
rect 42641 1923 42671 2123
rect 42713 1923 42743 2123
rect 43715 1923 43745 2123
rect 43787 1923 43817 2123
rect 44529 1923 44559 2123
rect 44601 1923 44631 2123
rect 45597 1923 45627 2123
rect 45669 1923 45699 2123
rect 46411 1923 46441 2123
rect 46483 1923 46513 2123
rect 47485 1923 47515 2123
rect 47557 1923 47587 2123
rect 48299 1923 48329 2123
rect 48371 1923 48401 2123
rect 49373 1923 49403 2123
rect 49445 1923 49475 2123
rect 50187 1923 50217 2123
rect 50259 1923 50289 2123
rect 51261 1923 51291 2123
rect 51333 1923 51363 2123
rect 52075 1923 52105 2123
rect 52147 1923 52177 2123
rect 53149 1923 53179 2123
rect 53221 1923 53251 2123
rect 53963 1923 53993 2123
rect 54035 1923 54065 2123
rect 55037 1923 55067 2123
rect 55109 1923 55139 2123
rect 55851 1923 55881 2123
rect 55923 1923 55953 2123
rect 56925 1923 56955 2123
rect 56997 1923 57027 2123
rect 57739 1923 57769 2123
rect 57811 1923 57841 2123
rect 58813 1923 58843 2123
rect 58885 1923 58915 2123
rect 59627 1923 59657 2123
rect 59699 1923 59729 2123
rect 160 869 190 1069
rect 1356 877 1386 1077
rect 1661 917 1691 1075
rect 1749 917 1779 1075
rect 2048 869 2078 1069
rect 3244 877 3274 1077
rect 3549 917 3579 1075
rect 3637 917 3667 1075
rect 3936 869 3966 1069
rect 5132 877 5162 1077
rect 5437 917 5467 1075
rect 5525 917 5555 1075
rect 5824 869 5854 1069
rect 7020 877 7050 1077
rect 7325 917 7355 1075
rect 7413 917 7443 1075
rect 7712 869 7742 1069
rect 8908 877 8938 1077
rect 9213 917 9243 1075
rect 9301 917 9331 1075
rect 9600 869 9630 1069
rect 10796 877 10826 1077
rect 11101 917 11131 1075
rect 11189 917 11219 1075
rect 11488 869 11518 1069
rect 12684 877 12714 1077
rect 12989 917 13019 1075
rect 13077 917 13107 1075
rect 13376 869 13406 1069
rect 14572 877 14602 1077
rect 14877 917 14907 1075
rect 14965 917 14995 1075
rect 15258 869 15288 1069
rect 16454 877 16484 1077
rect 16759 917 16789 1075
rect 16847 917 16877 1075
rect 17146 869 17176 1069
rect 18342 877 18372 1077
rect 18647 917 18677 1075
rect 18735 917 18765 1075
rect 19034 869 19064 1069
rect 20230 877 20260 1077
rect 20535 917 20565 1075
rect 20623 917 20653 1075
rect 20922 869 20952 1069
rect 22118 877 22148 1077
rect 22423 917 22453 1075
rect 22511 917 22541 1075
rect 22810 869 22840 1069
rect 24006 877 24036 1077
rect 24311 917 24341 1075
rect 24399 917 24429 1075
rect 24698 869 24728 1069
rect 25894 877 25924 1077
rect 26199 917 26229 1075
rect 26287 917 26317 1075
rect 26586 869 26616 1069
rect 27782 877 27812 1077
rect 28087 917 28117 1075
rect 28175 917 28205 1075
rect 28474 869 28504 1069
rect 29670 877 29700 1077
rect 29975 917 30005 1075
rect 30063 917 30093 1075
rect 30362 869 30392 1069
rect 31558 877 31588 1077
rect 31863 917 31893 1075
rect 31951 917 31981 1075
rect 32250 869 32280 1069
rect 33446 877 33476 1077
rect 33751 917 33781 1075
rect 33839 917 33869 1075
rect 34138 869 34168 1069
rect 35334 877 35364 1077
rect 35639 917 35669 1075
rect 35727 917 35757 1075
rect 36026 869 36056 1069
rect 37222 877 37252 1077
rect 37527 917 37557 1075
rect 37615 917 37645 1075
rect 37914 869 37944 1069
rect 39110 877 39140 1077
rect 39415 917 39445 1075
rect 39503 917 39533 1075
rect 39802 869 39832 1069
rect 40998 877 41028 1077
rect 41303 917 41333 1075
rect 41391 917 41421 1075
rect 41690 869 41720 1069
rect 42886 877 42916 1077
rect 43191 917 43221 1075
rect 43279 917 43309 1075
rect 43578 869 43608 1069
rect 44774 877 44804 1077
rect 45079 917 45109 1075
rect 45167 917 45197 1075
rect 45460 869 45490 1069
rect 46656 877 46686 1077
rect 46961 917 46991 1075
rect 47049 917 47079 1075
rect 47348 869 47378 1069
rect 48544 877 48574 1077
rect 48849 917 48879 1075
rect 48937 917 48967 1075
rect 49236 869 49266 1069
rect 50432 877 50462 1077
rect 50737 917 50767 1075
rect 50825 917 50855 1075
rect 51124 869 51154 1069
rect 52320 877 52350 1077
rect 52625 917 52655 1075
rect 52713 917 52743 1075
rect 53012 869 53042 1069
rect 54208 877 54238 1077
rect 54513 917 54543 1075
rect 54601 917 54631 1075
rect 54900 869 54930 1069
rect 56096 877 56126 1077
rect 56401 917 56431 1075
rect 56489 917 56519 1075
rect 56788 869 56818 1069
rect 57984 877 58014 1077
rect 58289 917 58319 1075
rect 58377 917 58407 1075
rect 58676 869 58706 1069
rect 59872 877 59902 1077
rect 60177 917 60207 1075
rect 60265 917 60295 1075
<< pmoshvt >>
rect 356 6378 386 6578
rect 686 6538 716 6738
rect 782 6538 812 6738
rect 1002 6378 1032 6578
rect 2244 6378 2274 6578
rect 2574 6538 2604 6738
rect 2670 6538 2700 6738
rect 2890 6378 2920 6578
rect 4132 6378 4162 6578
rect 4462 6538 4492 6738
rect 4558 6538 4588 6738
rect 4778 6378 4808 6578
rect 6020 6378 6050 6578
rect 6350 6538 6380 6738
rect 6446 6538 6476 6738
rect 6666 6378 6696 6578
rect 7908 6378 7938 6578
rect 8238 6538 8268 6738
rect 8334 6538 8364 6738
rect 8554 6378 8584 6578
rect 9796 6378 9826 6578
rect 10126 6538 10156 6738
rect 10222 6538 10252 6738
rect 10442 6378 10472 6578
rect 11684 6378 11714 6578
rect 12014 6538 12044 6738
rect 12110 6538 12140 6738
rect 12330 6378 12360 6578
rect 13572 6378 13602 6578
rect 13902 6538 13932 6738
rect 13998 6538 14028 6738
rect 14218 6378 14248 6578
rect 15454 6378 15484 6578
rect 15784 6538 15814 6738
rect 15880 6538 15910 6738
rect 16100 6378 16130 6578
rect 17342 6378 17372 6578
rect 17672 6538 17702 6738
rect 17768 6538 17798 6738
rect 17988 6378 18018 6578
rect 19230 6378 19260 6578
rect 19560 6538 19590 6738
rect 19656 6538 19686 6738
rect 19876 6378 19906 6578
rect 21118 6378 21148 6578
rect 21448 6538 21478 6738
rect 21544 6538 21574 6738
rect 21764 6378 21794 6578
rect 23006 6378 23036 6578
rect 23336 6538 23366 6738
rect 23432 6538 23462 6738
rect 23652 6378 23682 6578
rect 24894 6378 24924 6578
rect 25224 6538 25254 6738
rect 25320 6538 25350 6738
rect 25540 6378 25570 6578
rect 26782 6378 26812 6578
rect 27112 6538 27142 6738
rect 27208 6538 27238 6738
rect 27428 6378 27458 6578
rect 28670 6378 28700 6578
rect 29000 6538 29030 6738
rect 29096 6538 29126 6738
rect 29316 6378 29346 6578
rect 30558 6378 30588 6578
rect 30888 6538 30918 6738
rect 30984 6538 31014 6738
rect 31204 6378 31234 6578
rect 32446 6378 32476 6578
rect 32776 6538 32806 6738
rect 32872 6538 32902 6738
rect 33092 6378 33122 6578
rect 34334 6378 34364 6578
rect 34664 6538 34694 6738
rect 34760 6538 34790 6738
rect 34980 6378 35010 6578
rect 36222 6378 36252 6578
rect 36552 6538 36582 6738
rect 36648 6538 36678 6738
rect 36868 6378 36898 6578
rect 38110 6378 38140 6578
rect 38440 6538 38470 6738
rect 38536 6538 38566 6738
rect 38756 6378 38786 6578
rect 39998 6378 40028 6578
rect 40328 6538 40358 6738
rect 40424 6538 40454 6738
rect 40644 6378 40674 6578
rect 41886 6378 41916 6578
rect 42216 6538 42246 6738
rect 42312 6538 42342 6738
rect 42532 6378 42562 6578
rect 43774 6378 43804 6578
rect 44104 6538 44134 6738
rect 44200 6538 44230 6738
rect 44420 6378 44450 6578
rect 45656 6378 45686 6578
rect 45986 6538 46016 6738
rect 46082 6538 46112 6738
rect 46302 6378 46332 6578
rect 47544 6378 47574 6578
rect 47874 6538 47904 6738
rect 47970 6538 48000 6738
rect 48190 6378 48220 6578
rect 49432 6378 49462 6578
rect 49762 6538 49792 6738
rect 49858 6538 49888 6738
rect 50078 6378 50108 6578
rect 51320 6378 51350 6578
rect 51650 6538 51680 6738
rect 51746 6538 51776 6738
rect 51966 6378 51996 6578
rect 53208 6378 53238 6578
rect 53538 6538 53568 6738
rect 53634 6538 53664 6738
rect 53854 6378 53884 6578
rect 55096 6378 55126 6578
rect 55426 6538 55456 6738
rect 55522 6538 55552 6738
rect 55742 6378 55772 6578
rect 56984 6378 57014 6578
rect 57314 6538 57344 6738
rect 57410 6538 57440 6738
rect 57630 6378 57660 6578
rect 58872 6378 58902 6578
rect 59202 6538 59232 6738
rect 59298 6538 59328 6738
rect 59518 6378 59548 6578
rect 684 5482 714 5682
rect 780 5482 810 5682
rect 2572 5482 2602 5682
rect 2668 5482 2698 5682
rect 4460 5482 4490 5682
rect 4556 5482 4586 5682
rect 6348 5482 6378 5682
rect 6444 5482 6474 5682
rect 8236 5482 8266 5682
rect 8332 5482 8362 5682
rect 10124 5482 10154 5682
rect 10220 5482 10250 5682
rect 12012 5482 12042 5682
rect 12108 5482 12138 5682
rect 13900 5482 13930 5682
rect 13996 5482 14026 5682
rect 15782 5482 15812 5682
rect 15878 5482 15908 5682
rect 17670 5482 17700 5682
rect 17766 5482 17796 5682
rect 19558 5482 19588 5682
rect 19654 5482 19684 5682
rect 21446 5482 21476 5682
rect 21542 5482 21572 5682
rect 23334 5482 23364 5682
rect 23430 5482 23460 5682
rect 25222 5482 25252 5682
rect 25318 5482 25348 5682
rect 27110 5482 27140 5682
rect 27206 5482 27236 5682
rect 28998 5482 29028 5682
rect 29094 5482 29124 5682
rect 30886 5482 30916 5682
rect 30982 5482 31012 5682
rect 32774 5482 32804 5682
rect 32870 5482 32900 5682
rect 34662 5482 34692 5682
rect 34758 5482 34788 5682
rect 36550 5482 36580 5682
rect 36646 5482 36676 5682
rect 38438 5482 38468 5682
rect 38534 5482 38564 5682
rect 40326 5482 40356 5682
rect 40422 5482 40452 5682
rect 42214 5482 42244 5682
rect 42310 5482 42340 5682
rect 44102 5482 44132 5682
rect 44198 5482 44228 5682
rect 45984 5482 46014 5682
rect 46080 5482 46110 5682
rect 47872 5482 47902 5682
rect 47968 5482 47998 5682
rect 49760 5482 49790 5682
rect 49856 5482 49886 5682
rect 51648 5482 51678 5682
rect 51744 5482 51774 5682
rect 53536 5482 53566 5682
rect 53632 5482 53662 5682
rect 55424 5482 55454 5682
rect 55520 5482 55550 5682
rect 57312 5482 57342 5682
rect 57408 5482 57438 5682
rect 59200 5482 59230 5682
rect 59296 5482 59326 5682
rect 656 1758 686 1958
rect 752 1758 782 1958
rect 2544 1758 2574 1958
rect 2640 1758 2670 1958
rect 4432 1758 4462 1958
rect 4528 1758 4558 1958
rect 6320 1758 6350 1958
rect 6416 1758 6446 1958
rect 8208 1758 8238 1958
rect 8304 1758 8334 1958
rect 10096 1758 10126 1958
rect 10192 1758 10222 1958
rect 11984 1758 12014 1958
rect 12080 1758 12110 1958
rect 13872 1758 13902 1958
rect 13968 1758 13998 1958
rect 15754 1758 15784 1958
rect 15850 1758 15880 1958
rect 17642 1758 17672 1958
rect 17738 1758 17768 1958
rect 19530 1758 19560 1958
rect 19626 1758 19656 1958
rect 21418 1758 21448 1958
rect 21514 1758 21544 1958
rect 23306 1758 23336 1958
rect 23402 1758 23432 1958
rect 25194 1758 25224 1958
rect 25290 1758 25320 1958
rect 27082 1758 27112 1958
rect 27178 1758 27208 1958
rect 28970 1758 29000 1958
rect 29066 1758 29096 1958
rect 30858 1758 30888 1958
rect 30954 1758 30984 1958
rect 32746 1758 32776 1958
rect 32842 1758 32872 1958
rect 34634 1758 34664 1958
rect 34730 1758 34760 1958
rect 36522 1758 36552 1958
rect 36618 1758 36648 1958
rect 38410 1758 38440 1958
rect 38506 1758 38536 1958
rect 40298 1758 40328 1958
rect 40394 1758 40424 1958
rect 42186 1758 42216 1958
rect 42282 1758 42312 1958
rect 44074 1758 44104 1958
rect 44170 1758 44200 1958
rect 45956 1758 45986 1958
rect 46052 1758 46082 1958
rect 47844 1758 47874 1958
rect 47940 1758 47970 1958
rect 49732 1758 49762 1958
rect 49828 1758 49858 1958
rect 51620 1758 51650 1958
rect 51716 1758 51746 1958
rect 53508 1758 53538 1958
rect 53604 1758 53634 1958
rect 55396 1758 55426 1958
rect 55492 1758 55522 1958
rect 57284 1758 57314 1958
rect 57380 1758 57410 1958
rect 59172 1758 59202 1958
rect 59268 1758 59298 1958
rect 434 862 464 1062
rect 654 702 684 902
rect 750 702 780 902
rect 1080 862 1110 1062
rect 2322 862 2352 1062
rect 2542 702 2572 902
rect 2638 702 2668 902
rect 2968 862 2998 1062
rect 4210 862 4240 1062
rect 4430 702 4460 902
rect 4526 702 4556 902
rect 4856 862 4886 1062
rect 6098 862 6128 1062
rect 6318 702 6348 902
rect 6414 702 6444 902
rect 6744 862 6774 1062
rect 7986 862 8016 1062
rect 8206 702 8236 902
rect 8302 702 8332 902
rect 8632 862 8662 1062
rect 9874 862 9904 1062
rect 10094 702 10124 902
rect 10190 702 10220 902
rect 10520 862 10550 1062
rect 11762 862 11792 1062
rect 11982 702 12012 902
rect 12078 702 12108 902
rect 12408 862 12438 1062
rect 13650 862 13680 1062
rect 13870 702 13900 902
rect 13966 702 13996 902
rect 14296 862 14326 1062
rect 15532 862 15562 1062
rect 15752 702 15782 902
rect 15848 702 15878 902
rect 16178 862 16208 1062
rect 17420 862 17450 1062
rect 17640 702 17670 902
rect 17736 702 17766 902
rect 18066 862 18096 1062
rect 19308 862 19338 1062
rect 19528 702 19558 902
rect 19624 702 19654 902
rect 19954 862 19984 1062
rect 21196 862 21226 1062
rect 21416 702 21446 902
rect 21512 702 21542 902
rect 21842 862 21872 1062
rect 23084 862 23114 1062
rect 23304 702 23334 902
rect 23400 702 23430 902
rect 23730 862 23760 1062
rect 24972 862 25002 1062
rect 25192 702 25222 902
rect 25288 702 25318 902
rect 25618 862 25648 1062
rect 26860 862 26890 1062
rect 27080 702 27110 902
rect 27176 702 27206 902
rect 27506 862 27536 1062
rect 28748 862 28778 1062
rect 28968 702 28998 902
rect 29064 702 29094 902
rect 29394 862 29424 1062
rect 30636 862 30666 1062
rect 30856 702 30886 902
rect 30952 702 30982 902
rect 31282 862 31312 1062
rect 32524 862 32554 1062
rect 32744 702 32774 902
rect 32840 702 32870 902
rect 33170 862 33200 1062
rect 34412 862 34442 1062
rect 34632 702 34662 902
rect 34728 702 34758 902
rect 35058 862 35088 1062
rect 36300 862 36330 1062
rect 36520 702 36550 902
rect 36616 702 36646 902
rect 36946 862 36976 1062
rect 38188 862 38218 1062
rect 38408 702 38438 902
rect 38504 702 38534 902
rect 38834 862 38864 1062
rect 40076 862 40106 1062
rect 40296 702 40326 902
rect 40392 702 40422 902
rect 40722 862 40752 1062
rect 41964 862 41994 1062
rect 42184 702 42214 902
rect 42280 702 42310 902
rect 42610 862 42640 1062
rect 43852 862 43882 1062
rect 44072 702 44102 902
rect 44168 702 44198 902
rect 44498 862 44528 1062
rect 45734 862 45764 1062
rect 45954 702 45984 902
rect 46050 702 46080 902
rect 46380 862 46410 1062
rect 47622 862 47652 1062
rect 47842 702 47872 902
rect 47938 702 47968 902
rect 48268 862 48298 1062
rect 49510 862 49540 1062
rect 49730 702 49760 902
rect 49826 702 49856 902
rect 50156 862 50186 1062
rect 51398 862 51428 1062
rect 51618 702 51648 902
rect 51714 702 51744 902
rect 52044 862 52074 1062
rect 53286 862 53316 1062
rect 53506 702 53536 902
rect 53602 702 53632 902
rect 53932 862 53962 1062
rect 55174 862 55204 1062
rect 55394 702 55424 902
rect 55490 702 55520 902
rect 55820 862 55850 1062
rect 57062 862 57092 1062
rect 57282 702 57312 902
rect 57378 702 57408 902
rect 57708 862 57738 1062
rect 58950 862 58980 1062
rect 59170 702 59200 902
rect 59266 702 59296 902
rect 59596 862 59626 1062
<< ndiff >>
rect 608 7054 670 7068
rect 608 7020 620 7054
rect 654 7020 670 7054
rect 608 6986 670 7020
rect 608 6952 620 6986
rect 654 6952 670 6986
rect 608 6938 670 6952
rect 700 7054 766 7068
rect 700 7020 716 7054
rect 750 7020 766 7054
rect 700 6986 766 7020
rect 700 6952 716 6986
rect 750 6952 766 6986
rect 700 6938 766 6952
rect 796 7054 858 7068
rect 796 7020 812 7054
rect 846 7020 858 7054
rect 796 6986 858 7020
rect 796 6952 812 6986
rect 846 6952 858 6986
rect 796 6938 858 6952
rect 2496 7054 2558 7068
rect 2496 7020 2508 7054
rect 2542 7020 2558 7054
rect 2496 6986 2558 7020
rect 2496 6952 2508 6986
rect 2542 6952 2558 6986
rect 2496 6938 2558 6952
rect 2588 7054 2654 7068
rect 2588 7020 2604 7054
rect 2638 7020 2654 7054
rect 2588 6986 2654 7020
rect 2588 6952 2604 6986
rect 2638 6952 2654 6986
rect 2588 6938 2654 6952
rect 2684 7054 2746 7068
rect 2684 7020 2700 7054
rect 2734 7020 2746 7054
rect 2684 6986 2746 7020
rect 2684 6952 2700 6986
rect 2734 6952 2746 6986
rect 2684 6938 2746 6952
rect 4384 7054 4446 7068
rect 4384 7020 4396 7054
rect 4430 7020 4446 7054
rect 4384 6986 4446 7020
rect 4384 6952 4396 6986
rect 4430 6952 4446 6986
rect 4384 6938 4446 6952
rect 4476 7054 4542 7068
rect 4476 7020 4492 7054
rect 4526 7020 4542 7054
rect 4476 6986 4542 7020
rect 4476 6952 4492 6986
rect 4526 6952 4542 6986
rect 4476 6938 4542 6952
rect 4572 7054 4634 7068
rect 4572 7020 4588 7054
rect 4622 7020 4634 7054
rect 4572 6986 4634 7020
rect 4572 6952 4588 6986
rect 4622 6952 4634 6986
rect 4572 6938 4634 6952
rect 6272 7054 6334 7068
rect 6272 7020 6284 7054
rect 6318 7020 6334 7054
rect 6272 6986 6334 7020
rect 6272 6952 6284 6986
rect 6318 6952 6334 6986
rect 6272 6938 6334 6952
rect 6364 7054 6430 7068
rect 6364 7020 6380 7054
rect 6414 7020 6430 7054
rect 6364 6986 6430 7020
rect 6364 6952 6380 6986
rect 6414 6952 6430 6986
rect 6364 6938 6430 6952
rect 6460 7054 6522 7068
rect 6460 7020 6476 7054
rect 6510 7020 6522 7054
rect 6460 6986 6522 7020
rect 6460 6952 6476 6986
rect 6510 6952 6522 6986
rect 6460 6938 6522 6952
rect 8160 7054 8222 7068
rect 8160 7020 8172 7054
rect 8206 7020 8222 7054
rect 8160 6986 8222 7020
rect 8160 6952 8172 6986
rect 8206 6952 8222 6986
rect 8160 6938 8222 6952
rect 8252 7054 8318 7068
rect 8252 7020 8268 7054
rect 8302 7020 8318 7054
rect 8252 6986 8318 7020
rect 8252 6952 8268 6986
rect 8302 6952 8318 6986
rect 8252 6938 8318 6952
rect 8348 7054 8410 7068
rect 8348 7020 8364 7054
rect 8398 7020 8410 7054
rect 8348 6986 8410 7020
rect 8348 6952 8364 6986
rect 8398 6952 8410 6986
rect 8348 6938 8410 6952
rect 10048 7054 10110 7068
rect 10048 7020 10060 7054
rect 10094 7020 10110 7054
rect 10048 6986 10110 7020
rect 10048 6952 10060 6986
rect 10094 6952 10110 6986
rect 10048 6938 10110 6952
rect 10140 7054 10206 7068
rect 10140 7020 10156 7054
rect 10190 7020 10206 7054
rect 10140 6986 10206 7020
rect 10140 6952 10156 6986
rect 10190 6952 10206 6986
rect 10140 6938 10206 6952
rect 10236 7054 10298 7068
rect 10236 7020 10252 7054
rect 10286 7020 10298 7054
rect 10236 6986 10298 7020
rect 10236 6952 10252 6986
rect 10286 6952 10298 6986
rect 10236 6938 10298 6952
rect 11936 7054 11998 7068
rect 11936 7020 11948 7054
rect 11982 7020 11998 7054
rect 11936 6986 11998 7020
rect 11936 6952 11948 6986
rect 11982 6952 11998 6986
rect 11936 6938 11998 6952
rect 12028 7054 12094 7068
rect 12028 7020 12044 7054
rect 12078 7020 12094 7054
rect 12028 6986 12094 7020
rect 12028 6952 12044 6986
rect 12078 6952 12094 6986
rect 12028 6938 12094 6952
rect 12124 7054 12186 7068
rect 12124 7020 12140 7054
rect 12174 7020 12186 7054
rect 12124 6986 12186 7020
rect 12124 6952 12140 6986
rect 12174 6952 12186 6986
rect 12124 6938 12186 6952
rect 13824 7054 13886 7068
rect 13824 7020 13836 7054
rect 13870 7020 13886 7054
rect 13824 6986 13886 7020
rect 13824 6952 13836 6986
rect 13870 6952 13886 6986
rect 13824 6938 13886 6952
rect 13916 7054 13982 7068
rect 13916 7020 13932 7054
rect 13966 7020 13982 7054
rect 13916 6986 13982 7020
rect 13916 6952 13932 6986
rect 13966 6952 13982 6986
rect 13916 6938 13982 6952
rect 14012 7054 14074 7068
rect 14012 7020 14028 7054
rect 14062 7020 14074 7054
rect 14012 6986 14074 7020
rect 14012 6952 14028 6986
rect 14062 6952 14074 6986
rect 14012 6938 14074 6952
rect 15706 7054 15768 7068
rect 15706 7020 15718 7054
rect 15752 7020 15768 7054
rect 15706 6986 15768 7020
rect 15706 6952 15718 6986
rect 15752 6952 15768 6986
rect 15706 6938 15768 6952
rect 15798 7054 15864 7068
rect 15798 7020 15814 7054
rect 15848 7020 15864 7054
rect 15798 6986 15864 7020
rect 15798 6952 15814 6986
rect 15848 6952 15864 6986
rect 15798 6938 15864 6952
rect 15894 7054 15956 7068
rect 15894 7020 15910 7054
rect 15944 7020 15956 7054
rect 15894 6986 15956 7020
rect 15894 6952 15910 6986
rect 15944 6952 15956 6986
rect 15894 6938 15956 6952
rect 17594 7054 17656 7068
rect 17594 7020 17606 7054
rect 17640 7020 17656 7054
rect 17594 6986 17656 7020
rect 17594 6952 17606 6986
rect 17640 6952 17656 6986
rect 17594 6938 17656 6952
rect 17686 7054 17752 7068
rect 17686 7020 17702 7054
rect 17736 7020 17752 7054
rect 17686 6986 17752 7020
rect 17686 6952 17702 6986
rect 17736 6952 17752 6986
rect 17686 6938 17752 6952
rect 17782 7054 17844 7068
rect 17782 7020 17798 7054
rect 17832 7020 17844 7054
rect 17782 6986 17844 7020
rect 17782 6952 17798 6986
rect 17832 6952 17844 6986
rect 17782 6938 17844 6952
rect 19482 7054 19544 7068
rect 19482 7020 19494 7054
rect 19528 7020 19544 7054
rect 19482 6986 19544 7020
rect 19482 6952 19494 6986
rect 19528 6952 19544 6986
rect 19482 6938 19544 6952
rect 19574 7054 19640 7068
rect 19574 7020 19590 7054
rect 19624 7020 19640 7054
rect 19574 6986 19640 7020
rect 19574 6952 19590 6986
rect 19624 6952 19640 6986
rect 19574 6938 19640 6952
rect 19670 7054 19732 7068
rect 19670 7020 19686 7054
rect 19720 7020 19732 7054
rect 19670 6986 19732 7020
rect 19670 6952 19686 6986
rect 19720 6952 19732 6986
rect 19670 6938 19732 6952
rect 21370 7054 21432 7068
rect 21370 7020 21382 7054
rect 21416 7020 21432 7054
rect 21370 6986 21432 7020
rect 21370 6952 21382 6986
rect 21416 6952 21432 6986
rect 21370 6938 21432 6952
rect 21462 7054 21528 7068
rect 21462 7020 21478 7054
rect 21512 7020 21528 7054
rect 21462 6986 21528 7020
rect 21462 6952 21478 6986
rect 21512 6952 21528 6986
rect 21462 6938 21528 6952
rect 21558 7054 21620 7068
rect 21558 7020 21574 7054
rect 21608 7020 21620 7054
rect 21558 6986 21620 7020
rect 21558 6952 21574 6986
rect 21608 6952 21620 6986
rect 21558 6938 21620 6952
rect 23258 7054 23320 7068
rect 23258 7020 23270 7054
rect 23304 7020 23320 7054
rect 23258 6986 23320 7020
rect 23258 6952 23270 6986
rect 23304 6952 23320 6986
rect 23258 6938 23320 6952
rect 23350 7054 23416 7068
rect 23350 7020 23366 7054
rect 23400 7020 23416 7054
rect 23350 6986 23416 7020
rect 23350 6952 23366 6986
rect 23400 6952 23416 6986
rect 23350 6938 23416 6952
rect 23446 7054 23508 7068
rect 23446 7020 23462 7054
rect 23496 7020 23508 7054
rect 23446 6986 23508 7020
rect 23446 6952 23462 6986
rect 23496 6952 23508 6986
rect 23446 6938 23508 6952
rect 25146 7054 25208 7068
rect 25146 7020 25158 7054
rect 25192 7020 25208 7054
rect 25146 6986 25208 7020
rect 25146 6952 25158 6986
rect 25192 6952 25208 6986
rect 25146 6938 25208 6952
rect 25238 7054 25304 7068
rect 25238 7020 25254 7054
rect 25288 7020 25304 7054
rect 25238 6986 25304 7020
rect 25238 6952 25254 6986
rect 25288 6952 25304 6986
rect 25238 6938 25304 6952
rect 25334 7054 25396 7068
rect 25334 7020 25350 7054
rect 25384 7020 25396 7054
rect 25334 6986 25396 7020
rect 25334 6952 25350 6986
rect 25384 6952 25396 6986
rect 25334 6938 25396 6952
rect 27034 7054 27096 7068
rect 27034 7020 27046 7054
rect 27080 7020 27096 7054
rect 27034 6986 27096 7020
rect 27034 6952 27046 6986
rect 27080 6952 27096 6986
rect 27034 6938 27096 6952
rect 27126 7054 27192 7068
rect 27126 7020 27142 7054
rect 27176 7020 27192 7054
rect 27126 6986 27192 7020
rect 27126 6952 27142 6986
rect 27176 6952 27192 6986
rect 27126 6938 27192 6952
rect 27222 7054 27284 7068
rect 27222 7020 27238 7054
rect 27272 7020 27284 7054
rect 27222 6986 27284 7020
rect 27222 6952 27238 6986
rect 27272 6952 27284 6986
rect 27222 6938 27284 6952
rect 28922 7054 28984 7068
rect 28922 7020 28934 7054
rect 28968 7020 28984 7054
rect 28922 6986 28984 7020
rect 28922 6952 28934 6986
rect 28968 6952 28984 6986
rect 28922 6938 28984 6952
rect 29014 7054 29080 7068
rect 29014 7020 29030 7054
rect 29064 7020 29080 7054
rect 29014 6986 29080 7020
rect 29014 6952 29030 6986
rect 29064 6952 29080 6986
rect 29014 6938 29080 6952
rect 29110 7054 29172 7068
rect 29110 7020 29126 7054
rect 29160 7020 29172 7054
rect 29110 6986 29172 7020
rect 29110 6952 29126 6986
rect 29160 6952 29172 6986
rect 29110 6938 29172 6952
rect 30810 7054 30872 7068
rect 30810 7020 30822 7054
rect 30856 7020 30872 7054
rect 30810 6986 30872 7020
rect 30810 6952 30822 6986
rect 30856 6952 30872 6986
rect 30810 6938 30872 6952
rect 30902 7054 30968 7068
rect 30902 7020 30918 7054
rect 30952 7020 30968 7054
rect 30902 6986 30968 7020
rect 30902 6952 30918 6986
rect 30952 6952 30968 6986
rect 30902 6938 30968 6952
rect 30998 7054 31060 7068
rect 30998 7020 31014 7054
rect 31048 7020 31060 7054
rect 30998 6986 31060 7020
rect 30998 6952 31014 6986
rect 31048 6952 31060 6986
rect 30998 6938 31060 6952
rect 32698 7054 32760 7068
rect 32698 7020 32710 7054
rect 32744 7020 32760 7054
rect 32698 6986 32760 7020
rect 32698 6952 32710 6986
rect 32744 6952 32760 6986
rect 32698 6938 32760 6952
rect 32790 7054 32856 7068
rect 32790 7020 32806 7054
rect 32840 7020 32856 7054
rect 32790 6986 32856 7020
rect 32790 6952 32806 6986
rect 32840 6952 32856 6986
rect 32790 6938 32856 6952
rect 32886 7054 32948 7068
rect 32886 7020 32902 7054
rect 32936 7020 32948 7054
rect 32886 6986 32948 7020
rect 32886 6952 32902 6986
rect 32936 6952 32948 6986
rect 32886 6938 32948 6952
rect 34586 7054 34648 7068
rect 34586 7020 34598 7054
rect 34632 7020 34648 7054
rect 34586 6986 34648 7020
rect 34586 6952 34598 6986
rect 34632 6952 34648 6986
rect 34586 6938 34648 6952
rect 34678 7054 34744 7068
rect 34678 7020 34694 7054
rect 34728 7020 34744 7054
rect 34678 6986 34744 7020
rect 34678 6952 34694 6986
rect 34728 6952 34744 6986
rect 34678 6938 34744 6952
rect 34774 7054 34836 7068
rect 34774 7020 34790 7054
rect 34824 7020 34836 7054
rect 34774 6986 34836 7020
rect 34774 6952 34790 6986
rect 34824 6952 34836 6986
rect 34774 6938 34836 6952
rect 36474 7054 36536 7068
rect 36474 7020 36486 7054
rect 36520 7020 36536 7054
rect 36474 6986 36536 7020
rect 36474 6952 36486 6986
rect 36520 6952 36536 6986
rect 36474 6938 36536 6952
rect 36566 7054 36632 7068
rect 36566 7020 36582 7054
rect 36616 7020 36632 7054
rect 36566 6986 36632 7020
rect 36566 6952 36582 6986
rect 36616 6952 36632 6986
rect 36566 6938 36632 6952
rect 36662 7054 36724 7068
rect 36662 7020 36678 7054
rect 36712 7020 36724 7054
rect 36662 6986 36724 7020
rect 36662 6952 36678 6986
rect 36712 6952 36724 6986
rect 36662 6938 36724 6952
rect 38362 7054 38424 7068
rect 38362 7020 38374 7054
rect 38408 7020 38424 7054
rect 38362 6986 38424 7020
rect 38362 6952 38374 6986
rect 38408 6952 38424 6986
rect 38362 6938 38424 6952
rect 38454 7054 38520 7068
rect 38454 7020 38470 7054
rect 38504 7020 38520 7054
rect 38454 6986 38520 7020
rect 38454 6952 38470 6986
rect 38504 6952 38520 6986
rect 38454 6938 38520 6952
rect 38550 7054 38612 7068
rect 38550 7020 38566 7054
rect 38600 7020 38612 7054
rect 38550 6986 38612 7020
rect 38550 6952 38566 6986
rect 38600 6952 38612 6986
rect 38550 6938 38612 6952
rect 40250 7054 40312 7068
rect 40250 7020 40262 7054
rect 40296 7020 40312 7054
rect 40250 6986 40312 7020
rect 40250 6952 40262 6986
rect 40296 6952 40312 6986
rect 40250 6938 40312 6952
rect 40342 7054 40408 7068
rect 40342 7020 40358 7054
rect 40392 7020 40408 7054
rect 40342 6986 40408 7020
rect 40342 6952 40358 6986
rect 40392 6952 40408 6986
rect 40342 6938 40408 6952
rect 40438 7054 40500 7068
rect 40438 7020 40454 7054
rect 40488 7020 40500 7054
rect 40438 6986 40500 7020
rect 40438 6952 40454 6986
rect 40488 6952 40500 6986
rect 40438 6938 40500 6952
rect 42138 7054 42200 7068
rect 42138 7020 42150 7054
rect 42184 7020 42200 7054
rect 42138 6986 42200 7020
rect 42138 6952 42150 6986
rect 42184 6952 42200 6986
rect 42138 6938 42200 6952
rect 42230 7054 42296 7068
rect 42230 7020 42246 7054
rect 42280 7020 42296 7054
rect 42230 6986 42296 7020
rect 42230 6952 42246 6986
rect 42280 6952 42296 6986
rect 42230 6938 42296 6952
rect 42326 7054 42388 7068
rect 42326 7020 42342 7054
rect 42376 7020 42388 7054
rect 42326 6986 42388 7020
rect 42326 6952 42342 6986
rect 42376 6952 42388 6986
rect 42326 6938 42388 6952
rect 44026 7054 44088 7068
rect 44026 7020 44038 7054
rect 44072 7020 44088 7054
rect 44026 6986 44088 7020
rect 44026 6952 44038 6986
rect 44072 6952 44088 6986
rect 44026 6938 44088 6952
rect 44118 7054 44184 7068
rect 44118 7020 44134 7054
rect 44168 7020 44184 7054
rect 44118 6986 44184 7020
rect 44118 6952 44134 6986
rect 44168 6952 44184 6986
rect 44118 6938 44184 6952
rect 44214 7054 44276 7068
rect 44214 7020 44230 7054
rect 44264 7020 44276 7054
rect 44214 6986 44276 7020
rect 44214 6952 44230 6986
rect 44264 6952 44276 6986
rect 44214 6938 44276 6952
rect 45908 7054 45970 7068
rect 45908 7020 45920 7054
rect 45954 7020 45970 7054
rect 45908 6986 45970 7020
rect 45908 6952 45920 6986
rect 45954 6952 45970 6986
rect 45908 6938 45970 6952
rect 46000 7054 46066 7068
rect 46000 7020 46016 7054
rect 46050 7020 46066 7054
rect 46000 6986 46066 7020
rect 46000 6952 46016 6986
rect 46050 6952 46066 6986
rect 46000 6938 46066 6952
rect 46096 7054 46158 7068
rect 46096 7020 46112 7054
rect 46146 7020 46158 7054
rect 46096 6986 46158 7020
rect 46096 6952 46112 6986
rect 46146 6952 46158 6986
rect 46096 6938 46158 6952
rect 47796 7054 47858 7068
rect 47796 7020 47808 7054
rect 47842 7020 47858 7054
rect 47796 6986 47858 7020
rect 47796 6952 47808 6986
rect 47842 6952 47858 6986
rect 47796 6938 47858 6952
rect 47888 7054 47954 7068
rect 47888 7020 47904 7054
rect 47938 7020 47954 7054
rect 47888 6986 47954 7020
rect 47888 6952 47904 6986
rect 47938 6952 47954 6986
rect 47888 6938 47954 6952
rect 47984 7054 48046 7068
rect 47984 7020 48000 7054
rect 48034 7020 48046 7054
rect 47984 6986 48046 7020
rect 47984 6952 48000 6986
rect 48034 6952 48046 6986
rect 47984 6938 48046 6952
rect 49684 7054 49746 7068
rect 49684 7020 49696 7054
rect 49730 7020 49746 7054
rect 49684 6986 49746 7020
rect 49684 6952 49696 6986
rect 49730 6952 49746 6986
rect 49684 6938 49746 6952
rect 49776 7054 49842 7068
rect 49776 7020 49792 7054
rect 49826 7020 49842 7054
rect 49776 6986 49842 7020
rect 49776 6952 49792 6986
rect 49826 6952 49842 6986
rect 49776 6938 49842 6952
rect 49872 7054 49934 7068
rect 49872 7020 49888 7054
rect 49922 7020 49934 7054
rect 49872 6986 49934 7020
rect 49872 6952 49888 6986
rect 49922 6952 49934 6986
rect 49872 6938 49934 6952
rect 51572 7054 51634 7068
rect 51572 7020 51584 7054
rect 51618 7020 51634 7054
rect 51572 6986 51634 7020
rect 51572 6952 51584 6986
rect 51618 6952 51634 6986
rect 51572 6938 51634 6952
rect 51664 7054 51730 7068
rect 51664 7020 51680 7054
rect 51714 7020 51730 7054
rect 51664 6986 51730 7020
rect 51664 6952 51680 6986
rect 51714 6952 51730 6986
rect 51664 6938 51730 6952
rect 51760 7054 51822 7068
rect 51760 7020 51776 7054
rect 51810 7020 51822 7054
rect 51760 6986 51822 7020
rect 51760 6952 51776 6986
rect 51810 6952 51822 6986
rect 51760 6938 51822 6952
rect 53460 7054 53522 7068
rect 53460 7020 53472 7054
rect 53506 7020 53522 7054
rect 53460 6986 53522 7020
rect 53460 6952 53472 6986
rect 53506 6952 53522 6986
rect 53460 6938 53522 6952
rect 53552 7054 53618 7068
rect 53552 7020 53568 7054
rect 53602 7020 53618 7054
rect 53552 6986 53618 7020
rect 53552 6952 53568 6986
rect 53602 6952 53618 6986
rect 53552 6938 53618 6952
rect 53648 7054 53710 7068
rect 53648 7020 53664 7054
rect 53698 7020 53710 7054
rect 53648 6986 53710 7020
rect 53648 6952 53664 6986
rect 53698 6952 53710 6986
rect 53648 6938 53710 6952
rect 55348 7054 55410 7068
rect 55348 7020 55360 7054
rect 55394 7020 55410 7054
rect 55348 6986 55410 7020
rect 55348 6952 55360 6986
rect 55394 6952 55410 6986
rect 55348 6938 55410 6952
rect 55440 7054 55506 7068
rect 55440 7020 55456 7054
rect 55490 7020 55506 7054
rect 55440 6986 55506 7020
rect 55440 6952 55456 6986
rect 55490 6952 55506 6986
rect 55440 6938 55506 6952
rect 55536 7054 55598 7068
rect 55536 7020 55552 7054
rect 55586 7020 55598 7054
rect 55536 6986 55598 7020
rect 55536 6952 55552 6986
rect 55586 6952 55598 6986
rect 55536 6938 55598 6952
rect 57236 7054 57298 7068
rect 57236 7020 57248 7054
rect 57282 7020 57298 7054
rect 57236 6986 57298 7020
rect 57236 6952 57248 6986
rect 57282 6952 57298 6986
rect 57236 6938 57298 6952
rect 57328 7054 57394 7068
rect 57328 7020 57344 7054
rect 57378 7020 57394 7054
rect 57328 6986 57394 7020
rect 57328 6952 57344 6986
rect 57378 6952 57394 6986
rect 57328 6938 57394 6952
rect 57424 7054 57486 7068
rect 57424 7020 57440 7054
rect 57474 7020 57486 7054
rect 57424 6986 57486 7020
rect 57424 6952 57440 6986
rect 57474 6952 57486 6986
rect 57424 6938 57486 6952
rect 59124 7054 59186 7068
rect 59124 7020 59136 7054
rect 59170 7020 59186 7054
rect 59124 6986 59186 7020
rect 59124 6952 59136 6986
rect 59170 6952 59186 6986
rect 59124 6938 59186 6952
rect 59216 7054 59282 7068
rect 59216 7020 59232 7054
rect 59266 7020 59282 7054
rect 59216 6986 59282 7020
rect 59216 6952 59232 6986
rect 59266 6952 59282 6986
rect 59216 6938 59282 6952
rect 59312 7054 59374 7068
rect 59312 7020 59328 7054
rect 59362 7020 59374 7054
rect 59312 6986 59374 7020
rect 59312 6952 59328 6986
rect 59362 6952 59374 6986
rect 59312 6938 59374 6952
rect -365 6773 -313 6815
rect -365 6739 -357 6773
rect -323 6739 -313 6773
rect -365 6711 -313 6739
rect -283 6803 -225 6815
rect -283 6769 -271 6803
rect -237 6769 -225 6803
rect -283 6711 -225 6769
rect -195 6790 -143 6815
rect -195 6756 -185 6790
rect -151 6756 -143 6790
rect -195 6711 -143 6756
rect 28 6797 80 6813
rect 28 6763 36 6797
rect 70 6763 80 6797
rect 28 6729 80 6763
rect 28 6695 36 6729
rect 70 6695 80 6729
rect 28 6683 80 6695
rect 110 6797 162 6813
rect 110 6763 120 6797
rect 154 6763 162 6797
rect 1224 6805 1276 6821
rect 1224 6771 1232 6805
rect 1266 6771 1276 6805
rect 110 6729 162 6763
rect 110 6695 120 6729
rect 154 6695 162 6729
rect 110 6683 162 6695
rect 1224 6737 1276 6771
rect 1224 6703 1232 6737
rect 1266 6703 1276 6737
rect 1224 6691 1276 6703
rect 1306 6805 1358 6821
rect 1306 6771 1316 6805
rect 1350 6771 1358 6805
rect 1306 6737 1358 6771
rect 1306 6703 1316 6737
rect 1350 6703 1358 6737
rect 1523 6773 1575 6815
rect 1523 6739 1531 6773
rect 1565 6739 1575 6773
rect 1523 6711 1575 6739
rect 1605 6803 1663 6815
rect 1605 6769 1617 6803
rect 1651 6769 1663 6803
rect 1605 6711 1663 6769
rect 1693 6790 1745 6815
rect 1693 6756 1703 6790
rect 1737 6756 1745 6790
rect 1693 6711 1745 6756
rect 1916 6797 1968 6813
rect 1916 6763 1924 6797
rect 1958 6763 1968 6797
rect 1916 6729 1968 6763
rect 1306 6691 1358 6703
rect 1916 6695 1924 6729
rect 1958 6695 1968 6729
rect 1916 6683 1968 6695
rect 1998 6797 2050 6813
rect 1998 6763 2008 6797
rect 2042 6763 2050 6797
rect 3112 6805 3164 6821
rect 3112 6771 3120 6805
rect 3154 6771 3164 6805
rect 1998 6729 2050 6763
rect 1998 6695 2008 6729
rect 2042 6695 2050 6729
rect 1998 6683 2050 6695
rect 3112 6737 3164 6771
rect 3112 6703 3120 6737
rect 3154 6703 3164 6737
rect 3112 6691 3164 6703
rect 3194 6805 3246 6821
rect 3194 6771 3204 6805
rect 3238 6771 3246 6805
rect 3194 6737 3246 6771
rect 3194 6703 3204 6737
rect 3238 6703 3246 6737
rect 3411 6773 3463 6815
rect 3411 6739 3419 6773
rect 3453 6739 3463 6773
rect 3411 6711 3463 6739
rect 3493 6803 3551 6815
rect 3493 6769 3505 6803
rect 3539 6769 3551 6803
rect 3493 6711 3551 6769
rect 3581 6790 3633 6815
rect 3581 6756 3591 6790
rect 3625 6756 3633 6790
rect 3581 6711 3633 6756
rect 3804 6797 3856 6813
rect 3804 6763 3812 6797
rect 3846 6763 3856 6797
rect 3804 6729 3856 6763
rect 3194 6691 3246 6703
rect 3804 6695 3812 6729
rect 3846 6695 3856 6729
rect 3804 6683 3856 6695
rect 3886 6797 3938 6813
rect 3886 6763 3896 6797
rect 3930 6763 3938 6797
rect 5000 6805 5052 6821
rect 5000 6771 5008 6805
rect 5042 6771 5052 6805
rect 3886 6729 3938 6763
rect 3886 6695 3896 6729
rect 3930 6695 3938 6729
rect 3886 6683 3938 6695
rect 5000 6737 5052 6771
rect 5000 6703 5008 6737
rect 5042 6703 5052 6737
rect 5000 6691 5052 6703
rect 5082 6805 5134 6821
rect 5082 6771 5092 6805
rect 5126 6771 5134 6805
rect 5082 6737 5134 6771
rect 5082 6703 5092 6737
rect 5126 6703 5134 6737
rect 5299 6773 5351 6815
rect 5299 6739 5307 6773
rect 5341 6739 5351 6773
rect 5299 6711 5351 6739
rect 5381 6803 5439 6815
rect 5381 6769 5393 6803
rect 5427 6769 5439 6803
rect 5381 6711 5439 6769
rect 5469 6790 5521 6815
rect 5469 6756 5479 6790
rect 5513 6756 5521 6790
rect 5469 6711 5521 6756
rect 5692 6797 5744 6813
rect 5692 6763 5700 6797
rect 5734 6763 5744 6797
rect 5692 6729 5744 6763
rect 5082 6691 5134 6703
rect 5692 6695 5700 6729
rect 5734 6695 5744 6729
rect 5692 6683 5744 6695
rect 5774 6797 5826 6813
rect 5774 6763 5784 6797
rect 5818 6763 5826 6797
rect 6888 6805 6940 6821
rect 6888 6771 6896 6805
rect 6930 6771 6940 6805
rect 5774 6729 5826 6763
rect 5774 6695 5784 6729
rect 5818 6695 5826 6729
rect 5774 6683 5826 6695
rect 6888 6737 6940 6771
rect 6888 6703 6896 6737
rect 6930 6703 6940 6737
rect 6888 6691 6940 6703
rect 6970 6805 7022 6821
rect 6970 6771 6980 6805
rect 7014 6771 7022 6805
rect 6970 6737 7022 6771
rect 6970 6703 6980 6737
rect 7014 6703 7022 6737
rect 7187 6773 7239 6815
rect 7187 6739 7195 6773
rect 7229 6739 7239 6773
rect 7187 6711 7239 6739
rect 7269 6803 7327 6815
rect 7269 6769 7281 6803
rect 7315 6769 7327 6803
rect 7269 6711 7327 6769
rect 7357 6790 7409 6815
rect 7357 6756 7367 6790
rect 7401 6756 7409 6790
rect 7357 6711 7409 6756
rect 7580 6797 7632 6813
rect 7580 6763 7588 6797
rect 7622 6763 7632 6797
rect 7580 6729 7632 6763
rect 6970 6691 7022 6703
rect 7580 6695 7588 6729
rect 7622 6695 7632 6729
rect 7580 6683 7632 6695
rect 7662 6797 7714 6813
rect 7662 6763 7672 6797
rect 7706 6763 7714 6797
rect 8776 6805 8828 6821
rect 8776 6771 8784 6805
rect 8818 6771 8828 6805
rect 7662 6729 7714 6763
rect 7662 6695 7672 6729
rect 7706 6695 7714 6729
rect 7662 6683 7714 6695
rect 8776 6737 8828 6771
rect 8776 6703 8784 6737
rect 8818 6703 8828 6737
rect 8776 6691 8828 6703
rect 8858 6805 8910 6821
rect 8858 6771 8868 6805
rect 8902 6771 8910 6805
rect 8858 6737 8910 6771
rect 8858 6703 8868 6737
rect 8902 6703 8910 6737
rect 9075 6773 9127 6815
rect 9075 6739 9083 6773
rect 9117 6739 9127 6773
rect 9075 6711 9127 6739
rect 9157 6803 9215 6815
rect 9157 6769 9169 6803
rect 9203 6769 9215 6803
rect 9157 6711 9215 6769
rect 9245 6790 9297 6815
rect 9245 6756 9255 6790
rect 9289 6756 9297 6790
rect 9245 6711 9297 6756
rect 9468 6797 9520 6813
rect 9468 6763 9476 6797
rect 9510 6763 9520 6797
rect 9468 6729 9520 6763
rect 8858 6691 8910 6703
rect 9468 6695 9476 6729
rect 9510 6695 9520 6729
rect 9468 6683 9520 6695
rect 9550 6797 9602 6813
rect 9550 6763 9560 6797
rect 9594 6763 9602 6797
rect 10664 6805 10716 6821
rect 10664 6771 10672 6805
rect 10706 6771 10716 6805
rect 9550 6729 9602 6763
rect 9550 6695 9560 6729
rect 9594 6695 9602 6729
rect 9550 6683 9602 6695
rect 10664 6737 10716 6771
rect 10664 6703 10672 6737
rect 10706 6703 10716 6737
rect 10664 6691 10716 6703
rect 10746 6805 10798 6821
rect 10746 6771 10756 6805
rect 10790 6771 10798 6805
rect 10746 6737 10798 6771
rect 10746 6703 10756 6737
rect 10790 6703 10798 6737
rect 10963 6773 11015 6815
rect 10963 6739 10971 6773
rect 11005 6739 11015 6773
rect 10963 6711 11015 6739
rect 11045 6803 11103 6815
rect 11045 6769 11057 6803
rect 11091 6769 11103 6803
rect 11045 6711 11103 6769
rect 11133 6790 11185 6815
rect 11133 6756 11143 6790
rect 11177 6756 11185 6790
rect 11133 6711 11185 6756
rect 11356 6797 11408 6813
rect 11356 6763 11364 6797
rect 11398 6763 11408 6797
rect 11356 6729 11408 6763
rect 10746 6691 10798 6703
rect 11356 6695 11364 6729
rect 11398 6695 11408 6729
rect 11356 6683 11408 6695
rect 11438 6797 11490 6813
rect 11438 6763 11448 6797
rect 11482 6763 11490 6797
rect 12552 6805 12604 6821
rect 12552 6771 12560 6805
rect 12594 6771 12604 6805
rect 11438 6729 11490 6763
rect 11438 6695 11448 6729
rect 11482 6695 11490 6729
rect 11438 6683 11490 6695
rect 12552 6737 12604 6771
rect 12552 6703 12560 6737
rect 12594 6703 12604 6737
rect 12552 6691 12604 6703
rect 12634 6805 12686 6821
rect 12634 6771 12644 6805
rect 12678 6771 12686 6805
rect 12634 6737 12686 6771
rect 12634 6703 12644 6737
rect 12678 6703 12686 6737
rect 12851 6773 12903 6815
rect 12851 6739 12859 6773
rect 12893 6739 12903 6773
rect 12851 6711 12903 6739
rect 12933 6803 12991 6815
rect 12933 6769 12945 6803
rect 12979 6769 12991 6803
rect 12933 6711 12991 6769
rect 13021 6790 13073 6815
rect 13021 6756 13031 6790
rect 13065 6756 13073 6790
rect 13021 6711 13073 6756
rect 13244 6797 13296 6813
rect 13244 6763 13252 6797
rect 13286 6763 13296 6797
rect 13244 6729 13296 6763
rect 12634 6691 12686 6703
rect 13244 6695 13252 6729
rect 13286 6695 13296 6729
rect 13244 6683 13296 6695
rect 13326 6797 13378 6813
rect 13326 6763 13336 6797
rect 13370 6763 13378 6797
rect 14440 6805 14492 6821
rect 14440 6771 14448 6805
rect 14482 6771 14492 6805
rect 13326 6729 13378 6763
rect 13326 6695 13336 6729
rect 13370 6695 13378 6729
rect 13326 6683 13378 6695
rect 14440 6737 14492 6771
rect 14440 6703 14448 6737
rect 14482 6703 14492 6737
rect 14440 6691 14492 6703
rect 14522 6805 14574 6821
rect 14522 6771 14532 6805
rect 14566 6771 14574 6805
rect 14522 6737 14574 6771
rect 14522 6703 14532 6737
rect 14566 6703 14574 6737
rect 14733 6773 14785 6815
rect 14733 6739 14741 6773
rect 14775 6739 14785 6773
rect 14733 6711 14785 6739
rect 14815 6803 14873 6815
rect 14815 6769 14827 6803
rect 14861 6769 14873 6803
rect 14815 6711 14873 6769
rect 14903 6790 14955 6815
rect 14903 6756 14913 6790
rect 14947 6756 14955 6790
rect 14903 6711 14955 6756
rect 15126 6797 15178 6813
rect 15126 6763 15134 6797
rect 15168 6763 15178 6797
rect 15126 6729 15178 6763
rect 14522 6691 14574 6703
rect 15126 6695 15134 6729
rect 15168 6695 15178 6729
rect 15126 6683 15178 6695
rect 15208 6797 15260 6813
rect 15208 6763 15218 6797
rect 15252 6763 15260 6797
rect 16322 6805 16374 6821
rect 16322 6771 16330 6805
rect 16364 6771 16374 6805
rect 15208 6729 15260 6763
rect 15208 6695 15218 6729
rect 15252 6695 15260 6729
rect 15208 6683 15260 6695
rect 16322 6737 16374 6771
rect 16322 6703 16330 6737
rect 16364 6703 16374 6737
rect 16322 6691 16374 6703
rect 16404 6805 16456 6821
rect 16404 6771 16414 6805
rect 16448 6771 16456 6805
rect 16404 6737 16456 6771
rect 16404 6703 16414 6737
rect 16448 6703 16456 6737
rect 16621 6773 16673 6815
rect 16621 6739 16629 6773
rect 16663 6739 16673 6773
rect 16621 6711 16673 6739
rect 16703 6803 16761 6815
rect 16703 6769 16715 6803
rect 16749 6769 16761 6803
rect 16703 6711 16761 6769
rect 16791 6790 16843 6815
rect 16791 6756 16801 6790
rect 16835 6756 16843 6790
rect 16791 6711 16843 6756
rect 17014 6797 17066 6813
rect 17014 6763 17022 6797
rect 17056 6763 17066 6797
rect 17014 6729 17066 6763
rect 16404 6691 16456 6703
rect 17014 6695 17022 6729
rect 17056 6695 17066 6729
rect 17014 6683 17066 6695
rect 17096 6797 17148 6813
rect 17096 6763 17106 6797
rect 17140 6763 17148 6797
rect 18210 6805 18262 6821
rect 18210 6771 18218 6805
rect 18252 6771 18262 6805
rect 17096 6729 17148 6763
rect 17096 6695 17106 6729
rect 17140 6695 17148 6729
rect 17096 6683 17148 6695
rect 18210 6737 18262 6771
rect 18210 6703 18218 6737
rect 18252 6703 18262 6737
rect 18210 6691 18262 6703
rect 18292 6805 18344 6821
rect 18292 6771 18302 6805
rect 18336 6771 18344 6805
rect 18292 6737 18344 6771
rect 18292 6703 18302 6737
rect 18336 6703 18344 6737
rect 18509 6773 18561 6815
rect 18509 6739 18517 6773
rect 18551 6739 18561 6773
rect 18509 6711 18561 6739
rect 18591 6803 18649 6815
rect 18591 6769 18603 6803
rect 18637 6769 18649 6803
rect 18591 6711 18649 6769
rect 18679 6790 18731 6815
rect 18679 6756 18689 6790
rect 18723 6756 18731 6790
rect 18679 6711 18731 6756
rect 18902 6797 18954 6813
rect 18902 6763 18910 6797
rect 18944 6763 18954 6797
rect 18902 6729 18954 6763
rect 18292 6691 18344 6703
rect 18902 6695 18910 6729
rect 18944 6695 18954 6729
rect 18902 6683 18954 6695
rect 18984 6797 19036 6813
rect 18984 6763 18994 6797
rect 19028 6763 19036 6797
rect 20098 6805 20150 6821
rect 20098 6771 20106 6805
rect 20140 6771 20150 6805
rect 18984 6729 19036 6763
rect 18984 6695 18994 6729
rect 19028 6695 19036 6729
rect 18984 6683 19036 6695
rect 20098 6737 20150 6771
rect 20098 6703 20106 6737
rect 20140 6703 20150 6737
rect 20098 6691 20150 6703
rect 20180 6805 20232 6821
rect 20180 6771 20190 6805
rect 20224 6771 20232 6805
rect 20180 6737 20232 6771
rect 20180 6703 20190 6737
rect 20224 6703 20232 6737
rect 20397 6773 20449 6815
rect 20397 6739 20405 6773
rect 20439 6739 20449 6773
rect 20397 6711 20449 6739
rect 20479 6803 20537 6815
rect 20479 6769 20491 6803
rect 20525 6769 20537 6803
rect 20479 6711 20537 6769
rect 20567 6790 20619 6815
rect 20567 6756 20577 6790
rect 20611 6756 20619 6790
rect 20567 6711 20619 6756
rect 20790 6797 20842 6813
rect 20790 6763 20798 6797
rect 20832 6763 20842 6797
rect 20790 6729 20842 6763
rect 20180 6691 20232 6703
rect 20790 6695 20798 6729
rect 20832 6695 20842 6729
rect 20790 6683 20842 6695
rect 20872 6797 20924 6813
rect 20872 6763 20882 6797
rect 20916 6763 20924 6797
rect 21986 6805 22038 6821
rect 21986 6771 21994 6805
rect 22028 6771 22038 6805
rect 20872 6729 20924 6763
rect 20872 6695 20882 6729
rect 20916 6695 20924 6729
rect 20872 6683 20924 6695
rect 21986 6737 22038 6771
rect 21986 6703 21994 6737
rect 22028 6703 22038 6737
rect 21986 6691 22038 6703
rect 22068 6805 22120 6821
rect 22068 6771 22078 6805
rect 22112 6771 22120 6805
rect 22068 6737 22120 6771
rect 22068 6703 22078 6737
rect 22112 6703 22120 6737
rect 22285 6773 22337 6815
rect 22285 6739 22293 6773
rect 22327 6739 22337 6773
rect 22285 6711 22337 6739
rect 22367 6803 22425 6815
rect 22367 6769 22379 6803
rect 22413 6769 22425 6803
rect 22367 6711 22425 6769
rect 22455 6790 22507 6815
rect 22455 6756 22465 6790
rect 22499 6756 22507 6790
rect 22455 6711 22507 6756
rect 22678 6797 22730 6813
rect 22678 6763 22686 6797
rect 22720 6763 22730 6797
rect 22678 6729 22730 6763
rect 22068 6691 22120 6703
rect 22678 6695 22686 6729
rect 22720 6695 22730 6729
rect 22678 6683 22730 6695
rect 22760 6797 22812 6813
rect 22760 6763 22770 6797
rect 22804 6763 22812 6797
rect 23874 6805 23926 6821
rect 23874 6771 23882 6805
rect 23916 6771 23926 6805
rect 22760 6729 22812 6763
rect 22760 6695 22770 6729
rect 22804 6695 22812 6729
rect 22760 6683 22812 6695
rect 23874 6737 23926 6771
rect 23874 6703 23882 6737
rect 23916 6703 23926 6737
rect 23874 6691 23926 6703
rect 23956 6805 24008 6821
rect 23956 6771 23966 6805
rect 24000 6771 24008 6805
rect 23956 6737 24008 6771
rect 23956 6703 23966 6737
rect 24000 6703 24008 6737
rect 24173 6773 24225 6815
rect 24173 6739 24181 6773
rect 24215 6739 24225 6773
rect 24173 6711 24225 6739
rect 24255 6803 24313 6815
rect 24255 6769 24267 6803
rect 24301 6769 24313 6803
rect 24255 6711 24313 6769
rect 24343 6790 24395 6815
rect 24343 6756 24353 6790
rect 24387 6756 24395 6790
rect 24343 6711 24395 6756
rect 24566 6797 24618 6813
rect 24566 6763 24574 6797
rect 24608 6763 24618 6797
rect 24566 6729 24618 6763
rect 23956 6691 24008 6703
rect 24566 6695 24574 6729
rect 24608 6695 24618 6729
rect 24566 6683 24618 6695
rect 24648 6797 24700 6813
rect 24648 6763 24658 6797
rect 24692 6763 24700 6797
rect 25762 6805 25814 6821
rect 25762 6771 25770 6805
rect 25804 6771 25814 6805
rect 24648 6729 24700 6763
rect 24648 6695 24658 6729
rect 24692 6695 24700 6729
rect 24648 6683 24700 6695
rect 25762 6737 25814 6771
rect 25762 6703 25770 6737
rect 25804 6703 25814 6737
rect 25762 6691 25814 6703
rect 25844 6805 25896 6821
rect 25844 6771 25854 6805
rect 25888 6771 25896 6805
rect 25844 6737 25896 6771
rect 25844 6703 25854 6737
rect 25888 6703 25896 6737
rect 26061 6773 26113 6815
rect 26061 6739 26069 6773
rect 26103 6739 26113 6773
rect 26061 6711 26113 6739
rect 26143 6803 26201 6815
rect 26143 6769 26155 6803
rect 26189 6769 26201 6803
rect 26143 6711 26201 6769
rect 26231 6790 26283 6815
rect 26231 6756 26241 6790
rect 26275 6756 26283 6790
rect 26231 6711 26283 6756
rect 26454 6797 26506 6813
rect 26454 6763 26462 6797
rect 26496 6763 26506 6797
rect 26454 6729 26506 6763
rect 25844 6691 25896 6703
rect 26454 6695 26462 6729
rect 26496 6695 26506 6729
rect 26454 6683 26506 6695
rect 26536 6797 26588 6813
rect 26536 6763 26546 6797
rect 26580 6763 26588 6797
rect 27650 6805 27702 6821
rect 27650 6771 27658 6805
rect 27692 6771 27702 6805
rect 26536 6729 26588 6763
rect 26536 6695 26546 6729
rect 26580 6695 26588 6729
rect 26536 6683 26588 6695
rect 27650 6737 27702 6771
rect 27650 6703 27658 6737
rect 27692 6703 27702 6737
rect 27650 6691 27702 6703
rect 27732 6805 27784 6821
rect 27732 6771 27742 6805
rect 27776 6771 27784 6805
rect 27732 6737 27784 6771
rect 27732 6703 27742 6737
rect 27776 6703 27784 6737
rect 27949 6773 28001 6815
rect 27949 6739 27957 6773
rect 27991 6739 28001 6773
rect 27949 6711 28001 6739
rect 28031 6803 28089 6815
rect 28031 6769 28043 6803
rect 28077 6769 28089 6803
rect 28031 6711 28089 6769
rect 28119 6790 28171 6815
rect 28119 6756 28129 6790
rect 28163 6756 28171 6790
rect 28119 6711 28171 6756
rect 28342 6797 28394 6813
rect 28342 6763 28350 6797
rect 28384 6763 28394 6797
rect 28342 6729 28394 6763
rect 27732 6691 27784 6703
rect 28342 6695 28350 6729
rect 28384 6695 28394 6729
rect 28342 6683 28394 6695
rect 28424 6797 28476 6813
rect 28424 6763 28434 6797
rect 28468 6763 28476 6797
rect 29538 6805 29590 6821
rect 29538 6771 29546 6805
rect 29580 6771 29590 6805
rect 28424 6729 28476 6763
rect 28424 6695 28434 6729
rect 28468 6695 28476 6729
rect 28424 6683 28476 6695
rect 29538 6737 29590 6771
rect 29538 6703 29546 6737
rect 29580 6703 29590 6737
rect 29538 6691 29590 6703
rect 29620 6805 29672 6821
rect 29620 6771 29630 6805
rect 29664 6771 29672 6805
rect 29620 6737 29672 6771
rect 29620 6703 29630 6737
rect 29664 6703 29672 6737
rect 29837 6773 29889 6815
rect 29837 6739 29845 6773
rect 29879 6739 29889 6773
rect 29837 6711 29889 6739
rect 29919 6803 29977 6815
rect 29919 6769 29931 6803
rect 29965 6769 29977 6803
rect 29919 6711 29977 6769
rect 30007 6790 30059 6815
rect 30007 6756 30017 6790
rect 30051 6756 30059 6790
rect 30007 6711 30059 6756
rect 30230 6797 30282 6813
rect 30230 6763 30238 6797
rect 30272 6763 30282 6797
rect 30230 6729 30282 6763
rect 29620 6691 29672 6703
rect 30230 6695 30238 6729
rect 30272 6695 30282 6729
rect 30230 6683 30282 6695
rect 30312 6797 30364 6813
rect 30312 6763 30322 6797
rect 30356 6763 30364 6797
rect 31426 6805 31478 6821
rect 31426 6771 31434 6805
rect 31468 6771 31478 6805
rect 30312 6729 30364 6763
rect 30312 6695 30322 6729
rect 30356 6695 30364 6729
rect 30312 6683 30364 6695
rect 31426 6737 31478 6771
rect 31426 6703 31434 6737
rect 31468 6703 31478 6737
rect 31426 6691 31478 6703
rect 31508 6805 31560 6821
rect 31508 6771 31518 6805
rect 31552 6771 31560 6805
rect 31508 6737 31560 6771
rect 31508 6703 31518 6737
rect 31552 6703 31560 6737
rect 31725 6773 31777 6815
rect 31725 6739 31733 6773
rect 31767 6739 31777 6773
rect 31725 6711 31777 6739
rect 31807 6803 31865 6815
rect 31807 6769 31819 6803
rect 31853 6769 31865 6803
rect 31807 6711 31865 6769
rect 31895 6790 31947 6815
rect 31895 6756 31905 6790
rect 31939 6756 31947 6790
rect 31895 6711 31947 6756
rect 32118 6797 32170 6813
rect 32118 6763 32126 6797
rect 32160 6763 32170 6797
rect 32118 6729 32170 6763
rect 31508 6691 31560 6703
rect 32118 6695 32126 6729
rect 32160 6695 32170 6729
rect 32118 6683 32170 6695
rect 32200 6797 32252 6813
rect 32200 6763 32210 6797
rect 32244 6763 32252 6797
rect 33314 6805 33366 6821
rect 33314 6771 33322 6805
rect 33356 6771 33366 6805
rect 32200 6729 32252 6763
rect 32200 6695 32210 6729
rect 32244 6695 32252 6729
rect 32200 6683 32252 6695
rect 33314 6737 33366 6771
rect 33314 6703 33322 6737
rect 33356 6703 33366 6737
rect 33314 6691 33366 6703
rect 33396 6805 33448 6821
rect 33396 6771 33406 6805
rect 33440 6771 33448 6805
rect 33396 6737 33448 6771
rect 33396 6703 33406 6737
rect 33440 6703 33448 6737
rect 33613 6773 33665 6815
rect 33613 6739 33621 6773
rect 33655 6739 33665 6773
rect 33613 6711 33665 6739
rect 33695 6803 33753 6815
rect 33695 6769 33707 6803
rect 33741 6769 33753 6803
rect 33695 6711 33753 6769
rect 33783 6790 33835 6815
rect 33783 6756 33793 6790
rect 33827 6756 33835 6790
rect 33783 6711 33835 6756
rect 34006 6797 34058 6813
rect 34006 6763 34014 6797
rect 34048 6763 34058 6797
rect 34006 6729 34058 6763
rect 33396 6691 33448 6703
rect 34006 6695 34014 6729
rect 34048 6695 34058 6729
rect 34006 6683 34058 6695
rect 34088 6797 34140 6813
rect 34088 6763 34098 6797
rect 34132 6763 34140 6797
rect 35202 6805 35254 6821
rect 35202 6771 35210 6805
rect 35244 6771 35254 6805
rect 34088 6729 34140 6763
rect 34088 6695 34098 6729
rect 34132 6695 34140 6729
rect 34088 6683 34140 6695
rect 35202 6737 35254 6771
rect 35202 6703 35210 6737
rect 35244 6703 35254 6737
rect 35202 6691 35254 6703
rect 35284 6805 35336 6821
rect 35284 6771 35294 6805
rect 35328 6771 35336 6805
rect 35284 6737 35336 6771
rect 35284 6703 35294 6737
rect 35328 6703 35336 6737
rect 35501 6773 35553 6815
rect 35501 6739 35509 6773
rect 35543 6739 35553 6773
rect 35501 6711 35553 6739
rect 35583 6803 35641 6815
rect 35583 6769 35595 6803
rect 35629 6769 35641 6803
rect 35583 6711 35641 6769
rect 35671 6790 35723 6815
rect 35671 6756 35681 6790
rect 35715 6756 35723 6790
rect 35671 6711 35723 6756
rect 35894 6797 35946 6813
rect 35894 6763 35902 6797
rect 35936 6763 35946 6797
rect 35894 6729 35946 6763
rect 35284 6691 35336 6703
rect 35894 6695 35902 6729
rect 35936 6695 35946 6729
rect 35894 6683 35946 6695
rect 35976 6797 36028 6813
rect 35976 6763 35986 6797
rect 36020 6763 36028 6797
rect 37090 6805 37142 6821
rect 37090 6771 37098 6805
rect 37132 6771 37142 6805
rect 35976 6729 36028 6763
rect 35976 6695 35986 6729
rect 36020 6695 36028 6729
rect 35976 6683 36028 6695
rect 37090 6737 37142 6771
rect 37090 6703 37098 6737
rect 37132 6703 37142 6737
rect 37090 6691 37142 6703
rect 37172 6805 37224 6821
rect 37172 6771 37182 6805
rect 37216 6771 37224 6805
rect 37172 6737 37224 6771
rect 37172 6703 37182 6737
rect 37216 6703 37224 6737
rect 37389 6773 37441 6815
rect 37389 6739 37397 6773
rect 37431 6739 37441 6773
rect 37389 6711 37441 6739
rect 37471 6803 37529 6815
rect 37471 6769 37483 6803
rect 37517 6769 37529 6803
rect 37471 6711 37529 6769
rect 37559 6790 37611 6815
rect 37559 6756 37569 6790
rect 37603 6756 37611 6790
rect 37559 6711 37611 6756
rect 37782 6797 37834 6813
rect 37782 6763 37790 6797
rect 37824 6763 37834 6797
rect 37782 6729 37834 6763
rect 37172 6691 37224 6703
rect 37782 6695 37790 6729
rect 37824 6695 37834 6729
rect 37782 6683 37834 6695
rect 37864 6797 37916 6813
rect 37864 6763 37874 6797
rect 37908 6763 37916 6797
rect 38978 6805 39030 6821
rect 38978 6771 38986 6805
rect 39020 6771 39030 6805
rect 37864 6729 37916 6763
rect 37864 6695 37874 6729
rect 37908 6695 37916 6729
rect 37864 6683 37916 6695
rect 38978 6737 39030 6771
rect 38978 6703 38986 6737
rect 39020 6703 39030 6737
rect 38978 6691 39030 6703
rect 39060 6805 39112 6821
rect 39060 6771 39070 6805
rect 39104 6771 39112 6805
rect 39060 6737 39112 6771
rect 39060 6703 39070 6737
rect 39104 6703 39112 6737
rect 39277 6773 39329 6815
rect 39277 6739 39285 6773
rect 39319 6739 39329 6773
rect 39277 6711 39329 6739
rect 39359 6803 39417 6815
rect 39359 6769 39371 6803
rect 39405 6769 39417 6803
rect 39359 6711 39417 6769
rect 39447 6790 39499 6815
rect 39447 6756 39457 6790
rect 39491 6756 39499 6790
rect 39447 6711 39499 6756
rect 39670 6797 39722 6813
rect 39670 6763 39678 6797
rect 39712 6763 39722 6797
rect 39670 6729 39722 6763
rect 39060 6691 39112 6703
rect 39670 6695 39678 6729
rect 39712 6695 39722 6729
rect 39670 6683 39722 6695
rect 39752 6797 39804 6813
rect 39752 6763 39762 6797
rect 39796 6763 39804 6797
rect 40866 6805 40918 6821
rect 40866 6771 40874 6805
rect 40908 6771 40918 6805
rect 39752 6729 39804 6763
rect 39752 6695 39762 6729
rect 39796 6695 39804 6729
rect 39752 6683 39804 6695
rect 40866 6737 40918 6771
rect 40866 6703 40874 6737
rect 40908 6703 40918 6737
rect 40866 6691 40918 6703
rect 40948 6805 41000 6821
rect 40948 6771 40958 6805
rect 40992 6771 41000 6805
rect 40948 6737 41000 6771
rect 40948 6703 40958 6737
rect 40992 6703 41000 6737
rect 41165 6773 41217 6815
rect 41165 6739 41173 6773
rect 41207 6739 41217 6773
rect 41165 6711 41217 6739
rect 41247 6803 41305 6815
rect 41247 6769 41259 6803
rect 41293 6769 41305 6803
rect 41247 6711 41305 6769
rect 41335 6790 41387 6815
rect 41335 6756 41345 6790
rect 41379 6756 41387 6790
rect 41335 6711 41387 6756
rect 41558 6797 41610 6813
rect 41558 6763 41566 6797
rect 41600 6763 41610 6797
rect 41558 6729 41610 6763
rect 40948 6691 41000 6703
rect 41558 6695 41566 6729
rect 41600 6695 41610 6729
rect 41558 6683 41610 6695
rect 41640 6797 41692 6813
rect 41640 6763 41650 6797
rect 41684 6763 41692 6797
rect 42754 6805 42806 6821
rect 42754 6771 42762 6805
rect 42796 6771 42806 6805
rect 41640 6729 41692 6763
rect 41640 6695 41650 6729
rect 41684 6695 41692 6729
rect 41640 6683 41692 6695
rect 42754 6737 42806 6771
rect 42754 6703 42762 6737
rect 42796 6703 42806 6737
rect 42754 6691 42806 6703
rect 42836 6805 42888 6821
rect 42836 6771 42846 6805
rect 42880 6771 42888 6805
rect 42836 6737 42888 6771
rect 42836 6703 42846 6737
rect 42880 6703 42888 6737
rect 43053 6773 43105 6815
rect 43053 6739 43061 6773
rect 43095 6739 43105 6773
rect 43053 6711 43105 6739
rect 43135 6803 43193 6815
rect 43135 6769 43147 6803
rect 43181 6769 43193 6803
rect 43135 6711 43193 6769
rect 43223 6790 43275 6815
rect 43223 6756 43233 6790
rect 43267 6756 43275 6790
rect 43223 6711 43275 6756
rect 43446 6797 43498 6813
rect 43446 6763 43454 6797
rect 43488 6763 43498 6797
rect 43446 6729 43498 6763
rect 42836 6691 42888 6703
rect 43446 6695 43454 6729
rect 43488 6695 43498 6729
rect 43446 6683 43498 6695
rect 43528 6797 43580 6813
rect 43528 6763 43538 6797
rect 43572 6763 43580 6797
rect 44642 6805 44694 6821
rect 44642 6771 44650 6805
rect 44684 6771 44694 6805
rect 43528 6729 43580 6763
rect 43528 6695 43538 6729
rect 43572 6695 43580 6729
rect 43528 6683 43580 6695
rect 44642 6737 44694 6771
rect 44642 6703 44650 6737
rect 44684 6703 44694 6737
rect 44642 6691 44694 6703
rect 44724 6805 44776 6821
rect 44724 6771 44734 6805
rect 44768 6771 44776 6805
rect 44724 6737 44776 6771
rect 44724 6703 44734 6737
rect 44768 6703 44776 6737
rect 44935 6773 44987 6815
rect 44935 6739 44943 6773
rect 44977 6739 44987 6773
rect 44935 6711 44987 6739
rect 45017 6803 45075 6815
rect 45017 6769 45029 6803
rect 45063 6769 45075 6803
rect 45017 6711 45075 6769
rect 45105 6790 45157 6815
rect 45105 6756 45115 6790
rect 45149 6756 45157 6790
rect 45105 6711 45157 6756
rect 45328 6797 45380 6813
rect 45328 6763 45336 6797
rect 45370 6763 45380 6797
rect 45328 6729 45380 6763
rect 44724 6691 44776 6703
rect 45328 6695 45336 6729
rect 45370 6695 45380 6729
rect 45328 6683 45380 6695
rect 45410 6797 45462 6813
rect 45410 6763 45420 6797
rect 45454 6763 45462 6797
rect 46524 6805 46576 6821
rect 46524 6771 46532 6805
rect 46566 6771 46576 6805
rect 45410 6729 45462 6763
rect 45410 6695 45420 6729
rect 45454 6695 45462 6729
rect 45410 6683 45462 6695
rect 46524 6737 46576 6771
rect 46524 6703 46532 6737
rect 46566 6703 46576 6737
rect 46524 6691 46576 6703
rect 46606 6805 46658 6821
rect 46606 6771 46616 6805
rect 46650 6771 46658 6805
rect 46606 6737 46658 6771
rect 46606 6703 46616 6737
rect 46650 6703 46658 6737
rect 46823 6773 46875 6815
rect 46823 6739 46831 6773
rect 46865 6739 46875 6773
rect 46823 6711 46875 6739
rect 46905 6803 46963 6815
rect 46905 6769 46917 6803
rect 46951 6769 46963 6803
rect 46905 6711 46963 6769
rect 46993 6790 47045 6815
rect 46993 6756 47003 6790
rect 47037 6756 47045 6790
rect 46993 6711 47045 6756
rect 47216 6797 47268 6813
rect 47216 6763 47224 6797
rect 47258 6763 47268 6797
rect 47216 6729 47268 6763
rect 46606 6691 46658 6703
rect 47216 6695 47224 6729
rect 47258 6695 47268 6729
rect 47216 6683 47268 6695
rect 47298 6797 47350 6813
rect 47298 6763 47308 6797
rect 47342 6763 47350 6797
rect 48412 6805 48464 6821
rect 48412 6771 48420 6805
rect 48454 6771 48464 6805
rect 47298 6729 47350 6763
rect 47298 6695 47308 6729
rect 47342 6695 47350 6729
rect 47298 6683 47350 6695
rect 48412 6737 48464 6771
rect 48412 6703 48420 6737
rect 48454 6703 48464 6737
rect 48412 6691 48464 6703
rect 48494 6805 48546 6821
rect 48494 6771 48504 6805
rect 48538 6771 48546 6805
rect 48494 6737 48546 6771
rect 48494 6703 48504 6737
rect 48538 6703 48546 6737
rect 48711 6773 48763 6815
rect 48711 6739 48719 6773
rect 48753 6739 48763 6773
rect 48711 6711 48763 6739
rect 48793 6803 48851 6815
rect 48793 6769 48805 6803
rect 48839 6769 48851 6803
rect 48793 6711 48851 6769
rect 48881 6790 48933 6815
rect 48881 6756 48891 6790
rect 48925 6756 48933 6790
rect 48881 6711 48933 6756
rect 49104 6797 49156 6813
rect 49104 6763 49112 6797
rect 49146 6763 49156 6797
rect 49104 6729 49156 6763
rect 48494 6691 48546 6703
rect 49104 6695 49112 6729
rect 49146 6695 49156 6729
rect 49104 6683 49156 6695
rect 49186 6797 49238 6813
rect 49186 6763 49196 6797
rect 49230 6763 49238 6797
rect 50300 6805 50352 6821
rect 50300 6771 50308 6805
rect 50342 6771 50352 6805
rect 49186 6729 49238 6763
rect 49186 6695 49196 6729
rect 49230 6695 49238 6729
rect 49186 6683 49238 6695
rect 50300 6737 50352 6771
rect 50300 6703 50308 6737
rect 50342 6703 50352 6737
rect 50300 6691 50352 6703
rect 50382 6805 50434 6821
rect 50382 6771 50392 6805
rect 50426 6771 50434 6805
rect 50382 6737 50434 6771
rect 50382 6703 50392 6737
rect 50426 6703 50434 6737
rect 50599 6773 50651 6815
rect 50599 6739 50607 6773
rect 50641 6739 50651 6773
rect 50599 6711 50651 6739
rect 50681 6803 50739 6815
rect 50681 6769 50693 6803
rect 50727 6769 50739 6803
rect 50681 6711 50739 6769
rect 50769 6790 50821 6815
rect 50769 6756 50779 6790
rect 50813 6756 50821 6790
rect 50769 6711 50821 6756
rect 50992 6797 51044 6813
rect 50992 6763 51000 6797
rect 51034 6763 51044 6797
rect 50992 6729 51044 6763
rect 50382 6691 50434 6703
rect 50992 6695 51000 6729
rect 51034 6695 51044 6729
rect 50992 6683 51044 6695
rect 51074 6797 51126 6813
rect 51074 6763 51084 6797
rect 51118 6763 51126 6797
rect 52188 6805 52240 6821
rect 52188 6771 52196 6805
rect 52230 6771 52240 6805
rect 51074 6729 51126 6763
rect 51074 6695 51084 6729
rect 51118 6695 51126 6729
rect 51074 6683 51126 6695
rect 52188 6737 52240 6771
rect 52188 6703 52196 6737
rect 52230 6703 52240 6737
rect 52188 6691 52240 6703
rect 52270 6805 52322 6821
rect 52270 6771 52280 6805
rect 52314 6771 52322 6805
rect 52270 6737 52322 6771
rect 52270 6703 52280 6737
rect 52314 6703 52322 6737
rect 52487 6773 52539 6815
rect 52487 6739 52495 6773
rect 52529 6739 52539 6773
rect 52487 6711 52539 6739
rect 52569 6803 52627 6815
rect 52569 6769 52581 6803
rect 52615 6769 52627 6803
rect 52569 6711 52627 6769
rect 52657 6790 52709 6815
rect 52657 6756 52667 6790
rect 52701 6756 52709 6790
rect 52657 6711 52709 6756
rect 52880 6797 52932 6813
rect 52880 6763 52888 6797
rect 52922 6763 52932 6797
rect 52880 6729 52932 6763
rect 52270 6691 52322 6703
rect 52880 6695 52888 6729
rect 52922 6695 52932 6729
rect 52880 6683 52932 6695
rect 52962 6797 53014 6813
rect 52962 6763 52972 6797
rect 53006 6763 53014 6797
rect 54076 6805 54128 6821
rect 54076 6771 54084 6805
rect 54118 6771 54128 6805
rect 52962 6729 53014 6763
rect 52962 6695 52972 6729
rect 53006 6695 53014 6729
rect 52962 6683 53014 6695
rect 54076 6737 54128 6771
rect 54076 6703 54084 6737
rect 54118 6703 54128 6737
rect 54076 6691 54128 6703
rect 54158 6805 54210 6821
rect 54158 6771 54168 6805
rect 54202 6771 54210 6805
rect 54158 6737 54210 6771
rect 54158 6703 54168 6737
rect 54202 6703 54210 6737
rect 54375 6773 54427 6815
rect 54375 6739 54383 6773
rect 54417 6739 54427 6773
rect 54375 6711 54427 6739
rect 54457 6803 54515 6815
rect 54457 6769 54469 6803
rect 54503 6769 54515 6803
rect 54457 6711 54515 6769
rect 54545 6790 54597 6815
rect 54545 6756 54555 6790
rect 54589 6756 54597 6790
rect 54545 6711 54597 6756
rect 54768 6797 54820 6813
rect 54768 6763 54776 6797
rect 54810 6763 54820 6797
rect 54768 6729 54820 6763
rect 54158 6691 54210 6703
rect 54768 6695 54776 6729
rect 54810 6695 54820 6729
rect 54768 6683 54820 6695
rect 54850 6797 54902 6813
rect 54850 6763 54860 6797
rect 54894 6763 54902 6797
rect 55964 6805 56016 6821
rect 55964 6771 55972 6805
rect 56006 6771 56016 6805
rect 54850 6729 54902 6763
rect 54850 6695 54860 6729
rect 54894 6695 54902 6729
rect 54850 6683 54902 6695
rect 55964 6737 56016 6771
rect 55964 6703 55972 6737
rect 56006 6703 56016 6737
rect 55964 6691 56016 6703
rect 56046 6805 56098 6821
rect 56046 6771 56056 6805
rect 56090 6771 56098 6805
rect 56046 6737 56098 6771
rect 56046 6703 56056 6737
rect 56090 6703 56098 6737
rect 56263 6773 56315 6815
rect 56263 6739 56271 6773
rect 56305 6739 56315 6773
rect 56263 6711 56315 6739
rect 56345 6803 56403 6815
rect 56345 6769 56357 6803
rect 56391 6769 56403 6803
rect 56345 6711 56403 6769
rect 56433 6790 56485 6815
rect 56433 6756 56443 6790
rect 56477 6756 56485 6790
rect 56433 6711 56485 6756
rect 56656 6797 56708 6813
rect 56656 6763 56664 6797
rect 56698 6763 56708 6797
rect 56656 6729 56708 6763
rect 56046 6691 56098 6703
rect 56656 6695 56664 6729
rect 56698 6695 56708 6729
rect 56656 6683 56708 6695
rect 56738 6797 56790 6813
rect 56738 6763 56748 6797
rect 56782 6763 56790 6797
rect 57852 6805 57904 6821
rect 57852 6771 57860 6805
rect 57894 6771 57904 6805
rect 56738 6729 56790 6763
rect 56738 6695 56748 6729
rect 56782 6695 56790 6729
rect 56738 6683 56790 6695
rect 57852 6737 57904 6771
rect 57852 6703 57860 6737
rect 57894 6703 57904 6737
rect 57852 6691 57904 6703
rect 57934 6805 57986 6821
rect 57934 6771 57944 6805
rect 57978 6771 57986 6805
rect 57934 6737 57986 6771
rect 57934 6703 57944 6737
rect 57978 6703 57986 6737
rect 58151 6773 58203 6815
rect 58151 6739 58159 6773
rect 58193 6739 58203 6773
rect 58151 6711 58203 6739
rect 58233 6803 58291 6815
rect 58233 6769 58245 6803
rect 58279 6769 58291 6803
rect 58233 6711 58291 6769
rect 58321 6790 58373 6815
rect 58321 6756 58331 6790
rect 58365 6756 58373 6790
rect 58321 6711 58373 6756
rect 58544 6797 58596 6813
rect 58544 6763 58552 6797
rect 58586 6763 58596 6797
rect 58544 6729 58596 6763
rect 57934 6691 57986 6703
rect 58544 6695 58552 6729
rect 58586 6695 58596 6729
rect 58544 6683 58596 6695
rect 58626 6797 58678 6813
rect 58626 6763 58636 6797
rect 58670 6763 58678 6797
rect 59740 6805 59792 6821
rect 59740 6771 59748 6805
rect 59782 6771 59792 6805
rect 58626 6729 58678 6763
rect 58626 6695 58636 6729
rect 58670 6695 58678 6729
rect 58626 6683 58678 6695
rect 59740 6737 59792 6771
rect 59740 6703 59748 6737
rect 59782 6703 59792 6737
rect 59740 6691 59792 6703
rect 59822 6805 59874 6821
rect 59822 6771 59832 6805
rect 59866 6771 59874 6805
rect 59822 6737 59874 6771
rect 59822 6703 59832 6737
rect 59866 6703 59874 6737
rect 59822 6691 59874 6703
rect 606 5998 668 6012
rect 606 5964 618 5998
rect 652 5964 668 5998
rect 606 5930 668 5964
rect 606 5896 618 5930
rect 652 5896 668 5930
rect 606 5882 668 5896
rect 698 5998 764 6012
rect 698 5964 714 5998
rect 748 5964 764 5998
rect 698 5930 764 5964
rect 698 5896 714 5930
rect 748 5896 764 5930
rect 698 5882 764 5896
rect 794 5998 856 6012
rect 794 5964 810 5998
rect 844 5964 856 5998
rect 794 5930 856 5964
rect 794 5896 810 5930
rect 844 5896 856 5930
rect 794 5882 856 5896
rect 2494 5998 2556 6012
rect 2494 5964 2506 5998
rect 2540 5964 2556 5998
rect 2494 5930 2556 5964
rect 2494 5896 2506 5930
rect 2540 5896 2556 5930
rect 2494 5882 2556 5896
rect 2586 5998 2652 6012
rect 2586 5964 2602 5998
rect 2636 5964 2652 5998
rect 2586 5930 2652 5964
rect 2586 5896 2602 5930
rect 2636 5896 2652 5930
rect 2586 5882 2652 5896
rect 2682 5998 2744 6012
rect 2682 5964 2698 5998
rect 2732 5964 2744 5998
rect 2682 5930 2744 5964
rect 2682 5896 2698 5930
rect 2732 5896 2744 5930
rect 2682 5882 2744 5896
rect 4382 5998 4444 6012
rect 4382 5964 4394 5998
rect 4428 5964 4444 5998
rect 4382 5930 4444 5964
rect 4382 5896 4394 5930
rect 4428 5896 4444 5930
rect 4382 5882 4444 5896
rect 4474 5998 4540 6012
rect 4474 5964 4490 5998
rect 4524 5964 4540 5998
rect 4474 5930 4540 5964
rect 4474 5896 4490 5930
rect 4524 5896 4540 5930
rect 4474 5882 4540 5896
rect 4570 5998 4632 6012
rect 4570 5964 4586 5998
rect 4620 5964 4632 5998
rect 4570 5930 4632 5964
rect 4570 5896 4586 5930
rect 4620 5896 4632 5930
rect 4570 5882 4632 5896
rect 6270 5998 6332 6012
rect 6270 5964 6282 5998
rect 6316 5964 6332 5998
rect 6270 5930 6332 5964
rect 6270 5896 6282 5930
rect 6316 5896 6332 5930
rect 6270 5882 6332 5896
rect 6362 5998 6428 6012
rect 6362 5964 6378 5998
rect 6412 5964 6428 5998
rect 6362 5930 6428 5964
rect 6362 5896 6378 5930
rect 6412 5896 6428 5930
rect 6362 5882 6428 5896
rect 6458 5998 6520 6012
rect 6458 5964 6474 5998
rect 6508 5964 6520 5998
rect 6458 5930 6520 5964
rect 6458 5896 6474 5930
rect 6508 5896 6520 5930
rect 6458 5882 6520 5896
rect 8158 5998 8220 6012
rect 8158 5964 8170 5998
rect 8204 5964 8220 5998
rect 8158 5930 8220 5964
rect 8158 5896 8170 5930
rect 8204 5896 8220 5930
rect 8158 5882 8220 5896
rect 8250 5998 8316 6012
rect 8250 5964 8266 5998
rect 8300 5964 8316 5998
rect 8250 5930 8316 5964
rect 8250 5896 8266 5930
rect 8300 5896 8316 5930
rect 8250 5882 8316 5896
rect 8346 5998 8408 6012
rect 8346 5964 8362 5998
rect 8396 5964 8408 5998
rect 8346 5930 8408 5964
rect 8346 5896 8362 5930
rect 8396 5896 8408 5930
rect 8346 5882 8408 5896
rect 10046 5998 10108 6012
rect 10046 5964 10058 5998
rect 10092 5964 10108 5998
rect 10046 5930 10108 5964
rect 10046 5896 10058 5930
rect 10092 5896 10108 5930
rect 10046 5882 10108 5896
rect 10138 5998 10204 6012
rect 10138 5964 10154 5998
rect 10188 5964 10204 5998
rect 10138 5930 10204 5964
rect 10138 5896 10154 5930
rect 10188 5896 10204 5930
rect 10138 5882 10204 5896
rect 10234 5998 10296 6012
rect 10234 5964 10250 5998
rect 10284 5964 10296 5998
rect 10234 5930 10296 5964
rect 10234 5896 10250 5930
rect 10284 5896 10296 5930
rect 10234 5882 10296 5896
rect 11934 5998 11996 6012
rect 11934 5964 11946 5998
rect 11980 5964 11996 5998
rect 11934 5930 11996 5964
rect 11934 5896 11946 5930
rect 11980 5896 11996 5930
rect 11934 5882 11996 5896
rect 12026 5998 12092 6012
rect 12026 5964 12042 5998
rect 12076 5964 12092 5998
rect 12026 5930 12092 5964
rect 12026 5896 12042 5930
rect 12076 5896 12092 5930
rect 12026 5882 12092 5896
rect 12122 5998 12184 6012
rect 12122 5964 12138 5998
rect 12172 5964 12184 5998
rect 12122 5930 12184 5964
rect 12122 5896 12138 5930
rect 12172 5896 12184 5930
rect 12122 5882 12184 5896
rect 13822 5998 13884 6012
rect 13822 5964 13834 5998
rect 13868 5964 13884 5998
rect 13822 5930 13884 5964
rect 13822 5896 13834 5930
rect 13868 5896 13884 5930
rect 13822 5882 13884 5896
rect 13914 5998 13980 6012
rect 13914 5964 13930 5998
rect 13964 5964 13980 5998
rect 13914 5930 13980 5964
rect 13914 5896 13930 5930
rect 13964 5896 13980 5930
rect 13914 5882 13980 5896
rect 14010 5998 14072 6012
rect 14010 5964 14026 5998
rect 14060 5964 14072 5998
rect 14010 5930 14072 5964
rect 14010 5896 14026 5930
rect 14060 5896 14072 5930
rect 14010 5882 14072 5896
rect 15704 5998 15766 6012
rect 15704 5964 15716 5998
rect 15750 5964 15766 5998
rect 15704 5930 15766 5964
rect 15704 5896 15716 5930
rect 15750 5896 15766 5930
rect 15704 5882 15766 5896
rect 15796 5998 15862 6012
rect 15796 5964 15812 5998
rect 15846 5964 15862 5998
rect 15796 5930 15862 5964
rect 15796 5896 15812 5930
rect 15846 5896 15862 5930
rect 15796 5882 15862 5896
rect 15892 5998 15954 6012
rect 15892 5964 15908 5998
rect 15942 5964 15954 5998
rect 15892 5930 15954 5964
rect 15892 5896 15908 5930
rect 15942 5896 15954 5930
rect 15892 5882 15954 5896
rect 17592 5998 17654 6012
rect 17592 5964 17604 5998
rect 17638 5964 17654 5998
rect 17592 5930 17654 5964
rect 17592 5896 17604 5930
rect 17638 5896 17654 5930
rect 17592 5882 17654 5896
rect 17684 5998 17750 6012
rect 17684 5964 17700 5998
rect 17734 5964 17750 5998
rect 17684 5930 17750 5964
rect 17684 5896 17700 5930
rect 17734 5896 17750 5930
rect 17684 5882 17750 5896
rect 17780 5998 17842 6012
rect 17780 5964 17796 5998
rect 17830 5964 17842 5998
rect 17780 5930 17842 5964
rect 17780 5896 17796 5930
rect 17830 5896 17842 5930
rect 17780 5882 17842 5896
rect 19480 5998 19542 6012
rect 19480 5964 19492 5998
rect 19526 5964 19542 5998
rect 19480 5930 19542 5964
rect 19480 5896 19492 5930
rect 19526 5896 19542 5930
rect 19480 5882 19542 5896
rect 19572 5998 19638 6012
rect 19572 5964 19588 5998
rect 19622 5964 19638 5998
rect 19572 5930 19638 5964
rect 19572 5896 19588 5930
rect 19622 5896 19638 5930
rect 19572 5882 19638 5896
rect 19668 5998 19730 6012
rect 19668 5964 19684 5998
rect 19718 5964 19730 5998
rect 19668 5930 19730 5964
rect 19668 5896 19684 5930
rect 19718 5896 19730 5930
rect 19668 5882 19730 5896
rect 21368 5998 21430 6012
rect 21368 5964 21380 5998
rect 21414 5964 21430 5998
rect 21368 5930 21430 5964
rect 21368 5896 21380 5930
rect 21414 5896 21430 5930
rect 21368 5882 21430 5896
rect 21460 5998 21526 6012
rect 21460 5964 21476 5998
rect 21510 5964 21526 5998
rect 21460 5930 21526 5964
rect 21460 5896 21476 5930
rect 21510 5896 21526 5930
rect 21460 5882 21526 5896
rect 21556 5998 21618 6012
rect 21556 5964 21572 5998
rect 21606 5964 21618 5998
rect 21556 5930 21618 5964
rect 21556 5896 21572 5930
rect 21606 5896 21618 5930
rect 21556 5882 21618 5896
rect 23256 5998 23318 6012
rect 23256 5964 23268 5998
rect 23302 5964 23318 5998
rect 23256 5930 23318 5964
rect 23256 5896 23268 5930
rect 23302 5896 23318 5930
rect 23256 5882 23318 5896
rect 23348 5998 23414 6012
rect 23348 5964 23364 5998
rect 23398 5964 23414 5998
rect 23348 5930 23414 5964
rect 23348 5896 23364 5930
rect 23398 5896 23414 5930
rect 23348 5882 23414 5896
rect 23444 5998 23506 6012
rect 23444 5964 23460 5998
rect 23494 5964 23506 5998
rect 23444 5930 23506 5964
rect 23444 5896 23460 5930
rect 23494 5896 23506 5930
rect 23444 5882 23506 5896
rect 25144 5998 25206 6012
rect 25144 5964 25156 5998
rect 25190 5964 25206 5998
rect 25144 5930 25206 5964
rect 25144 5896 25156 5930
rect 25190 5896 25206 5930
rect 25144 5882 25206 5896
rect 25236 5998 25302 6012
rect 25236 5964 25252 5998
rect 25286 5964 25302 5998
rect 25236 5930 25302 5964
rect 25236 5896 25252 5930
rect 25286 5896 25302 5930
rect 25236 5882 25302 5896
rect 25332 5998 25394 6012
rect 25332 5964 25348 5998
rect 25382 5964 25394 5998
rect 25332 5930 25394 5964
rect 25332 5896 25348 5930
rect 25382 5896 25394 5930
rect 25332 5882 25394 5896
rect 27032 5998 27094 6012
rect 27032 5964 27044 5998
rect 27078 5964 27094 5998
rect 27032 5930 27094 5964
rect 27032 5896 27044 5930
rect 27078 5896 27094 5930
rect 27032 5882 27094 5896
rect 27124 5998 27190 6012
rect 27124 5964 27140 5998
rect 27174 5964 27190 5998
rect 27124 5930 27190 5964
rect 27124 5896 27140 5930
rect 27174 5896 27190 5930
rect 27124 5882 27190 5896
rect 27220 5998 27282 6012
rect 27220 5964 27236 5998
rect 27270 5964 27282 5998
rect 27220 5930 27282 5964
rect 27220 5896 27236 5930
rect 27270 5896 27282 5930
rect 27220 5882 27282 5896
rect 28920 5998 28982 6012
rect 28920 5964 28932 5998
rect 28966 5964 28982 5998
rect 28920 5930 28982 5964
rect 28920 5896 28932 5930
rect 28966 5896 28982 5930
rect 28920 5882 28982 5896
rect 29012 5998 29078 6012
rect 29012 5964 29028 5998
rect 29062 5964 29078 5998
rect 29012 5930 29078 5964
rect 29012 5896 29028 5930
rect 29062 5896 29078 5930
rect 29012 5882 29078 5896
rect 29108 5998 29170 6012
rect 29108 5964 29124 5998
rect 29158 5964 29170 5998
rect 29108 5930 29170 5964
rect 29108 5896 29124 5930
rect 29158 5896 29170 5930
rect 29108 5882 29170 5896
rect 30808 5998 30870 6012
rect 30808 5964 30820 5998
rect 30854 5964 30870 5998
rect 30808 5930 30870 5964
rect 30808 5896 30820 5930
rect 30854 5896 30870 5930
rect 30808 5882 30870 5896
rect 30900 5998 30966 6012
rect 30900 5964 30916 5998
rect 30950 5964 30966 5998
rect 30900 5930 30966 5964
rect 30900 5896 30916 5930
rect 30950 5896 30966 5930
rect 30900 5882 30966 5896
rect 30996 5998 31058 6012
rect 30996 5964 31012 5998
rect 31046 5964 31058 5998
rect 30996 5930 31058 5964
rect 30996 5896 31012 5930
rect 31046 5896 31058 5930
rect 30996 5882 31058 5896
rect 32696 5998 32758 6012
rect 32696 5964 32708 5998
rect 32742 5964 32758 5998
rect 32696 5930 32758 5964
rect 32696 5896 32708 5930
rect 32742 5896 32758 5930
rect 32696 5882 32758 5896
rect 32788 5998 32854 6012
rect 32788 5964 32804 5998
rect 32838 5964 32854 5998
rect 32788 5930 32854 5964
rect 32788 5896 32804 5930
rect 32838 5896 32854 5930
rect 32788 5882 32854 5896
rect 32884 5998 32946 6012
rect 32884 5964 32900 5998
rect 32934 5964 32946 5998
rect 32884 5930 32946 5964
rect 32884 5896 32900 5930
rect 32934 5896 32946 5930
rect 32884 5882 32946 5896
rect 34584 5998 34646 6012
rect 34584 5964 34596 5998
rect 34630 5964 34646 5998
rect 34584 5930 34646 5964
rect 34584 5896 34596 5930
rect 34630 5896 34646 5930
rect 34584 5882 34646 5896
rect 34676 5998 34742 6012
rect 34676 5964 34692 5998
rect 34726 5964 34742 5998
rect 34676 5930 34742 5964
rect 34676 5896 34692 5930
rect 34726 5896 34742 5930
rect 34676 5882 34742 5896
rect 34772 5998 34834 6012
rect 34772 5964 34788 5998
rect 34822 5964 34834 5998
rect 34772 5930 34834 5964
rect 34772 5896 34788 5930
rect 34822 5896 34834 5930
rect 34772 5882 34834 5896
rect 36472 5998 36534 6012
rect 36472 5964 36484 5998
rect 36518 5964 36534 5998
rect 36472 5930 36534 5964
rect 36472 5896 36484 5930
rect 36518 5896 36534 5930
rect 36472 5882 36534 5896
rect 36564 5998 36630 6012
rect 36564 5964 36580 5998
rect 36614 5964 36630 5998
rect 36564 5930 36630 5964
rect 36564 5896 36580 5930
rect 36614 5896 36630 5930
rect 36564 5882 36630 5896
rect 36660 5998 36722 6012
rect 36660 5964 36676 5998
rect 36710 5964 36722 5998
rect 36660 5930 36722 5964
rect 36660 5896 36676 5930
rect 36710 5896 36722 5930
rect 36660 5882 36722 5896
rect 38360 5998 38422 6012
rect 38360 5964 38372 5998
rect 38406 5964 38422 5998
rect 38360 5930 38422 5964
rect 38360 5896 38372 5930
rect 38406 5896 38422 5930
rect 38360 5882 38422 5896
rect 38452 5998 38518 6012
rect 38452 5964 38468 5998
rect 38502 5964 38518 5998
rect 38452 5930 38518 5964
rect 38452 5896 38468 5930
rect 38502 5896 38518 5930
rect 38452 5882 38518 5896
rect 38548 5998 38610 6012
rect 38548 5964 38564 5998
rect 38598 5964 38610 5998
rect 38548 5930 38610 5964
rect 38548 5896 38564 5930
rect 38598 5896 38610 5930
rect 38548 5882 38610 5896
rect 40248 5998 40310 6012
rect 40248 5964 40260 5998
rect 40294 5964 40310 5998
rect 40248 5930 40310 5964
rect 40248 5896 40260 5930
rect 40294 5896 40310 5930
rect 40248 5882 40310 5896
rect 40340 5998 40406 6012
rect 40340 5964 40356 5998
rect 40390 5964 40406 5998
rect 40340 5930 40406 5964
rect 40340 5896 40356 5930
rect 40390 5896 40406 5930
rect 40340 5882 40406 5896
rect 40436 5998 40498 6012
rect 40436 5964 40452 5998
rect 40486 5964 40498 5998
rect 40436 5930 40498 5964
rect 40436 5896 40452 5930
rect 40486 5896 40498 5930
rect 40436 5882 40498 5896
rect 42136 5998 42198 6012
rect 42136 5964 42148 5998
rect 42182 5964 42198 5998
rect 42136 5930 42198 5964
rect 42136 5896 42148 5930
rect 42182 5896 42198 5930
rect 42136 5882 42198 5896
rect 42228 5998 42294 6012
rect 42228 5964 42244 5998
rect 42278 5964 42294 5998
rect 42228 5930 42294 5964
rect 42228 5896 42244 5930
rect 42278 5896 42294 5930
rect 42228 5882 42294 5896
rect 42324 5998 42386 6012
rect 42324 5964 42340 5998
rect 42374 5964 42386 5998
rect 42324 5930 42386 5964
rect 42324 5896 42340 5930
rect 42374 5896 42386 5930
rect 42324 5882 42386 5896
rect 44024 5998 44086 6012
rect 44024 5964 44036 5998
rect 44070 5964 44086 5998
rect 44024 5930 44086 5964
rect 44024 5896 44036 5930
rect 44070 5896 44086 5930
rect 44024 5882 44086 5896
rect 44116 5998 44182 6012
rect 44116 5964 44132 5998
rect 44166 5964 44182 5998
rect 44116 5930 44182 5964
rect 44116 5896 44132 5930
rect 44166 5896 44182 5930
rect 44116 5882 44182 5896
rect 44212 5998 44274 6012
rect 44212 5964 44228 5998
rect 44262 5964 44274 5998
rect 44212 5930 44274 5964
rect 44212 5896 44228 5930
rect 44262 5896 44274 5930
rect 44212 5882 44274 5896
rect 45906 5998 45968 6012
rect 45906 5964 45918 5998
rect 45952 5964 45968 5998
rect 45906 5930 45968 5964
rect 45906 5896 45918 5930
rect 45952 5896 45968 5930
rect 45906 5882 45968 5896
rect 45998 5998 46064 6012
rect 45998 5964 46014 5998
rect 46048 5964 46064 5998
rect 45998 5930 46064 5964
rect 45998 5896 46014 5930
rect 46048 5896 46064 5930
rect 45998 5882 46064 5896
rect 46094 5998 46156 6012
rect 46094 5964 46110 5998
rect 46144 5964 46156 5998
rect 46094 5930 46156 5964
rect 46094 5896 46110 5930
rect 46144 5896 46156 5930
rect 46094 5882 46156 5896
rect 47794 5998 47856 6012
rect 47794 5964 47806 5998
rect 47840 5964 47856 5998
rect 47794 5930 47856 5964
rect 47794 5896 47806 5930
rect 47840 5896 47856 5930
rect 47794 5882 47856 5896
rect 47886 5998 47952 6012
rect 47886 5964 47902 5998
rect 47936 5964 47952 5998
rect 47886 5930 47952 5964
rect 47886 5896 47902 5930
rect 47936 5896 47952 5930
rect 47886 5882 47952 5896
rect 47982 5998 48044 6012
rect 47982 5964 47998 5998
rect 48032 5964 48044 5998
rect 47982 5930 48044 5964
rect 47982 5896 47998 5930
rect 48032 5896 48044 5930
rect 47982 5882 48044 5896
rect 49682 5998 49744 6012
rect 49682 5964 49694 5998
rect 49728 5964 49744 5998
rect 49682 5930 49744 5964
rect 49682 5896 49694 5930
rect 49728 5896 49744 5930
rect 49682 5882 49744 5896
rect 49774 5998 49840 6012
rect 49774 5964 49790 5998
rect 49824 5964 49840 5998
rect 49774 5930 49840 5964
rect 49774 5896 49790 5930
rect 49824 5896 49840 5930
rect 49774 5882 49840 5896
rect 49870 5998 49932 6012
rect 49870 5964 49886 5998
rect 49920 5964 49932 5998
rect 49870 5930 49932 5964
rect 49870 5896 49886 5930
rect 49920 5896 49932 5930
rect 49870 5882 49932 5896
rect 51570 5998 51632 6012
rect 51570 5964 51582 5998
rect 51616 5964 51632 5998
rect 51570 5930 51632 5964
rect 51570 5896 51582 5930
rect 51616 5896 51632 5930
rect 51570 5882 51632 5896
rect 51662 5998 51728 6012
rect 51662 5964 51678 5998
rect 51712 5964 51728 5998
rect 51662 5930 51728 5964
rect 51662 5896 51678 5930
rect 51712 5896 51728 5930
rect 51662 5882 51728 5896
rect 51758 5998 51820 6012
rect 51758 5964 51774 5998
rect 51808 5964 51820 5998
rect 51758 5930 51820 5964
rect 51758 5896 51774 5930
rect 51808 5896 51820 5930
rect 51758 5882 51820 5896
rect 53458 5998 53520 6012
rect 53458 5964 53470 5998
rect 53504 5964 53520 5998
rect 53458 5930 53520 5964
rect 53458 5896 53470 5930
rect 53504 5896 53520 5930
rect 53458 5882 53520 5896
rect 53550 5998 53616 6012
rect 53550 5964 53566 5998
rect 53600 5964 53616 5998
rect 53550 5930 53616 5964
rect 53550 5896 53566 5930
rect 53600 5896 53616 5930
rect 53550 5882 53616 5896
rect 53646 5998 53708 6012
rect 53646 5964 53662 5998
rect 53696 5964 53708 5998
rect 53646 5930 53708 5964
rect 53646 5896 53662 5930
rect 53696 5896 53708 5930
rect 53646 5882 53708 5896
rect 55346 5998 55408 6012
rect 55346 5964 55358 5998
rect 55392 5964 55408 5998
rect 55346 5930 55408 5964
rect 55346 5896 55358 5930
rect 55392 5896 55408 5930
rect 55346 5882 55408 5896
rect 55438 5998 55504 6012
rect 55438 5964 55454 5998
rect 55488 5964 55504 5998
rect 55438 5930 55504 5964
rect 55438 5896 55454 5930
rect 55488 5896 55504 5930
rect 55438 5882 55504 5896
rect 55534 5998 55596 6012
rect 55534 5964 55550 5998
rect 55584 5964 55596 5998
rect 55534 5930 55596 5964
rect 55534 5896 55550 5930
rect 55584 5896 55596 5930
rect 55534 5882 55596 5896
rect 57234 5998 57296 6012
rect 57234 5964 57246 5998
rect 57280 5964 57296 5998
rect 57234 5930 57296 5964
rect 57234 5896 57246 5930
rect 57280 5896 57296 5930
rect 57234 5882 57296 5896
rect 57326 5998 57392 6012
rect 57326 5964 57342 5998
rect 57376 5964 57392 5998
rect 57326 5930 57392 5964
rect 57326 5896 57342 5930
rect 57376 5896 57392 5930
rect 57326 5882 57392 5896
rect 57422 5998 57484 6012
rect 57422 5964 57438 5998
rect 57472 5964 57484 5998
rect 57422 5930 57484 5964
rect 57422 5896 57438 5930
rect 57472 5896 57484 5930
rect 57422 5882 57484 5896
rect 59122 5998 59184 6012
rect 59122 5964 59134 5998
rect 59168 5964 59184 5998
rect 59122 5930 59184 5964
rect 59122 5896 59134 5930
rect 59168 5896 59184 5930
rect 59122 5882 59184 5896
rect 59214 5998 59280 6012
rect 59214 5964 59230 5998
rect 59264 5964 59280 5998
rect 59214 5930 59280 5964
rect 59214 5896 59230 5930
rect 59264 5896 59280 5930
rect 59214 5882 59280 5896
rect 59310 5998 59372 6012
rect 59310 5964 59326 5998
rect 59360 5964 59372 5998
rect 59310 5930 59372 5964
rect 59310 5896 59326 5930
rect 59360 5896 59372 5930
rect 59310 5882 59372 5896
rect 189 5753 241 5767
rect 189 5719 197 5753
rect 231 5719 241 5753
rect 189 5685 241 5719
rect 189 5651 197 5685
rect 231 5651 241 5685
rect 189 5637 241 5651
rect 271 5753 325 5767
rect 271 5719 281 5753
rect 315 5719 325 5753
rect 271 5685 325 5719
rect 271 5651 281 5685
rect 315 5651 325 5685
rect 271 5637 325 5651
rect 355 5753 407 5767
rect 355 5719 365 5753
rect 399 5719 407 5753
rect 355 5685 407 5719
rect 1003 5753 1055 5767
rect 1003 5719 1011 5753
rect 1045 5719 1055 5753
rect 355 5651 365 5685
rect 399 5651 407 5685
rect 1003 5685 1055 5719
rect 355 5637 407 5651
rect 1003 5651 1011 5685
rect 1045 5651 1055 5685
rect 1003 5637 1055 5651
rect 1085 5753 1139 5767
rect 1085 5719 1095 5753
rect 1129 5719 1139 5753
rect 1085 5685 1139 5719
rect 1085 5651 1095 5685
rect 1129 5651 1139 5685
rect 1085 5637 1139 5651
rect 1169 5753 1221 5767
rect 1169 5719 1179 5753
rect 1213 5719 1221 5753
rect 1169 5685 1221 5719
rect 1169 5651 1179 5685
rect 1213 5651 1221 5685
rect 1169 5637 1221 5651
rect 2077 5753 2129 5767
rect 2077 5719 2085 5753
rect 2119 5719 2129 5753
rect 2077 5685 2129 5719
rect 2077 5651 2085 5685
rect 2119 5651 2129 5685
rect 2077 5637 2129 5651
rect 2159 5753 2213 5767
rect 2159 5719 2169 5753
rect 2203 5719 2213 5753
rect 2159 5685 2213 5719
rect 2159 5651 2169 5685
rect 2203 5651 2213 5685
rect 2159 5637 2213 5651
rect 2243 5753 2295 5767
rect 2243 5719 2253 5753
rect 2287 5719 2295 5753
rect 2243 5685 2295 5719
rect 2891 5753 2943 5767
rect 2891 5719 2899 5753
rect 2933 5719 2943 5753
rect 2243 5651 2253 5685
rect 2287 5651 2295 5685
rect 2891 5685 2943 5719
rect 2243 5637 2295 5651
rect 2891 5651 2899 5685
rect 2933 5651 2943 5685
rect 2891 5637 2943 5651
rect 2973 5753 3027 5767
rect 2973 5719 2983 5753
rect 3017 5719 3027 5753
rect 2973 5685 3027 5719
rect 2973 5651 2983 5685
rect 3017 5651 3027 5685
rect 2973 5637 3027 5651
rect 3057 5753 3109 5767
rect 3057 5719 3067 5753
rect 3101 5719 3109 5753
rect 3057 5685 3109 5719
rect 3057 5651 3067 5685
rect 3101 5651 3109 5685
rect 3057 5637 3109 5651
rect 3965 5753 4017 5767
rect 3965 5719 3973 5753
rect 4007 5719 4017 5753
rect 3965 5685 4017 5719
rect 3965 5651 3973 5685
rect 4007 5651 4017 5685
rect 3965 5637 4017 5651
rect 4047 5753 4101 5767
rect 4047 5719 4057 5753
rect 4091 5719 4101 5753
rect 4047 5685 4101 5719
rect 4047 5651 4057 5685
rect 4091 5651 4101 5685
rect 4047 5637 4101 5651
rect 4131 5753 4183 5767
rect 4131 5719 4141 5753
rect 4175 5719 4183 5753
rect 4131 5685 4183 5719
rect 4779 5753 4831 5767
rect 4779 5719 4787 5753
rect 4821 5719 4831 5753
rect 4131 5651 4141 5685
rect 4175 5651 4183 5685
rect 4779 5685 4831 5719
rect 4131 5637 4183 5651
rect 4779 5651 4787 5685
rect 4821 5651 4831 5685
rect 4779 5637 4831 5651
rect 4861 5753 4915 5767
rect 4861 5719 4871 5753
rect 4905 5719 4915 5753
rect 4861 5685 4915 5719
rect 4861 5651 4871 5685
rect 4905 5651 4915 5685
rect 4861 5637 4915 5651
rect 4945 5753 4997 5767
rect 4945 5719 4955 5753
rect 4989 5719 4997 5753
rect 4945 5685 4997 5719
rect 4945 5651 4955 5685
rect 4989 5651 4997 5685
rect 4945 5637 4997 5651
rect 5853 5753 5905 5767
rect 5853 5719 5861 5753
rect 5895 5719 5905 5753
rect 5853 5685 5905 5719
rect 5853 5651 5861 5685
rect 5895 5651 5905 5685
rect 5853 5637 5905 5651
rect 5935 5753 5989 5767
rect 5935 5719 5945 5753
rect 5979 5719 5989 5753
rect 5935 5685 5989 5719
rect 5935 5651 5945 5685
rect 5979 5651 5989 5685
rect 5935 5637 5989 5651
rect 6019 5753 6071 5767
rect 6019 5719 6029 5753
rect 6063 5719 6071 5753
rect 6019 5685 6071 5719
rect 6667 5753 6719 5767
rect 6667 5719 6675 5753
rect 6709 5719 6719 5753
rect 6019 5651 6029 5685
rect 6063 5651 6071 5685
rect 6667 5685 6719 5719
rect 6019 5637 6071 5651
rect 6667 5651 6675 5685
rect 6709 5651 6719 5685
rect 6667 5637 6719 5651
rect 6749 5753 6803 5767
rect 6749 5719 6759 5753
rect 6793 5719 6803 5753
rect 6749 5685 6803 5719
rect 6749 5651 6759 5685
rect 6793 5651 6803 5685
rect 6749 5637 6803 5651
rect 6833 5753 6885 5767
rect 6833 5719 6843 5753
rect 6877 5719 6885 5753
rect 6833 5685 6885 5719
rect 6833 5651 6843 5685
rect 6877 5651 6885 5685
rect 6833 5637 6885 5651
rect 7741 5753 7793 5767
rect 7741 5719 7749 5753
rect 7783 5719 7793 5753
rect 7741 5685 7793 5719
rect 7741 5651 7749 5685
rect 7783 5651 7793 5685
rect 7741 5637 7793 5651
rect 7823 5753 7877 5767
rect 7823 5719 7833 5753
rect 7867 5719 7877 5753
rect 7823 5685 7877 5719
rect 7823 5651 7833 5685
rect 7867 5651 7877 5685
rect 7823 5637 7877 5651
rect 7907 5753 7959 5767
rect 7907 5719 7917 5753
rect 7951 5719 7959 5753
rect 7907 5685 7959 5719
rect 8555 5753 8607 5767
rect 8555 5719 8563 5753
rect 8597 5719 8607 5753
rect 7907 5651 7917 5685
rect 7951 5651 7959 5685
rect 8555 5685 8607 5719
rect 7907 5637 7959 5651
rect 8555 5651 8563 5685
rect 8597 5651 8607 5685
rect 8555 5637 8607 5651
rect 8637 5753 8691 5767
rect 8637 5719 8647 5753
rect 8681 5719 8691 5753
rect 8637 5685 8691 5719
rect 8637 5651 8647 5685
rect 8681 5651 8691 5685
rect 8637 5637 8691 5651
rect 8721 5753 8773 5767
rect 8721 5719 8731 5753
rect 8765 5719 8773 5753
rect 8721 5685 8773 5719
rect 8721 5651 8731 5685
rect 8765 5651 8773 5685
rect 8721 5637 8773 5651
rect 9629 5753 9681 5767
rect 9629 5719 9637 5753
rect 9671 5719 9681 5753
rect 9629 5685 9681 5719
rect 9629 5651 9637 5685
rect 9671 5651 9681 5685
rect 9629 5637 9681 5651
rect 9711 5753 9765 5767
rect 9711 5719 9721 5753
rect 9755 5719 9765 5753
rect 9711 5685 9765 5719
rect 9711 5651 9721 5685
rect 9755 5651 9765 5685
rect 9711 5637 9765 5651
rect 9795 5753 9847 5767
rect 9795 5719 9805 5753
rect 9839 5719 9847 5753
rect 9795 5685 9847 5719
rect 10443 5753 10495 5767
rect 10443 5719 10451 5753
rect 10485 5719 10495 5753
rect 9795 5651 9805 5685
rect 9839 5651 9847 5685
rect 10443 5685 10495 5719
rect 9795 5637 9847 5651
rect 10443 5651 10451 5685
rect 10485 5651 10495 5685
rect 10443 5637 10495 5651
rect 10525 5753 10579 5767
rect 10525 5719 10535 5753
rect 10569 5719 10579 5753
rect 10525 5685 10579 5719
rect 10525 5651 10535 5685
rect 10569 5651 10579 5685
rect 10525 5637 10579 5651
rect 10609 5753 10661 5767
rect 10609 5719 10619 5753
rect 10653 5719 10661 5753
rect 10609 5685 10661 5719
rect 10609 5651 10619 5685
rect 10653 5651 10661 5685
rect 10609 5637 10661 5651
rect 11517 5753 11569 5767
rect 11517 5719 11525 5753
rect 11559 5719 11569 5753
rect 11517 5685 11569 5719
rect 11517 5651 11525 5685
rect 11559 5651 11569 5685
rect 11517 5637 11569 5651
rect 11599 5753 11653 5767
rect 11599 5719 11609 5753
rect 11643 5719 11653 5753
rect 11599 5685 11653 5719
rect 11599 5651 11609 5685
rect 11643 5651 11653 5685
rect 11599 5637 11653 5651
rect 11683 5753 11735 5767
rect 11683 5719 11693 5753
rect 11727 5719 11735 5753
rect 11683 5685 11735 5719
rect 12331 5753 12383 5767
rect 12331 5719 12339 5753
rect 12373 5719 12383 5753
rect 11683 5651 11693 5685
rect 11727 5651 11735 5685
rect 12331 5685 12383 5719
rect 11683 5637 11735 5651
rect 12331 5651 12339 5685
rect 12373 5651 12383 5685
rect 12331 5637 12383 5651
rect 12413 5753 12467 5767
rect 12413 5719 12423 5753
rect 12457 5719 12467 5753
rect 12413 5685 12467 5719
rect 12413 5651 12423 5685
rect 12457 5651 12467 5685
rect 12413 5637 12467 5651
rect 12497 5753 12549 5767
rect 12497 5719 12507 5753
rect 12541 5719 12549 5753
rect 12497 5685 12549 5719
rect 12497 5651 12507 5685
rect 12541 5651 12549 5685
rect 12497 5637 12549 5651
rect 13405 5753 13457 5767
rect 13405 5719 13413 5753
rect 13447 5719 13457 5753
rect 13405 5685 13457 5719
rect 13405 5651 13413 5685
rect 13447 5651 13457 5685
rect 13405 5637 13457 5651
rect 13487 5753 13541 5767
rect 13487 5719 13497 5753
rect 13531 5719 13541 5753
rect 13487 5685 13541 5719
rect 13487 5651 13497 5685
rect 13531 5651 13541 5685
rect 13487 5637 13541 5651
rect 13571 5753 13623 5767
rect 13571 5719 13581 5753
rect 13615 5719 13623 5753
rect 13571 5685 13623 5719
rect 14219 5753 14271 5767
rect 14219 5719 14227 5753
rect 14261 5719 14271 5753
rect 13571 5651 13581 5685
rect 13615 5651 13623 5685
rect 14219 5685 14271 5719
rect 13571 5637 13623 5651
rect 14219 5651 14227 5685
rect 14261 5651 14271 5685
rect 14219 5637 14271 5651
rect 14301 5753 14355 5767
rect 14301 5719 14311 5753
rect 14345 5719 14355 5753
rect 14301 5685 14355 5719
rect 14301 5651 14311 5685
rect 14345 5651 14355 5685
rect 14301 5637 14355 5651
rect 14385 5753 14437 5767
rect 14385 5719 14395 5753
rect 14429 5719 14437 5753
rect 14385 5685 14437 5719
rect 14385 5651 14395 5685
rect 14429 5651 14437 5685
rect 14385 5637 14437 5651
rect 15287 5753 15339 5767
rect 15287 5719 15295 5753
rect 15329 5719 15339 5753
rect 15287 5685 15339 5719
rect 15287 5651 15295 5685
rect 15329 5651 15339 5685
rect 15287 5637 15339 5651
rect 15369 5753 15423 5767
rect 15369 5719 15379 5753
rect 15413 5719 15423 5753
rect 15369 5685 15423 5719
rect 15369 5651 15379 5685
rect 15413 5651 15423 5685
rect 15369 5637 15423 5651
rect 15453 5753 15505 5767
rect 15453 5719 15463 5753
rect 15497 5719 15505 5753
rect 15453 5685 15505 5719
rect 16101 5753 16153 5767
rect 16101 5719 16109 5753
rect 16143 5719 16153 5753
rect 15453 5651 15463 5685
rect 15497 5651 15505 5685
rect 16101 5685 16153 5719
rect 15453 5637 15505 5651
rect 16101 5651 16109 5685
rect 16143 5651 16153 5685
rect 16101 5637 16153 5651
rect 16183 5753 16237 5767
rect 16183 5719 16193 5753
rect 16227 5719 16237 5753
rect 16183 5685 16237 5719
rect 16183 5651 16193 5685
rect 16227 5651 16237 5685
rect 16183 5637 16237 5651
rect 16267 5753 16319 5767
rect 16267 5719 16277 5753
rect 16311 5719 16319 5753
rect 16267 5685 16319 5719
rect 16267 5651 16277 5685
rect 16311 5651 16319 5685
rect 16267 5637 16319 5651
rect 17175 5753 17227 5767
rect 17175 5719 17183 5753
rect 17217 5719 17227 5753
rect 17175 5685 17227 5719
rect 17175 5651 17183 5685
rect 17217 5651 17227 5685
rect 17175 5637 17227 5651
rect 17257 5753 17311 5767
rect 17257 5719 17267 5753
rect 17301 5719 17311 5753
rect 17257 5685 17311 5719
rect 17257 5651 17267 5685
rect 17301 5651 17311 5685
rect 17257 5637 17311 5651
rect 17341 5753 17393 5767
rect 17341 5719 17351 5753
rect 17385 5719 17393 5753
rect 17341 5685 17393 5719
rect 17989 5753 18041 5767
rect 17989 5719 17997 5753
rect 18031 5719 18041 5753
rect 17341 5651 17351 5685
rect 17385 5651 17393 5685
rect 17989 5685 18041 5719
rect 17341 5637 17393 5651
rect 17989 5651 17997 5685
rect 18031 5651 18041 5685
rect 17989 5637 18041 5651
rect 18071 5753 18125 5767
rect 18071 5719 18081 5753
rect 18115 5719 18125 5753
rect 18071 5685 18125 5719
rect 18071 5651 18081 5685
rect 18115 5651 18125 5685
rect 18071 5637 18125 5651
rect 18155 5753 18207 5767
rect 18155 5719 18165 5753
rect 18199 5719 18207 5753
rect 18155 5685 18207 5719
rect 18155 5651 18165 5685
rect 18199 5651 18207 5685
rect 18155 5637 18207 5651
rect 19063 5753 19115 5767
rect 19063 5719 19071 5753
rect 19105 5719 19115 5753
rect 19063 5685 19115 5719
rect 19063 5651 19071 5685
rect 19105 5651 19115 5685
rect 19063 5637 19115 5651
rect 19145 5753 19199 5767
rect 19145 5719 19155 5753
rect 19189 5719 19199 5753
rect 19145 5685 19199 5719
rect 19145 5651 19155 5685
rect 19189 5651 19199 5685
rect 19145 5637 19199 5651
rect 19229 5753 19281 5767
rect 19229 5719 19239 5753
rect 19273 5719 19281 5753
rect 19229 5685 19281 5719
rect 19877 5753 19929 5767
rect 19877 5719 19885 5753
rect 19919 5719 19929 5753
rect 19229 5651 19239 5685
rect 19273 5651 19281 5685
rect 19877 5685 19929 5719
rect 19229 5637 19281 5651
rect 19877 5651 19885 5685
rect 19919 5651 19929 5685
rect 19877 5637 19929 5651
rect 19959 5753 20013 5767
rect 19959 5719 19969 5753
rect 20003 5719 20013 5753
rect 19959 5685 20013 5719
rect 19959 5651 19969 5685
rect 20003 5651 20013 5685
rect 19959 5637 20013 5651
rect 20043 5753 20095 5767
rect 20043 5719 20053 5753
rect 20087 5719 20095 5753
rect 20043 5685 20095 5719
rect 20043 5651 20053 5685
rect 20087 5651 20095 5685
rect 20043 5637 20095 5651
rect 20951 5753 21003 5767
rect 20951 5719 20959 5753
rect 20993 5719 21003 5753
rect 20951 5685 21003 5719
rect 20951 5651 20959 5685
rect 20993 5651 21003 5685
rect 20951 5637 21003 5651
rect 21033 5753 21087 5767
rect 21033 5719 21043 5753
rect 21077 5719 21087 5753
rect 21033 5685 21087 5719
rect 21033 5651 21043 5685
rect 21077 5651 21087 5685
rect 21033 5637 21087 5651
rect 21117 5753 21169 5767
rect 21117 5719 21127 5753
rect 21161 5719 21169 5753
rect 21117 5685 21169 5719
rect 21765 5753 21817 5767
rect 21765 5719 21773 5753
rect 21807 5719 21817 5753
rect 21117 5651 21127 5685
rect 21161 5651 21169 5685
rect 21765 5685 21817 5719
rect 21117 5637 21169 5651
rect 21765 5651 21773 5685
rect 21807 5651 21817 5685
rect 21765 5637 21817 5651
rect 21847 5753 21901 5767
rect 21847 5719 21857 5753
rect 21891 5719 21901 5753
rect 21847 5685 21901 5719
rect 21847 5651 21857 5685
rect 21891 5651 21901 5685
rect 21847 5637 21901 5651
rect 21931 5753 21983 5767
rect 21931 5719 21941 5753
rect 21975 5719 21983 5753
rect 21931 5685 21983 5719
rect 21931 5651 21941 5685
rect 21975 5651 21983 5685
rect 21931 5637 21983 5651
rect 22839 5753 22891 5767
rect 22839 5719 22847 5753
rect 22881 5719 22891 5753
rect 22839 5685 22891 5719
rect 22839 5651 22847 5685
rect 22881 5651 22891 5685
rect 22839 5637 22891 5651
rect 22921 5753 22975 5767
rect 22921 5719 22931 5753
rect 22965 5719 22975 5753
rect 22921 5685 22975 5719
rect 22921 5651 22931 5685
rect 22965 5651 22975 5685
rect 22921 5637 22975 5651
rect 23005 5753 23057 5767
rect 23005 5719 23015 5753
rect 23049 5719 23057 5753
rect 23005 5685 23057 5719
rect 23653 5753 23705 5767
rect 23653 5719 23661 5753
rect 23695 5719 23705 5753
rect 23005 5651 23015 5685
rect 23049 5651 23057 5685
rect 23653 5685 23705 5719
rect 23005 5637 23057 5651
rect 23653 5651 23661 5685
rect 23695 5651 23705 5685
rect 23653 5637 23705 5651
rect 23735 5753 23789 5767
rect 23735 5719 23745 5753
rect 23779 5719 23789 5753
rect 23735 5685 23789 5719
rect 23735 5651 23745 5685
rect 23779 5651 23789 5685
rect 23735 5637 23789 5651
rect 23819 5753 23871 5767
rect 23819 5719 23829 5753
rect 23863 5719 23871 5753
rect 23819 5685 23871 5719
rect 23819 5651 23829 5685
rect 23863 5651 23871 5685
rect 23819 5637 23871 5651
rect 24727 5753 24779 5767
rect 24727 5719 24735 5753
rect 24769 5719 24779 5753
rect 24727 5685 24779 5719
rect 24727 5651 24735 5685
rect 24769 5651 24779 5685
rect 24727 5637 24779 5651
rect 24809 5753 24863 5767
rect 24809 5719 24819 5753
rect 24853 5719 24863 5753
rect 24809 5685 24863 5719
rect 24809 5651 24819 5685
rect 24853 5651 24863 5685
rect 24809 5637 24863 5651
rect 24893 5753 24945 5767
rect 24893 5719 24903 5753
rect 24937 5719 24945 5753
rect 24893 5685 24945 5719
rect 25541 5753 25593 5767
rect 25541 5719 25549 5753
rect 25583 5719 25593 5753
rect 24893 5651 24903 5685
rect 24937 5651 24945 5685
rect 25541 5685 25593 5719
rect 24893 5637 24945 5651
rect 25541 5651 25549 5685
rect 25583 5651 25593 5685
rect 25541 5637 25593 5651
rect 25623 5753 25677 5767
rect 25623 5719 25633 5753
rect 25667 5719 25677 5753
rect 25623 5685 25677 5719
rect 25623 5651 25633 5685
rect 25667 5651 25677 5685
rect 25623 5637 25677 5651
rect 25707 5753 25759 5767
rect 25707 5719 25717 5753
rect 25751 5719 25759 5753
rect 25707 5685 25759 5719
rect 25707 5651 25717 5685
rect 25751 5651 25759 5685
rect 25707 5637 25759 5651
rect 26615 5753 26667 5767
rect 26615 5719 26623 5753
rect 26657 5719 26667 5753
rect 26615 5685 26667 5719
rect 26615 5651 26623 5685
rect 26657 5651 26667 5685
rect 26615 5637 26667 5651
rect 26697 5753 26751 5767
rect 26697 5719 26707 5753
rect 26741 5719 26751 5753
rect 26697 5685 26751 5719
rect 26697 5651 26707 5685
rect 26741 5651 26751 5685
rect 26697 5637 26751 5651
rect 26781 5753 26833 5767
rect 26781 5719 26791 5753
rect 26825 5719 26833 5753
rect 26781 5685 26833 5719
rect 27429 5753 27481 5767
rect 27429 5719 27437 5753
rect 27471 5719 27481 5753
rect 26781 5651 26791 5685
rect 26825 5651 26833 5685
rect 27429 5685 27481 5719
rect 26781 5637 26833 5651
rect 27429 5651 27437 5685
rect 27471 5651 27481 5685
rect 27429 5637 27481 5651
rect 27511 5753 27565 5767
rect 27511 5719 27521 5753
rect 27555 5719 27565 5753
rect 27511 5685 27565 5719
rect 27511 5651 27521 5685
rect 27555 5651 27565 5685
rect 27511 5637 27565 5651
rect 27595 5753 27647 5767
rect 27595 5719 27605 5753
rect 27639 5719 27647 5753
rect 27595 5685 27647 5719
rect 27595 5651 27605 5685
rect 27639 5651 27647 5685
rect 27595 5637 27647 5651
rect 28503 5753 28555 5767
rect 28503 5719 28511 5753
rect 28545 5719 28555 5753
rect 28503 5685 28555 5719
rect 28503 5651 28511 5685
rect 28545 5651 28555 5685
rect 28503 5637 28555 5651
rect 28585 5753 28639 5767
rect 28585 5719 28595 5753
rect 28629 5719 28639 5753
rect 28585 5685 28639 5719
rect 28585 5651 28595 5685
rect 28629 5651 28639 5685
rect 28585 5637 28639 5651
rect 28669 5753 28721 5767
rect 28669 5719 28679 5753
rect 28713 5719 28721 5753
rect 28669 5685 28721 5719
rect 29317 5753 29369 5767
rect 29317 5719 29325 5753
rect 29359 5719 29369 5753
rect 28669 5651 28679 5685
rect 28713 5651 28721 5685
rect 29317 5685 29369 5719
rect 28669 5637 28721 5651
rect 29317 5651 29325 5685
rect 29359 5651 29369 5685
rect 29317 5637 29369 5651
rect 29399 5753 29453 5767
rect 29399 5719 29409 5753
rect 29443 5719 29453 5753
rect 29399 5685 29453 5719
rect 29399 5651 29409 5685
rect 29443 5651 29453 5685
rect 29399 5637 29453 5651
rect 29483 5753 29535 5767
rect 29483 5719 29493 5753
rect 29527 5719 29535 5753
rect 29483 5685 29535 5719
rect 29483 5651 29493 5685
rect 29527 5651 29535 5685
rect 29483 5637 29535 5651
rect 30391 5753 30443 5767
rect 30391 5719 30399 5753
rect 30433 5719 30443 5753
rect 30391 5685 30443 5719
rect 30391 5651 30399 5685
rect 30433 5651 30443 5685
rect 30391 5637 30443 5651
rect 30473 5753 30527 5767
rect 30473 5719 30483 5753
rect 30517 5719 30527 5753
rect 30473 5685 30527 5719
rect 30473 5651 30483 5685
rect 30517 5651 30527 5685
rect 30473 5637 30527 5651
rect 30557 5753 30609 5767
rect 30557 5719 30567 5753
rect 30601 5719 30609 5753
rect 30557 5685 30609 5719
rect 31205 5753 31257 5767
rect 31205 5719 31213 5753
rect 31247 5719 31257 5753
rect 30557 5651 30567 5685
rect 30601 5651 30609 5685
rect 31205 5685 31257 5719
rect 30557 5637 30609 5651
rect 31205 5651 31213 5685
rect 31247 5651 31257 5685
rect 31205 5637 31257 5651
rect 31287 5753 31341 5767
rect 31287 5719 31297 5753
rect 31331 5719 31341 5753
rect 31287 5685 31341 5719
rect 31287 5651 31297 5685
rect 31331 5651 31341 5685
rect 31287 5637 31341 5651
rect 31371 5753 31423 5767
rect 31371 5719 31381 5753
rect 31415 5719 31423 5753
rect 31371 5685 31423 5719
rect 31371 5651 31381 5685
rect 31415 5651 31423 5685
rect 31371 5637 31423 5651
rect 32279 5753 32331 5767
rect 32279 5719 32287 5753
rect 32321 5719 32331 5753
rect 32279 5685 32331 5719
rect 32279 5651 32287 5685
rect 32321 5651 32331 5685
rect 32279 5637 32331 5651
rect 32361 5753 32415 5767
rect 32361 5719 32371 5753
rect 32405 5719 32415 5753
rect 32361 5685 32415 5719
rect 32361 5651 32371 5685
rect 32405 5651 32415 5685
rect 32361 5637 32415 5651
rect 32445 5753 32497 5767
rect 32445 5719 32455 5753
rect 32489 5719 32497 5753
rect 32445 5685 32497 5719
rect 33093 5753 33145 5767
rect 33093 5719 33101 5753
rect 33135 5719 33145 5753
rect 32445 5651 32455 5685
rect 32489 5651 32497 5685
rect 33093 5685 33145 5719
rect 32445 5637 32497 5651
rect 33093 5651 33101 5685
rect 33135 5651 33145 5685
rect 33093 5637 33145 5651
rect 33175 5753 33229 5767
rect 33175 5719 33185 5753
rect 33219 5719 33229 5753
rect 33175 5685 33229 5719
rect 33175 5651 33185 5685
rect 33219 5651 33229 5685
rect 33175 5637 33229 5651
rect 33259 5753 33311 5767
rect 33259 5719 33269 5753
rect 33303 5719 33311 5753
rect 33259 5685 33311 5719
rect 33259 5651 33269 5685
rect 33303 5651 33311 5685
rect 33259 5637 33311 5651
rect 34167 5753 34219 5767
rect 34167 5719 34175 5753
rect 34209 5719 34219 5753
rect 34167 5685 34219 5719
rect 34167 5651 34175 5685
rect 34209 5651 34219 5685
rect 34167 5637 34219 5651
rect 34249 5753 34303 5767
rect 34249 5719 34259 5753
rect 34293 5719 34303 5753
rect 34249 5685 34303 5719
rect 34249 5651 34259 5685
rect 34293 5651 34303 5685
rect 34249 5637 34303 5651
rect 34333 5753 34385 5767
rect 34333 5719 34343 5753
rect 34377 5719 34385 5753
rect 34333 5685 34385 5719
rect 34981 5753 35033 5767
rect 34981 5719 34989 5753
rect 35023 5719 35033 5753
rect 34333 5651 34343 5685
rect 34377 5651 34385 5685
rect 34981 5685 35033 5719
rect 34333 5637 34385 5651
rect 34981 5651 34989 5685
rect 35023 5651 35033 5685
rect 34981 5637 35033 5651
rect 35063 5753 35117 5767
rect 35063 5719 35073 5753
rect 35107 5719 35117 5753
rect 35063 5685 35117 5719
rect 35063 5651 35073 5685
rect 35107 5651 35117 5685
rect 35063 5637 35117 5651
rect 35147 5753 35199 5767
rect 35147 5719 35157 5753
rect 35191 5719 35199 5753
rect 35147 5685 35199 5719
rect 35147 5651 35157 5685
rect 35191 5651 35199 5685
rect 35147 5637 35199 5651
rect 36055 5753 36107 5767
rect 36055 5719 36063 5753
rect 36097 5719 36107 5753
rect 36055 5685 36107 5719
rect 36055 5651 36063 5685
rect 36097 5651 36107 5685
rect 36055 5637 36107 5651
rect 36137 5753 36191 5767
rect 36137 5719 36147 5753
rect 36181 5719 36191 5753
rect 36137 5685 36191 5719
rect 36137 5651 36147 5685
rect 36181 5651 36191 5685
rect 36137 5637 36191 5651
rect 36221 5753 36273 5767
rect 36221 5719 36231 5753
rect 36265 5719 36273 5753
rect 36221 5685 36273 5719
rect 36869 5753 36921 5767
rect 36869 5719 36877 5753
rect 36911 5719 36921 5753
rect 36221 5651 36231 5685
rect 36265 5651 36273 5685
rect 36869 5685 36921 5719
rect 36221 5637 36273 5651
rect 36869 5651 36877 5685
rect 36911 5651 36921 5685
rect 36869 5637 36921 5651
rect 36951 5753 37005 5767
rect 36951 5719 36961 5753
rect 36995 5719 37005 5753
rect 36951 5685 37005 5719
rect 36951 5651 36961 5685
rect 36995 5651 37005 5685
rect 36951 5637 37005 5651
rect 37035 5753 37087 5767
rect 37035 5719 37045 5753
rect 37079 5719 37087 5753
rect 37035 5685 37087 5719
rect 37035 5651 37045 5685
rect 37079 5651 37087 5685
rect 37035 5637 37087 5651
rect 37943 5753 37995 5767
rect 37943 5719 37951 5753
rect 37985 5719 37995 5753
rect 37943 5685 37995 5719
rect 37943 5651 37951 5685
rect 37985 5651 37995 5685
rect 37943 5637 37995 5651
rect 38025 5753 38079 5767
rect 38025 5719 38035 5753
rect 38069 5719 38079 5753
rect 38025 5685 38079 5719
rect 38025 5651 38035 5685
rect 38069 5651 38079 5685
rect 38025 5637 38079 5651
rect 38109 5753 38161 5767
rect 38109 5719 38119 5753
rect 38153 5719 38161 5753
rect 38109 5685 38161 5719
rect 38757 5753 38809 5767
rect 38757 5719 38765 5753
rect 38799 5719 38809 5753
rect 38109 5651 38119 5685
rect 38153 5651 38161 5685
rect 38757 5685 38809 5719
rect 38109 5637 38161 5651
rect 38757 5651 38765 5685
rect 38799 5651 38809 5685
rect 38757 5637 38809 5651
rect 38839 5753 38893 5767
rect 38839 5719 38849 5753
rect 38883 5719 38893 5753
rect 38839 5685 38893 5719
rect 38839 5651 38849 5685
rect 38883 5651 38893 5685
rect 38839 5637 38893 5651
rect 38923 5753 38975 5767
rect 38923 5719 38933 5753
rect 38967 5719 38975 5753
rect 38923 5685 38975 5719
rect 38923 5651 38933 5685
rect 38967 5651 38975 5685
rect 38923 5637 38975 5651
rect 39831 5753 39883 5767
rect 39831 5719 39839 5753
rect 39873 5719 39883 5753
rect 39831 5685 39883 5719
rect 39831 5651 39839 5685
rect 39873 5651 39883 5685
rect 39831 5637 39883 5651
rect 39913 5753 39967 5767
rect 39913 5719 39923 5753
rect 39957 5719 39967 5753
rect 39913 5685 39967 5719
rect 39913 5651 39923 5685
rect 39957 5651 39967 5685
rect 39913 5637 39967 5651
rect 39997 5753 40049 5767
rect 39997 5719 40007 5753
rect 40041 5719 40049 5753
rect 39997 5685 40049 5719
rect 40645 5753 40697 5767
rect 40645 5719 40653 5753
rect 40687 5719 40697 5753
rect 39997 5651 40007 5685
rect 40041 5651 40049 5685
rect 40645 5685 40697 5719
rect 39997 5637 40049 5651
rect 40645 5651 40653 5685
rect 40687 5651 40697 5685
rect 40645 5637 40697 5651
rect 40727 5753 40781 5767
rect 40727 5719 40737 5753
rect 40771 5719 40781 5753
rect 40727 5685 40781 5719
rect 40727 5651 40737 5685
rect 40771 5651 40781 5685
rect 40727 5637 40781 5651
rect 40811 5753 40863 5767
rect 40811 5719 40821 5753
rect 40855 5719 40863 5753
rect 40811 5685 40863 5719
rect 40811 5651 40821 5685
rect 40855 5651 40863 5685
rect 40811 5637 40863 5651
rect 41719 5753 41771 5767
rect 41719 5719 41727 5753
rect 41761 5719 41771 5753
rect 41719 5685 41771 5719
rect 41719 5651 41727 5685
rect 41761 5651 41771 5685
rect 41719 5637 41771 5651
rect 41801 5753 41855 5767
rect 41801 5719 41811 5753
rect 41845 5719 41855 5753
rect 41801 5685 41855 5719
rect 41801 5651 41811 5685
rect 41845 5651 41855 5685
rect 41801 5637 41855 5651
rect 41885 5753 41937 5767
rect 41885 5719 41895 5753
rect 41929 5719 41937 5753
rect 41885 5685 41937 5719
rect 42533 5753 42585 5767
rect 42533 5719 42541 5753
rect 42575 5719 42585 5753
rect 41885 5651 41895 5685
rect 41929 5651 41937 5685
rect 42533 5685 42585 5719
rect 41885 5637 41937 5651
rect 42533 5651 42541 5685
rect 42575 5651 42585 5685
rect 42533 5637 42585 5651
rect 42615 5753 42669 5767
rect 42615 5719 42625 5753
rect 42659 5719 42669 5753
rect 42615 5685 42669 5719
rect 42615 5651 42625 5685
rect 42659 5651 42669 5685
rect 42615 5637 42669 5651
rect 42699 5753 42751 5767
rect 42699 5719 42709 5753
rect 42743 5719 42751 5753
rect 42699 5685 42751 5719
rect 42699 5651 42709 5685
rect 42743 5651 42751 5685
rect 42699 5637 42751 5651
rect 43607 5753 43659 5767
rect 43607 5719 43615 5753
rect 43649 5719 43659 5753
rect 43607 5685 43659 5719
rect 43607 5651 43615 5685
rect 43649 5651 43659 5685
rect 43607 5637 43659 5651
rect 43689 5753 43743 5767
rect 43689 5719 43699 5753
rect 43733 5719 43743 5753
rect 43689 5685 43743 5719
rect 43689 5651 43699 5685
rect 43733 5651 43743 5685
rect 43689 5637 43743 5651
rect 43773 5753 43825 5767
rect 43773 5719 43783 5753
rect 43817 5719 43825 5753
rect 43773 5685 43825 5719
rect 44421 5753 44473 5767
rect 44421 5719 44429 5753
rect 44463 5719 44473 5753
rect 43773 5651 43783 5685
rect 43817 5651 43825 5685
rect 44421 5685 44473 5719
rect 43773 5637 43825 5651
rect 44421 5651 44429 5685
rect 44463 5651 44473 5685
rect 44421 5637 44473 5651
rect 44503 5753 44557 5767
rect 44503 5719 44513 5753
rect 44547 5719 44557 5753
rect 44503 5685 44557 5719
rect 44503 5651 44513 5685
rect 44547 5651 44557 5685
rect 44503 5637 44557 5651
rect 44587 5753 44639 5767
rect 44587 5719 44597 5753
rect 44631 5719 44639 5753
rect 44587 5685 44639 5719
rect 44587 5651 44597 5685
rect 44631 5651 44639 5685
rect 44587 5637 44639 5651
rect 45489 5753 45541 5767
rect 45489 5719 45497 5753
rect 45531 5719 45541 5753
rect 45489 5685 45541 5719
rect 45489 5651 45497 5685
rect 45531 5651 45541 5685
rect 45489 5637 45541 5651
rect 45571 5753 45625 5767
rect 45571 5719 45581 5753
rect 45615 5719 45625 5753
rect 45571 5685 45625 5719
rect 45571 5651 45581 5685
rect 45615 5651 45625 5685
rect 45571 5637 45625 5651
rect 45655 5753 45707 5767
rect 45655 5719 45665 5753
rect 45699 5719 45707 5753
rect 45655 5685 45707 5719
rect 46303 5753 46355 5767
rect 46303 5719 46311 5753
rect 46345 5719 46355 5753
rect 45655 5651 45665 5685
rect 45699 5651 45707 5685
rect 46303 5685 46355 5719
rect 45655 5637 45707 5651
rect 46303 5651 46311 5685
rect 46345 5651 46355 5685
rect 46303 5637 46355 5651
rect 46385 5753 46439 5767
rect 46385 5719 46395 5753
rect 46429 5719 46439 5753
rect 46385 5685 46439 5719
rect 46385 5651 46395 5685
rect 46429 5651 46439 5685
rect 46385 5637 46439 5651
rect 46469 5753 46521 5767
rect 46469 5719 46479 5753
rect 46513 5719 46521 5753
rect 46469 5685 46521 5719
rect 46469 5651 46479 5685
rect 46513 5651 46521 5685
rect 46469 5637 46521 5651
rect 47377 5753 47429 5767
rect 47377 5719 47385 5753
rect 47419 5719 47429 5753
rect 47377 5685 47429 5719
rect 47377 5651 47385 5685
rect 47419 5651 47429 5685
rect 47377 5637 47429 5651
rect 47459 5753 47513 5767
rect 47459 5719 47469 5753
rect 47503 5719 47513 5753
rect 47459 5685 47513 5719
rect 47459 5651 47469 5685
rect 47503 5651 47513 5685
rect 47459 5637 47513 5651
rect 47543 5753 47595 5767
rect 47543 5719 47553 5753
rect 47587 5719 47595 5753
rect 47543 5685 47595 5719
rect 48191 5753 48243 5767
rect 48191 5719 48199 5753
rect 48233 5719 48243 5753
rect 47543 5651 47553 5685
rect 47587 5651 47595 5685
rect 48191 5685 48243 5719
rect 47543 5637 47595 5651
rect 48191 5651 48199 5685
rect 48233 5651 48243 5685
rect 48191 5637 48243 5651
rect 48273 5753 48327 5767
rect 48273 5719 48283 5753
rect 48317 5719 48327 5753
rect 48273 5685 48327 5719
rect 48273 5651 48283 5685
rect 48317 5651 48327 5685
rect 48273 5637 48327 5651
rect 48357 5753 48409 5767
rect 48357 5719 48367 5753
rect 48401 5719 48409 5753
rect 48357 5685 48409 5719
rect 48357 5651 48367 5685
rect 48401 5651 48409 5685
rect 48357 5637 48409 5651
rect 49265 5753 49317 5767
rect 49265 5719 49273 5753
rect 49307 5719 49317 5753
rect 49265 5685 49317 5719
rect 49265 5651 49273 5685
rect 49307 5651 49317 5685
rect 49265 5637 49317 5651
rect 49347 5753 49401 5767
rect 49347 5719 49357 5753
rect 49391 5719 49401 5753
rect 49347 5685 49401 5719
rect 49347 5651 49357 5685
rect 49391 5651 49401 5685
rect 49347 5637 49401 5651
rect 49431 5753 49483 5767
rect 49431 5719 49441 5753
rect 49475 5719 49483 5753
rect 49431 5685 49483 5719
rect 50079 5753 50131 5767
rect 50079 5719 50087 5753
rect 50121 5719 50131 5753
rect 49431 5651 49441 5685
rect 49475 5651 49483 5685
rect 50079 5685 50131 5719
rect 49431 5637 49483 5651
rect 50079 5651 50087 5685
rect 50121 5651 50131 5685
rect 50079 5637 50131 5651
rect 50161 5753 50215 5767
rect 50161 5719 50171 5753
rect 50205 5719 50215 5753
rect 50161 5685 50215 5719
rect 50161 5651 50171 5685
rect 50205 5651 50215 5685
rect 50161 5637 50215 5651
rect 50245 5753 50297 5767
rect 50245 5719 50255 5753
rect 50289 5719 50297 5753
rect 50245 5685 50297 5719
rect 50245 5651 50255 5685
rect 50289 5651 50297 5685
rect 50245 5637 50297 5651
rect 51153 5753 51205 5767
rect 51153 5719 51161 5753
rect 51195 5719 51205 5753
rect 51153 5685 51205 5719
rect 51153 5651 51161 5685
rect 51195 5651 51205 5685
rect 51153 5637 51205 5651
rect 51235 5753 51289 5767
rect 51235 5719 51245 5753
rect 51279 5719 51289 5753
rect 51235 5685 51289 5719
rect 51235 5651 51245 5685
rect 51279 5651 51289 5685
rect 51235 5637 51289 5651
rect 51319 5753 51371 5767
rect 51319 5719 51329 5753
rect 51363 5719 51371 5753
rect 51319 5685 51371 5719
rect 51967 5753 52019 5767
rect 51967 5719 51975 5753
rect 52009 5719 52019 5753
rect 51319 5651 51329 5685
rect 51363 5651 51371 5685
rect 51967 5685 52019 5719
rect 51319 5637 51371 5651
rect 51967 5651 51975 5685
rect 52009 5651 52019 5685
rect 51967 5637 52019 5651
rect 52049 5753 52103 5767
rect 52049 5719 52059 5753
rect 52093 5719 52103 5753
rect 52049 5685 52103 5719
rect 52049 5651 52059 5685
rect 52093 5651 52103 5685
rect 52049 5637 52103 5651
rect 52133 5753 52185 5767
rect 52133 5719 52143 5753
rect 52177 5719 52185 5753
rect 52133 5685 52185 5719
rect 52133 5651 52143 5685
rect 52177 5651 52185 5685
rect 52133 5637 52185 5651
rect 53041 5753 53093 5767
rect 53041 5719 53049 5753
rect 53083 5719 53093 5753
rect 53041 5685 53093 5719
rect 53041 5651 53049 5685
rect 53083 5651 53093 5685
rect 53041 5637 53093 5651
rect 53123 5753 53177 5767
rect 53123 5719 53133 5753
rect 53167 5719 53177 5753
rect 53123 5685 53177 5719
rect 53123 5651 53133 5685
rect 53167 5651 53177 5685
rect 53123 5637 53177 5651
rect 53207 5753 53259 5767
rect 53207 5719 53217 5753
rect 53251 5719 53259 5753
rect 53207 5685 53259 5719
rect 53855 5753 53907 5767
rect 53855 5719 53863 5753
rect 53897 5719 53907 5753
rect 53207 5651 53217 5685
rect 53251 5651 53259 5685
rect 53855 5685 53907 5719
rect 53207 5637 53259 5651
rect 53855 5651 53863 5685
rect 53897 5651 53907 5685
rect 53855 5637 53907 5651
rect 53937 5753 53991 5767
rect 53937 5719 53947 5753
rect 53981 5719 53991 5753
rect 53937 5685 53991 5719
rect 53937 5651 53947 5685
rect 53981 5651 53991 5685
rect 53937 5637 53991 5651
rect 54021 5753 54073 5767
rect 54021 5719 54031 5753
rect 54065 5719 54073 5753
rect 54021 5685 54073 5719
rect 54021 5651 54031 5685
rect 54065 5651 54073 5685
rect 54021 5637 54073 5651
rect 54929 5753 54981 5767
rect 54929 5719 54937 5753
rect 54971 5719 54981 5753
rect 54929 5685 54981 5719
rect 54929 5651 54937 5685
rect 54971 5651 54981 5685
rect 54929 5637 54981 5651
rect 55011 5753 55065 5767
rect 55011 5719 55021 5753
rect 55055 5719 55065 5753
rect 55011 5685 55065 5719
rect 55011 5651 55021 5685
rect 55055 5651 55065 5685
rect 55011 5637 55065 5651
rect 55095 5753 55147 5767
rect 55095 5719 55105 5753
rect 55139 5719 55147 5753
rect 55095 5685 55147 5719
rect 55743 5753 55795 5767
rect 55743 5719 55751 5753
rect 55785 5719 55795 5753
rect 55095 5651 55105 5685
rect 55139 5651 55147 5685
rect 55743 5685 55795 5719
rect 55095 5637 55147 5651
rect 55743 5651 55751 5685
rect 55785 5651 55795 5685
rect 55743 5637 55795 5651
rect 55825 5753 55879 5767
rect 55825 5719 55835 5753
rect 55869 5719 55879 5753
rect 55825 5685 55879 5719
rect 55825 5651 55835 5685
rect 55869 5651 55879 5685
rect 55825 5637 55879 5651
rect 55909 5753 55961 5767
rect 55909 5719 55919 5753
rect 55953 5719 55961 5753
rect 55909 5685 55961 5719
rect 55909 5651 55919 5685
rect 55953 5651 55961 5685
rect 55909 5637 55961 5651
rect 56817 5753 56869 5767
rect 56817 5719 56825 5753
rect 56859 5719 56869 5753
rect 56817 5685 56869 5719
rect 56817 5651 56825 5685
rect 56859 5651 56869 5685
rect 56817 5637 56869 5651
rect 56899 5753 56953 5767
rect 56899 5719 56909 5753
rect 56943 5719 56953 5753
rect 56899 5685 56953 5719
rect 56899 5651 56909 5685
rect 56943 5651 56953 5685
rect 56899 5637 56953 5651
rect 56983 5753 57035 5767
rect 56983 5719 56993 5753
rect 57027 5719 57035 5753
rect 56983 5685 57035 5719
rect 57631 5753 57683 5767
rect 57631 5719 57639 5753
rect 57673 5719 57683 5753
rect 56983 5651 56993 5685
rect 57027 5651 57035 5685
rect 57631 5685 57683 5719
rect 56983 5637 57035 5651
rect 57631 5651 57639 5685
rect 57673 5651 57683 5685
rect 57631 5637 57683 5651
rect 57713 5753 57767 5767
rect 57713 5719 57723 5753
rect 57757 5719 57767 5753
rect 57713 5685 57767 5719
rect 57713 5651 57723 5685
rect 57757 5651 57767 5685
rect 57713 5637 57767 5651
rect 57797 5753 57849 5767
rect 57797 5719 57807 5753
rect 57841 5719 57849 5753
rect 57797 5685 57849 5719
rect 57797 5651 57807 5685
rect 57841 5651 57849 5685
rect 57797 5637 57849 5651
rect 58705 5753 58757 5767
rect 58705 5719 58713 5753
rect 58747 5719 58757 5753
rect 58705 5685 58757 5719
rect 58705 5651 58713 5685
rect 58747 5651 58757 5685
rect 58705 5637 58757 5651
rect 58787 5753 58841 5767
rect 58787 5719 58797 5753
rect 58831 5719 58841 5753
rect 58787 5685 58841 5719
rect 58787 5651 58797 5685
rect 58831 5651 58841 5685
rect 58787 5637 58841 5651
rect 58871 5753 58923 5767
rect 58871 5719 58881 5753
rect 58915 5719 58923 5753
rect 58871 5685 58923 5719
rect 59519 5753 59571 5767
rect 59519 5719 59527 5753
rect 59561 5719 59571 5753
rect 58871 5651 58881 5685
rect 58915 5651 58923 5685
rect 59519 5685 59571 5719
rect 58871 5637 58923 5651
rect 59519 5651 59527 5685
rect 59561 5651 59571 5685
rect 59519 5637 59571 5651
rect 59601 5753 59655 5767
rect 59601 5719 59611 5753
rect 59645 5719 59655 5753
rect 59601 5685 59655 5719
rect 59601 5651 59611 5685
rect 59645 5651 59655 5685
rect 59601 5637 59655 5651
rect 59685 5753 59737 5767
rect 59685 5719 59695 5753
rect 59729 5719 59737 5753
rect 59685 5685 59737 5719
rect 59685 5651 59695 5685
rect 59729 5651 59737 5685
rect 59685 5637 59737 5651
rect 5702 4809 5754 4825
rect 5702 4775 5710 4809
rect 5744 4775 5754 4809
rect 5702 4741 5754 4775
rect 5702 4707 5710 4741
rect 5744 4707 5754 4741
rect 5702 4695 5754 4707
rect 5784 4809 5838 4825
rect 5784 4775 5794 4809
rect 5828 4775 5838 4809
rect 5784 4741 5838 4775
rect 5784 4707 5794 4741
rect 5828 4707 5838 4741
rect 5784 4695 5838 4707
rect 5868 4741 5922 4825
rect 5868 4707 5878 4741
rect 5912 4707 5922 4741
rect 5868 4695 5922 4707
rect 5952 4809 6006 4825
rect 5952 4775 5962 4809
rect 5996 4775 6006 4809
rect 5952 4741 6006 4775
rect 5952 4707 5962 4741
rect 5996 4707 6006 4741
rect 5952 4695 6006 4707
rect 6036 4741 6090 4825
rect 6036 4707 6046 4741
rect 6080 4707 6090 4741
rect 6036 4695 6090 4707
rect 6120 4809 6174 4825
rect 6120 4775 6130 4809
rect 6164 4775 6174 4809
rect 6120 4741 6174 4775
rect 6120 4707 6130 4741
rect 6164 4707 6174 4741
rect 6120 4695 6174 4707
rect 6204 4741 6258 4825
rect 6204 4707 6214 4741
rect 6248 4707 6258 4741
rect 6204 4695 6258 4707
rect 6288 4809 6342 4825
rect 6288 4775 6298 4809
rect 6332 4775 6342 4809
rect 6288 4741 6342 4775
rect 6288 4707 6298 4741
rect 6332 4707 6342 4741
rect 6288 4695 6342 4707
rect 6372 4741 6426 4825
rect 6372 4707 6382 4741
rect 6416 4707 6426 4741
rect 6372 4695 6426 4707
rect 6456 4809 6510 4825
rect 6456 4775 6466 4809
rect 6500 4775 6510 4809
rect 6456 4741 6510 4775
rect 6456 4707 6466 4741
rect 6500 4707 6510 4741
rect 6456 4695 6510 4707
rect 6540 4741 6594 4825
rect 6540 4707 6550 4741
rect 6584 4707 6594 4741
rect 6540 4695 6594 4707
rect 6624 4809 6678 4825
rect 6624 4775 6634 4809
rect 6668 4775 6678 4809
rect 6624 4741 6678 4775
rect 6624 4707 6634 4741
rect 6668 4707 6678 4741
rect 6624 4695 6678 4707
rect 6708 4741 6762 4825
rect 6708 4707 6718 4741
rect 6752 4707 6762 4741
rect 6708 4695 6762 4707
rect 6792 4809 6846 4825
rect 6792 4775 6802 4809
rect 6836 4775 6846 4809
rect 6792 4741 6846 4775
rect 6792 4707 6802 4741
rect 6836 4707 6846 4741
rect 6792 4695 6846 4707
rect 6876 4741 6930 4825
rect 6876 4707 6886 4741
rect 6920 4707 6930 4741
rect 6876 4695 6930 4707
rect 6960 4809 7014 4825
rect 6960 4775 6970 4809
rect 7004 4775 7014 4809
rect 6960 4741 7014 4775
rect 6960 4707 6970 4741
rect 7004 4707 7014 4741
rect 6960 4695 7014 4707
rect 7044 4809 7096 4825
rect 7044 4775 7054 4809
rect 7088 4775 7096 4809
rect 7044 4741 7096 4775
rect 7044 4707 7054 4741
rect 7088 4707 7096 4741
rect 7044 4695 7096 4707
rect 7584 4807 7636 4823
rect 7584 4773 7592 4807
rect 7626 4773 7636 4807
rect 7584 4739 7636 4773
rect 7584 4705 7592 4739
rect 7626 4705 7636 4739
rect 7584 4693 7636 4705
rect 7666 4807 7720 4823
rect 7666 4773 7676 4807
rect 7710 4773 7720 4807
rect 7666 4739 7720 4773
rect 7666 4705 7676 4739
rect 7710 4705 7720 4739
rect 7666 4693 7720 4705
rect 7750 4739 7804 4823
rect 7750 4705 7760 4739
rect 7794 4705 7804 4739
rect 7750 4693 7804 4705
rect 7834 4807 7888 4823
rect 7834 4773 7844 4807
rect 7878 4773 7888 4807
rect 7834 4739 7888 4773
rect 7834 4705 7844 4739
rect 7878 4705 7888 4739
rect 7834 4693 7888 4705
rect 7918 4739 7972 4823
rect 7918 4705 7928 4739
rect 7962 4705 7972 4739
rect 7918 4693 7972 4705
rect 8002 4807 8056 4823
rect 8002 4773 8012 4807
rect 8046 4773 8056 4807
rect 8002 4739 8056 4773
rect 8002 4705 8012 4739
rect 8046 4705 8056 4739
rect 8002 4693 8056 4705
rect 8086 4739 8140 4823
rect 8086 4705 8096 4739
rect 8130 4705 8140 4739
rect 8086 4693 8140 4705
rect 8170 4807 8224 4823
rect 8170 4773 8180 4807
rect 8214 4773 8224 4807
rect 8170 4739 8224 4773
rect 8170 4705 8180 4739
rect 8214 4705 8224 4739
rect 8170 4693 8224 4705
rect 8254 4739 8308 4823
rect 8254 4705 8264 4739
rect 8298 4705 8308 4739
rect 8254 4693 8308 4705
rect 8338 4807 8392 4823
rect 8338 4773 8348 4807
rect 8382 4773 8392 4807
rect 8338 4739 8392 4773
rect 8338 4705 8348 4739
rect 8382 4705 8392 4739
rect 8338 4693 8392 4705
rect 8422 4739 8476 4823
rect 8422 4705 8432 4739
rect 8466 4705 8476 4739
rect 8422 4693 8476 4705
rect 8506 4807 8560 4823
rect 8506 4773 8516 4807
rect 8550 4773 8560 4807
rect 8506 4739 8560 4773
rect 8506 4705 8516 4739
rect 8550 4705 8560 4739
rect 8506 4693 8560 4705
rect 8590 4739 8644 4823
rect 8590 4705 8600 4739
rect 8634 4705 8644 4739
rect 8590 4693 8644 4705
rect 8674 4807 8728 4823
rect 8674 4773 8684 4807
rect 8718 4773 8728 4807
rect 8674 4739 8728 4773
rect 8674 4705 8684 4739
rect 8718 4705 8728 4739
rect 8674 4693 8728 4705
rect 8758 4739 8812 4823
rect 8758 4705 8768 4739
rect 8802 4705 8812 4739
rect 8758 4693 8812 4705
rect 8842 4807 8896 4823
rect 8842 4773 8852 4807
rect 8886 4773 8896 4807
rect 8842 4739 8896 4773
rect 8842 4705 8852 4739
rect 8886 4705 8896 4739
rect 8842 4693 8896 4705
rect 8926 4807 8978 4823
rect 8926 4773 8936 4807
rect 8970 4773 8978 4807
rect 8926 4739 8978 4773
rect 8926 4705 8936 4739
rect 8970 4705 8978 4739
rect 8926 4693 8978 4705
rect 20800 4809 20852 4825
rect 20800 4775 20808 4809
rect 20842 4775 20852 4809
rect 20800 4741 20852 4775
rect 20800 4707 20808 4741
rect 20842 4707 20852 4741
rect 20800 4695 20852 4707
rect 20882 4809 20936 4825
rect 20882 4775 20892 4809
rect 20926 4775 20936 4809
rect 20882 4741 20936 4775
rect 20882 4707 20892 4741
rect 20926 4707 20936 4741
rect 20882 4695 20936 4707
rect 20966 4741 21020 4825
rect 20966 4707 20976 4741
rect 21010 4707 21020 4741
rect 20966 4695 21020 4707
rect 21050 4809 21104 4825
rect 21050 4775 21060 4809
rect 21094 4775 21104 4809
rect 21050 4741 21104 4775
rect 21050 4707 21060 4741
rect 21094 4707 21104 4741
rect 21050 4695 21104 4707
rect 21134 4741 21188 4825
rect 21134 4707 21144 4741
rect 21178 4707 21188 4741
rect 21134 4695 21188 4707
rect 21218 4809 21272 4825
rect 21218 4775 21228 4809
rect 21262 4775 21272 4809
rect 21218 4741 21272 4775
rect 21218 4707 21228 4741
rect 21262 4707 21272 4741
rect 21218 4695 21272 4707
rect 21302 4741 21356 4825
rect 21302 4707 21312 4741
rect 21346 4707 21356 4741
rect 21302 4695 21356 4707
rect 21386 4809 21440 4825
rect 21386 4775 21396 4809
rect 21430 4775 21440 4809
rect 21386 4741 21440 4775
rect 21386 4707 21396 4741
rect 21430 4707 21440 4741
rect 21386 4695 21440 4707
rect 21470 4741 21524 4825
rect 21470 4707 21480 4741
rect 21514 4707 21524 4741
rect 21470 4695 21524 4707
rect 21554 4809 21608 4825
rect 21554 4775 21564 4809
rect 21598 4775 21608 4809
rect 21554 4741 21608 4775
rect 21554 4707 21564 4741
rect 21598 4707 21608 4741
rect 21554 4695 21608 4707
rect 21638 4741 21692 4825
rect 21638 4707 21648 4741
rect 21682 4707 21692 4741
rect 21638 4695 21692 4707
rect 21722 4809 21776 4825
rect 21722 4775 21732 4809
rect 21766 4775 21776 4809
rect 21722 4741 21776 4775
rect 21722 4707 21732 4741
rect 21766 4707 21776 4741
rect 21722 4695 21776 4707
rect 21806 4741 21860 4825
rect 21806 4707 21816 4741
rect 21850 4707 21860 4741
rect 21806 4695 21860 4707
rect 21890 4809 21944 4825
rect 21890 4775 21900 4809
rect 21934 4775 21944 4809
rect 21890 4741 21944 4775
rect 21890 4707 21900 4741
rect 21934 4707 21944 4741
rect 21890 4695 21944 4707
rect 21974 4741 22028 4825
rect 21974 4707 21984 4741
rect 22018 4707 22028 4741
rect 21974 4695 22028 4707
rect 22058 4809 22112 4825
rect 22058 4775 22068 4809
rect 22102 4775 22112 4809
rect 22058 4741 22112 4775
rect 22058 4707 22068 4741
rect 22102 4707 22112 4741
rect 22058 4695 22112 4707
rect 22142 4809 22194 4825
rect 22142 4775 22152 4809
rect 22186 4775 22194 4809
rect 22142 4741 22194 4775
rect 22142 4707 22152 4741
rect 22186 4707 22194 4741
rect 22142 4695 22194 4707
rect 22682 4807 22734 4823
rect 22682 4773 22690 4807
rect 22724 4773 22734 4807
rect 22682 4739 22734 4773
rect 22682 4705 22690 4739
rect 22724 4705 22734 4739
rect 22682 4693 22734 4705
rect 22764 4807 22818 4823
rect 22764 4773 22774 4807
rect 22808 4773 22818 4807
rect 22764 4739 22818 4773
rect 22764 4705 22774 4739
rect 22808 4705 22818 4739
rect 22764 4693 22818 4705
rect 22848 4739 22902 4823
rect 22848 4705 22858 4739
rect 22892 4705 22902 4739
rect 22848 4693 22902 4705
rect 22932 4807 22986 4823
rect 22932 4773 22942 4807
rect 22976 4773 22986 4807
rect 22932 4739 22986 4773
rect 22932 4705 22942 4739
rect 22976 4705 22986 4739
rect 22932 4693 22986 4705
rect 23016 4739 23070 4823
rect 23016 4705 23026 4739
rect 23060 4705 23070 4739
rect 23016 4693 23070 4705
rect 23100 4807 23154 4823
rect 23100 4773 23110 4807
rect 23144 4773 23154 4807
rect 23100 4739 23154 4773
rect 23100 4705 23110 4739
rect 23144 4705 23154 4739
rect 23100 4693 23154 4705
rect 23184 4739 23238 4823
rect 23184 4705 23194 4739
rect 23228 4705 23238 4739
rect 23184 4693 23238 4705
rect 23268 4807 23322 4823
rect 23268 4773 23278 4807
rect 23312 4773 23322 4807
rect 23268 4739 23322 4773
rect 23268 4705 23278 4739
rect 23312 4705 23322 4739
rect 23268 4693 23322 4705
rect 23352 4739 23406 4823
rect 23352 4705 23362 4739
rect 23396 4705 23406 4739
rect 23352 4693 23406 4705
rect 23436 4807 23490 4823
rect 23436 4773 23446 4807
rect 23480 4773 23490 4807
rect 23436 4739 23490 4773
rect 23436 4705 23446 4739
rect 23480 4705 23490 4739
rect 23436 4693 23490 4705
rect 23520 4739 23574 4823
rect 23520 4705 23530 4739
rect 23564 4705 23574 4739
rect 23520 4693 23574 4705
rect 23604 4807 23658 4823
rect 23604 4773 23614 4807
rect 23648 4773 23658 4807
rect 23604 4739 23658 4773
rect 23604 4705 23614 4739
rect 23648 4705 23658 4739
rect 23604 4693 23658 4705
rect 23688 4739 23742 4823
rect 23688 4705 23698 4739
rect 23732 4705 23742 4739
rect 23688 4693 23742 4705
rect 23772 4807 23826 4823
rect 23772 4773 23782 4807
rect 23816 4773 23826 4807
rect 23772 4739 23826 4773
rect 23772 4705 23782 4739
rect 23816 4705 23826 4739
rect 23772 4693 23826 4705
rect 23856 4739 23910 4823
rect 23856 4705 23866 4739
rect 23900 4705 23910 4739
rect 23856 4693 23910 4705
rect 23940 4807 23994 4823
rect 23940 4773 23950 4807
rect 23984 4773 23994 4807
rect 23940 4739 23994 4773
rect 23940 4705 23950 4739
rect 23984 4705 23994 4739
rect 23940 4693 23994 4705
rect 24024 4807 24076 4823
rect 24024 4773 24034 4807
rect 24068 4773 24076 4807
rect 24024 4739 24076 4773
rect 24024 4705 24034 4739
rect 24068 4705 24076 4739
rect 24024 4693 24076 4705
rect 35904 4809 35956 4825
rect 35904 4775 35912 4809
rect 35946 4775 35956 4809
rect 35904 4741 35956 4775
rect 35904 4707 35912 4741
rect 35946 4707 35956 4741
rect 35904 4695 35956 4707
rect 35986 4809 36040 4825
rect 35986 4775 35996 4809
rect 36030 4775 36040 4809
rect 35986 4741 36040 4775
rect 35986 4707 35996 4741
rect 36030 4707 36040 4741
rect 35986 4695 36040 4707
rect 36070 4741 36124 4825
rect 36070 4707 36080 4741
rect 36114 4707 36124 4741
rect 36070 4695 36124 4707
rect 36154 4809 36208 4825
rect 36154 4775 36164 4809
rect 36198 4775 36208 4809
rect 36154 4741 36208 4775
rect 36154 4707 36164 4741
rect 36198 4707 36208 4741
rect 36154 4695 36208 4707
rect 36238 4741 36292 4825
rect 36238 4707 36248 4741
rect 36282 4707 36292 4741
rect 36238 4695 36292 4707
rect 36322 4809 36376 4825
rect 36322 4775 36332 4809
rect 36366 4775 36376 4809
rect 36322 4741 36376 4775
rect 36322 4707 36332 4741
rect 36366 4707 36376 4741
rect 36322 4695 36376 4707
rect 36406 4741 36460 4825
rect 36406 4707 36416 4741
rect 36450 4707 36460 4741
rect 36406 4695 36460 4707
rect 36490 4809 36544 4825
rect 36490 4775 36500 4809
rect 36534 4775 36544 4809
rect 36490 4741 36544 4775
rect 36490 4707 36500 4741
rect 36534 4707 36544 4741
rect 36490 4695 36544 4707
rect 36574 4741 36628 4825
rect 36574 4707 36584 4741
rect 36618 4707 36628 4741
rect 36574 4695 36628 4707
rect 36658 4809 36712 4825
rect 36658 4775 36668 4809
rect 36702 4775 36712 4809
rect 36658 4741 36712 4775
rect 36658 4707 36668 4741
rect 36702 4707 36712 4741
rect 36658 4695 36712 4707
rect 36742 4741 36796 4825
rect 36742 4707 36752 4741
rect 36786 4707 36796 4741
rect 36742 4695 36796 4707
rect 36826 4809 36880 4825
rect 36826 4775 36836 4809
rect 36870 4775 36880 4809
rect 36826 4741 36880 4775
rect 36826 4707 36836 4741
rect 36870 4707 36880 4741
rect 36826 4695 36880 4707
rect 36910 4741 36964 4825
rect 36910 4707 36920 4741
rect 36954 4707 36964 4741
rect 36910 4695 36964 4707
rect 36994 4809 37048 4825
rect 36994 4775 37004 4809
rect 37038 4775 37048 4809
rect 36994 4741 37048 4775
rect 36994 4707 37004 4741
rect 37038 4707 37048 4741
rect 36994 4695 37048 4707
rect 37078 4741 37132 4825
rect 37078 4707 37088 4741
rect 37122 4707 37132 4741
rect 37078 4695 37132 4707
rect 37162 4809 37216 4825
rect 37162 4775 37172 4809
rect 37206 4775 37216 4809
rect 37162 4741 37216 4775
rect 37162 4707 37172 4741
rect 37206 4707 37216 4741
rect 37162 4695 37216 4707
rect 37246 4809 37298 4825
rect 37246 4775 37256 4809
rect 37290 4775 37298 4809
rect 37246 4741 37298 4775
rect 37246 4707 37256 4741
rect 37290 4707 37298 4741
rect 37246 4695 37298 4707
rect 37786 4807 37838 4823
rect 37786 4773 37794 4807
rect 37828 4773 37838 4807
rect 37786 4739 37838 4773
rect 37786 4705 37794 4739
rect 37828 4705 37838 4739
rect 37786 4693 37838 4705
rect 37868 4807 37922 4823
rect 37868 4773 37878 4807
rect 37912 4773 37922 4807
rect 37868 4739 37922 4773
rect 37868 4705 37878 4739
rect 37912 4705 37922 4739
rect 37868 4693 37922 4705
rect 37952 4739 38006 4823
rect 37952 4705 37962 4739
rect 37996 4705 38006 4739
rect 37952 4693 38006 4705
rect 38036 4807 38090 4823
rect 38036 4773 38046 4807
rect 38080 4773 38090 4807
rect 38036 4739 38090 4773
rect 38036 4705 38046 4739
rect 38080 4705 38090 4739
rect 38036 4693 38090 4705
rect 38120 4739 38174 4823
rect 38120 4705 38130 4739
rect 38164 4705 38174 4739
rect 38120 4693 38174 4705
rect 38204 4807 38258 4823
rect 38204 4773 38214 4807
rect 38248 4773 38258 4807
rect 38204 4739 38258 4773
rect 38204 4705 38214 4739
rect 38248 4705 38258 4739
rect 38204 4693 38258 4705
rect 38288 4739 38342 4823
rect 38288 4705 38298 4739
rect 38332 4705 38342 4739
rect 38288 4693 38342 4705
rect 38372 4807 38426 4823
rect 38372 4773 38382 4807
rect 38416 4773 38426 4807
rect 38372 4739 38426 4773
rect 38372 4705 38382 4739
rect 38416 4705 38426 4739
rect 38372 4693 38426 4705
rect 38456 4739 38510 4823
rect 38456 4705 38466 4739
rect 38500 4705 38510 4739
rect 38456 4693 38510 4705
rect 38540 4807 38594 4823
rect 38540 4773 38550 4807
rect 38584 4773 38594 4807
rect 38540 4739 38594 4773
rect 38540 4705 38550 4739
rect 38584 4705 38594 4739
rect 38540 4693 38594 4705
rect 38624 4739 38678 4823
rect 38624 4705 38634 4739
rect 38668 4705 38678 4739
rect 38624 4693 38678 4705
rect 38708 4807 38762 4823
rect 38708 4773 38718 4807
rect 38752 4773 38762 4807
rect 38708 4739 38762 4773
rect 38708 4705 38718 4739
rect 38752 4705 38762 4739
rect 38708 4693 38762 4705
rect 38792 4739 38846 4823
rect 38792 4705 38802 4739
rect 38836 4705 38846 4739
rect 38792 4693 38846 4705
rect 38876 4807 38930 4823
rect 38876 4773 38886 4807
rect 38920 4773 38930 4807
rect 38876 4739 38930 4773
rect 38876 4705 38886 4739
rect 38920 4705 38930 4739
rect 38876 4693 38930 4705
rect 38960 4739 39014 4823
rect 38960 4705 38970 4739
rect 39004 4705 39014 4739
rect 38960 4693 39014 4705
rect 39044 4807 39098 4823
rect 39044 4773 39054 4807
rect 39088 4773 39098 4807
rect 39044 4739 39098 4773
rect 39044 4705 39054 4739
rect 39088 4705 39098 4739
rect 39044 4693 39098 4705
rect 39128 4807 39180 4823
rect 39128 4773 39138 4807
rect 39172 4773 39180 4807
rect 39128 4739 39180 4773
rect 39128 4705 39138 4739
rect 39172 4705 39180 4739
rect 39128 4693 39180 4705
rect 51002 4809 51054 4825
rect 51002 4775 51010 4809
rect 51044 4775 51054 4809
rect 51002 4741 51054 4775
rect 51002 4707 51010 4741
rect 51044 4707 51054 4741
rect 51002 4695 51054 4707
rect 51084 4809 51138 4825
rect 51084 4775 51094 4809
rect 51128 4775 51138 4809
rect 51084 4741 51138 4775
rect 51084 4707 51094 4741
rect 51128 4707 51138 4741
rect 51084 4695 51138 4707
rect 51168 4741 51222 4825
rect 51168 4707 51178 4741
rect 51212 4707 51222 4741
rect 51168 4695 51222 4707
rect 51252 4809 51306 4825
rect 51252 4775 51262 4809
rect 51296 4775 51306 4809
rect 51252 4741 51306 4775
rect 51252 4707 51262 4741
rect 51296 4707 51306 4741
rect 51252 4695 51306 4707
rect 51336 4741 51390 4825
rect 51336 4707 51346 4741
rect 51380 4707 51390 4741
rect 51336 4695 51390 4707
rect 51420 4809 51474 4825
rect 51420 4775 51430 4809
rect 51464 4775 51474 4809
rect 51420 4741 51474 4775
rect 51420 4707 51430 4741
rect 51464 4707 51474 4741
rect 51420 4695 51474 4707
rect 51504 4741 51558 4825
rect 51504 4707 51514 4741
rect 51548 4707 51558 4741
rect 51504 4695 51558 4707
rect 51588 4809 51642 4825
rect 51588 4775 51598 4809
rect 51632 4775 51642 4809
rect 51588 4741 51642 4775
rect 51588 4707 51598 4741
rect 51632 4707 51642 4741
rect 51588 4695 51642 4707
rect 51672 4741 51726 4825
rect 51672 4707 51682 4741
rect 51716 4707 51726 4741
rect 51672 4695 51726 4707
rect 51756 4809 51810 4825
rect 51756 4775 51766 4809
rect 51800 4775 51810 4809
rect 51756 4741 51810 4775
rect 51756 4707 51766 4741
rect 51800 4707 51810 4741
rect 51756 4695 51810 4707
rect 51840 4741 51894 4825
rect 51840 4707 51850 4741
rect 51884 4707 51894 4741
rect 51840 4695 51894 4707
rect 51924 4809 51978 4825
rect 51924 4775 51934 4809
rect 51968 4775 51978 4809
rect 51924 4741 51978 4775
rect 51924 4707 51934 4741
rect 51968 4707 51978 4741
rect 51924 4695 51978 4707
rect 52008 4741 52062 4825
rect 52008 4707 52018 4741
rect 52052 4707 52062 4741
rect 52008 4695 52062 4707
rect 52092 4809 52146 4825
rect 52092 4775 52102 4809
rect 52136 4775 52146 4809
rect 52092 4741 52146 4775
rect 52092 4707 52102 4741
rect 52136 4707 52146 4741
rect 52092 4695 52146 4707
rect 52176 4741 52230 4825
rect 52176 4707 52186 4741
rect 52220 4707 52230 4741
rect 52176 4695 52230 4707
rect 52260 4809 52314 4825
rect 52260 4775 52270 4809
rect 52304 4775 52314 4809
rect 52260 4741 52314 4775
rect 52260 4707 52270 4741
rect 52304 4707 52314 4741
rect 52260 4695 52314 4707
rect 52344 4809 52396 4825
rect 52344 4775 52354 4809
rect 52388 4775 52396 4809
rect 52344 4741 52396 4775
rect 52344 4707 52354 4741
rect 52388 4707 52396 4741
rect 52344 4695 52396 4707
rect 52884 4807 52936 4823
rect 52884 4773 52892 4807
rect 52926 4773 52936 4807
rect 52884 4739 52936 4773
rect 52884 4705 52892 4739
rect 52926 4705 52936 4739
rect 52884 4693 52936 4705
rect 52966 4807 53020 4823
rect 52966 4773 52976 4807
rect 53010 4773 53020 4807
rect 52966 4739 53020 4773
rect 52966 4705 52976 4739
rect 53010 4705 53020 4739
rect 52966 4693 53020 4705
rect 53050 4739 53104 4823
rect 53050 4705 53060 4739
rect 53094 4705 53104 4739
rect 53050 4693 53104 4705
rect 53134 4807 53188 4823
rect 53134 4773 53144 4807
rect 53178 4773 53188 4807
rect 53134 4739 53188 4773
rect 53134 4705 53144 4739
rect 53178 4705 53188 4739
rect 53134 4693 53188 4705
rect 53218 4739 53272 4823
rect 53218 4705 53228 4739
rect 53262 4705 53272 4739
rect 53218 4693 53272 4705
rect 53302 4807 53356 4823
rect 53302 4773 53312 4807
rect 53346 4773 53356 4807
rect 53302 4739 53356 4773
rect 53302 4705 53312 4739
rect 53346 4705 53356 4739
rect 53302 4693 53356 4705
rect 53386 4739 53440 4823
rect 53386 4705 53396 4739
rect 53430 4705 53440 4739
rect 53386 4693 53440 4705
rect 53470 4807 53524 4823
rect 53470 4773 53480 4807
rect 53514 4773 53524 4807
rect 53470 4739 53524 4773
rect 53470 4705 53480 4739
rect 53514 4705 53524 4739
rect 53470 4693 53524 4705
rect 53554 4739 53608 4823
rect 53554 4705 53564 4739
rect 53598 4705 53608 4739
rect 53554 4693 53608 4705
rect 53638 4807 53692 4823
rect 53638 4773 53648 4807
rect 53682 4773 53692 4807
rect 53638 4739 53692 4773
rect 53638 4705 53648 4739
rect 53682 4705 53692 4739
rect 53638 4693 53692 4705
rect 53722 4739 53776 4823
rect 53722 4705 53732 4739
rect 53766 4705 53776 4739
rect 53722 4693 53776 4705
rect 53806 4807 53860 4823
rect 53806 4773 53816 4807
rect 53850 4773 53860 4807
rect 53806 4739 53860 4773
rect 53806 4705 53816 4739
rect 53850 4705 53860 4739
rect 53806 4693 53860 4705
rect 53890 4739 53944 4823
rect 53890 4705 53900 4739
rect 53934 4705 53944 4739
rect 53890 4693 53944 4705
rect 53974 4807 54028 4823
rect 53974 4773 53984 4807
rect 54018 4773 54028 4807
rect 53974 4739 54028 4773
rect 53974 4705 53984 4739
rect 54018 4705 54028 4739
rect 53974 4693 54028 4705
rect 54058 4739 54112 4823
rect 54058 4705 54068 4739
rect 54102 4705 54112 4739
rect 54058 4693 54112 4705
rect 54142 4807 54196 4823
rect 54142 4773 54152 4807
rect 54186 4773 54196 4807
rect 54142 4739 54196 4773
rect 54142 4705 54152 4739
rect 54186 4705 54196 4739
rect 54142 4693 54196 4705
rect 54226 4807 54278 4823
rect 54226 4773 54236 4807
rect 54270 4773 54278 4807
rect 54226 4739 54278 4773
rect 54226 4705 54236 4739
rect 54270 4705 54278 4739
rect 54226 4693 54278 4705
rect 30064 3664 30116 3748
rect 30064 3630 30072 3664
rect 30106 3630 30116 3664
rect 30064 3618 30116 3630
rect 30146 3672 30200 3748
rect 30146 3638 30156 3672
rect 30190 3638 30200 3672
rect 30146 3618 30200 3638
rect 30230 3664 30284 3748
rect 30230 3630 30240 3664
rect 30274 3630 30284 3664
rect 30230 3618 30284 3630
rect 30314 3672 30368 3748
rect 30314 3638 30324 3672
rect 30358 3638 30368 3672
rect 30314 3618 30368 3638
rect 30398 3665 30450 3748
rect 30398 3631 30408 3665
rect 30442 3631 30450 3665
rect 30398 3618 30450 3631
rect 30595 3732 30647 3748
rect 30595 3698 30603 3732
rect 30637 3698 30647 3732
rect 30595 3664 30647 3698
rect 30595 3630 30603 3664
rect 30637 3630 30647 3664
rect 30595 3618 30647 3630
rect 30677 3732 30731 3748
rect 30677 3698 30687 3732
rect 30721 3698 30731 3732
rect 30677 3664 30731 3698
rect 30677 3630 30687 3664
rect 30721 3630 30731 3664
rect 30677 3618 30731 3630
rect 30761 3664 30815 3748
rect 30761 3630 30771 3664
rect 30805 3630 30815 3664
rect 30761 3618 30815 3630
rect 30845 3732 30899 3748
rect 30845 3698 30855 3732
rect 30889 3698 30899 3732
rect 30845 3664 30899 3698
rect 30845 3630 30855 3664
rect 30889 3630 30899 3664
rect 30845 3618 30899 3630
rect 30929 3664 30983 3748
rect 30929 3630 30939 3664
rect 30973 3630 30983 3664
rect 30929 3618 30983 3630
rect 31013 3732 31067 3748
rect 31013 3698 31023 3732
rect 31057 3698 31067 3732
rect 31013 3664 31067 3698
rect 31013 3630 31023 3664
rect 31057 3630 31067 3664
rect 31013 3618 31067 3630
rect 31097 3664 31151 3748
rect 31097 3630 31107 3664
rect 31141 3630 31151 3664
rect 31097 3618 31151 3630
rect 31181 3732 31235 3748
rect 31181 3698 31191 3732
rect 31225 3698 31235 3732
rect 31181 3664 31235 3698
rect 31181 3630 31191 3664
rect 31225 3630 31235 3664
rect 31181 3618 31235 3630
rect 31265 3664 31319 3748
rect 31265 3630 31275 3664
rect 31309 3630 31319 3664
rect 31265 3618 31319 3630
rect 31349 3732 31403 3748
rect 31349 3698 31359 3732
rect 31393 3698 31403 3732
rect 31349 3664 31403 3698
rect 31349 3630 31359 3664
rect 31393 3630 31403 3664
rect 31349 3618 31403 3630
rect 31433 3664 31487 3748
rect 31433 3630 31443 3664
rect 31477 3630 31487 3664
rect 31433 3618 31487 3630
rect 31517 3732 31571 3748
rect 31517 3698 31527 3732
rect 31561 3698 31571 3732
rect 31517 3664 31571 3698
rect 31517 3630 31527 3664
rect 31561 3630 31571 3664
rect 31517 3618 31571 3630
rect 31601 3664 31655 3748
rect 31601 3630 31611 3664
rect 31645 3630 31655 3664
rect 31601 3618 31655 3630
rect 31685 3732 31739 3748
rect 31685 3698 31695 3732
rect 31729 3698 31739 3732
rect 31685 3664 31739 3698
rect 31685 3630 31695 3664
rect 31729 3630 31739 3664
rect 31685 3618 31739 3630
rect 31769 3664 31823 3748
rect 31769 3630 31779 3664
rect 31813 3630 31823 3664
rect 31769 3618 31823 3630
rect 31853 3732 31907 3748
rect 31853 3698 31863 3732
rect 31897 3698 31907 3732
rect 31853 3664 31907 3698
rect 31853 3630 31863 3664
rect 31897 3630 31907 3664
rect 31853 3618 31907 3630
rect 31937 3732 31989 3748
rect 31937 3698 31947 3732
rect 31981 3698 31989 3732
rect 31937 3664 31989 3698
rect 31937 3630 31947 3664
rect 31981 3630 31989 3664
rect 31937 3618 31989 3630
rect 43421 3516 43473 3532
rect 43421 3482 43429 3516
rect 43463 3482 43473 3516
rect 43421 3448 43473 3482
rect 43421 3414 43429 3448
rect 43463 3414 43473 3448
rect 43421 3402 43473 3414
rect 43503 3516 43557 3532
rect 43503 3482 43513 3516
rect 43547 3482 43557 3516
rect 43503 3448 43557 3482
rect 43503 3414 43513 3448
rect 43547 3414 43557 3448
rect 43503 3402 43557 3414
rect 43587 3448 43641 3532
rect 43587 3414 43597 3448
rect 43631 3414 43641 3448
rect 43587 3402 43641 3414
rect 43671 3516 43725 3532
rect 43671 3482 43681 3516
rect 43715 3482 43725 3516
rect 43671 3448 43725 3482
rect 43671 3414 43681 3448
rect 43715 3414 43725 3448
rect 43671 3402 43725 3414
rect 43755 3448 43809 3532
rect 43755 3414 43765 3448
rect 43799 3414 43809 3448
rect 43755 3402 43809 3414
rect 43839 3516 43893 3532
rect 43839 3482 43849 3516
rect 43883 3482 43893 3516
rect 43839 3448 43893 3482
rect 43839 3414 43849 3448
rect 43883 3414 43893 3448
rect 43839 3402 43893 3414
rect 43923 3448 43977 3532
rect 43923 3414 43933 3448
rect 43967 3414 43977 3448
rect 43923 3402 43977 3414
rect 44007 3516 44061 3532
rect 44007 3482 44017 3516
rect 44051 3482 44061 3516
rect 44007 3448 44061 3482
rect 44007 3414 44017 3448
rect 44051 3414 44061 3448
rect 44007 3402 44061 3414
rect 44091 3448 44145 3532
rect 44091 3414 44101 3448
rect 44135 3414 44145 3448
rect 44091 3402 44145 3414
rect 44175 3516 44229 3532
rect 44175 3482 44185 3516
rect 44219 3482 44229 3516
rect 44175 3448 44229 3482
rect 44175 3414 44185 3448
rect 44219 3414 44229 3448
rect 44175 3402 44229 3414
rect 44259 3448 44313 3532
rect 44259 3414 44269 3448
rect 44303 3414 44313 3448
rect 44259 3402 44313 3414
rect 44343 3516 44397 3532
rect 44343 3482 44353 3516
rect 44387 3482 44397 3516
rect 44343 3448 44397 3482
rect 44343 3414 44353 3448
rect 44387 3414 44397 3448
rect 44343 3402 44397 3414
rect 44427 3448 44481 3532
rect 44427 3414 44437 3448
rect 44471 3414 44481 3448
rect 44427 3402 44481 3414
rect 44511 3516 44565 3532
rect 44511 3482 44521 3516
rect 44555 3482 44565 3516
rect 44511 3448 44565 3482
rect 44511 3414 44521 3448
rect 44555 3414 44565 3448
rect 44511 3402 44565 3414
rect 44595 3448 44649 3532
rect 44595 3414 44605 3448
rect 44639 3414 44649 3448
rect 44595 3402 44649 3414
rect 44679 3516 44733 3532
rect 44679 3482 44689 3516
rect 44723 3482 44733 3516
rect 44679 3448 44733 3482
rect 44679 3414 44689 3448
rect 44723 3414 44733 3448
rect 44679 3402 44733 3414
rect 44763 3516 44815 3532
rect 44763 3482 44773 3516
rect 44807 3482 44815 3516
rect 44763 3448 44815 3482
rect 44763 3414 44773 3448
rect 44807 3414 44815 3448
rect 44763 3402 44815 3414
rect 45351 3516 45403 3532
rect 45351 3482 45359 3516
rect 45393 3482 45403 3516
rect 45351 3448 45403 3482
rect 45351 3414 45359 3448
rect 45393 3414 45403 3448
rect 45351 3402 45403 3414
rect 45433 3516 45487 3532
rect 45433 3482 45443 3516
rect 45477 3482 45487 3516
rect 45433 3448 45487 3482
rect 45433 3414 45443 3448
rect 45477 3414 45487 3448
rect 45433 3402 45487 3414
rect 45517 3448 45571 3532
rect 45517 3414 45527 3448
rect 45561 3414 45571 3448
rect 45517 3402 45571 3414
rect 45601 3516 45655 3532
rect 45601 3482 45611 3516
rect 45645 3482 45655 3516
rect 45601 3448 45655 3482
rect 45601 3414 45611 3448
rect 45645 3414 45655 3448
rect 45601 3402 45655 3414
rect 45685 3448 45739 3532
rect 45685 3414 45695 3448
rect 45729 3414 45739 3448
rect 45685 3402 45739 3414
rect 45769 3516 45823 3532
rect 45769 3482 45779 3516
rect 45813 3482 45823 3516
rect 45769 3448 45823 3482
rect 45769 3414 45779 3448
rect 45813 3414 45823 3448
rect 45769 3402 45823 3414
rect 45853 3448 45907 3532
rect 45853 3414 45863 3448
rect 45897 3414 45907 3448
rect 45853 3402 45907 3414
rect 45937 3516 45991 3532
rect 45937 3482 45947 3516
rect 45981 3482 45991 3516
rect 45937 3448 45991 3482
rect 45937 3414 45947 3448
rect 45981 3414 45991 3448
rect 45937 3402 45991 3414
rect 46021 3448 46075 3532
rect 46021 3414 46031 3448
rect 46065 3414 46075 3448
rect 46021 3402 46075 3414
rect 46105 3516 46159 3532
rect 46105 3482 46115 3516
rect 46149 3482 46159 3516
rect 46105 3448 46159 3482
rect 46105 3414 46115 3448
rect 46149 3414 46159 3448
rect 46105 3402 46159 3414
rect 46189 3448 46243 3532
rect 46189 3414 46199 3448
rect 46233 3414 46243 3448
rect 46189 3402 46243 3414
rect 46273 3516 46327 3532
rect 46273 3482 46283 3516
rect 46317 3482 46327 3516
rect 46273 3448 46327 3482
rect 46273 3414 46283 3448
rect 46317 3414 46327 3448
rect 46273 3402 46327 3414
rect 46357 3448 46411 3532
rect 46357 3414 46367 3448
rect 46401 3414 46411 3448
rect 46357 3402 46411 3414
rect 46441 3516 46495 3532
rect 46441 3482 46451 3516
rect 46485 3482 46495 3516
rect 46441 3448 46495 3482
rect 46441 3414 46451 3448
rect 46485 3414 46495 3448
rect 46441 3402 46495 3414
rect 46525 3448 46579 3532
rect 46525 3414 46535 3448
rect 46569 3414 46579 3448
rect 46525 3402 46579 3414
rect 46609 3516 46663 3532
rect 46609 3482 46619 3516
rect 46653 3482 46663 3516
rect 46609 3448 46663 3482
rect 46609 3414 46619 3448
rect 46653 3414 46663 3448
rect 46609 3402 46663 3414
rect 46693 3516 46745 3532
rect 46693 3482 46703 3516
rect 46737 3482 46745 3516
rect 46693 3448 46745 3482
rect 46693 3414 46703 3448
rect 46737 3414 46745 3448
rect 46693 3402 46745 3414
rect 13279 3356 13331 3372
rect 13279 3322 13287 3356
rect 13321 3322 13331 3356
rect 13279 3288 13331 3322
rect 13279 3254 13287 3288
rect 13321 3254 13331 3288
rect 13279 3242 13331 3254
rect 13361 3356 13415 3372
rect 13361 3322 13371 3356
rect 13405 3322 13415 3356
rect 13361 3288 13415 3322
rect 13361 3254 13371 3288
rect 13405 3254 13415 3288
rect 13361 3242 13415 3254
rect 13445 3288 13499 3372
rect 13445 3254 13455 3288
rect 13489 3254 13499 3288
rect 13445 3242 13499 3254
rect 13529 3356 13583 3372
rect 13529 3322 13539 3356
rect 13573 3322 13583 3356
rect 13529 3288 13583 3322
rect 13529 3254 13539 3288
rect 13573 3254 13583 3288
rect 13529 3242 13583 3254
rect 13613 3288 13667 3372
rect 13613 3254 13623 3288
rect 13657 3254 13667 3288
rect 13613 3242 13667 3254
rect 13697 3356 13751 3372
rect 13697 3322 13707 3356
rect 13741 3322 13751 3356
rect 13697 3288 13751 3322
rect 13697 3254 13707 3288
rect 13741 3254 13751 3288
rect 13697 3242 13751 3254
rect 13781 3288 13835 3372
rect 13781 3254 13791 3288
rect 13825 3254 13835 3288
rect 13781 3242 13835 3254
rect 13865 3356 13919 3372
rect 13865 3322 13875 3356
rect 13909 3322 13919 3356
rect 13865 3288 13919 3322
rect 13865 3254 13875 3288
rect 13909 3254 13919 3288
rect 13865 3242 13919 3254
rect 13949 3288 14003 3372
rect 13949 3254 13959 3288
rect 13993 3254 14003 3288
rect 13949 3242 14003 3254
rect 14033 3356 14087 3372
rect 14033 3322 14043 3356
rect 14077 3322 14087 3356
rect 14033 3288 14087 3322
rect 14033 3254 14043 3288
rect 14077 3254 14087 3288
rect 14033 3242 14087 3254
rect 14117 3288 14171 3372
rect 14117 3254 14127 3288
rect 14161 3254 14171 3288
rect 14117 3242 14171 3254
rect 14201 3356 14255 3372
rect 14201 3322 14211 3356
rect 14245 3322 14255 3356
rect 14201 3288 14255 3322
rect 14201 3254 14211 3288
rect 14245 3254 14255 3288
rect 14201 3242 14255 3254
rect 14285 3288 14339 3372
rect 14285 3254 14295 3288
rect 14329 3254 14339 3288
rect 14285 3242 14339 3254
rect 14369 3356 14423 3372
rect 14369 3322 14379 3356
rect 14413 3322 14423 3356
rect 14369 3288 14423 3322
rect 14369 3254 14379 3288
rect 14413 3254 14423 3288
rect 14369 3242 14423 3254
rect 14453 3288 14507 3372
rect 14453 3254 14463 3288
rect 14497 3254 14507 3288
rect 14453 3242 14507 3254
rect 14537 3356 14591 3372
rect 14537 3322 14547 3356
rect 14581 3322 14591 3356
rect 14537 3288 14591 3322
rect 14537 3254 14547 3288
rect 14581 3254 14591 3288
rect 14537 3242 14591 3254
rect 14621 3356 14673 3372
rect 14621 3322 14631 3356
rect 14665 3322 14673 3356
rect 14621 3288 14673 3322
rect 14621 3254 14631 3288
rect 14665 3254 14673 3288
rect 14621 3242 14673 3254
rect 15209 3356 15261 3372
rect 15209 3322 15217 3356
rect 15251 3322 15261 3356
rect 15209 3288 15261 3322
rect 15209 3254 15217 3288
rect 15251 3254 15261 3288
rect 15209 3242 15261 3254
rect 15291 3356 15345 3372
rect 15291 3322 15301 3356
rect 15335 3322 15345 3356
rect 15291 3288 15345 3322
rect 15291 3254 15301 3288
rect 15335 3254 15345 3288
rect 15291 3242 15345 3254
rect 15375 3288 15429 3372
rect 15375 3254 15385 3288
rect 15419 3254 15429 3288
rect 15375 3242 15429 3254
rect 15459 3356 15513 3372
rect 15459 3322 15469 3356
rect 15503 3322 15513 3356
rect 15459 3288 15513 3322
rect 15459 3254 15469 3288
rect 15503 3254 15513 3288
rect 15459 3242 15513 3254
rect 15543 3288 15597 3372
rect 15543 3254 15553 3288
rect 15587 3254 15597 3288
rect 15543 3242 15597 3254
rect 15627 3356 15681 3372
rect 15627 3322 15637 3356
rect 15671 3322 15681 3356
rect 15627 3288 15681 3322
rect 15627 3254 15637 3288
rect 15671 3254 15681 3288
rect 15627 3242 15681 3254
rect 15711 3288 15765 3372
rect 15711 3254 15721 3288
rect 15755 3254 15765 3288
rect 15711 3242 15765 3254
rect 15795 3356 15849 3372
rect 15795 3322 15805 3356
rect 15839 3322 15849 3356
rect 15795 3288 15849 3322
rect 15795 3254 15805 3288
rect 15839 3254 15849 3288
rect 15795 3242 15849 3254
rect 15879 3288 15933 3372
rect 15879 3254 15889 3288
rect 15923 3254 15933 3288
rect 15879 3242 15933 3254
rect 15963 3356 16017 3372
rect 15963 3322 15973 3356
rect 16007 3322 16017 3356
rect 15963 3288 16017 3322
rect 15963 3254 15973 3288
rect 16007 3254 16017 3288
rect 15963 3242 16017 3254
rect 16047 3288 16101 3372
rect 16047 3254 16057 3288
rect 16091 3254 16101 3288
rect 16047 3242 16101 3254
rect 16131 3356 16185 3372
rect 16131 3322 16141 3356
rect 16175 3322 16185 3356
rect 16131 3288 16185 3322
rect 16131 3254 16141 3288
rect 16175 3254 16185 3288
rect 16131 3242 16185 3254
rect 16215 3288 16269 3372
rect 16215 3254 16225 3288
rect 16259 3254 16269 3288
rect 16215 3242 16269 3254
rect 16299 3356 16353 3372
rect 16299 3322 16309 3356
rect 16343 3322 16353 3356
rect 16299 3288 16353 3322
rect 16299 3254 16309 3288
rect 16343 3254 16353 3288
rect 16299 3242 16353 3254
rect 16383 3288 16437 3372
rect 16383 3254 16393 3288
rect 16427 3254 16437 3288
rect 16383 3242 16437 3254
rect 16467 3356 16521 3372
rect 16467 3322 16477 3356
rect 16511 3322 16521 3356
rect 16467 3288 16521 3322
rect 16467 3254 16477 3288
rect 16511 3254 16521 3288
rect 16467 3242 16521 3254
rect 16551 3356 16603 3372
rect 16551 3322 16561 3356
rect 16595 3322 16603 3356
rect 16551 3288 16603 3322
rect 16551 3254 16561 3288
rect 16595 3254 16603 3288
rect 16551 3242 16603 3254
rect 5704 2735 5756 2747
rect 5704 2701 5712 2735
rect 5746 2701 5756 2735
rect 5704 2667 5756 2701
rect 5704 2633 5712 2667
rect 5746 2633 5756 2667
rect 5704 2617 5756 2633
rect 5786 2735 5840 2747
rect 5786 2701 5796 2735
rect 5830 2701 5840 2735
rect 5786 2667 5840 2701
rect 5786 2633 5796 2667
rect 5830 2633 5840 2667
rect 5786 2617 5840 2633
rect 5870 2735 5924 2747
rect 5870 2701 5880 2735
rect 5914 2701 5924 2735
rect 5870 2617 5924 2701
rect 5954 2735 6008 2747
rect 5954 2701 5964 2735
rect 5998 2701 6008 2735
rect 5954 2667 6008 2701
rect 5954 2633 5964 2667
rect 5998 2633 6008 2667
rect 5954 2617 6008 2633
rect 6038 2735 6092 2747
rect 6038 2701 6048 2735
rect 6082 2701 6092 2735
rect 6038 2617 6092 2701
rect 6122 2735 6176 2747
rect 6122 2701 6132 2735
rect 6166 2701 6176 2735
rect 6122 2667 6176 2701
rect 6122 2633 6132 2667
rect 6166 2633 6176 2667
rect 6122 2617 6176 2633
rect 6206 2735 6260 2747
rect 6206 2701 6216 2735
rect 6250 2701 6260 2735
rect 6206 2617 6260 2701
rect 6290 2735 6344 2747
rect 6290 2701 6300 2735
rect 6334 2701 6344 2735
rect 6290 2667 6344 2701
rect 6290 2633 6300 2667
rect 6334 2633 6344 2667
rect 6290 2617 6344 2633
rect 6374 2735 6428 2747
rect 6374 2701 6384 2735
rect 6418 2701 6428 2735
rect 6374 2617 6428 2701
rect 6458 2735 6512 2747
rect 6458 2701 6468 2735
rect 6502 2701 6512 2735
rect 6458 2667 6512 2701
rect 6458 2633 6468 2667
rect 6502 2633 6512 2667
rect 6458 2617 6512 2633
rect 6542 2735 6596 2747
rect 6542 2701 6552 2735
rect 6586 2701 6596 2735
rect 6542 2617 6596 2701
rect 6626 2735 6680 2747
rect 6626 2701 6636 2735
rect 6670 2701 6680 2735
rect 6626 2667 6680 2701
rect 6626 2633 6636 2667
rect 6670 2633 6680 2667
rect 6626 2617 6680 2633
rect 6710 2735 6764 2747
rect 6710 2701 6720 2735
rect 6754 2701 6764 2735
rect 6710 2617 6764 2701
rect 6794 2735 6848 2747
rect 6794 2701 6804 2735
rect 6838 2701 6848 2735
rect 6794 2667 6848 2701
rect 6794 2633 6804 2667
rect 6838 2633 6848 2667
rect 6794 2617 6848 2633
rect 6878 2735 6932 2747
rect 6878 2701 6888 2735
rect 6922 2701 6932 2735
rect 6878 2617 6932 2701
rect 6962 2735 7016 2747
rect 6962 2701 6972 2735
rect 7006 2701 7016 2735
rect 6962 2667 7016 2701
rect 6962 2633 6972 2667
rect 7006 2633 7016 2667
rect 6962 2617 7016 2633
rect 7046 2735 7098 2747
rect 7046 2701 7056 2735
rect 7090 2701 7098 2735
rect 7046 2667 7098 2701
rect 7046 2633 7056 2667
rect 7090 2633 7098 2667
rect 7046 2617 7098 2633
rect 7586 2733 7638 2745
rect 7586 2699 7594 2733
rect 7628 2699 7638 2733
rect 7586 2665 7638 2699
rect 7586 2631 7594 2665
rect 7628 2631 7638 2665
rect 7586 2615 7638 2631
rect 7668 2733 7722 2745
rect 7668 2699 7678 2733
rect 7712 2699 7722 2733
rect 7668 2665 7722 2699
rect 7668 2631 7678 2665
rect 7712 2631 7722 2665
rect 7668 2615 7722 2631
rect 7752 2733 7806 2745
rect 7752 2699 7762 2733
rect 7796 2699 7806 2733
rect 7752 2615 7806 2699
rect 7836 2733 7890 2745
rect 7836 2699 7846 2733
rect 7880 2699 7890 2733
rect 7836 2665 7890 2699
rect 7836 2631 7846 2665
rect 7880 2631 7890 2665
rect 7836 2615 7890 2631
rect 7920 2733 7974 2745
rect 7920 2699 7930 2733
rect 7964 2699 7974 2733
rect 7920 2615 7974 2699
rect 8004 2733 8058 2745
rect 8004 2699 8014 2733
rect 8048 2699 8058 2733
rect 8004 2665 8058 2699
rect 8004 2631 8014 2665
rect 8048 2631 8058 2665
rect 8004 2615 8058 2631
rect 8088 2733 8142 2745
rect 8088 2699 8098 2733
rect 8132 2699 8142 2733
rect 8088 2615 8142 2699
rect 8172 2733 8226 2745
rect 8172 2699 8182 2733
rect 8216 2699 8226 2733
rect 8172 2665 8226 2699
rect 8172 2631 8182 2665
rect 8216 2631 8226 2665
rect 8172 2615 8226 2631
rect 8256 2733 8310 2745
rect 8256 2699 8266 2733
rect 8300 2699 8310 2733
rect 8256 2615 8310 2699
rect 8340 2733 8394 2745
rect 8340 2699 8350 2733
rect 8384 2699 8394 2733
rect 8340 2665 8394 2699
rect 8340 2631 8350 2665
rect 8384 2631 8394 2665
rect 8340 2615 8394 2631
rect 8424 2733 8478 2745
rect 8424 2699 8434 2733
rect 8468 2699 8478 2733
rect 8424 2615 8478 2699
rect 8508 2733 8562 2745
rect 8508 2699 8518 2733
rect 8552 2699 8562 2733
rect 8508 2665 8562 2699
rect 8508 2631 8518 2665
rect 8552 2631 8562 2665
rect 8508 2615 8562 2631
rect 8592 2733 8646 2745
rect 8592 2699 8602 2733
rect 8636 2699 8646 2733
rect 8592 2615 8646 2699
rect 8676 2733 8730 2745
rect 8676 2699 8686 2733
rect 8720 2699 8730 2733
rect 8676 2665 8730 2699
rect 8676 2631 8686 2665
rect 8720 2631 8730 2665
rect 8676 2615 8730 2631
rect 8760 2733 8814 2745
rect 8760 2699 8770 2733
rect 8804 2699 8814 2733
rect 8760 2615 8814 2699
rect 8844 2733 8898 2745
rect 8844 2699 8854 2733
rect 8888 2699 8898 2733
rect 8844 2665 8898 2699
rect 8844 2631 8854 2665
rect 8888 2631 8898 2665
rect 8844 2615 8898 2631
rect 8928 2733 8980 2745
rect 8928 2699 8938 2733
rect 8972 2699 8980 2733
rect 8928 2665 8980 2699
rect 8928 2631 8938 2665
rect 8972 2631 8980 2665
rect 8928 2615 8980 2631
rect 20802 2735 20854 2747
rect 20802 2701 20810 2735
rect 20844 2701 20854 2735
rect 20802 2667 20854 2701
rect 20802 2633 20810 2667
rect 20844 2633 20854 2667
rect 20802 2617 20854 2633
rect 20884 2735 20938 2747
rect 20884 2701 20894 2735
rect 20928 2701 20938 2735
rect 20884 2667 20938 2701
rect 20884 2633 20894 2667
rect 20928 2633 20938 2667
rect 20884 2617 20938 2633
rect 20968 2735 21022 2747
rect 20968 2701 20978 2735
rect 21012 2701 21022 2735
rect 20968 2617 21022 2701
rect 21052 2735 21106 2747
rect 21052 2701 21062 2735
rect 21096 2701 21106 2735
rect 21052 2667 21106 2701
rect 21052 2633 21062 2667
rect 21096 2633 21106 2667
rect 21052 2617 21106 2633
rect 21136 2735 21190 2747
rect 21136 2701 21146 2735
rect 21180 2701 21190 2735
rect 21136 2617 21190 2701
rect 21220 2735 21274 2747
rect 21220 2701 21230 2735
rect 21264 2701 21274 2735
rect 21220 2667 21274 2701
rect 21220 2633 21230 2667
rect 21264 2633 21274 2667
rect 21220 2617 21274 2633
rect 21304 2735 21358 2747
rect 21304 2701 21314 2735
rect 21348 2701 21358 2735
rect 21304 2617 21358 2701
rect 21388 2735 21442 2747
rect 21388 2701 21398 2735
rect 21432 2701 21442 2735
rect 21388 2667 21442 2701
rect 21388 2633 21398 2667
rect 21432 2633 21442 2667
rect 21388 2617 21442 2633
rect 21472 2735 21526 2747
rect 21472 2701 21482 2735
rect 21516 2701 21526 2735
rect 21472 2617 21526 2701
rect 21556 2735 21610 2747
rect 21556 2701 21566 2735
rect 21600 2701 21610 2735
rect 21556 2667 21610 2701
rect 21556 2633 21566 2667
rect 21600 2633 21610 2667
rect 21556 2617 21610 2633
rect 21640 2735 21694 2747
rect 21640 2701 21650 2735
rect 21684 2701 21694 2735
rect 21640 2617 21694 2701
rect 21724 2735 21778 2747
rect 21724 2701 21734 2735
rect 21768 2701 21778 2735
rect 21724 2667 21778 2701
rect 21724 2633 21734 2667
rect 21768 2633 21778 2667
rect 21724 2617 21778 2633
rect 21808 2735 21862 2747
rect 21808 2701 21818 2735
rect 21852 2701 21862 2735
rect 21808 2617 21862 2701
rect 21892 2735 21946 2747
rect 21892 2701 21902 2735
rect 21936 2701 21946 2735
rect 21892 2667 21946 2701
rect 21892 2633 21902 2667
rect 21936 2633 21946 2667
rect 21892 2617 21946 2633
rect 21976 2735 22030 2747
rect 21976 2701 21986 2735
rect 22020 2701 22030 2735
rect 21976 2617 22030 2701
rect 22060 2735 22114 2747
rect 22060 2701 22070 2735
rect 22104 2701 22114 2735
rect 22060 2667 22114 2701
rect 22060 2633 22070 2667
rect 22104 2633 22114 2667
rect 22060 2617 22114 2633
rect 22144 2735 22196 2747
rect 22144 2701 22154 2735
rect 22188 2701 22196 2735
rect 22144 2667 22196 2701
rect 22144 2633 22154 2667
rect 22188 2633 22196 2667
rect 22144 2617 22196 2633
rect 22684 2733 22736 2745
rect 22684 2699 22692 2733
rect 22726 2699 22736 2733
rect 22684 2665 22736 2699
rect 22684 2631 22692 2665
rect 22726 2631 22736 2665
rect 22684 2615 22736 2631
rect 22766 2733 22820 2745
rect 22766 2699 22776 2733
rect 22810 2699 22820 2733
rect 22766 2665 22820 2699
rect 22766 2631 22776 2665
rect 22810 2631 22820 2665
rect 22766 2615 22820 2631
rect 22850 2733 22904 2745
rect 22850 2699 22860 2733
rect 22894 2699 22904 2733
rect 22850 2615 22904 2699
rect 22934 2733 22988 2745
rect 22934 2699 22944 2733
rect 22978 2699 22988 2733
rect 22934 2665 22988 2699
rect 22934 2631 22944 2665
rect 22978 2631 22988 2665
rect 22934 2615 22988 2631
rect 23018 2733 23072 2745
rect 23018 2699 23028 2733
rect 23062 2699 23072 2733
rect 23018 2615 23072 2699
rect 23102 2733 23156 2745
rect 23102 2699 23112 2733
rect 23146 2699 23156 2733
rect 23102 2665 23156 2699
rect 23102 2631 23112 2665
rect 23146 2631 23156 2665
rect 23102 2615 23156 2631
rect 23186 2733 23240 2745
rect 23186 2699 23196 2733
rect 23230 2699 23240 2733
rect 23186 2615 23240 2699
rect 23270 2733 23324 2745
rect 23270 2699 23280 2733
rect 23314 2699 23324 2733
rect 23270 2665 23324 2699
rect 23270 2631 23280 2665
rect 23314 2631 23324 2665
rect 23270 2615 23324 2631
rect 23354 2733 23408 2745
rect 23354 2699 23364 2733
rect 23398 2699 23408 2733
rect 23354 2615 23408 2699
rect 23438 2733 23492 2745
rect 23438 2699 23448 2733
rect 23482 2699 23492 2733
rect 23438 2665 23492 2699
rect 23438 2631 23448 2665
rect 23482 2631 23492 2665
rect 23438 2615 23492 2631
rect 23522 2733 23576 2745
rect 23522 2699 23532 2733
rect 23566 2699 23576 2733
rect 23522 2615 23576 2699
rect 23606 2733 23660 2745
rect 23606 2699 23616 2733
rect 23650 2699 23660 2733
rect 23606 2665 23660 2699
rect 23606 2631 23616 2665
rect 23650 2631 23660 2665
rect 23606 2615 23660 2631
rect 23690 2733 23744 2745
rect 23690 2699 23700 2733
rect 23734 2699 23744 2733
rect 23690 2615 23744 2699
rect 23774 2733 23828 2745
rect 23774 2699 23784 2733
rect 23818 2699 23828 2733
rect 23774 2665 23828 2699
rect 23774 2631 23784 2665
rect 23818 2631 23828 2665
rect 23774 2615 23828 2631
rect 23858 2733 23912 2745
rect 23858 2699 23868 2733
rect 23902 2699 23912 2733
rect 23858 2615 23912 2699
rect 23942 2733 23996 2745
rect 23942 2699 23952 2733
rect 23986 2699 23996 2733
rect 23942 2665 23996 2699
rect 23942 2631 23952 2665
rect 23986 2631 23996 2665
rect 23942 2615 23996 2631
rect 24026 2733 24078 2745
rect 24026 2699 24036 2733
rect 24070 2699 24078 2733
rect 24026 2665 24078 2699
rect 24026 2631 24036 2665
rect 24070 2631 24078 2665
rect 24026 2615 24078 2631
rect 35906 2735 35958 2747
rect 35906 2701 35914 2735
rect 35948 2701 35958 2735
rect 35906 2667 35958 2701
rect 35906 2633 35914 2667
rect 35948 2633 35958 2667
rect 35906 2617 35958 2633
rect 35988 2735 36042 2747
rect 35988 2701 35998 2735
rect 36032 2701 36042 2735
rect 35988 2667 36042 2701
rect 35988 2633 35998 2667
rect 36032 2633 36042 2667
rect 35988 2617 36042 2633
rect 36072 2735 36126 2747
rect 36072 2701 36082 2735
rect 36116 2701 36126 2735
rect 36072 2617 36126 2701
rect 36156 2735 36210 2747
rect 36156 2701 36166 2735
rect 36200 2701 36210 2735
rect 36156 2667 36210 2701
rect 36156 2633 36166 2667
rect 36200 2633 36210 2667
rect 36156 2617 36210 2633
rect 36240 2735 36294 2747
rect 36240 2701 36250 2735
rect 36284 2701 36294 2735
rect 36240 2617 36294 2701
rect 36324 2735 36378 2747
rect 36324 2701 36334 2735
rect 36368 2701 36378 2735
rect 36324 2667 36378 2701
rect 36324 2633 36334 2667
rect 36368 2633 36378 2667
rect 36324 2617 36378 2633
rect 36408 2735 36462 2747
rect 36408 2701 36418 2735
rect 36452 2701 36462 2735
rect 36408 2617 36462 2701
rect 36492 2735 36546 2747
rect 36492 2701 36502 2735
rect 36536 2701 36546 2735
rect 36492 2667 36546 2701
rect 36492 2633 36502 2667
rect 36536 2633 36546 2667
rect 36492 2617 36546 2633
rect 36576 2735 36630 2747
rect 36576 2701 36586 2735
rect 36620 2701 36630 2735
rect 36576 2617 36630 2701
rect 36660 2735 36714 2747
rect 36660 2701 36670 2735
rect 36704 2701 36714 2735
rect 36660 2667 36714 2701
rect 36660 2633 36670 2667
rect 36704 2633 36714 2667
rect 36660 2617 36714 2633
rect 36744 2735 36798 2747
rect 36744 2701 36754 2735
rect 36788 2701 36798 2735
rect 36744 2617 36798 2701
rect 36828 2735 36882 2747
rect 36828 2701 36838 2735
rect 36872 2701 36882 2735
rect 36828 2667 36882 2701
rect 36828 2633 36838 2667
rect 36872 2633 36882 2667
rect 36828 2617 36882 2633
rect 36912 2735 36966 2747
rect 36912 2701 36922 2735
rect 36956 2701 36966 2735
rect 36912 2617 36966 2701
rect 36996 2735 37050 2747
rect 36996 2701 37006 2735
rect 37040 2701 37050 2735
rect 36996 2667 37050 2701
rect 36996 2633 37006 2667
rect 37040 2633 37050 2667
rect 36996 2617 37050 2633
rect 37080 2735 37134 2747
rect 37080 2701 37090 2735
rect 37124 2701 37134 2735
rect 37080 2617 37134 2701
rect 37164 2735 37218 2747
rect 37164 2701 37174 2735
rect 37208 2701 37218 2735
rect 37164 2667 37218 2701
rect 37164 2633 37174 2667
rect 37208 2633 37218 2667
rect 37164 2617 37218 2633
rect 37248 2735 37300 2747
rect 37248 2701 37258 2735
rect 37292 2701 37300 2735
rect 37248 2667 37300 2701
rect 37248 2633 37258 2667
rect 37292 2633 37300 2667
rect 37248 2617 37300 2633
rect 37788 2733 37840 2745
rect 37788 2699 37796 2733
rect 37830 2699 37840 2733
rect 37788 2665 37840 2699
rect 37788 2631 37796 2665
rect 37830 2631 37840 2665
rect 37788 2615 37840 2631
rect 37870 2733 37924 2745
rect 37870 2699 37880 2733
rect 37914 2699 37924 2733
rect 37870 2665 37924 2699
rect 37870 2631 37880 2665
rect 37914 2631 37924 2665
rect 37870 2615 37924 2631
rect 37954 2733 38008 2745
rect 37954 2699 37964 2733
rect 37998 2699 38008 2733
rect 37954 2615 38008 2699
rect 38038 2733 38092 2745
rect 38038 2699 38048 2733
rect 38082 2699 38092 2733
rect 38038 2665 38092 2699
rect 38038 2631 38048 2665
rect 38082 2631 38092 2665
rect 38038 2615 38092 2631
rect 38122 2733 38176 2745
rect 38122 2699 38132 2733
rect 38166 2699 38176 2733
rect 38122 2615 38176 2699
rect 38206 2733 38260 2745
rect 38206 2699 38216 2733
rect 38250 2699 38260 2733
rect 38206 2665 38260 2699
rect 38206 2631 38216 2665
rect 38250 2631 38260 2665
rect 38206 2615 38260 2631
rect 38290 2733 38344 2745
rect 38290 2699 38300 2733
rect 38334 2699 38344 2733
rect 38290 2615 38344 2699
rect 38374 2733 38428 2745
rect 38374 2699 38384 2733
rect 38418 2699 38428 2733
rect 38374 2665 38428 2699
rect 38374 2631 38384 2665
rect 38418 2631 38428 2665
rect 38374 2615 38428 2631
rect 38458 2733 38512 2745
rect 38458 2699 38468 2733
rect 38502 2699 38512 2733
rect 38458 2615 38512 2699
rect 38542 2733 38596 2745
rect 38542 2699 38552 2733
rect 38586 2699 38596 2733
rect 38542 2665 38596 2699
rect 38542 2631 38552 2665
rect 38586 2631 38596 2665
rect 38542 2615 38596 2631
rect 38626 2733 38680 2745
rect 38626 2699 38636 2733
rect 38670 2699 38680 2733
rect 38626 2615 38680 2699
rect 38710 2733 38764 2745
rect 38710 2699 38720 2733
rect 38754 2699 38764 2733
rect 38710 2665 38764 2699
rect 38710 2631 38720 2665
rect 38754 2631 38764 2665
rect 38710 2615 38764 2631
rect 38794 2733 38848 2745
rect 38794 2699 38804 2733
rect 38838 2699 38848 2733
rect 38794 2615 38848 2699
rect 38878 2733 38932 2745
rect 38878 2699 38888 2733
rect 38922 2699 38932 2733
rect 38878 2665 38932 2699
rect 38878 2631 38888 2665
rect 38922 2631 38932 2665
rect 38878 2615 38932 2631
rect 38962 2733 39016 2745
rect 38962 2699 38972 2733
rect 39006 2699 39016 2733
rect 38962 2615 39016 2699
rect 39046 2733 39100 2745
rect 39046 2699 39056 2733
rect 39090 2699 39100 2733
rect 39046 2665 39100 2699
rect 39046 2631 39056 2665
rect 39090 2631 39100 2665
rect 39046 2615 39100 2631
rect 39130 2733 39182 2745
rect 39130 2699 39140 2733
rect 39174 2699 39182 2733
rect 39130 2665 39182 2699
rect 39130 2631 39140 2665
rect 39174 2631 39182 2665
rect 39130 2615 39182 2631
rect 51004 2735 51056 2747
rect 51004 2701 51012 2735
rect 51046 2701 51056 2735
rect 51004 2667 51056 2701
rect 51004 2633 51012 2667
rect 51046 2633 51056 2667
rect 51004 2617 51056 2633
rect 51086 2735 51140 2747
rect 51086 2701 51096 2735
rect 51130 2701 51140 2735
rect 51086 2667 51140 2701
rect 51086 2633 51096 2667
rect 51130 2633 51140 2667
rect 51086 2617 51140 2633
rect 51170 2735 51224 2747
rect 51170 2701 51180 2735
rect 51214 2701 51224 2735
rect 51170 2617 51224 2701
rect 51254 2735 51308 2747
rect 51254 2701 51264 2735
rect 51298 2701 51308 2735
rect 51254 2667 51308 2701
rect 51254 2633 51264 2667
rect 51298 2633 51308 2667
rect 51254 2617 51308 2633
rect 51338 2735 51392 2747
rect 51338 2701 51348 2735
rect 51382 2701 51392 2735
rect 51338 2617 51392 2701
rect 51422 2735 51476 2747
rect 51422 2701 51432 2735
rect 51466 2701 51476 2735
rect 51422 2667 51476 2701
rect 51422 2633 51432 2667
rect 51466 2633 51476 2667
rect 51422 2617 51476 2633
rect 51506 2735 51560 2747
rect 51506 2701 51516 2735
rect 51550 2701 51560 2735
rect 51506 2617 51560 2701
rect 51590 2735 51644 2747
rect 51590 2701 51600 2735
rect 51634 2701 51644 2735
rect 51590 2667 51644 2701
rect 51590 2633 51600 2667
rect 51634 2633 51644 2667
rect 51590 2617 51644 2633
rect 51674 2735 51728 2747
rect 51674 2701 51684 2735
rect 51718 2701 51728 2735
rect 51674 2617 51728 2701
rect 51758 2735 51812 2747
rect 51758 2701 51768 2735
rect 51802 2701 51812 2735
rect 51758 2667 51812 2701
rect 51758 2633 51768 2667
rect 51802 2633 51812 2667
rect 51758 2617 51812 2633
rect 51842 2735 51896 2747
rect 51842 2701 51852 2735
rect 51886 2701 51896 2735
rect 51842 2617 51896 2701
rect 51926 2735 51980 2747
rect 51926 2701 51936 2735
rect 51970 2701 51980 2735
rect 51926 2667 51980 2701
rect 51926 2633 51936 2667
rect 51970 2633 51980 2667
rect 51926 2617 51980 2633
rect 52010 2735 52064 2747
rect 52010 2701 52020 2735
rect 52054 2701 52064 2735
rect 52010 2617 52064 2701
rect 52094 2735 52148 2747
rect 52094 2701 52104 2735
rect 52138 2701 52148 2735
rect 52094 2667 52148 2701
rect 52094 2633 52104 2667
rect 52138 2633 52148 2667
rect 52094 2617 52148 2633
rect 52178 2735 52232 2747
rect 52178 2701 52188 2735
rect 52222 2701 52232 2735
rect 52178 2617 52232 2701
rect 52262 2735 52316 2747
rect 52262 2701 52272 2735
rect 52306 2701 52316 2735
rect 52262 2667 52316 2701
rect 52262 2633 52272 2667
rect 52306 2633 52316 2667
rect 52262 2617 52316 2633
rect 52346 2735 52398 2747
rect 52346 2701 52356 2735
rect 52390 2701 52398 2735
rect 52346 2667 52398 2701
rect 52346 2633 52356 2667
rect 52390 2633 52398 2667
rect 52346 2617 52398 2633
rect 52886 2733 52938 2745
rect 52886 2699 52894 2733
rect 52928 2699 52938 2733
rect 52886 2665 52938 2699
rect 52886 2631 52894 2665
rect 52928 2631 52938 2665
rect 52886 2615 52938 2631
rect 52968 2733 53022 2745
rect 52968 2699 52978 2733
rect 53012 2699 53022 2733
rect 52968 2665 53022 2699
rect 52968 2631 52978 2665
rect 53012 2631 53022 2665
rect 52968 2615 53022 2631
rect 53052 2733 53106 2745
rect 53052 2699 53062 2733
rect 53096 2699 53106 2733
rect 53052 2615 53106 2699
rect 53136 2733 53190 2745
rect 53136 2699 53146 2733
rect 53180 2699 53190 2733
rect 53136 2665 53190 2699
rect 53136 2631 53146 2665
rect 53180 2631 53190 2665
rect 53136 2615 53190 2631
rect 53220 2733 53274 2745
rect 53220 2699 53230 2733
rect 53264 2699 53274 2733
rect 53220 2615 53274 2699
rect 53304 2733 53358 2745
rect 53304 2699 53314 2733
rect 53348 2699 53358 2733
rect 53304 2665 53358 2699
rect 53304 2631 53314 2665
rect 53348 2631 53358 2665
rect 53304 2615 53358 2631
rect 53388 2733 53442 2745
rect 53388 2699 53398 2733
rect 53432 2699 53442 2733
rect 53388 2615 53442 2699
rect 53472 2733 53526 2745
rect 53472 2699 53482 2733
rect 53516 2699 53526 2733
rect 53472 2665 53526 2699
rect 53472 2631 53482 2665
rect 53516 2631 53526 2665
rect 53472 2615 53526 2631
rect 53556 2733 53610 2745
rect 53556 2699 53566 2733
rect 53600 2699 53610 2733
rect 53556 2615 53610 2699
rect 53640 2733 53694 2745
rect 53640 2699 53650 2733
rect 53684 2699 53694 2733
rect 53640 2665 53694 2699
rect 53640 2631 53650 2665
rect 53684 2631 53694 2665
rect 53640 2615 53694 2631
rect 53724 2733 53778 2745
rect 53724 2699 53734 2733
rect 53768 2699 53778 2733
rect 53724 2615 53778 2699
rect 53808 2733 53862 2745
rect 53808 2699 53818 2733
rect 53852 2699 53862 2733
rect 53808 2665 53862 2699
rect 53808 2631 53818 2665
rect 53852 2631 53862 2665
rect 53808 2615 53862 2631
rect 53892 2733 53946 2745
rect 53892 2699 53902 2733
rect 53936 2699 53946 2733
rect 53892 2615 53946 2699
rect 53976 2733 54030 2745
rect 53976 2699 53986 2733
rect 54020 2699 54030 2733
rect 53976 2665 54030 2699
rect 53976 2631 53986 2665
rect 54020 2631 54030 2665
rect 53976 2615 54030 2631
rect 54060 2733 54114 2745
rect 54060 2699 54070 2733
rect 54104 2699 54114 2733
rect 54060 2615 54114 2699
rect 54144 2733 54198 2745
rect 54144 2699 54154 2733
rect 54188 2699 54198 2733
rect 54144 2665 54198 2699
rect 54144 2631 54154 2665
rect 54188 2631 54198 2665
rect 54144 2615 54198 2631
rect 54228 2733 54280 2745
rect 54228 2699 54238 2733
rect 54272 2699 54280 2733
rect 54228 2665 54280 2699
rect 54228 2631 54238 2665
rect 54272 2631 54280 2665
rect 54228 2615 54280 2631
rect 245 1789 297 1803
rect 245 1755 253 1789
rect 287 1755 297 1789
rect 245 1721 297 1755
rect 245 1687 253 1721
rect 287 1687 297 1721
rect 245 1673 297 1687
rect 327 1789 381 1803
rect 327 1755 337 1789
rect 371 1755 381 1789
rect 327 1721 381 1755
rect 327 1687 337 1721
rect 371 1687 381 1721
rect 327 1673 381 1687
rect 411 1789 463 1803
rect 411 1755 421 1789
rect 455 1755 463 1789
rect 1059 1789 1111 1803
rect 411 1721 463 1755
rect 1059 1755 1067 1789
rect 1101 1755 1111 1789
rect 411 1687 421 1721
rect 455 1687 463 1721
rect 411 1673 463 1687
rect 1059 1721 1111 1755
rect 1059 1687 1067 1721
rect 1101 1687 1111 1721
rect 1059 1673 1111 1687
rect 1141 1789 1195 1803
rect 1141 1755 1151 1789
rect 1185 1755 1195 1789
rect 1141 1721 1195 1755
rect 1141 1687 1151 1721
rect 1185 1687 1195 1721
rect 1141 1673 1195 1687
rect 1225 1789 1277 1803
rect 1225 1755 1235 1789
rect 1269 1755 1277 1789
rect 1225 1721 1277 1755
rect 1225 1687 1235 1721
rect 1269 1687 1277 1721
rect 1225 1673 1277 1687
rect 2133 1789 2185 1803
rect 2133 1755 2141 1789
rect 2175 1755 2185 1789
rect 2133 1721 2185 1755
rect 2133 1687 2141 1721
rect 2175 1687 2185 1721
rect 2133 1673 2185 1687
rect 2215 1789 2269 1803
rect 2215 1755 2225 1789
rect 2259 1755 2269 1789
rect 2215 1721 2269 1755
rect 2215 1687 2225 1721
rect 2259 1687 2269 1721
rect 2215 1673 2269 1687
rect 2299 1789 2351 1803
rect 2299 1755 2309 1789
rect 2343 1755 2351 1789
rect 2947 1789 2999 1803
rect 2299 1721 2351 1755
rect 2947 1755 2955 1789
rect 2989 1755 2999 1789
rect 2299 1687 2309 1721
rect 2343 1687 2351 1721
rect 2299 1673 2351 1687
rect 2947 1721 2999 1755
rect 2947 1687 2955 1721
rect 2989 1687 2999 1721
rect 2947 1673 2999 1687
rect 3029 1789 3083 1803
rect 3029 1755 3039 1789
rect 3073 1755 3083 1789
rect 3029 1721 3083 1755
rect 3029 1687 3039 1721
rect 3073 1687 3083 1721
rect 3029 1673 3083 1687
rect 3113 1789 3165 1803
rect 3113 1755 3123 1789
rect 3157 1755 3165 1789
rect 3113 1721 3165 1755
rect 3113 1687 3123 1721
rect 3157 1687 3165 1721
rect 3113 1673 3165 1687
rect 4021 1789 4073 1803
rect 4021 1755 4029 1789
rect 4063 1755 4073 1789
rect 4021 1721 4073 1755
rect 4021 1687 4029 1721
rect 4063 1687 4073 1721
rect 4021 1673 4073 1687
rect 4103 1789 4157 1803
rect 4103 1755 4113 1789
rect 4147 1755 4157 1789
rect 4103 1721 4157 1755
rect 4103 1687 4113 1721
rect 4147 1687 4157 1721
rect 4103 1673 4157 1687
rect 4187 1789 4239 1803
rect 4187 1755 4197 1789
rect 4231 1755 4239 1789
rect 4835 1789 4887 1803
rect 4187 1721 4239 1755
rect 4835 1755 4843 1789
rect 4877 1755 4887 1789
rect 4187 1687 4197 1721
rect 4231 1687 4239 1721
rect 4187 1673 4239 1687
rect 4835 1721 4887 1755
rect 4835 1687 4843 1721
rect 4877 1687 4887 1721
rect 4835 1673 4887 1687
rect 4917 1789 4971 1803
rect 4917 1755 4927 1789
rect 4961 1755 4971 1789
rect 4917 1721 4971 1755
rect 4917 1687 4927 1721
rect 4961 1687 4971 1721
rect 4917 1673 4971 1687
rect 5001 1789 5053 1803
rect 5001 1755 5011 1789
rect 5045 1755 5053 1789
rect 5001 1721 5053 1755
rect 5001 1687 5011 1721
rect 5045 1687 5053 1721
rect 5001 1673 5053 1687
rect 5909 1789 5961 1803
rect 5909 1755 5917 1789
rect 5951 1755 5961 1789
rect 5909 1721 5961 1755
rect 5909 1687 5917 1721
rect 5951 1687 5961 1721
rect 5909 1673 5961 1687
rect 5991 1789 6045 1803
rect 5991 1755 6001 1789
rect 6035 1755 6045 1789
rect 5991 1721 6045 1755
rect 5991 1687 6001 1721
rect 6035 1687 6045 1721
rect 5991 1673 6045 1687
rect 6075 1789 6127 1803
rect 6075 1755 6085 1789
rect 6119 1755 6127 1789
rect 6723 1789 6775 1803
rect 6075 1721 6127 1755
rect 6723 1755 6731 1789
rect 6765 1755 6775 1789
rect 6075 1687 6085 1721
rect 6119 1687 6127 1721
rect 6075 1673 6127 1687
rect 6723 1721 6775 1755
rect 6723 1687 6731 1721
rect 6765 1687 6775 1721
rect 6723 1673 6775 1687
rect 6805 1789 6859 1803
rect 6805 1755 6815 1789
rect 6849 1755 6859 1789
rect 6805 1721 6859 1755
rect 6805 1687 6815 1721
rect 6849 1687 6859 1721
rect 6805 1673 6859 1687
rect 6889 1789 6941 1803
rect 6889 1755 6899 1789
rect 6933 1755 6941 1789
rect 6889 1721 6941 1755
rect 6889 1687 6899 1721
rect 6933 1687 6941 1721
rect 6889 1673 6941 1687
rect 7797 1789 7849 1803
rect 7797 1755 7805 1789
rect 7839 1755 7849 1789
rect 7797 1721 7849 1755
rect 7797 1687 7805 1721
rect 7839 1687 7849 1721
rect 7797 1673 7849 1687
rect 7879 1789 7933 1803
rect 7879 1755 7889 1789
rect 7923 1755 7933 1789
rect 7879 1721 7933 1755
rect 7879 1687 7889 1721
rect 7923 1687 7933 1721
rect 7879 1673 7933 1687
rect 7963 1789 8015 1803
rect 7963 1755 7973 1789
rect 8007 1755 8015 1789
rect 8611 1789 8663 1803
rect 7963 1721 8015 1755
rect 8611 1755 8619 1789
rect 8653 1755 8663 1789
rect 7963 1687 7973 1721
rect 8007 1687 8015 1721
rect 7963 1673 8015 1687
rect 8611 1721 8663 1755
rect 8611 1687 8619 1721
rect 8653 1687 8663 1721
rect 8611 1673 8663 1687
rect 8693 1789 8747 1803
rect 8693 1755 8703 1789
rect 8737 1755 8747 1789
rect 8693 1721 8747 1755
rect 8693 1687 8703 1721
rect 8737 1687 8747 1721
rect 8693 1673 8747 1687
rect 8777 1789 8829 1803
rect 8777 1755 8787 1789
rect 8821 1755 8829 1789
rect 8777 1721 8829 1755
rect 8777 1687 8787 1721
rect 8821 1687 8829 1721
rect 8777 1673 8829 1687
rect 9685 1789 9737 1803
rect 9685 1755 9693 1789
rect 9727 1755 9737 1789
rect 9685 1721 9737 1755
rect 9685 1687 9693 1721
rect 9727 1687 9737 1721
rect 9685 1673 9737 1687
rect 9767 1789 9821 1803
rect 9767 1755 9777 1789
rect 9811 1755 9821 1789
rect 9767 1721 9821 1755
rect 9767 1687 9777 1721
rect 9811 1687 9821 1721
rect 9767 1673 9821 1687
rect 9851 1789 9903 1803
rect 9851 1755 9861 1789
rect 9895 1755 9903 1789
rect 10499 1789 10551 1803
rect 9851 1721 9903 1755
rect 10499 1755 10507 1789
rect 10541 1755 10551 1789
rect 9851 1687 9861 1721
rect 9895 1687 9903 1721
rect 9851 1673 9903 1687
rect 10499 1721 10551 1755
rect 10499 1687 10507 1721
rect 10541 1687 10551 1721
rect 10499 1673 10551 1687
rect 10581 1789 10635 1803
rect 10581 1755 10591 1789
rect 10625 1755 10635 1789
rect 10581 1721 10635 1755
rect 10581 1687 10591 1721
rect 10625 1687 10635 1721
rect 10581 1673 10635 1687
rect 10665 1789 10717 1803
rect 10665 1755 10675 1789
rect 10709 1755 10717 1789
rect 10665 1721 10717 1755
rect 10665 1687 10675 1721
rect 10709 1687 10717 1721
rect 10665 1673 10717 1687
rect 11573 1789 11625 1803
rect 11573 1755 11581 1789
rect 11615 1755 11625 1789
rect 11573 1721 11625 1755
rect 11573 1687 11581 1721
rect 11615 1687 11625 1721
rect 11573 1673 11625 1687
rect 11655 1789 11709 1803
rect 11655 1755 11665 1789
rect 11699 1755 11709 1789
rect 11655 1721 11709 1755
rect 11655 1687 11665 1721
rect 11699 1687 11709 1721
rect 11655 1673 11709 1687
rect 11739 1789 11791 1803
rect 11739 1755 11749 1789
rect 11783 1755 11791 1789
rect 12387 1789 12439 1803
rect 11739 1721 11791 1755
rect 12387 1755 12395 1789
rect 12429 1755 12439 1789
rect 11739 1687 11749 1721
rect 11783 1687 11791 1721
rect 11739 1673 11791 1687
rect 12387 1721 12439 1755
rect 12387 1687 12395 1721
rect 12429 1687 12439 1721
rect 12387 1673 12439 1687
rect 12469 1789 12523 1803
rect 12469 1755 12479 1789
rect 12513 1755 12523 1789
rect 12469 1721 12523 1755
rect 12469 1687 12479 1721
rect 12513 1687 12523 1721
rect 12469 1673 12523 1687
rect 12553 1789 12605 1803
rect 12553 1755 12563 1789
rect 12597 1755 12605 1789
rect 12553 1721 12605 1755
rect 12553 1687 12563 1721
rect 12597 1687 12605 1721
rect 12553 1673 12605 1687
rect 13461 1789 13513 1803
rect 13461 1755 13469 1789
rect 13503 1755 13513 1789
rect 13461 1721 13513 1755
rect 13461 1687 13469 1721
rect 13503 1687 13513 1721
rect 13461 1673 13513 1687
rect 13543 1789 13597 1803
rect 13543 1755 13553 1789
rect 13587 1755 13597 1789
rect 13543 1721 13597 1755
rect 13543 1687 13553 1721
rect 13587 1687 13597 1721
rect 13543 1673 13597 1687
rect 13627 1789 13679 1803
rect 13627 1755 13637 1789
rect 13671 1755 13679 1789
rect 14275 1789 14327 1803
rect 13627 1721 13679 1755
rect 14275 1755 14283 1789
rect 14317 1755 14327 1789
rect 13627 1687 13637 1721
rect 13671 1687 13679 1721
rect 13627 1673 13679 1687
rect 14275 1721 14327 1755
rect 14275 1687 14283 1721
rect 14317 1687 14327 1721
rect 14275 1673 14327 1687
rect 14357 1789 14411 1803
rect 14357 1755 14367 1789
rect 14401 1755 14411 1789
rect 14357 1721 14411 1755
rect 14357 1687 14367 1721
rect 14401 1687 14411 1721
rect 14357 1673 14411 1687
rect 14441 1789 14493 1803
rect 14441 1755 14451 1789
rect 14485 1755 14493 1789
rect 14441 1721 14493 1755
rect 14441 1687 14451 1721
rect 14485 1687 14493 1721
rect 14441 1673 14493 1687
rect 15343 1789 15395 1803
rect 15343 1755 15351 1789
rect 15385 1755 15395 1789
rect 15343 1721 15395 1755
rect 15343 1687 15351 1721
rect 15385 1687 15395 1721
rect 15343 1673 15395 1687
rect 15425 1789 15479 1803
rect 15425 1755 15435 1789
rect 15469 1755 15479 1789
rect 15425 1721 15479 1755
rect 15425 1687 15435 1721
rect 15469 1687 15479 1721
rect 15425 1673 15479 1687
rect 15509 1789 15561 1803
rect 15509 1755 15519 1789
rect 15553 1755 15561 1789
rect 16157 1789 16209 1803
rect 15509 1721 15561 1755
rect 16157 1755 16165 1789
rect 16199 1755 16209 1789
rect 15509 1687 15519 1721
rect 15553 1687 15561 1721
rect 15509 1673 15561 1687
rect 16157 1721 16209 1755
rect 16157 1687 16165 1721
rect 16199 1687 16209 1721
rect 16157 1673 16209 1687
rect 16239 1789 16293 1803
rect 16239 1755 16249 1789
rect 16283 1755 16293 1789
rect 16239 1721 16293 1755
rect 16239 1687 16249 1721
rect 16283 1687 16293 1721
rect 16239 1673 16293 1687
rect 16323 1789 16375 1803
rect 16323 1755 16333 1789
rect 16367 1755 16375 1789
rect 16323 1721 16375 1755
rect 16323 1687 16333 1721
rect 16367 1687 16375 1721
rect 16323 1673 16375 1687
rect 17231 1789 17283 1803
rect 17231 1755 17239 1789
rect 17273 1755 17283 1789
rect 17231 1721 17283 1755
rect 17231 1687 17239 1721
rect 17273 1687 17283 1721
rect 17231 1673 17283 1687
rect 17313 1789 17367 1803
rect 17313 1755 17323 1789
rect 17357 1755 17367 1789
rect 17313 1721 17367 1755
rect 17313 1687 17323 1721
rect 17357 1687 17367 1721
rect 17313 1673 17367 1687
rect 17397 1789 17449 1803
rect 17397 1755 17407 1789
rect 17441 1755 17449 1789
rect 18045 1789 18097 1803
rect 17397 1721 17449 1755
rect 18045 1755 18053 1789
rect 18087 1755 18097 1789
rect 17397 1687 17407 1721
rect 17441 1687 17449 1721
rect 17397 1673 17449 1687
rect 18045 1721 18097 1755
rect 18045 1687 18053 1721
rect 18087 1687 18097 1721
rect 18045 1673 18097 1687
rect 18127 1789 18181 1803
rect 18127 1755 18137 1789
rect 18171 1755 18181 1789
rect 18127 1721 18181 1755
rect 18127 1687 18137 1721
rect 18171 1687 18181 1721
rect 18127 1673 18181 1687
rect 18211 1789 18263 1803
rect 18211 1755 18221 1789
rect 18255 1755 18263 1789
rect 18211 1721 18263 1755
rect 18211 1687 18221 1721
rect 18255 1687 18263 1721
rect 18211 1673 18263 1687
rect 19119 1789 19171 1803
rect 19119 1755 19127 1789
rect 19161 1755 19171 1789
rect 19119 1721 19171 1755
rect 19119 1687 19127 1721
rect 19161 1687 19171 1721
rect 19119 1673 19171 1687
rect 19201 1789 19255 1803
rect 19201 1755 19211 1789
rect 19245 1755 19255 1789
rect 19201 1721 19255 1755
rect 19201 1687 19211 1721
rect 19245 1687 19255 1721
rect 19201 1673 19255 1687
rect 19285 1789 19337 1803
rect 19285 1755 19295 1789
rect 19329 1755 19337 1789
rect 19933 1789 19985 1803
rect 19285 1721 19337 1755
rect 19933 1755 19941 1789
rect 19975 1755 19985 1789
rect 19285 1687 19295 1721
rect 19329 1687 19337 1721
rect 19285 1673 19337 1687
rect 19933 1721 19985 1755
rect 19933 1687 19941 1721
rect 19975 1687 19985 1721
rect 19933 1673 19985 1687
rect 20015 1789 20069 1803
rect 20015 1755 20025 1789
rect 20059 1755 20069 1789
rect 20015 1721 20069 1755
rect 20015 1687 20025 1721
rect 20059 1687 20069 1721
rect 20015 1673 20069 1687
rect 20099 1789 20151 1803
rect 20099 1755 20109 1789
rect 20143 1755 20151 1789
rect 20099 1721 20151 1755
rect 20099 1687 20109 1721
rect 20143 1687 20151 1721
rect 20099 1673 20151 1687
rect 21007 1789 21059 1803
rect 21007 1755 21015 1789
rect 21049 1755 21059 1789
rect 21007 1721 21059 1755
rect 21007 1687 21015 1721
rect 21049 1687 21059 1721
rect 21007 1673 21059 1687
rect 21089 1789 21143 1803
rect 21089 1755 21099 1789
rect 21133 1755 21143 1789
rect 21089 1721 21143 1755
rect 21089 1687 21099 1721
rect 21133 1687 21143 1721
rect 21089 1673 21143 1687
rect 21173 1789 21225 1803
rect 21173 1755 21183 1789
rect 21217 1755 21225 1789
rect 21821 1789 21873 1803
rect 21173 1721 21225 1755
rect 21821 1755 21829 1789
rect 21863 1755 21873 1789
rect 21173 1687 21183 1721
rect 21217 1687 21225 1721
rect 21173 1673 21225 1687
rect 21821 1721 21873 1755
rect 21821 1687 21829 1721
rect 21863 1687 21873 1721
rect 21821 1673 21873 1687
rect 21903 1789 21957 1803
rect 21903 1755 21913 1789
rect 21947 1755 21957 1789
rect 21903 1721 21957 1755
rect 21903 1687 21913 1721
rect 21947 1687 21957 1721
rect 21903 1673 21957 1687
rect 21987 1789 22039 1803
rect 21987 1755 21997 1789
rect 22031 1755 22039 1789
rect 21987 1721 22039 1755
rect 21987 1687 21997 1721
rect 22031 1687 22039 1721
rect 21987 1673 22039 1687
rect 22895 1789 22947 1803
rect 22895 1755 22903 1789
rect 22937 1755 22947 1789
rect 22895 1721 22947 1755
rect 22895 1687 22903 1721
rect 22937 1687 22947 1721
rect 22895 1673 22947 1687
rect 22977 1789 23031 1803
rect 22977 1755 22987 1789
rect 23021 1755 23031 1789
rect 22977 1721 23031 1755
rect 22977 1687 22987 1721
rect 23021 1687 23031 1721
rect 22977 1673 23031 1687
rect 23061 1789 23113 1803
rect 23061 1755 23071 1789
rect 23105 1755 23113 1789
rect 23709 1789 23761 1803
rect 23061 1721 23113 1755
rect 23709 1755 23717 1789
rect 23751 1755 23761 1789
rect 23061 1687 23071 1721
rect 23105 1687 23113 1721
rect 23061 1673 23113 1687
rect 23709 1721 23761 1755
rect 23709 1687 23717 1721
rect 23751 1687 23761 1721
rect 23709 1673 23761 1687
rect 23791 1789 23845 1803
rect 23791 1755 23801 1789
rect 23835 1755 23845 1789
rect 23791 1721 23845 1755
rect 23791 1687 23801 1721
rect 23835 1687 23845 1721
rect 23791 1673 23845 1687
rect 23875 1789 23927 1803
rect 23875 1755 23885 1789
rect 23919 1755 23927 1789
rect 23875 1721 23927 1755
rect 23875 1687 23885 1721
rect 23919 1687 23927 1721
rect 23875 1673 23927 1687
rect 24783 1789 24835 1803
rect 24783 1755 24791 1789
rect 24825 1755 24835 1789
rect 24783 1721 24835 1755
rect 24783 1687 24791 1721
rect 24825 1687 24835 1721
rect 24783 1673 24835 1687
rect 24865 1789 24919 1803
rect 24865 1755 24875 1789
rect 24909 1755 24919 1789
rect 24865 1721 24919 1755
rect 24865 1687 24875 1721
rect 24909 1687 24919 1721
rect 24865 1673 24919 1687
rect 24949 1789 25001 1803
rect 24949 1755 24959 1789
rect 24993 1755 25001 1789
rect 25597 1789 25649 1803
rect 24949 1721 25001 1755
rect 25597 1755 25605 1789
rect 25639 1755 25649 1789
rect 24949 1687 24959 1721
rect 24993 1687 25001 1721
rect 24949 1673 25001 1687
rect 25597 1721 25649 1755
rect 25597 1687 25605 1721
rect 25639 1687 25649 1721
rect 25597 1673 25649 1687
rect 25679 1789 25733 1803
rect 25679 1755 25689 1789
rect 25723 1755 25733 1789
rect 25679 1721 25733 1755
rect 25679 1687 25689 1721
rect 25723 1687 25733 1721
rect 25679 1673 25733 1687
rect 25763 1789 25815 1803
rect 25763 1755 25773 1789
rect 25807 1755 25815 1789
rect 25763 1721 25815 1755
rect 25763 1687 25773 1721
rect 25807 1687 25815 1721
rect 25763 1673 25815 1687
rect 26671 1789 26723 1803
rect 26671 1755 26679 1789
rect 26713 1755 26723 1789
rect 26671 1721 26723 1755
rect 26671 1687 26679 1721
rect 26713 1687 26723 1721
rect 26671 1673 26723 1687
rect 26753 1789 26807 1803
rect 26753 1755 26763 1789
rect 26797 1755 26807 1789
rect 26753 1721 26807 1755
rect 26753 1687 26763 1721
rect 26797 1687 26807 1721
rect 26753 1673 26807 1687
rect 26837 1789 26889 1803
rect 26837 1755 26847 1789
rect 26881 1755 26889 1789
rect 27485 1789 27537 1803
rect 26837 1721 26889 1755
rect 27485 1755 27493 1789
rect 27527 1755 27537 1789
rect 26837 1687 26847 1721
rect 26881 1687 26889 1721
rect 26837 1673 26889 1687
rect 27485 1721 27537 1755
rect 27485 1687 27493 1721
rect 27527 1687 27537 1721
rect 27485 1673 27537 1687
rect 27567 1789 27621 1803
rect 27567 1755 27577 1789
rect 27611 1755 27621 1789
rect 27567 1721 27621 1755
rect 27567 1687 27577 1721
rect 27611 1687 27621 1721
rect 27567 1673 27621 1687
rect 27651 1789 27703 1803
rect 27651 1755 27661 1789
rect 27695 1755 27703 1789
rect 27651 1721 27703 1755
rect 27651 1687 27661 1721
rect 27695 1687 27703 1721
rect 27651 1673 27703 1687
rect 28559 1789 28611 1803
rect 28559 1755 28567 1789
rect 28601 1755 28611 1789
rect 28559 1721 28611 1755
rect 28559 1687 28567 1721
rect 28601 1687 28611 1721
rect 28559 1673 28611 1687
rect 28641 1789 28695 1803
rect 28641 1755 28651 1789
rect 28685 1755 28695 1789
rect 28641 1721 28695 1755
rect 28641 1687 28651 1721
rect 28685 1687 28695 1721
rect 28641 1673 28695 1687
rect 28725 1789 28777 1803
rect 28725 1755 28735 1789
rect 28769 1755 28777 1789
rect 29373 1789 29425 1803
rect 28725 1721 28777 1755
rect 29373 1755 29381 1789
rect 29415 1755 29425 1789
rect 28725 1687 28735 1721
rect 28769 1687 28777 1721
rect 28725 1673 28777 1687
rect 29373 1721 29425 1755
rect 29373 1687 29381 1721
rect 29415 1687 29425 1721
rect 29373 1673 29425 1687
rect 29455 1789 29509 1803
rect 29455 1755 29465 1789
rect 29499 1755 29509 1789
rect 29455 1721 29509 1755
rect 29455 1687 29465 1721
rect 29499 1687 29509 1721
rect 29455 1673 29509 1687
rect 29539 1789 29591 1803
rect 29539 1755 29549 1789
rect 29583 1755 29591 1789
rect 29539 1721 29591 1755
rect 29539 1687 29549 1721
rect 29583 1687 29591 1721
rect 29539 1673 29591 1687
rect 30447 1789 30499 1803
rect 30447 1755 30455 1789
rect 30489 1755 30499 1789
rect 30447 1721 30499 1755
rect 30447 1687 30455 1721
rect 30489 1687 30499 1721
rect 30447 1673 30499 1687
rect 30529 1789 30583 1803
rect 30529 1755 30539 1789
rect 30573 1755 30583 1789
rect 30529 1721 30583 1755
rect 30529 1687 30539 1721
rect 30573 1687 30583 1721
rect 30529 1673 30583 1687
rect 30613 1789 30665 1803
rect 30613 1755 30623 1789
rect 30657 1755 30665 1789
rect 31261 1789 31313 1803
rect 30613 1721 30665 1755
rect 31261 1755 31269 1789
rect 31303 1755 31313 1789
rect 30613 1687 30623 1721
rect 30657 1687 30665 1721
rect 30613 1673 30665 1687
rect 31261 1721 31313 1755
rect 31261 1687 31269 1721
rect 31303 1687 31313 1721
rect 31261 1673 31313 1687
rect 31343 1789 31397 1803
rect 31343 1755 31353 1789
rect 31387 1755 31397 1789
rect 31343 1721 31397 1755
rect 31343 1687 31353 1721
rect 31387 1687 31397 1721
rect 31343 1673 31397 1687
rect 31427 1789 31479 1803
rect 31427 1755 31437 1789
rect 31471 1755 31479 1789
rect 31427 1721 31479 1755
rect 31427 1687 31437 1721
rect 31471 1687 31479 1721
rect 31427 1673 31479 1687
rect 32335 1789 32387 1803
rect 32335 1755 32343 1789
rect 32377 1755 32387 1789
rect 32335 1721 32387 1755
rect 32335 1687 32343 1721
rect 32377 1687 32387 1721
rect 32335 1673 32387 1687
rect 32417 1789 32471 1803
rect 32417 1755 32427 1789
rect 32461 1755 32471 1789
rect 32417 1721 32471 1755
rect 32417 1687 32427 1721
rect 32461 1687 32471 1721
rect 32417 1673 32471 1687
rect 32501 1789 32553 1803
rect 32501 1755 32511 1789
rect 32545 1755 32553 1789
rect 33149 1789 33201 1803
rect 32501 1721 32553 1755
rect 33149 1755 33157 1789
rect 33191 1755 33201 1789
rect 32501 1687 32511 1721
rect 32545 1687 32553 1721
rect 32501 1673 32553 1687
rect 33149 1721 33201 1755
rect 33149 1687 33157 1721
rect 33191 1687 33201 1721
rect 33149 1673 33201 1687
rect 33231 1789 33285 1803
rect 33231 1755 33241 1789
rect 33275 1755 33285 1789
rect 33231 1721 33285 1755
rect 33231 1687 33241 1721
rect 33275 1687 33285 1721
rect 33231 1673 33285 1687
rect 33315 1789 33367 1803
rect 33315 1755 33325 1789
rect 33359 1755 33367 1789
rect 33315 1721 33367 1755
rect 33315 1687 33325 1721
rect 33359 1687 33367 1721
rect 33315 1673 33367 1687
rect 34223 1789 34275 1803
rect 34223 1755 34231 1789
rect 34265 1755 34275 1789
rect 34223 1721 34275 1755
rect 34223 1687 34231 1721
rect 34265 1687 34275 1721
rect 34223 1673 34275 1687
rect 34305 1789 34359 1803
rect 34305 1755 34315 1789
rect 34349 1755 34359 1789
rect 34305 1721 34359 1755
rect 34305 1687 34315 1721
rect 34349 1687 34359 1721
rect 34305 1673 34359 1687
rect 34389 1789 34441 1803
rect 34389 1755 34399 1789
rect 34433 1755 34441 1789
rect 35037 1789 35089 1803
rect 34389 1721 34441 1755
rect 35037 1755 35045 1789
rect 35079 1755 35089 1789
rect 34389 1687 34399 1721
rect 34433 1687 34441 1721
rect 34389 1673 34441 1687
rect 35037 1721 35089 1755
rect 35037 1687 35045 1721
rect 35079 1687 35089 1721
rect 35037 1673 35089 1687
rect 35119 1789 35173 1803
rect 35119 1755 35129 1789
rect 35163 1755 35173 1789
rect 35119 1721 35173 1755
rect 35119 1687 35129 1721
rect 35163 1687 35173 1721
rect 35119 1673 35173 1687
rect 35203 1789 35255 1803
rect 35203 1755 35213 1789
rect 35247 1755 35255 1789
rect 35203 1721 35255 1755
rect 35203 1687 35213 1721
rect 35247 1687 35255 1721
rect 35203 1673 35255 1687
rect 36111 1789 36163 1803
rect 36111 1755 36119 1789
rect 36153 1755 36163 1789
rect 36111 1721 36163 1755
rect 36111 1687 36119 1721
rect 36153 1687 36163 1721
rect 36111 1673 36163 1687
rect 36193 1789 36247 1803
rect 36193 1755 36203 1789
rect 36237 1755 36247 1789
rect 36193 1721 36247 1755
rect 36193 1687 36203 1721
rect 36237 1687 36247 1721
rect 36193 1673 36247 1687
rect 36277 1789 36329 1803
rect 36277 1755 36287 1789
rect 36321 1755 36329 1789
rect 36925 1789 36977 1803
rect 36277 1721 36329 1755
rect 36925 1755 36933 1789
rect 36967 1755 36977 1789
rect 36277 1687 36287 1721
rect 36321 1687 36329 1721
rect 36277 1673 36329 1687
rect 36925 1721 36977 1755
rect 36925 1687 36933 1721
rect 36967 1687 36977 1721
rect 36925 1673 36977 1687
rect 37007 1789 37061 1803
rect 37007 1755 37017 1789
rect 37051 1755 37061 1789
rect 37007 1721 37061 1755
rect 37007 1687 37017 1721
rect 37051 1687 37061 1721
rect 37007 1673 37061 1687
rect 37091 1789 37143 1803
rect 37091 1755 37101 1789
rect 37135 1755 37143 1789
rect 37091 1721 37143 1755
rect 37091 1687 37101 1721
rect 37135 1687 37143 1721
rect 37091 1673 37143 1687
rect 37999 1789 38051 1803
rect 37999 1755 38007 1789
rect 38041 1755 38051 1789
rect 37999 1721 38051 1755
rect 37999 1687 38007 1721
rect 38041 1687 38051 1721
rect 37999 1673 38051 1687
rect 38081 1789 38135 1803
rect 38081 1755 38091 1789
rect 38125 1755 38135 1789
rect 38081 1721 38135 1755
rect 38081 1687 38091 1721
rect 38125 1687 38135 1721
rect 38081 1673 38135 1687
rect 38165 1789 38217 1803
rect 38165 1755 38175 1789
rect 38209 1755 38217 1789
rect 38813 1789 38865 1803
rect 38165 1721 38217 1755
rect 38813 1755 38821 1789
rect 38855 1755 38865 1789
rect 38165 1687 38175 1721
rect 38209 1687 38217 1721
rect 38165 1673 38217 1687
rect 38813 1721 38865 1755
rect 38813 1687 38821 1721
rect 38855 1687 38865 1721
rect 38813 1673 38865 1687
rect 38895 1789 38949 1803
rect 38895 1755 38905 1789
rect 38939 1755 38949 1789
rect 38895 1721 38949 1755
rect 38895 1687 38905 1721
rect 38939 1687 38949 1721
rect 38895 1673 38949 1687
rect 38979 1789 39031 1803
rect 38979 1755 38989 1789
rect 39023 1755 39031 1789
rect 38979 1721 39031 1755
rect 38979 1687 38989 1721
rect 39023 1687 39031 1721
rect 38979 1673 39031 1687
rect 39887 1789 39939 1803
rect 39887 1755 39895 1789
rect 39929 1755 39939 1789
rect 39887 1721 39939 1755
rect 39887 1687 39895 1721
rect 39929 1687 39939 1721
rect 39887 1673 39939 1687
rect 39969 1789 40023 1803
rect 39969 1755 39979 1789
rect 40013 1755 40023 1789
rect 39969 1721 40023 1755
rect 39969 1687 39979 1721
rect 40013 1687 40023 1721
rect 39969 1673 40023 1687
rect 40053 1789 40105 1803
rect 40053 1755 40063 1789
rect 40097 1755 40105 1789
rect 40701 1789 40753 1803
rect 40053 1721 40105 1755
rect 40701 1755 40709 1789
rect 40743 1755 40753 1789
rect 40053 1687 40063 1721
rect 40097 1687 40105 1721
rect 40053 1673 40105 1687
rect 40701 1721 40753 1755
rect 40701 1687 40709 1721
rect 40743 1687 40753 1721
rect 40701 1673 40753 1687
rect 40783 1789 40837 1803
rect 40783 1755 40793 1789
rect 40827 1755 40837 1789
rect 40783 1721 40837 1755
rect 40783 1687 40793 1721
rect 40827 1687 40837 1721
rect 40783 1673 40837 1687
rect 40867 1789 40919 1803
rect 40867 1755 40877 1789
rect 40911 1755 40919 1789
rect 40867 1721 40919 1755
rect 40867 1687 40877 1721
rect 40911 1687 40919 1721
rect 40867 1673 40919 1687
rect 41775 1789 41827 1803
rect 41775 1755 41783 1789
rect 41817 1755 41827 1789
rect 41775 1721 41827 1755
rect 41775 1687 41783 1721
rect 41817 1687 41827 1721
rect 41775 1673 41827 1687
rect 41857 1789 41911 1803
rect 41857 1755 41867 1789
rect 41901 1755 41911 1789
rect 41857 1721 41911 1755
rect 41857 1687 41867 1721
rect 41901 1687 41911 1721
rect 41857 1673 41911 1687
rect 41941 1789 41993 1803
rect 41941 1755 41951 1789
rect 41985 1755 41993 1789
rect 42589 1789 42641 1803
rect 41941 1721 41993 1755
rect 42589 1755 42597 1789
rect 42631 1755 42641 1789
rect 41941 1687 41951 1721
rect 41985 1687 41993 1721
rect 41941 1673 41993 1687
rect 42589 1721 42641 1755
rect 42589 1687 42597 1721
rect 42631 1687 42641 1721
rect 42589 1673 42641 1687
rect 42671 1789 42725 1803
rect 42671 1755 42681 1789
rect 42715 1755 42725 1789
rect 42671 1721 42725 1755
rect 42671 1687 42681 1721
rect 42715 1687 42725 1721
rect 42671 1673 42725 1687
rect 42755 1789 42807 1803
rect 42755 1755 42765 1789
rect 42799 1755 42807 1789
rect 42755 1721 42807 1755
rect 42755 1687 42765 1721
rect 42799 1687 42807 1721
rect 42755 1673 42807 1687
rect 43663 1789 43715 1803
rect 43663 1755 43671 1789
rect 43705 1755 43715 1789
rect 43663 1721 43715 1755
rect 43663 1687 43671 1721
rect 43705 1687 43715 1721
rect 43663 1673 43715 1687
rect 43745 1789 43799 1803
rect 43745 1755 43755 1789
rect 43789 1755 43799 1789
rect 43745 1721 43799 1755
rect 43745 1687 43755 1721
rect 43789 1687 43799 1721
rect 43745 1673 43799 1687
rect 43829 1789 43881 1803
rect 43829 1755 43839 1789
rect 43873 1755 43881 1789
rect 44477 1789 44529 1803
rect 43829 1721 43881 1755
rect 44477 1755 44485 1789
rect 44519 1755 44529 1789
rect 43829 1687 43839 1721
rect 43873 1687 43881 1721
rect 43829 1673 43881 1687
rect 44477 1721 44529 1755
rect 44477 1687 44485 1721
rect 44519 1687 44529 1721
rect 44477 1673 44529 1687
rect 44559 1789 44613 1803
rect 44559 1755 44569 1789
rect 44603 1755 44613 1789
rect 44559 1721 44613 1755
rect 44559 1687 44569 1721
rect 44603 1687 44613 1721
rect 44559 1673 44613 1687
rect 44643 1789 44695 1803
rect 44643 1755 44653 1789
rect 44687 1755 44695 1789
rect 44643 1721 44695 1755
rect 44643 1687 44653 1721
rect 44687 1687 44695 1721
rect 44643 1673 44695 1687
rect 45545 1789 45597 1803
rect 45545 1755 45553 1789
rect 45587 1755 45597 1789
rect 45545 1721 45597 1755
rect 45545 1687 45553 1721
rect 45587 1687 45597 1721
rect 45545 1673 45597 1687
rect 45627 1789 45681 1803
rect 45627 1755 45637 1789
rect 45671 1755 45681 1789
rect 45627 1721 45681 1755
rect 45627 1687 45637 1721
rect 45671 1687 45681 1721
rect 45627 1673 45681 1687
rect 45711 1789 45763 1803
rect 45711 1755 45721 1789
rect 45755 1755 45763 1789
rect 46359 1789 46411 1803
rect 45711 1721 45763 1755
rect 46359 1755 46367 1789
rect 46401 1755 46411 1789
rect 45711 1687 45721 1721
rect 45755 1687 45763 1721
rect 45711 1673 45763 1687
rect 46359 1721 46411 1755
rect 46359 1687 46367 1721
rect 46401 1687 46411 1721
rect 46359 1673 46411 1687
rect 46441 1789 46495 1803
rect 46441 1755 46451 1789
rect 46485 1755 46495 1789
rect 46441 1721 46495 1755
rect 46441 1687 46451 1721
rect 46485 1687 46495 1721
rect 46441 1673 46495 1687
rect 46525 1789 46577 1803
rect 46525 1755 46535 1789
rect 46569 1755 46577 1789
rect 46525 1721 46577 1755
rect 46525 1687 46535 1721
rect 46569 1687 46577 1721
rect 46525 1673 46577 1687
rect 47433 1789 47485 1803
rect 47433 1755 47441 1789
rect 47475 1755 47485 1789
rect 47433 1721 47485 1755
rect 47433 1687 47441 1721
rect 47475 1687 47485 1721
rect 47433 1673 47485 1687
rect 47515 1789 47569 1803
rect 47515 1755 47525 1789
rect 47559 1755 47569 1789
rect 47515 1721 47569 1755
rect 47515 1687 47525 1721
rect 47559 1687 47569 1721
rect 47515 1673 47569 1687
rect 47599 1789 47651 1803
rect 47599 1755 47609 1789
rect 47643 1755 47651 1789
rect 48247 1789 48299 1803
rect 47599 1721 47651 1755
rect 48247 1755 48255 1789
rect 48289 1755 48299 1789
rect 47599 1687 47609 1721
rect 47643 1687 47651 1721
rect 47599 1673 47651 1687
rect 48247 1721 48299 1755
rect 48247 1687 48255 1721
rect 48289 1687 48299 1721
rect 48247 1673 48299 1687
rect 48329 1789 48383 1803
rect 48329 1755 48339 1789
rect 48373 1755 48383 1789
rect 48329 1721 48383 1755
rect 48329 1687 48339 1721
rect 48373 1687 48383 1721
rect 48329 1673 48383 1687
rect 48413 1789 48465 1803
rect 48413 1755 48423 1789
rect 48457 1755 48465 1789
rect 48413 1721 48465 1755
rect 48413 1687 48423 1721
rect 48457 1687 48465 1721
rect 48413 1673 48465 1687
rect 49321 1789 49373 1803
rect 49321 1755 49329 1789
rect 49363 1755 49373 1789
rect 49321 1721 49373 1755
rect 49321 1687 49329 1721
rect 49363 1687 49373 1721
rect 49321 1673 49373 1687
rect 49403 1789 49457 1803
rect 49403 1755 49413 1789
rect 49447 1755 49457 1789
rect 49403 1721 49457 1755
rect 49403 1687 49413 1721
rect 49447 1687 49457 1721
rect 49403 1673 49457 1687
rect 49487 1789 49539 1803
rect 49487 1755 49497 1789
rect 49531 1755 49539 1789
rect 50135 1789 50187 1803
rect 49487 1721 49539 1755
rect 50135 1755 50143 1789
rect 50177 1755 50187 1789
rect 49487 1687 49497 1721
rect 49531 1687 49539 1721
rect 49487 1673 49539 1687
rect 50135 1721 50187 1755
rect 50135 1687 50143 1721
rect 50177 1687 50187 1721
rect 50135 1673 50187 1687
rect 50217 1789 50271 1803
rect 50217 1755 50227 1789
rect 50261 1755 50271 1789
rect 50217 1721 50271 1755
rect 50217 1687 50227 1721
rect 50261 1687 50271 1721
rect 50217 1673 50271 1687
rect 50301 1789 50353 1803
rect 50301 1755 50311 1789
rect 50345 1755 50353 1789
rect 50301 1721 50353 1755
rect 50301 1687 50311 1721
rect 50345 1687 50353 1721
rect 50301 1673 50353 1687
rect 51209 1789 51261 1803
rect 51209 1755 51217 1789
rect 51251 1755 51261 1789
rect 51209 1721 51261 1755
rect 51209 1687 51217 1721
rect 51251 1687 51261 1721
rect 51209 1673 51261 1687
rect 51291 1789 51345 1803
rect 51291 1755 51301 1789
rect 51335 1755 51345 1789
rect 51291 1721 51345 1755
rect 51291 1687 51301 1721
rect 51335 1687 51345 1721
rect 51291 1673 51345 1687
rect 51375 1789 51427 1803
rect 51375 1755 51385 1789
rect 51419 1755 51427 1789
rect 52023 1789 52075 1803
rect 51375 1721 51427 1755
rect 52023 1755 52031 1789
rect 52065 1755 52075 1789
rect 51375 1687 51385 1721
rect 51419 1687 51427 1721
rect 51375 1673 51427 1687
rect 52023 1721 52075 1755
rect 52023 1687 52031 1721
rect 52065 1687 52075 1721
rect 52023 1673 52075 1687
rect 52105 1789 52159 1803
rect 52105 1755 52115 1789
rect 52149 1755 52159 1789
rect 52105 1721 52159 1755
rect 52105 1687 52115 1721
rect 52149 1687 52159 1721
rect 52105 1673 52159 1687
rect 52189 1789 52241 1803
rect 52189 1755 52199 1789
rect 52233 1755 52241 1789
rect 52189 1721 52241 1755
rect 52189 1687 52199 1721
rect 52233 1687 52241 1721
rect 52189 1673 52241 1687
rect 53097 1789 53149 1803
rect 53097 1755 53105 1789
rect 53139 1755 53149 1789
rect 53097 1721 53149 1755
rect 53097 1687 53105 1721
rect 53139 1687 53149 1721
rect 53097 1673 53149 1687
rect 53179 1789 53233 1803
rect 53179 1755 53189 1789
rect 53223 1755 53233 1789
rect 53179 1721 53233 1755
rect 53179 1687 53189 1721
rect 53223 1687 53233 1721
rect 53179 1673 53233 1687
rect 53263 1789 53315 1803
rect 53263 1755 53273 1789
rect 53307 1755 53315 1789
rect 53911 1789 53963 1803
rect 53263 1721 53315 1755
rect 53911 1755 53919 1789
rect 53953 1755 53963 1789
rect 53263 1687 53273 1721
rect 53307 1687 53315 1721
rect 53263 1673 53315 1687
rect 53911 1721 53963 1755
rect 53911 1687 53919 1721
rect 53953 1687 53963 1721
rect 53911 1673 53963 1687
rect 53993 1789 54047 1803
rect 53993 1755 54003 1789
rect 54037 1755 54047 1789
rect 53993 1721 54047 1755
rect 53993 1687 54003 1721
rect 54037 1687 54047 1721
rect 53993 1673 54047 1687
rect 54077 1789 54129 1803
rect 54077 1755 54087 1789
rect 54121 1755 54129 1789
rect 54077 1721 54129 1755
rect 54077 1687 54087 1721
rect 54121 1687 54129 1721
rect 54077 1673 54129 1687
rect 54985 1789 55037 1803
rect 54985 1755 54993 1789
rect 55027 1755 55037 1789
rect 54985 1721 55037 1755
rect 54985 1687 54993 1721
rect 55027 1687 55037 1721
rect 54985 1673 55037 1687
rect 55067 1789 55121 1803
rect 55067 1755 55077 1789
rect 55111 1755 55121 1789
rect 55067 1721 55121 1755
rect 55067 1687 55077 1721
rect 55111 1687 55121 1721
rect 55067 1673 55121 1687
rect 55151 1789 55203 1803
rect 55151 1755 55161 1789
rect 55195 1755 55203 1789
rect 55799 1789 55851 1803
rect 55151 1721 55203 1755
rect 55799 1755 55807 1789
rect 55841 1755 55851 1789
rect 55151 1687 55161 1721
rect 55195 1687 55203 1721
rect 55151 1673 55203 1687
rect 55799 1721 55851 1755
rect 55799 1687 55807 1721
rect 55841 1687 55851 1721
rect 55799 1673 55851 1687
rect 55881 1789 55935 1803
rect 55881 1755 55891 1789
rect 55925 1755 55935 1789
rect 55881 1721 55935 1755
rect 55881 1687 55891 1721
rect 55925 1687 55935 1721
rect 55881 1673 55935 1687
rect 55965 1789 56017 1803
rect 55965 1755 55975 1789
rect 56009 1755 56017 1789
rect 55965 1721 56017 1755
rect 55965 1687 55975 1721
rect 56009 1687 56017 1721
rect 55965 1673 56017 1687
rect 56873 1789 56925 1803
rect 56873 1755 56881 1789
rect 56915 1755 56925 1789
rect 56873 1721 56925 1755
rect 56873 1687 56881 1721
rect 56915 1687 56925 1721
rect 56873 1673 56925 1687
rect 56955 1789 57009 1803
rect 56955 1755 56965 1789
rect 56999 1755 57009 1789
rect 56955 1721 57009 1755
rect 56955 1687 56965 1721
rect 56999 1687 57009 1721
rect 56955 1673 57009 1687
rect 57039 1789 57091 1803
rect 57039 1755 57049 1789
rect 57083 1755 57091 1789
rect 57687 1789 57739 1803
rect 57039 1721 57091 1755
rect 57687 1755 57695 1789
rect 57729 1755 57739 1789
rect 57039 1687 57049 1721
rect 57083 1687 57091 1721
rect 57039 1673 57091 1687
rect 57687 1721 57739 1755
rect 57687 1687 57695 1721
rect 57729 1687 57739 1721
rect 57687 1673 57739 1687
rect 57769 1789 57823 1803
rect 57769 1755 57779 1789
rect 57813 1755 57823 1789
rect 57769 1721 57823 1755
rect 57769 1687 57779 1721
rect 57813 1687 57823 1721
rect 57769 1673 57823 1687
rect 57853 1789 57905 1803
rect 57853 1755 57863 1789
rect 57897 1755 57905 1789
rect 57853 1721 57905 1755
rect 57853 1687 57863 1721
rect 57897 1687 57905 1721
rect 57853 1673 57905 1687
rect 58761 1789 58813 1803
rect 58761 1755 58769 1789
rect 58803 1755 58813 1789
rect 58761 1721 58813 1755
rect 58761 1687 58769 1721
rect 58803 1687 58813 1721
rect 58761 1673 58813 1687
rect 58843 1789 58897 1803
rect 58843 1755 58853 1789
rect 58887 1755 58897 1789
rect 58843 1721 58897 1755
rect 58843 1687 58853 1721
rect 58887 1687 58897 1721
rect 58843 1673 58897 1687
rect 58927 1789 58979 1803
rect 58927 1755 58937 1789
rect 58971 1755 58979 1789
rect 59575 1789 59627 1803
rect 58927 1721 58979 1755
rect 59575 1755 59583 1789
rect 59617 1755 59627 1789
rect 58927 1687 58937 1721
rect 58971 1687 58979 1721
rect 58927 1673 58979 1687
rect 59575 1721 59627 1755
rect 59575 1687 59583 1721
rect 59617 1687 59627 1721
rect 59575 1673 59627 1687
rect 59657 1789 59711 1803
rect 59657 1755 59667 1789
rect 59701 1755 59711 1789
rect 59657 1721 59711 1755
rect 59657 1687 59667 1721
rect 59701 1687 59711 1721
rect 59657 1673 59711 1687
rect 59741 1789 59793 1803
rect 59741 1755 59751 1789
rect 59785 1755 59793 1789
rect 59741 1721 59793 1755
rect 59741 1687 59751 1721
rect 59785 1687 59793 1721
rect 59741 1673 59793 1687
rect 610 1544 672 1558
rect 610 1510 622 1544
rect 656 1510 672 1544
rect 610 1476 672 1510
rect 610 1442 622 1476
rect 656 1442 672 1476
rect 610 1428 672 1442
rect 702 1544 768 1558
rect 702 1510 718 1544
rect 752 1510 768 1544
rect 702 1476 768 1510
rect 702 1442 718 1476
rect 752 1442 768 1476
rect 702 1428 768 1442
rect 798 1544 860 1558
rect 798 1510 814 1544
rect 848 1510 860 1544
rect 798 1476 860 1510
rect 798 1442 814 1476
rect 848 1442 860 1476
rect 798 1428 860 1442
rect 2498 1544 2560 1558
rect 2498 1510 2510 1544
rect 2544 1510 2560 1544
rect 2498 1476 2560 1510
rect 2498 1442 2510 1476
rect 2544 1442 2560 1476
rect 2498 1428 2560 1442
rect 2590 1544 2656 1558
rect 2590 1510 2606 1544
rect 2640 1510 2656 1544
rect 2590 1476 2656 1510
rect 2590 1442 2606 1476
rect 2640 1442 2656 1476
rect 2590 1428 2656 1442
rect 2686 1544 2748 1558
rect 2686 1510 2702 1544
rect 2736 1510 2748 1544
rect 2686 1476 2748 1510
rect 2686 1442 2702 1476
rect 2736 1442 2748 1476
rect 2686 1428 2748 1442
rect 4386 1544 4448 1558
rect 4386 1510 4398 1544
rect 4432 1510 4448 1544
rect 4386 1476 4448 1510
rect 4386 1442 4398 1476
rect 4432 1442 4448 1476
rect 4386 1428 4448 1442
rect 4478 1544 4544 1558
rect 4478 1510 4494 1544
rect 4528 1510 4544 1544
rect 4478 1476 4544 1510
rect 4478 1442 4494 1476
rect 4528 1442 4544 1476
rect 4478 1428 4544 1442
rect 4574 1544 4636 1558
rect 4574 1510 4590 1544
rect 4624 1510 4636 1544
rect 4574 1476 4636 1510
rect 4574 1442 4590 1476
rect 4624 1442 4636 1476
rect 4574 1428 4636 1442
rect 6274 1544 6336 1558
rect 6274 1510 6286 1544
rect 6320 1510 6336 1544
rect 6274 1476 6336 1510
rect 6274 1442 6286 1476
rect 6320 1442 6336 1476
rect 6274 1428 6336 1442
rect 6366 1544 6432 1558
rect 6366 1510 6382 1544
rect 6416 1510 6432 1544
rect 6366 1476 6432 1510
rect 6366 1442 6382 1476
rect 6416 1442 6432 1476
rect 6366 1428 6432 1442
rect 6462 1544 6524 1558
rect 6462 1510 6478 1544
rect 6512 1510 6524 1544
rect 6462 1476 6524 1510
rect 6462 1442 6478 1476
rect 6512 1442 6524 1476
rect 6462 1428 6524 1442
rect 8162 1544 8224 1558
rect 8162 1510 8174 1544
rect 8208 1510 8224 1544
rect 8162 1476 8224 1510
rect 8162 1442 8174 1476
rect 8208 1442 8224 1476
rect 8162 1428 8224 1442
rect 8254 1544 8320 1558
rect 8254 1510 8270 1544
rect 8304 1510 8320 1544
rect 8254 1476 8320 1510
rect 8254 1442 8270 1476
rect 8304 1442 8320 1476
rect 8254 1428 8320 1442
rect 8350 1544 8412 1558
rect 8350 1510 8366 1544
rect 8400 1510 8412 1544
rect 8350 1476 8412 1510
rect 8350 1442 8366 1476
rect 8400 1442 8412 1476
rect 8350 1428 8412 1442
rect 10050 1544 10112 1558
rect 10050 1510 10062 1544
rect 10096 1510 10112 1544
rect 10050 1476 10112 1510
rect 10050 1442 10062 1476
rect 10096 1442 10112 1476
rect 10050 1428 10112 1442
rect 10142 1544 10208 1558
rect 10142 1510 10158 1544
rect 10192 1510 10208 1544
rect 10142 1476 10208 1510
rect 10142 1442 10158 1476
rect 10192 1442 10208 1476
rect 10142 1428 10208 1442
rect 10238 1544 10300 1558
rect 10238 1510 10254 1544
rect 10288 1510 10300 1544
rect 10238 1476 10300 1510
rect 10238 1442 10254 1476
rect 10288 1442 10300 1476
rect 10238 1428 10300 1442
rect 11938 1544 12000 1558
rect 11938 1510 11950 1544
rect 11984 1510 12000 1544
rect 11938 1476 12000 1510
rect 11938 1442 11950 1476
rect 11984 1442 12000 1476
rect 11938 1428 12000 1442
rect 12030 1544 12096 1558
rect 12030 1510 12046 1544
rect 12080 1510 12096 1544
rect 12030 1476 12096 1510
rect 12030 1442 12046 1476
rect 12080 1442 12096 1476
rect 12030 1428 12096 1442
rect 12126 1544 12188 1558
rect 12126 1510 12142 1544
rect 12176 1510 12188 1544
rect 12126 1476 12188 1510
rect 12126 1442 12142 1476
rect 12176 1442 12188 1476
rect 12126 1428 12188 1442
rect 13826 1544 13888 1558
rect 13826 1510 13838 1544
rect 13872 1510 13888 1544
rect 13826 1476 13888 1510
rect 13826 1442 13838 1476
rect 13872 1442 13888 1476
rect 13826 1428 13888 1442
rect 13918 1544 13984 1558
rect 13918 1510 13934 1544
rect 13968 1510 13984 1544
rect 13918 1476 13984 1510
rect 13918 1442 13934 1476
rect 13968 1442 13984 1476
rect 13918 1428 13984 1442
rect 14014 1544 14076 1558
rect 14014 1510 14030 1544
rect 14064 1510 14076 1544
rect 14014 1476 14076 1510
rect 14014 1442 14030 1476
rect 14064 1442 14076 1476
rect 14014 1428 14076 1442
rect 15708 1544 15770 1558
rect 15708 1510 15720 1544
rect 15754 1510 15770 1544
rect 15708 1476 15770 1510
rect 15708 1442 15720 1476
rect 15754 1442 15770 1476
rect 15708 1428 15770 1442
rect 15800 1544 15866 1558
rect 15800 1510 15816 1544
rect 15850 1510 15866 1544
rect 15800 1476 15866 1510
rect 15800 1442 15816 1476
rect 15850 1442 15866 1476
rect 15800 1428 15866 1442
rect 15896 1544 15958 1558
rect 15896 1510 15912 1544
rect 15946 1510 15958 1544
rect 15896 1476 15958 1510
rect 15896 1442 15912 1476
rect 15946 1442 15958 1476
rect 15896 1428 15958 1442
rect 17596 1544 17658 1558
rect 17596 1510 17608 1544
rect 17642 1510 17658 1544
rect 17596 1476 17658 1510
rect 17596 1442 17608 1476
rect 17642 1442 17658 1476
rect 17596 1428 17658 1442
rect 17688 1544 17754 1558
rect 17688 1510 17704 1544
rect 17738 1510 17754 1544
rect 17688 1476 17754 1510
rect 17688 1442 17704 1476
rect 17738 1442 17754 1476
rect 17688 1428 17754 1442
rect 17784 1544 17846 1558
rect 17784 1510 17800 1544
rect 17834 1510 17846 1544
rect 17784 1476 17846 1510
rect 17784 1442 17800 1476
rect 17834 1442 17846 1476
rect 17784 1428 17846 1442
rect 19484 1544 19546 1558
rect 19484 1510 19496 1544
rect 19530 1510 19546 1544
rect 19484 1476 19546 1510
rect 19484 1442 19496 1476
rect 19530 1442 19546 1476
rect 19484 1428 19546 1442
rect 19576 1544 19642 1558
rect 19576 1510 19592 1544
rect 19626 1510 19642 1544
rect 19576 1476 19642 1510
rect 19576 1442 19592 1476
rect 19626 1442 19642 1476
rect 19576 1428 19642 1442
rect 19672 1544 19734 1558
rect 19672 1510 19688 1544
rect 19722 1510 19734 1544
rect 19672 1476 19734 1510
rect 19672 1442 19688 1476
rect 19722 1442 19734 1476
rect 19672 1428 19734 1442
rect 21372 1544 21434 1558
rect 21372 1510 21384 1544
rect 21418 1510 21434 1544
rect 21372 1476 21434 1510
rect 21372 1442 21384 1476
rect 21418 1442 21434 1476
rect 21372 1428 21434 1442
rect 21464 1544 21530 1558
rect 21464 1510 21480 1544
rect 21514 1510 21530 1544
rect 21464 1476 21530 1510
rect 21464 1442 21480 1476
rect 21514 1442 21530 1476
rect 21464 1428 21530 1442
rect 21560 1544 21622 1558
rect 21560 1510 21576 1544
rect 21610 1510 21622 1544
rect 21560 1476 21622 1510
rect 21560 1442 21576 1476
rect 21610 1442 21622 1476
rect 21560 1428 21622 1442
rect 23260 1544 23322 1558
rect 23260 1510 23272 1544
rect 23306 1510 23322 1544
rect 23260 1476 23322 1510
rect 23260 1442 23272 1476
rect 23306 1442 23322 1476
rect 23260 1428 23322 1442
rect 23352 1544 23418 1558
rect 23352 1510 23368 1544
rect 23402 1510 23418 1544
rect 23352 1476 23418 1510
rect 23352 1442 23368 1476
rect 23402 1442 23418 1476
rect 23352 1428 23418 1442
rect 23448 1544 23510 1558
rect 23448 1510 23464 1544
rect 23498 1510 23510 1544
rect 23448 1476 23510 1510
rect 23448 1442 23464 1476
rect 23498 1442 23510 1476
rect 23448 1428 23510 1442
rect 25148 1544 25210 1558
rect 25148 1510 25160 1544
rect 25194 1510 25210 1544
rect 25148 1476 25210 1510
rect 25148 1442 25160 1476
rect 25194 1442 25210 1476
rect 25148 1428 25210 1442
rect 25240 1544 25306 1558
rect 25240 1510 25256 1544
rect 25290 1510 25306 1544
rect 25240 1476 25306 1510
rect 25240 1442 25256 1476
rect 25290 1442 25306 1476
rect 25240 1428 25306 1442
rect 25336 1544 25398 1558
rect 25336 1510 25352 1544
rect 25386 1510 25398 1544
rect 25336 1476 25398 1510
rect 25336 1442 25352 1476
rect 25386 1442 25398 1476
rect 25336 1428 25398 1442
rect 27036 1544 27098 1558
rect 27036 1510 27048 1544
rect 27082 1510 27098 1544
rect 27036 1476 27098 1510
rect 27036 1442 27048 1476
rect 27082 1442 27098 1476
rect 27036 1428 27098 1442
rect 27128 1544 27194 1558
rect 27128 1510 27144 1544
rect 27178 1510 27194 1544
rect 27128 1476 27194 1510
rect 27128 1442 27144 1476
rect 27178 1442 27194 1476
rect 27128 1428 27194 1442
rect 27224 1544 27286 1558
rect 27224 1510 27240 1544
rect 27274 1510 27286 1544
rect 27224 1476 27286 1510
rect 27224 1442 27240 1476
rect 27274 1442 27286 1476
rect 27224 1428 27286 1442
rect 28924 1544 28986 1558
rect 28924 1510 28936 1544
rect 28970 1510 28986 1544
rect 28924 1476 28986 1510
rect 28924 1442 28936 1476
rect 28970 1442 28986 1476
rect 28924 1428 28986 1442
rect 29016 1544 29082 1558
rect 29016 1510 29032 1544
rect 29066 1510 29082 1544
rect 29016 1476 29082 1510
rect 29016 1442 29032 1476
rect 29066 1442 29082 1476
rect 29016 1428 29082 1442
rect 29112 1544 29174 1558
rect 29112 1510 29128 1544
rect 29162 1510 29174 1544
rect 29112 1476 29174 1510
rect 29112 1442 29128 1476
rect 29162 1442 29174 1476
rect 29112 1428 29174 1442
rect 30812 1544 30874 1558
rect 30812 1510 30824 1544
rect 30858 1510 30874 1544
rect 30812 1476 30874 1510
rect 30812 1442 30824 1476
rect 30858 1442 30874 1476
rect 30812 1428 30874 1442
rect 30904 1544 30970 1558
rect 30904 1510 30920 1544
rect 30954 1510 30970 1544
rect 30904 1476 30970 1510
rect 30904 1442 30920 1476
rect 30954 1442 30970 1476
rect 30904 1428 30970 1442
rect 31000 1544 31062 1558
rect 31000 1510 31016 1544
rect 31050 1510 31062 1544
rect 31000 1476 31062 1510
rect 31000 1442 31016 1476
rect 31050 1442 31062 1476
rect 31000 1428 31062 1442
rect 32700 1544 32762 1558
rect 32700 1510 32712 1544
rect 32746 1510 32762 1544
rect 32700 1476 32762 1510
rect 32700 1442 32712 1476
rect 32746 1442 32762 1476
rect 32700 1428 32762 1442
rect 32792 1544 32858 1558
rect 32792 1510 32808 1544
rect 32842 1510 32858 1544
rect 32792 1476 32858 1510
rect 32792 1442 32808 1476
rect 32842 1442 32858 1476
rect 32792 1428 32858 1442
rect 32888 1544 32950 1558
rect 32888 1510 32904 1544
rect 32938 1510 32950 1544
rect 32888 1476 32950 1510
rect 32888 1442 32904 1476
rect 32938 1442 32950 1476
rect 32888 1428 32950 1442
rect 34588 1544 34650 1558
rect 34588 1510 34600 1544
rect 34634 1510 34650 1544
rect 34588 1476 34650 1510
rect 34588 1442 34600 1476
rect 34634 1442 34650 1476
rect 34588 1428 34650 1442
rect 34680 1544 34746 1558
rect 34680 1510 34696 1544
rect 34730 1510 34746 1544
rect 34680 1476 34746 1510
rect 34680 1442 34696 1476
rect 34730 1442 34746 1476
rect 34680 1428 34746 1442
rect 34776 1544 34838 1558
rect 34776 1510 34792 1544
rect 34826 1510 34838 1544
rect 34776 1476 34838 1510
rect 34776 1442 34792 1476
rect 34826 1442 34838 1476
rect 34776 1428 34838 1442
rect 36476 1544 36538 1558
rect 36476 1510 36488 1544
rect 36522 1510 36538 1544
rect 36476 1476 36538 1510
rect 36476 1442 36488 1476
rect 36522 1442 36538 1476
rect 36476 1428 36538 1442
rect 36568 1544 36634 1558
rect 36568 1510 36584 1544
rect 36618 1510 36634 1544
rect 36568 1476 36634 1510
rect 36568 1442 36584 1476
rect 36618 1442 36634 1476
rect 36568 1428 36634 1442
rect 36664 1544 36726 1558
rect 36664 1510 36680 1544
rect 36714 1510 36726 1544
rect 36664 1476 36726 1510
rect 36664 1442 36680 1476
rect 36714 1442 36726 1476
rect 36664 1428 36726 1442
rect 38364 1544 38426 1558
rect 38364 1510 38376 1544
rect 38410 1510 38426 1544
rect 38364 1476 38426 1510
rect 38364 1442 38376 1476
rect 38410 1442 38426 1476
rect 38364 1428 38426 1442
rect 38456 1544 38522 1558
rect 38456 1510 38472 1544
rect 38506 1510 38522 1544
rect 38456 1476 38522 1510
rect 38456 1442 38472 1476
rect 38506 1442 38522 1476
rect 38456 1428 38522 1442
rect 38552 1544 38614 1558
rect 38552 1510 38568 1544
rect 38602 1510 38614 1544
rect 38552 1476 38614 1510
rect 38552 1442 38568 1476
rect 38602 1442 38614 1476
rect 38552 1428 38614 1442
rect 40252 1544 40314 1558
rect 40252 1510 40264 1544
rect 40298 1510 40314 1544
rect 40252 1476 40314 1510
rect 40252 1442 40264 1476
rect 40298 1442 40314 1476
rect 40252 1428 40314 1442
rect 40344 1544 40410 1558
rect 40344 1510 40360 1544
rect 40394 1510 40410 1544
rect 40344 1476 40410 1510
rect 40344 1442 40360 1476
rect 40394 1442 40410 1476
rect 40344 1428 40410 1442
rect 40440 1544 40502 1558
rect 40440 1510 40456 1544
rect 40490 1510 40502 1544
rect 40440 1476 40502 1510
rect 40440 1442 40456 1476
rect 40490 1442 40502 1476
rect 40440 1428 40502 1442
rect 42140 1544 42202 1558
rect 42140 1510 42152 1544
rect 42186 1510 42202 1544
rect 42140 1476 42202 1510
rect 42140 1442 42152 1476
rect 42186 1442 42202 1476
rect 42140 1428 42202 1442
rect 42232 1544 42298 1558
rect 42232 1510 42248 1544
rect 42282 1510 42298 1544
rect 42232 1476 42298 1510
rect 42232 1442 42248 1476
rect 42282 1442 42298 1476
rect 42232 1428 42298 1442
rect 42328 1544 42390 1558
rect 42328 1510 42344 1544
rect 42378 1510 42390 1544
rect 42328 1476 42390 1510
rect 42328 1442 42344 1476
rect 42378 1442 42390 1476
rect 42328 1428 42390 1442
rect 44028 1544 44090 1558
rect 44028 1510 44040 1544
rect 44074 1510 44090 1544
rect 44028 1476 44090 1510
rect 44028 1442 44040 1476
rect 44074 1442 44090 1476
rect 44028 1428 44090 1442
rect 44120 1544 44186 1558
rect 44120 1510 44136 1544
rect 44170 1510 44186 1544
rect 44120 1476 44186 1510
rect 44120 1442 44136 1476
rect 44170 1442 44186 1476
rect 44120 1428 44186 1442
rect 44216 1544 44278 1558
rect 44216 1510 44232 1544
rect 44266 1510 44278 1544
rect 44216 1476 44278 1510
rect 44216 1442 44232 1476
rect 44266 1442 44278 1476
rect 44216 1428 44278 1442
rect 45910 1544 45972 1558
rect 45910 1510 45922 1544
rect 45956 1510 45972 1544
rect 45910 1476 45972 1510
rect 45910 1442 45922 1476
rect 45956 1442 45972 1476
rect 45910 1428 45972 1442
rect 46002 1544 46068 1558
rect 46002 1510 46018 1544
rect 46052 1510 46068 1544
rect 46002 1476 46068 1510
rect 46002 1442 46018 1476
rect 46052 1442 46068 1476
rect 46002 1428 46068 1442
rect 46098 1544 46160 1558
rect 46098 1510 46114 1544
rect 46148 1510 46160 1544
rect 46098 1476 46160 1510
rect 46098 1442 46114 1476
rect 46148 1442 46160 1476
rect 46098 1428 46160 1442
rect 47798 1544 47860 1558
rect 47798 1510 47810 1544
rect 47844 1510 47860 1544
rect 47798 1476 47860 1510
rect 47798 1442 47810 1476
rect 47844 1442 47860 1476
rect 47798 1428 47860 1442
rect 47890 1544 47956 1558
rect 47890 1510 47906 1544
rect 47940 1510 47956 1544
rect 47890 1476 47956 1510
rect 47890 1442 47906 1476
rect 47940 1442 47956 1476
rect 47890 1428 47956 1442
rect 47986 1544 48048 1558
rect 47986 1510 48002 1544
rect 48036 1510 48048 1544
rect 47986 1476 48048 1510
rect 47986 1442 48002 1476
rect 48036 1442 48048 1476
rect 47986 1428 48048 1442
rect 49686 1544 49748 1558
rect 49686 1510 49698 1544
rect 49732 1510 49748 1544
rect 49686 1476 49748 1510
rect 49686 1442 49698 1476
rect 49732 1442 49748 1476
rect 49686 1428 49748 1442
rect 49778 1544 49844 1558
rect 49778 1510 49794 1544
rect 49828 1510 49844 1544
rect 49778 1476 49844 1510
rect 49778 1442 49794 1476
rect 49828 1442 49844 1476
rect 49778 1428 49844 1442
rect 49874 1544 49936 1558
rect 49874 1510 49890 1544
rect 49924 1510 49936 1544
rect 49874 1476 49936 1510
rect 49874 1442 49890 1476
rect 49924 1442 49936 1476
rect 49874 1428 49936 1442
rect 51574 1544 51636 1558
rect 51574 1510 51586 1544
rect 51620 1510 51636 1544
rect 51574 1476 51636 1510
rect 51574 1442 51586 1476
rect 51620 1442 51636 1476
rect 51574 1428 51636 1442
rect 51666 1544 51732 1558
rect 51666 1510 51682 1544
rect 51716 1510 51732 1544
rect 51666 1476 51732 1510
rect 51666 1442 51682 1476
rect 51716 1442 51732 1476
rect 51666 1428 51732 1442
rect 51762 1544 51824 1558
rect 51762 1510 51778 1544
rect 51812 1510 51824 1544
rect 51762 1476 51824 1510
rect 51762 1442 51778 1476
rect 51812 1442 51824 1476
rect 51762 1428 51824 1442
rect 53462 1544 53524 1558
rect 53462 1510 53474 1544
rect 53508 1510 53524 1544
rect 53462 1476 53524 1510
rect 53462 1442 53474 1476
rect 53508 1442 53524 1476
rect 53462 1428 53524 1442
rect 53554 1544 53620 1558
rect 53554 1510 53570 1544
rect 53604 1510 53620 1544
rect 53554 1476 53620 1510
rect 53554 1442 53570 1476
rect 53604 1442 53620 1476
rect 53554 1428 53620 1442
rect 53650 1544 53712 1558
rect 53650 1510 53666 1544
rect 53700 1510 53712 1544
rect 53650 1476 53712 1510
rect 53650 1442 53666 1476
rect 53700 1442 53712 1476
rect 53650 1428 53712 1442
rect 55350 1544 55412 1558
rect 55350 1510 55362 1544
rect 55396 1510 55412 1544
rect 55350 1476 55412 1510
rect 55350 1442 55362 1476
rect 55396 1442 55412 1476
rect 55350 1428 55412 1442
rect 55442 1544 55508 1558
rect 55442 1510 55458 1544
rect 55492 1510 55508 1544
rect 55442 1476 55508 1510
rect 55442 1442 55458 1476
rect 55492 1442 55508 1476
rect 55442 1428 55508 1442
rect 55538 1544 55600 1558
rect 55538 1510 55554 1544
rect 55588 1510 55600 1544
rect 55538 1476 55600 1510
rect 55538 1442 55554 1476
rect 55588 1442 55600 1476
rect 55538 1428 55600 1442
rect 57238 1544 57300 1558
rect 57238 1510 57250 1544
rect 57284 1510 57300 1544
rect 57238 1476 57300 1510
rect 57238 1442 57250 1476
rect 57284 1442 57300 1476
rect 57238 1428 57300 1442
rect 57330 1544 57396 1558
rect 57330 1510 57346 1544
rect 57380 1510 57396 1544
rect 57330 1476 57396 1510
rect 57330 1442 57346 1476
rect 57380 1442 57396 1476
rect 57330 1428 57396 1442
rect 57426 1544 57488 1558
rect 57426 1510 57442 1544
rect 57476 1510 57488 1544
rect 57426 1476 57488 1510
rect 57426 1442 57442 1476
rect 57476 1442 57488 1476
rect 57426 1428 57488 1442
rect 59126 1544 59188 1558
rect 59126 1510 59138 1544
rect 59172 1510 59188 1544
rect 59126 1476 59188 1510
rect 59126 1442 59138 1476
rect 59172 1442 59188 1476
rect 59126 1428 59188 1442
rect 59218 1544 59284 1558
rect 59218 1510 59234 1544
rect 59268 1510 59284 1544
rect 59218 1476 59284 1510
rect 59218 1442 59234 1476
rect 59268 1442 59284 1476
rect 59218 1428 59284 1442
rect 59314 1544 59376 1558
rect 59314 1510 59330 1544
rect 59364 1510 59376 1544
rect 59314 1476 59376 1510
rect 59314 1442 59330 1476
rect 59364 1442 59376 1476
rect 59314 1428 59376 1442
rect 108 737 160 749
rect 108 703 116 737
rect 150 703 160 737
rect 108 669 160 703
rect 108 635 116 669
rect 150 635 160 669
rect 108 619 160 635
rect 190 737 242 749
rect 190 703 200 737
rect 234 703 242 737
rect 190 669 242 703
rect 1304 745 1356 757
rect 1304 711 1312 745
rect 1346 711 1356 745
rect 1304 677 1356 711
rect 190 635 200 669
rect 234 635 242 669
rect 190 619 242 635
rect 1304 643 1312 677
rect 1346 643 1356 677
rect 1304 627 1356 643
rect 1386 745 1438 757
rect 1386 711 1396 745
rect 1430 711 1438 745
rect 1996 737 2048 749
rect 1386 677 1438 711
rect 1386 643 1396 677
rect 1430 643 1438 677
rect 1386 627 1438 643
rect 1609 684 1661 729
rect 1609 650 1617 684
rect 1651 650 1661 684
rect 1609 625 1661 650
rect 1691 671 1749 729
rect 1691 637 1703 671
rect 1737 637 1749 671
rect 1691 625 1749 637
rect 1779 701 1831 729
rect 1779 667 1789 701
rect 1823 667 1831 701
rect 1779 625 1831 667
rect 1996 703 2004 737
rect 2038 703 2048 737
rect 1996 669 2048 703
rect 1996 635 2004 669
rect 2038 635 2048 669
rect 1996 619 2048 635
rect 2078 737 2130 749
rect 2078 703 2088 737
rect 2122 703 2130 737
rect 2078 669 2130 703
rect 3192 745 3244 757
rect 3192 711 3200 745
rect 3234 711 3244 745
rect 3192 677 3244 711
rect 2078 635 2088 669
rect 2122 635 2130 669
rect 2078 619 2130 635
rect 3192 643 3200 677
rect 3234 643 3244 677
rect 3192 627 3244 643
rect 3274 745 3326 757
rect 3274 711 3284 745
rect 3318 711 3326 745
rect 3884 737 3936 749
rect 3274 677 3326 711
rect 3274 643 3284 677
rect 3318 643 3326 677
rect 3274 627 3326 643
rect 3497 684 3549 729
rect 3497 650 3505 684
rect 3539 650 3549 684
rect 3497 625 3549 650
rect 3579 671 3637 729
rect 3579 637 3591 671
rect 3625 637 3637 671
rect 3579 625 3637 637
rect 3667 701 3719 729
rect 3667 667 3677 701
rect 3711 667 3719 701
rect 3667 625 3719 667
rect 3884 703 3892 737
rect 3926 703 3936 737
rect 3884 669 3936 703
rect 3884 635 3892 669
rect 3926 635 3936 669
rect 3884 619 3936 635
rect 3966 737 4018 749
rect 3966 703 3976 737
rect 4010 703 4018 737
rect 3966 669 4018 703
rect 5080 745 5132 757
rect 5080 711 5088 745
rect 5122 711 5132 745
rect 5080 677 5132 711
rect 3966 635 3976 669
rect 4010 635 4018 669
rect 3966 619 4018 635
rect 5080 643 5088 677
rect 5122 643 5132 677
rect 5080 627 5132 643
rect 5162 745 5214 757
rect 5162 711 5172 745
rect 5206 711 5214 745
rect 5772 737 5824 749
rect 5162 677 5214 711
rect 5162 643 5172 677
rect 5206 643 5214 677
rect 5162 627 5214 643
rect 5385 684 5437 729
rect 5385 650 5393 684
rect 5427 650 5437 684
rect 5385 625 5437 650
rect 5467 671 5525 729
rect 5467 637 5479 671
rect 5513 637 5525 671
rect 5467 625 5525 637
rect 5555 701 5607 729
rect 5555 667 5565 701
rect 5599 667 5607 701
rect 5555 625 5607 667
rect 5772 703 5780 737
rect 5814 703 5824 737
rect 5772 669 5824 703
rect 5772 635 5780 669
rect 5814 635 5824 669
rect 5772 619 5824 635
rect 5854 737 5906 749
rect 5854 703 5864 737
rect 5898 703 5906 737
rect 5854 669 5906 703
rect 6968 745 7020 757
rect 6968 711 6976 745
rect 7010 711 7020 745
rect 6968 677 7020 711
rect 5854 635 5864 669
rect 5898 635 5906 669
rect 5854 619 5906 635
rect 6968 643 6976 677
rect 7010 643 7020 677
rect 6968 627 7020 643
rect 7050 745 7102 757
rect 7050 711 7060 745
rect 7094 711 7102 745
rect 7660 737 7712 749
rect 7050 677 7102 711
rect 7050 643 7060 677
rect 7094 643 7102 677
rect 7050 627 7102 643
rect 7273 684 7325 729
rect 7273 650 7281 684
rect 7315 650 7325 684
rect 7273 625 7325 650
rect 7355 671 7413 729
rect 7355 637 7367 671
rect 7401 637 7413 671
rect 7355 625 7413 637
rect 7443 701 7495 729
rect 7443 667 7453 701
rect 7487 667 7495 701
rect 7443 625 7495 667
rect 7660 703 7668 737
rect 7702 703 7712 737
rect 7660 669 7712 703
rect 7660 635 7668 669
rect 7702 635 7712 669
rect 7660 619 7712 635
rect 7742 737 7794 749
rect 7742 703 7752 737
rect 7786 703 7794 737
rect 7742 669 7794 703
rect 8856 745 8908 757
rect 8856 711 8864 745
rect 8898 711 8908 745
rect 8856 677 8908 711
rect 7742 635 7752 669
rect 7786 635 7794 669
rect 7742 619 7794 635
rect 8856 643 8864 677
rect 8898 643 8908 677
rect 8856 627 8908 643
rect 8938 745 8990 757
rect 8938 711 8948 745
rect 8982 711 8990 745
rect 9548 737 9600 749
rect 8938 677 8990 711
rect 8938 643 8948 677
rect 8982 643 8990 677
rect 8938 627 8990 643
rect 9161 684 9213 729
rect 9161 650 9169 684
rect 9203 650 9213 684
rect 9161 625 9213 650
rect 9243 671 9301 729
rect 9243 637 9255 671
rect 9289 637 9301 671
rect 9243 625 9301 637
rect 9331 701 9383 729
rect 9331 667 9341 701
rect 9375 667 9383 701
rect 9331 625 9383 667
rect 9548 703 9556 737
rect 9590 703 9600 737
rect 9548 669 9600 703
rect 9548 635 9556 669
rect 9590 635 9600 669
rect 9548 619 9600 635
rect 9630 737 9682 749
rect 9630 703 9640 737
rect 9674 703 9682 737
rect 9630 669 9682 703
rect 10744 745 10796 757
rect 10744 711 10752 745
rect 10786 711 10796 745
rect 10744 677 10796 711
rect 9630 635 9640 669
rect 9674 635 9682 669
rect 9630 619 9682 635
rect 10744 643 10752 677
rect 10786 643 10796 677
rect 10744 627 10796 643
rect 10826 745 10878 757
rect 10826 711 10836 745
rect 10870 711 10878 745
rect 11436 737 11488 749
rect 10826 677 10878 711
rect 10826 643 10836 677
rect 10870 643 10878 677
rect 10826 627 10878 643
rect 11049 684 11101 729
rect 11049 650 11057 684
rect 11091 650 11101 684
rect 11049 625 11101 650
rect 11131 671 11189 729
rect 11131 637 11143 671
rect 11177 637 11189 671
rect 11131 625 11189 637
rect 11219 701 11271 729
rect 11219 667 11229 701
rect 11263 667 11271 701
rect 11219 625 11271 667
rect 11436 703 11444 737
rect 11478 703 11488 737
rect 11436 669 11488 703
rect 11436 635 11444 669
rect 11478 635 11488 669
rect 11436 619 11488 635
rect 11518 737 11570 749
rect 11518 703 11528 737
rect 11562 703 11570 737
rect 11518 669 11570 703
rect 12632 745 12684 757
rect 12632 711 12640 745
rect 12674 711 12684 745
rect 12632 677 12684 711
rect 11518 635 11528 669
rect 11562 635 11570 669
rect 11518 619 11570 635
rect 12632 643 12640 677
rect 12674 643 12684 677
rect 12632 627 12684 643
rect 12714 745 12766 757
rect 12714 711 12724 745
rect 12758 711 12766 745
rect 13324 737 13376 749
rect 12714 677 12766 711
rect 12714 643 12724 677
rect 12758 643 12766 677
rect 12714 627 12766 643
rect 12937 684 12989 729
rect 12937 650 12945 684
rect 12979 650 12989 684
rect 12937 625 12989 650
rect 13019 671 13077 729
rect 13019 637 13031 671
rect 13065 637 13077 671
rect 13019 625 13077 637
rect 13107 701 13159 729
rect 13107 667 13117 701
rect 13151 667 13159 701
rect 13107 625 13159 667
rect 13324 703 13332 737
rect 13366 703 13376 737
rect 13324 669 13376 703
rect 13324 635 13332 669
rect 13366 635 13376 669
rect 13324 619 13376 635
rect 13406 737 13458 749
rect 13406 703 13416 737
rect 13450 703 13458 737
rect 13406 669 13458 703
rect 14520 745 14572 757
rect 14520 711 14528 745
rect 14562 711 14572 745
rect 14520 677 14572 711
rect 13406 635 13416 669
rect 13450 635 13458 669
rect 13406 619 13458 635
rect 14520 643 14528 677
rect 14562 643 14572 677
rect 14520 627 14572 643
rect 14602 745 14654 757
rect 14602 711 14612 745
rect 14646 711 14654 745
rect 15206 737 15258 749
rect 14602 677 14654 711
rect 14602 643 14612 677
rect 14646 643 14654 677
rect 14602 627 14654 643
rect 14825 684 14877 729
rect 14825 650 14833 684
rect 14867 650 14877 684
rect 14825 625 14877 650
rect 14907 671 14965 729
rect 14907 637 14919 671
rect 14953 637 14965 671
rect 14907 625 14965 637
rect 14995 701 15047 729
rect 14995 667 15005 701
rect 15039 667 15047 701
rect 14995 625 15047 667
rect 15206 703 15214 737
rect 15248 703 15258 737
rect 15206 669 15258 703
rect 15206 635 15214 669
rect 15248 635 15258 669
rect 15206 619 15258 635
rect 15288 737 15340 749
rect 15288 703 15298 737
rect 15332 703 15340 737
rect 15288 669 15340 703
rect 16402 745 16454 757
rect 16402 711 16410 745
rect 16444 711 16454 745
rect 16402 677 16454 711
rect 15288 635 15298 669
rect 15332 635 15340 669
rect 15288 619 15340 635
rect 16402 643 16410 677
rect 16444 643 16454 677
rect 16402 627 16454 643
rect 16484 745 16536 757
rect 16484 711 16494 745
rect 16528 711 16536 745
rect 17094 737 17146 749
rect 16484 677 16536 711
rect 16484 643 16494 677
rect 16528 643 16536 677
rect 16484 627 16536 643
rect 16707 684 16759 729
rect 16707 650 16715 684
rect 16749 650 16759 684
rect 16707 625 16759 650
rect 16789 671 16847 729
rect 16789 637 16801 671
rect 16835 637 16847 671
rect 16789 625 16847 637
rect 16877 701 16929 729
rect 16877 667 16887 701
rect 16921 667 16929 701
rect 16877 625 16929 667
rect 17094 703 17102 737
rect 17136 703 17146 737
rect 17094 669 17146 703
rect 17094 635 17102 669
rect 17136 635 17146 669
rect 17094 619 17146 635
rect 17176 737 17228 749
rect 17176 703 17186 737
rect 17220 703 17228 737
rect 17176 669 17228 703
rect 18290 745 18342 757
rect 18290 711 18298 745
rect 18332 711 18342 745
rect 18290 677 18342 711
rect 17176 635 17186 669
rect 17220 635 17228 669
rect 17176 619 17228 635
rect 18290 643 18298 677
rect 18332 643 18342 677
rect 18290 627 18342 643
rect 18372 745 18424 757
rect 18372 711 18382 745
rect 18416 711 18424 745
rect 18982 737 19034 749
rect 18372 677 18424 711
rect 18372 643 18382 677
rect 18416 643 18424 677
rect 18372 627 18424 643
rect 18595 684 18647 729
rect 18595 650 18603 684
rect 18637 650 18647 684
rect 18595 625 18647 650
rect 18677 671 18735 729
rect 18677 637 18689 671
rect 18723 637 18735 671
rect 18677 625 18735 637
rect 18765 701 18817 729
rect 18765 667 18775 701
rect 18809 667 18817 701
rect 18765 625 18817 667
rect 18982 703 18990 737
rect 19024 703 19034 737
rect 18982 669 19034 703
rect 18982 635 18990 669
rect 19024 635 19034 669
rect 18982 619 19034 635
rect 19064 737 19116 749
rect 19064 703 19074 737
rect 19108 703 19116 737
rect 19064 669 19116 703
rect 20178 745 20230 757
rect 20178 711 20186 745
rect 20220 711 20230 745
rect 20178 677 20230 711
rect 19064 635 19074 669
rect 19108 635 19116 669
rect 19064 619 19116 635
rect 20178 643 20186 677
rect 20220 643 20230 677
rect 20178 627 20230 643
rect 20260 745 20312 757
rect 20260 711 20270 745
rect 20304 711 20312 745
rect 20870 737 20922 749
rect 20260 677 20312 711
rect 20260 643 20270 677
rect 20304 643 20312 677
rect 20260 627 20312 643
rect 20483 684 20535 729
rect 20483 650 20491 684
rect 20525 650 20535 684
rect 20483 625 20535 650
rect 20565 671 20623 729
rect 20565 637 20577 671
rect 20611 637 20623 671
rect 20565 625 20623 637
rect 20653 701 20705 729
rect 20653 667 20663 701
rect 20697 667 20705 701
rect 20653 625 20705 667
rect 20870 703 20878 737
rect 20912 703 20922 737
rect 20870 669 20922 703
rect 20870 635 20878 669
rect 20912 635 20922 669
rect 20870 619 20922 635
rect 20952 737 21004 749
rect 20952 703 20962 737
rect 20996 703 21004 737
rect 20952 669 21004 703
rect 22066 745 22118 757
rect 22066 711 22074 745
rect 22108 711 22118 745
rect 22066 677 22118 711
rect 20952 635 20962 669
rect 20996 635 21004 669
rect 20952 619 21004 635
rect 22066 643 22074 677
rect 22108 643 22118 677
rect 22066 627 22118 643
rect 22148 745 22200 757
rect 22148 711 22158 745
rect 22192 711 22200 745
rect 22758 737 22810 749
rect 22148 677 22200 711
rect 22148 643 22158 677
rect 22192 643 22200 677
rect 22148 627 22200 643
rect 22371 684 22423 729
rect 22371 650 22379 684
rect 22413 650 22423 684
rect 22371 625 22423 650
rect 22453 671 22511 729
rect 22453 637 22465 671
rect 22499 637 22511 671
rect 22453 625 22511 637
rect 22541 701 22593 729
rect 22541 667 22551 701
rect 22585 667 22593 701
rect 22541 625 22593 667
rect 22758 703 22766 737
rect 22800 703 22810 737
rect 22758 669 22810 703
rect 22758 635 22766 669
rect 22800 635 22810 669
rect 22758 619 22810 635
rect 22840 737 22892 749
rect 22840 703 22850 737
rect 22884 703 22892 737
rect 22840 669 22892 703
rect 23954 745 24006 757
rect 23954 711 23962 745
rect 23996 711 24006 745
rect 23954 677 24006 711
rect 22840 635 22850 669
rect 22884 635 22892 669
rect 22840 619 22892 635
rect 23954 643 23962 677
rect 23996 643 24006 677
rect 23954 627 24006 643
rect 24036 745 24088 757
rect 24036 711 24046 745
rect 24080 711 24088 745
rect 24646 737 24698 749
rect 24036 677 24088 711
rect 24036 643 24046 677
rect 24080 643 24088 677
rect 24036 627 24088 643
rect 24259 684 24311 729
rect 24259 650 24267 684
rect 24301 650 24311 684
rect 24259 625 24311 650
rect 24341 671 24399 729
rect 24341 637 24353 671
rect 24387 637 24399 671
rect 24341 625 24399 637
rect 24429 701 24481 729
rect 24429 667 24439 701
rect 24473 667 24481 701
rect 24429 625 24481 667
rect 24646 703 24654 737
rect 24688 703 24698 737
rect 24646 669 24698 703
rect 24646 635 24654 669
rect 24688 635 24698 669
rect 24646 619 24698 635
rect 24728 737 24780 749
rect 24728 703 24738 737
rect 24772 703 24780 737
rect 24728 669 24780 703
rect 25842 745 25894 757
rect 25842 711 25850 745
rect 25884 711 25894 745
rect 25842 677 25894 711
rect 24728 635 24738 669
rect 24772 635 24780 669
rect 24728 619 24780 635
rect 25842 643 25850 677
rect 25884 643 25894 677
rect 25842 627 25894 643
rect 25924 745 25976 757
rect 25924 711 25934 745
rect 25968 711 25976 745
rect 26534 737 26586 749
rect 25924 677 25976 711
rect 25924 643 25934 677
rect 25968 643 25976 677
rect 25924 627 25976 643
rect 26147 684 26199 729
rect 26147 650 26155 684
rect 26189 650 26199 684
rect 26147 625 26199 650
rect 26229 671 26287 729
rect 26229 637 26241 671
rect 26275 637 26287 671
rect 26229 625 26287 637
rect 26317 701 26369 729
rect 26317 667 26327 701
rect 26361 667 26369 701
rect 26317 625 26369 667
rect 26534 703 26542 737
rect 26576 703 26586 737
rect 26534 669 26586 703
rect 26534 635 26542 669
rect 26576 635 26586 669
rect 26534 619 26586 635
rect 26616 737 26668 749
rect 26616 703 26626 737
rect 26660 703 26668 737
rect 26616 669 26668 703
rect 27730 745 27782 757
rect 27730 711 27738 745
rect 27772 711 27782 745
rect 27730 677 27782 711
rect 26616 635 26626 669
rect 26660 635 26668 669
rect 26616 619 26668 635
rect 27730 643 27738 677
rect 27772 643 27782 677
rect 27730 627 27782 643
rect 27812 745 27864 757
rect 27812 711 27822 745
rect 27856 711 27864 745
rect 28422 737 28474 749
rect 27812 677 27864 711
rect 27812 643 27822 677
rect 27856 643 27864 677
rect 27812 627 27864 643
rect 28035 684 28087 729
rect 28035 650 28043 684
rect 28077 650 28087 684
rect 28035 625 28087 650
rect 28117 671 28175 729
rect 28117 637 28129 671
rect 28163 637 28175 671
rect 28117 625 28175 637
rect 28205 701 28257 729
rect 28205 667 28215 701
rect 28249 667 28257 701
rect 28205 625 28257 667
rect 28422 703 28430 737
rect 28464 703 28474 737
rect 28422 669 28474 703
rect 28422 635 28430 669
rect 28464 635 28474 669
rect 28422 619 28474 635
rect 28504 737 28556 749
rect 28504 703 28514 737
rect 28548 703 28556 737
rect 28504 669 28556 703
rect 29618 745 29670 757
rect 29618 711 29626 745
rect 29660 711 29670 745
rect 29618 677 29670 711
rect 28504 635 28514 669
rect 28548 635 28556 669
rect 28504 619 28556 635
rect 29618 643 29626 677
rect 29660 643 29670 677
rect 29618 627 29670 643
rect 29700 745 29752 757
rect 29700 711 29710 745
rect 29744 711 29752 745
rect 30310 737 30362 749
rect 29700 677 29752 711
rect 29700 643 29710 677
rect 29744 643 29752 677
rect 29700 627 29752 643
rect 29923 684 29975 729
rect 29923 650 29931 684
rect 29965 650 29975 684
rect 29923 625 29975 650
rect 30005 671 30063 729
rect 30005 637 30017 671
rect 30051 637 30063 671
rect 30005 625 30063 637
rect 30093 701 30145 729
rect 30093 667 30103 701
rect 30137 667 30145 701
rect 30093 625 30145 667
rect 30310 703 30318 737
rect 30352 703 30362 737
rect 30310 669 30362 703
rect 30310 635 30318 669
rect 30352 635 30362 669
rect 30310 619 30362 635
rect 30392 737 30444 749
rect 30392 703 30402 737
rect 30436 703 30444 737
rect 30392 669 30444 703
rect 31506 745 31558 757
rect 31506 711 31514 745
rect 31548 711 31558 745
rect 31506 677 31558 711
rect 30392 635 30402 669
rect 30436 635 30444 669
rect 30392 619 30444 635
rect 31506 643 31514 677
rect 31548 643 31558 677
rect 31506 627 31558 643
rect 31588 745 31640 757
rect 31588 711 31598 745
rect 31632 711 31640 745
rect 32198 737 32250 749
rect 31588 677 31640 711
rect 31588 643 31598 677
rect 31632 643 31640 677
rect 31588 627 31640 643
rect 31811 684 31863 729
rect 31811 650 31819 684
rect 31853 650 31863 684
rect 31811 625 31863 650
rect 31893 671 31951 729
rect 31893 637 31905 671
rect 31939 637 31951 671
rect 31893 625 31951 637
rect 31981 701 32033 729
rect 31981 667 31991 701
rect 32025 667 32033 701
rect 31981 625 32033 667
rect 32198 703 32206 737
rect 32240 703 32250 737
rect 32198 669 32250 703
rect 32198 635 32206 669
rect 32240 635 32250 669
rect 32198 619 32250 635
rect 32280 737 32332 749
rect 32280 703 32290 737
rect 32324 703 32332 737
rect 32280 669 32332 703
rect 33394 745 33446 757
rect 33394 711 33402 745
rect 33436 711 33446 745
rect 33394 677 33446 711
rect 32280 635 32290 669
rect 32324 635 32332 669
rect 32280 619 32332 635
rect 33394 643 33402 677
rect 33436 643 33446 677
rect 33394 627 33446 643
rect 33476 745 33528 757
rect 33476 711 33486 745
rect 33520 711 33528 745
rect 34086 737 34138 749
rect 33476 677 33528 711
rect 33476 643 33486 677
rect 33520 643 33528 677
rect 33476 627 33528 643
rect 33699 684 33751 729
rect 33699 650 33707 684
rect 33741 650 33751 684
rect 33699 625 33751 650
rect 33781 671 33839 729
rect 33781 637 33793 671
rect 33827 637 33839 671
rect 33781 625 33839 637
rect 33869 701 33921 729
rect 33869 667 33879 701
rect 33913 667 33921 701
rect 33869 625 33921 667
rect 34086 703 34094 737
rect 34128 703 34138 737
rect 34086 669 34138 703
rect 34086 635 34094 669
rect 34128 635 34138 669
rect 34086 619 34138 635
rect 34168 737 34220 749
rect 34168 703 34178 737
rect 34212 703 34220 737
rect 34168 669 34220 703
rect 35282 745 35334 757
rect 35282 711 35290 745
rect 35324 711 35334 745
rect 35282 677 35334 711
rect 34168 635 34178 669
rect 34212 635 34220 669
rect 34168 619 34220 635
rect 35282 643 35290 677
rect 35324 643 35334 677
rect 35282 627 35334 643
rect 35364 745 35416 757
rect 35364 711 35374 745
rect 35408 711 35416 745
rect 35974 737 36026 749
rect 35364 677 35416 711
rect 35364 643 35374 677
rect 35408 643 35416 677
rect 35364 627 35416 643
rect 35587 684 35639 729
rect 35587 650 35595 684
rect 35629 650 35639 684
rect 35587 625 35639 650
rect 35669 671 35727 729
rect 35669 637 35681 671
rect 35715 637 35727 671
rect 35669 625 35727 637
rect 35757 701 35809 729
rect 35757 667 35767 701
rect 35801 667 35809 701
rect 35757 625 35809 667
rect 35974 703 35982 737
rect 36016 703 36026 737
rect 35974 669 36026 703
rect 35974 635 35982 669
rect 36016 635 36026 669
rect 35974 619 36026 635
rect 36056 737 36108 749
rect 36056 703 36066 737
rect 36100 703 36108 737
rect 36056 669 36108 703
rect 37170 745 37222 757
rect 37170 711 37178 745
rect 37212 711 37222 745
rect 37170 677 37222 711
rect 36056 635 36066 669
rect 36100 635 36108 669
rect 36056 619 36108 635
rect 37170 643 37178 677
rect 37212 643 37222 677
rect 37170 627 37222 643
rect 37252 745 37304 757
rect 37252 711 37262 745
rect 37296 711 37304 745
rect 37862 737 37914 749
rect 37252 677 37304 711
rect 37252 643 37262 677
rect 37296 643 37304 677
rect 37252 627 37304 643
rect 37475 684 37527 729
rect 37475 650 37483 684
rect 37517 650 37527 684
rect 37475 625 37527 650
rect 37557 671 37615 729
rect 37557 637 37569 671
rect 37603 637 37615 671
rect 37557 625 37615 637
rect 37645 701 37697 729
rect 37645 667 37655 701
rect 37689 667 37697 701
rect 37645 625 37697 667
rect 37862 703 37870 737
rect 37904 703 37914 737
rect 37862 669 37914 703
rect 37862 635 37870 669
rect 37904 635 37914 669
rect 37862 619 37914 635
rect 37944 737 37996 749
rect 37944 703 37954 737
rect 37988 703 37996 737
rect 37944 669 37996 703
rect 39058 745 39110 757
rect 39058 711 39066 745
rect 39100 711 39110 745
rect 39058 677 39110 711
rect 37944 635 37954 669
rect 37988 635 37996 669
rect 37944 619 37996 635
rect 39058 643 39066 677
rect 39100 643 39110 677
rect 39058 627 39110 643
rect 39140 745 39192 757
rect 39140 711 39150 745
rect 39184 711 39192 745
rect 39750 737 39802 749
rect 39140 677 39192 711
rect 39140 643 39150 677
rect 39184 643 39192 677
rect 39140 627 39192 643
rect 39363 684 39415 729
rect 39363 650 39371 684
rect 39405 650 39415 684
rect 39363 625 39415 650
rect 39445 671 39503 729
rect 39445 637 39457 671
rect 39491 637 39503 671
rect 39445 625 39503 637
rect 39533 701 39585 729
rect 39533 667 39543 701
rect 39577 667 39585 701
rect 39533 625 39585 667
rect 39750 703 39758 737
rect 39792 703 39802 737
rect 39750 669 39802 703
rect 39750 635 39758 669
rect 39792 635 39802 669
rect 39750 619 39802 635
rect 39832 737 39884 749
rect 39832 703 39842 737
rect 39876 703 39884 737
rect 39832 669 39884 703
rect 40946 745 40998 757
rect 40946 711 40954 745
rect 40988 711 40998 745
rect 40946 677 40998 711
rect 39832 635 39842 669
rect 39876 635 39884 669
rect 39832 619 39884 635
rect 40946 643 40954 677
rect 40988 643 40998 677
rect 40946 627 40998 643
rect 41028 745 41080 757
rect 41028 711 41038 745
rect 41072 711 41080 745
rect 41638 737 41690 749
rect 41028 677 41080 711
rect 41028 643 41038 677
rect 41072 643 41080 677
rect 41028 627 41080 643
rect 41251 684 41303 729
rect 41251 650 41259 684
rect 41293 650 41303 684
rect 41251 625 41303 650
rect 41333 671 41391 729
rect 41333 637 41345 671
rect 41379 637 41391 671
rect 41333 625 41391 637
rect 41421 701 41473 729
rect 41421 667 41431 701
rect 41465 667 41473 701
rect 41421 625 41473 667
rect 41638 703 41646 737
rect 41680 703 41690 737
rect 41638 669 41690 703
rect 41638 635 41646 669
rect 41680 635 41690 669
rect 41638 619 41690 635
rect 41720 737 41772 749
rect 41720 703 41730 737
rect 41764 703 41772 737
rect 41720 669 41772 703
rect 42834 745 42886 757
rect 42834 711 42842 745
rect 42876 711 42886 745
rect 42834 677 42886 711
rect 41720 635 41730 669
rect 41764 635 41772 669
rect 41720 619 41772 635
rect 42834 643 42842 677
rect 42876 643 42886 677
rect 42834 627 42886 643
rect 42916 745 42968 757
rect 42916 711 42926 745
rect 42960 711 42968 745
rect 43526 737 43578 749
rect 42916 677 42968 711
rect 42916 643 42926 677
rect 42960 643 42968 677
rect 42916 627 42968 643
rect 43139 684 43191 729
rect 43139 650 43147 684
rect 43181 650 43191 684
rect 43139 625 43191 650
rect 43221 671 43279 729
rect 43221 637 43233 671
rect 43267 637 43279 671
rect 43221 625 43279 637
rect 43309 701 43361 729
rect 43309 667 43319 701
rect 43353 667 43361 701
rect 43309 625 43361 667
rect 43526 703 43534 737
rect 43568 703 43578 737
rect 43526 669 43578 703
rect 43526 635 43534 669
rect 43568 635 43578 669
rect 43526 619 43578 635
rect 43608 737 43660 749
rect 43608 703 43618 737
rect 43652 703 43660 737
rect 43608 669 43660 703
rect 44722 745 44774 757
rect 44722 711 44730 745
rect 44764 711 44774 745
rect 44722 677 44774 711
rect 43608 635 43618 669
rect 43652 635 43660 669
rect 43608 619 43660 635
rect 44722 643 44730 677
rect 44764 643 44774 677
rect 44722 627 44774 643
rect 44804 745 44856 757
rect 44804 711 44814 745
rect 44848 711 44856 745
rect 45408 737 45460 749
rect 44804 677 44856 711
rect 44804 643 44814 677
rect 44848 643 44856 677
rect 44804 627 44856 643
rect 45027 684 45079 729
rect 45027 650 45035 684
rect 45069 650 45079 684
rect 45027 625 45079 650
rect 45109 671 45167 729
rect 45109 637 45121 671
rect 45155 637 45167 671
rect 45109 625 45167 637
rect 45197 701 45249 729
rect 45197 667 45207 701
rect 45241 667 45249 701
rect 45197 625 45249 667
rect 45408 703 45416 737
rect 45450 703 45460 737
rect 45408 669 45460 703
rect 45408 635 45416 669
rect 45450 635 45460 669
rect 45408 619 45460 635
rect 45490 737 45542 749
rect 45490 703 45500 737
rect 45534 703 45542 737
rect 45490 669 45542 703
rect 46604 745 46656 757
rect 46604 711 46612 745
rect 46646 711 46656 745
rect 46604 677 46656 711
rect 45490 635 45500 669
rect 45534 635 45542 669
rect 45490 619 45542 635
rect 46604 643 46612 677
rect 46646 643 46656 677
rect 46604 627 46656 643
rect 46686 745 46738 757
rect 46686 711 46696 745
rect 46730 711 46738 745
rect 47296 737 47348 749
rect 46686 677 46738 711
rect 46686 643 46696 677
rect 46730 643 46738 677
rect 46686 627 46738 643
rect 46909 684 46961 729
rect 46909 650 46917 684
rect 46951 650 46961 684
rect 46909 625 46961 650
rect 46991 671 47049 729
rect 46991 637 47003 671
rect 47037 637 47049 671
rect 46991 625 47049 637
rect 47079 701 47131 729
rect 47079 667 47089 701
rect 47123 667 47131 701
rect 47079 625 47131 667
rect 47296 703 47304 737
rect 47338 703 47348 737
rect 47296 669 47348 703
rect 47296 635 47304 669
rect 47338 635 47348 669
rect 47296 619 47348 635
rect 47378 737 47430 749
rect 47378 703 47388 737
rect 47422 703 47430 737
rect 47378 669 47430 703
rect 48492 745 48544 757
rect 48492 711 48500 745
rect 48534 711 48544 745
rect 48492 677 48544 711
rect 47378 635 47388 669
rect 47422 635 47430 669
rect 47378 619 47430 635
rect 48492 643 48500 677
rect 48534 643 48544 677
rect 48492 627 48544 643
rect 48574 745 48626 757
rect 48574 711 48584 745
rect 48618 711 48626 745
rect 49184 737 49236 749
rect 48574 677 48626 711
rect 48574 643 48584 677
rect 48618 643 48626 677
rect 48574 627 48626 643
rect 48797 684 48849 729
rect 48797 650 48805 684
rect 48839 650 48849 684
rect 48797 625 48849 650
rect 48879 671 48937 729
rect 48879 637 48891 671
rect 48925 637 48937 671
rect 48879 625 48937 637
rect 48967 701 49019 729
rect 48967 667 48977 701
rect 49011 667 49019 701
rect 48967 625 49019 667
rect 49184 703 49192 737
rect 49226 703 49236 737
rect 49184 669 49236 703
rect 49184 635 49192 669
rect 49226 635 49236 669
rect 49184 619 49236 635
rect 49266 737 49318 749
rect 49266 703 49276 737
rect 49310 703 49318 737
rect 49266 669 49318 703
rect 50380 745 50432 757
rect 50380 711 50388 745
rect 50422 711 50432 745
rect 50380 677 50432 711
rect 49266 635 49276 669
rect 49310 635 49318 669
rect 49266 619 49318 635
rect 50380 643 50388 677
rect 50422 643 50432 677
rect 50380 627 50432 643
rect 50462 745 50514 757
rect 50462 711 50472 745
rect 50506 711 50514 745
rect 51072 737 51124 749
rect 50462 677 50514 711
rect 50462 643 50472 677
rect 50506 643 50514 677
rect 50462 627 50514 643
rect 50685 684 50737 729
rect 50685 650 50693 684
rect 50727 650 50737 684
rect 50685 625 50737 650
rect 50767 671 50825 729
rect 50767 637 50779 671
rect 50813 637 50825 671
rect 50767 625 50825 637
rect 50855 701 50907 729
rect 50855 667 50865 701
rect 50899 667 50907 701
rect 50855 625 50907 667
rect 51072 703 51080 737
rect 51114 703 51124 737
rect 51072 669 51124 703
rect 51072 635 51080 669
rect 51114 635 51124 669
rect 51072 619 51124 635
rect 51154 737 51206 749
rect 51154 703 51164 737
rect 51198 703 51206 737
rect 51154 669 51206 703
rect 52268 745 52320 757
rect 52268 711 52276 745
rect 52310 711 52320 745
rect 52268 677 52320 711
rect 51154 635 51164 669
rect 51198 635 51206 669
rect 51154 619 51206 635
rect 52268 643 52276 677
rect 52310 643 52320 677
rect 52268 627 52320 643
rect 52350 745 52402 757
rect 52350 711 52360 745
rect 52394 711 52402 745
rect 52960 737 53012 749
rect 52350 677 52402 711
rect 52350 643 52360 677
rect 52394 643 52402 677
rect 52350 627 52402 643
rect 52573 684 52625 729
rect 52573 650 52581 684
rect 52615 650 52625 684
rect 52573 625 52625 650
rect 52655 671 52713 729
rect 52655 637 52667 671
rect 52701 637 52713 671
rect 52655 625 52713 637
rect 52743 701 52795 729
rect 52743 667 52753 701
rect 52787 667 52795 701
rect 52743 625 52795 667
rect 52960 703 52968 737
rect 53002 703 53012 737
rect 52960 669 53012 703
rect 52960 635 52968 669
rect 53002 635 53012 669
rect 52960 619 53012 635
rect 53042 737 53094 749
rect 53042 703 53052 737
rect 53086 703 53094 737
rect 53042 669 53094 703
rect 54156 745 54208 757
rect 54156 711 54164 745
rect 54198 711 54208 745
rect 54156 677 54208 711
rect 53042 635 53052 669
rect 53086 635 53094 669
rect 53042 619 53094 635
rect 54156 643 54164 677
rect 54198 643 54208 677
rect 54156 627 54208 643
rect 54238 745 54290 757
rect 54238 711 54248 745
rect 54282 711 54290 745
rect 54848 737 54900 749
rect 54238 677 54290 711
rect 54238 643 54248 677
rect 54282 643 54290 677
rect 54238 627 54290 643
rect 54461 684 54513 729
rect 54461 650 54469 684
rect 54503 650 54513 684
rect 54461 625 54513 650
rect 54543 671 54601 729
rect 54543 637 54555 671
rect 54589 637 54601 671
rect 54543 625 54601 637
rect 54631 701 54683 729
rect 54631 667 54641 701
rect 54675 667 54683 701
rect 54631 625 54683 667
rect 54848 703 54856 737
rect 54890 703 54900 737
rect 54848 669 54900 703
rect 54848 635 54856 669
rect 54890 635 54900 669
rect 54848 619 54900 635
rect 54930 737 54982 749
rect 54930 703 54940 737
rect 54974 703 54982 737
rect 54930 669 54982 703
rect 56044 745 56096 757
rect 56044 711 56052 745
rect 56086 711 56096 745
rect 56044 677 56096 711
rect 54930 635 54940 669
rect 54974 635 54982 669
rect 54930 619 54982 635
rect 56044 643 56052 677
rect 56086 643 56096 677
rect 56044 627 56096 643
rect 56126 745 56178 757
rect 56126 711 56136 745
rect 56170 711 56178 745
rect 56736 737 56788 749
rect 56126 677 56178 711
rect 56126 643 56136 677
rect 56170 643 56178 677
rect 56126 627 56178 643
rect 56349 684 56401 729
rect 56349 650 56357 684
rect 56391 650 56401 684
rect 56349 625 56401 650
rect 56431 671 56489 729
rect 56431 637 56443 671
rect 56477 637 56489 671
rect 56431 625 56489 637
rect 56519 701 56571 729
rect 56519 667 56529 701
rect 56563 667 56571 701
rect 56519 625 56571 667
rect 56736 703 56744 737
rect 56778 703 56788 737
rect 56736 669 56788 703
rect 56736 635 56744 669
rect 56778 635 56788 669
rect 56736 619 56788 635
rect 56818 737 56870 749
rect 56818 703 56828 737
rect 56862 703 56870 737
rect 56818 669 56870 703
rect 57932 745 57984 757
rect 57932 711 57940 745
rect 57974 711 57984 745
rect 57932 677 57984 711
rect 56818 635 56828 669
rect 56862 635 56870 669
rect 56818 619 56870 635
rect 57932 643 57940 677
rect 57974 643 57984 677
rect 57932 627 57984 643
rect 58014 745 58066 757
rect 58014 711 58024 745
rect 58058 711 58066 745
rect 58624 737 58676 749
rect 58014 677 58066 711
rect 58014 643 58024 677
rect 58058 643 58066 677
rect 58014 627 58066 643
rect 58237 684 58289 729
rect 58237 650 58245 684
rect 58279 650 58289 684
rect 58237 625 58289 650
rect 58319 671 58377 729
rect 58319 637 58331 671
rect 58365 637 58377 671
rect 58319 625 58377 637
rect 58407 701 58459 729
rect 58407 667 58417 701
rect 58451 667 58459 701
rect 58407 625 58459 667
rect 58624 703 58632 737
rect 58666 703 58676 737
rect 58624 669 58676 703
rect 58624 635 58632 669
rect 58666 635 58676 669
rect 58624 619 58676 635
rect 58706 737 58758 749
rect 58706 703 58716 737
rect 58750 703 58758 737
rect 58706 669 58758 703
rect 59820 745 59872 757
rect 59820 711 59828 745
rect 59862 711 59872 745
rect 59820 677 59872 711
rect 58706 635 58716 669
rect 58750 635 58758 669
rect 58706 619 58758 635
rect 59820 643 59828 677
rect 59862 643 59872 677
rect 59820 627 59872 643
rect 59902 745 59954 757
rect 59902 711 59912 745
rect 59946 711 59954 745
rect 59902 677 59954 711
rect 59902 643 59912 677
rect 59946 643 59954 677
rect 59902 627 59954 643
rect 60125 684 60177 729
rect 60125 650 60133 684
rect 60167 650 60177 684
rect 60125 625 60177 650
rect 60207 671 60265 729
rect 60207 637 60219 671
rect 60253 637 60265 671
rect 60207 625 60265 637
rect 60295 701 60347 729
rect 60295 667 60305 701
rect 60339 667 60347 701
rect 60295 625 60347 667
rect 608 488 670 502
rect 608 454 620 488
rect 654 454 670 488
rect 608 420 670 454
rect 608 386 620 420
rect 654 386 670 420
rect 608 372 670 386
rect 700 488 766 502
rect 700 454 716 488
rect 750 454 766 488
rect 700 420 766 454
rect 700 386 716 420
rect 750 386 766 420
rect 700 372 766 386
rect 796 488 858 502
rect 796 454 812 488
rect 846 454 858 488
rect 796 420 858 454
rect 796 386 812 420
rect 846 386 858 420
rect 796 372 858 386
rect 2496 488 2558 502
rect 2496 454 2508 488
rect 2542 454 2558 488
rect 2496 420 2558 454
rect 2496 386 2508 420
rect 2542 386 2558 420
rect 2496 372 2558 386
rect 2588 488 2654 502
rect 2588 454 2604 488
rect 2638 454 2654 488
rect 2588 420 2654 454
rect 2588 386 2604 420
rect 2638 386 2654 420
rect 2588 372 2654 386
rect 2684 488 2746 502
rect 2684 454 2700 488
rect 2734 454 2746 488
rect 2684 420 2746 454
rect 2684 386 2700 420
rect 2734 386 2746 420
rect 2684 372 2746 386
rect 4384 488 4446 502
rect 4384 454 4396 488
rect 4430 454 4446 488
rect 4384 420 4446 454
rect 4384 386 4396 420
rect 4430 386 4446 420
rect 4384 372 4446 386
rect 4476 488 4542 502
rect 4476 454 4492 488
rect 4526 454 4542 488
rect 4476 420 4542 454
rect 4476 386 4492 420
rect 4526 386 4542 420
rect 4476 372 4542 386
rect 4572 488 4634 502
rect 4572 454 4588 488
rect 4622 454 4634 488
rect 4572 420 4634 454
rect 4572 386 4588 420
rect 4622 386 4634 420
rect 4572 372 4634 386
rect 6272 488 6334 502
rect 6272 454 6284 488
rect 6318 454 6334 488
rect 6272 420 6334 454
rect 6272 386 6284 420
rect 6318 386 6334 420
rect 6272 372 6334 386
rect 6364 488 6430 502
rect 6364 454 6380 488
rect 6414 454 6430 488
rect 6364 420 6430 454
rect 6364 386 6380 420
rect 6414 386 6430 420
rect 6364 372 6430 386
rect 6460 488 6522 502
rect 6460 454 6476 488
rect 6510 454 6522 488
rect 6460 420 6522 454
rect 6460 386 6476 420
rect 6510 386 6522 420
rect 6460 372 6522 386
rect 8160 488 8222 502
rect 8160 454 8172 488
rect 8206 454 8222 488
rect 8160 420 8222 454
rect 8160 386 8172 420
rect 8206 386 8222 420
rect 8160 372 8222 386
rect 8252 488 8318 502
rect 8252 454 8268 488
rect 8302 454 8318 488
rect 8252 420 8318 454
rect 8252 386 8268 420
rect 8302 386 8318 420
rect 8252 372 8318 386
rect 8348 488 8410 502
rect 8348 454 8364 488
rect 8398 454 8410 488
rect 8348 420 8410 454
rect 8348 386 8364 420
rect 8398 386 8410 420
rect 8348 372 8410 386
rect 10048 488 10110 502
rect 10048 454 10060 488
rect 10094 454 10110 488
rect 10048 420 10110 454
rect 10048 386 10060 420
rect 10094 386 10110 420
rect 10048 372 10110 386
rect 10140 488 10206 502
rect 10140 454 10156 488
rect 10190 454 10206 488
rect 10140 420 10206 454
rect 10140 386 10156 420
rect 10190 386 10206 420
rect 10140 372 10206 386
rect 10236 488 10298 502
rect 10236 454 10252 488
rect 10286 454 10298 488
rect 10236 420 10298 454
rect 10236 386 10252 420
rect 10286 386 10298 420
rect 10236 372 10298 386
rect 11936 488 11998 502
rect 11936 454 11948 488
rect 11982 454 11998 488
rect 11936 420 11998 454
rect 11936 386 11948 420
rect 11982 386 11998 420
rect 11936 372 11998 386
rect 12028 488 12094 502
rect 12028 454 12044 488
rect 12078 454 12094 488
rect 12028 420 12094 454
rect 12028 386 12044 420
rect 12078 386 12094 420
rect 12028 372 12094 386
rect 12124 488 12186 502
rect 12124 454 12140 488
rect 12174 454 12186 488
rect 12124 420 12186 454
rect 12124 386 12140 420
rect 12174 386 12186 420
rect 12124 372 12186 386
rect 13824 488 13886 502
rect 13824 454 13836 488
rect 13870 454 13886 488
rect 13824 420 13886 454
rect 13824 386 13836 420
rect 13870 386 13886 420
rect 13824 372 13886 386
rect 13916 488 13982 502
rect 13916 454 13932 488
rect 13966 454 13982 488
rect 13916 420 13982 454
rect 13916 386 13932 420
rect 13966 386 13982 420
rect 13916 372 13982 386
rect 14012 488 14074 502
rect 14012 454 14028 488
rect 14062 454 14074 488
rect 14012 420 14074 454
rect 14012 386 14028 420
rect 14062 386 14074 420
rect 14012 372 14074 386
rect 15706 488 15768 502
rect 15706 454 15718 488
rect 15752 454 15768 488
rect 15706 420 15768 454
rect 15706 386 15718 420
rect 15752 386 15768 420
rect 15706 372 15768 386
rect 15798 488 15864 502
rect 15798 454 15814 488
rect 15848 454 15864 488
rect 15798 420 15864 454
rect 15798 386 15814 420
rect 15848 386 15864 420
rect 15798 372 15864 386
rect 15894 488 15956 502
rect 15894 454 15910 488
rect 15944 454 15956 488
rect 15894 420 15956 454
rect 15894 386 15910 420
rect 15944 386 15956 420
rect 15894 372 15956 386
rect 17594 488 17656 502
rect 17594 454 17606 488
rect 17640 454 17656 488
rect 17594 420 17656 454
rect 17594 386 17606 420
rect 17640 386 17656 420
rect 17594 372 17656 386
rect 17686 488 17752 502
rect 17686 454 17702 488
rect 17736 454 17752 488
rect 17686 420 17752 454
rect 17686 386 17702 420
rect 17736 386 17752 420
rect 17686 372 17752 386
rect 17782 488 17844 502
rect 17782 454 17798 488
rect 17832 454 17844 488
rect 17782 420 17844 454
rect 17782 386 17798 420
rect 17832 386 17844 420
rect 17782 372 17844 386
rect 19482 488 19544 502
rect 19482 454 19494 488
rect 19528 454 19544 488
rect 19482 420 19544 454
rect 19482 386 19494 420
rect 19528 386 19544 420
rect 19482 372 19544 386
rect 19574 488 19640 502
rect 19574 454 19590 488
rect 19624 454 19640 488
rect 19574 420 19640 454
rect 19574 386 19590 420
rect 19624 386 19640 420
rect 19574 372 19640 386
rect 19670 488 19732 502
rect 19670 454 19686 488
rect 19720 454 19732 488
rect 19670 420 19732 454
rect 19670 386 19686 420
rect 19720 386 19732 420
rect 19670 372 19732 386
rect 21370 488 21432 502
rect 21370 454 21382 488
rect 21416 454 21432 488
rect 21370 420 21432 454
rect 21370 386 21382 420
rect 21416 386 21432 420
rect 21370 372 21432 386
rect 21462 488 21528 502
rect 21462 454 21478 488
rect 21512 454 21528 488
rect 21462 420 21528 454
rect 21462 386 21478 420
rect 21512 386 21528 420
rect 21462 372 21528 386
rect 21558 488 21620 502
rect 21558 454 21574 488
rect 21608 454 21620 488
rect 21558 420 21620 454
rect 21558 386 21574 420
rect 21608 386 21620 420
rect 21558 372 21620 386
rect 23258 488 23320 502
rect 23258 454 23270 488
rect 23304 454 23320 488
rect 23258 420 23320 454
rect 23258 386 23270 420
rect 23304 386 23320 420
rect 23258 372 23320 386
rect 23350 488 23416 502
rect 23350 454 23366 488
rect 23400 454 23416 488
rect 23350 420 23416 454
rect 23350 386 23366 420
rect 23400 386 23416 420
rect 23350 372 23416 386
rect 23446 488 23508 502
rect 23446 454 23462 488
rect 23496 454 23508 488
rect 23446 420 23508 454
rect 23446 386 23462 420
rect 23496 386 23508 420
rect 23446 372 23508 386
rect 25146 488 25208 502
rect 25146 454 25158 488
rect 25192 454 25208 488
rect 25146 420 25208 454
rect 25146 386 25158 420
rect 25192 386 25208 420
rect 25146 372 25208 386
rect 25238 488 25304 502
rect 25238 454 25254 488
rect 25288 454 25304 488
rect 25238 420 25304 454
rect 25238 386 25254 420
rect 25288 386 25304 420
rect 25238 372 25304 386
rect 25334 488 25396 502
rect 25334 454 25350 488
rect 25384 454 25396 488
rect 25334 420 25396 454
rect 25334 386 25350 420
rect 25384 386 25396 420
rect 25334 372 25396 386
rect 27034 488 27096 502
rect 27034 454 27046 488
rect 27080 454 27096 488
rect 27034 420 27096 454
rect 27034 386 27046 420
rect 27080 386 27096 420
rect 27034 372 27096 386
rect 27126 488 27192 502
rect 27126 454 27142 488
rect 27176 454 27192 488
rect 27126 420 27192 454
rect 27126 386 27142 420
rect 27176 386 27192 420
rect 27126 372 27192 386
rect 27222 488 27284 502
rect 27222 454 27238 488
rect 27272 454 27284 488
rect 27222 420 27284 454
rect 27222 386 27238 420
rect 27272 386 27284 420
rect 27222 372 27284 386
rect 28922 488 28984 502
rect 28922 454 28934 488
rect 28968 454 28984 488
rect 28922 420 28984 454
rect 28922 386 28934 420
rect 28968 386 28984 420
rect 28922 372 28984 386
rect 29014 488 29080 502
rect 29014 454 29030 488
rect 29064 454 29080 488
rect 29014 420 29080 454
rect 29014 386 29030 420
rect 29064 386 29080 420
rect 29014 372 29080 386
rect 29110 488 29172 502
rect 29110 454 29126 488
rect 29160 454 29172 488
rect 29110 420 29172 454
rect 29110 386 29126 420
rect 29160 386 29172 420
rect 29110 372 29172 386
rect 30810 488 30872 502
rect 30810 454 30822 488
rect 30856 454 30872 488
rect 30810 420 30872 454
rect 30810 386 30822 420
rect 30856 386 30872 420
rect 30810 372 30872 386
rect 30902 488 30968 502
rect 30902 454 30918 488
rect 30952 454 30968 488
rect 30902 420 30968 454
rect 30902 386 30918 420
rect 30952 386 30968 420
rect 30902 372 30968 386
rect 30998 488 31060 502
rect 30998 454 31014 488
rect 31048 454 31060 488
rect 30998 420 31060 454
rect 30998 386 31014 420
rect 31048 386 31060 420
rect 30998 372 31060 386
rect 32698 488 32760 502
rect 32698 454 32710 488
rect 32744 454 32760 488
rect 32698 420 32760 454
rect 32698 386 32710 420
rect 32744 386 32760 420
rect 32698 372 32760 386
rect 32790 488 32856 502
rect 32790 454 32806 488
rect 32840 454 32856 488
rect 32790 420 32856 454
rect 32790 386 32806 420
rect 32840 386 32856 420
rect 32790 372 32856 386
rect 32886 488 32948 502
rect 32886 454 32902 488
rect 32936 454 32948 488
rect 32886 420 32948 454
rect 32886 386 32902 420
rect 32936 386 32948 420
rect 32886 372 32948 386
rect 34586 488 34648 502
rect 34586 454 34598 488
rect 34632 454 34648 488
rect 34586 420 34648 454
rect 34586 386 34598 420
rect 34632 386 34648 420
rect 34586 372 34648 386
rect 34678 488 34744 502
rect 34678 454 34694 488
rect 34728 454 34744 488
rect 34678 420 34744 454
rect 34678 386 34694 420
rect 34728 386 34744 420
rect 34678 372 34744 386
rect 34774 488 34836 502
rect 34774 454 34790 488
rect 34824 454 34836 488
rect 34774 420 34836 454
rect 34774 386 34790 420
rect 34824 386 34836 420
rect 34774 372 34836 386
rect 36474 488 36536 502
rect 36474 454 36486 488
rect 36520 454 36536 488
rect 36474 420 36536 454
rect 36474 386 36486 420
rect 36520 386 36536 420
rect 36474 372 36536 386
rect 36566 488 36632 502
rect 36566 454 36582 488
rect 36616 454 36632 488
rect 36566 420 36632 454
rect 36566 386 36582 420
rect 36616 386 36632 420
rect 36566 372 36632 386
rect 36662 488 36724 502
rect 36662 454 36678 488
rect 36712 454 36724 488
rect 36662 420 36724 454
rect 36662 386 36678 420
rect 36712 386 36724 420
rect 36662 372 36724 386
rect 38362 488 38424 502
rect 38362 454 38374 488
rect 38408 454 38424 488
rect 38362 420 38424 454
rect 38362 386 38374 420
rect 38408 386 38424 420
rect 38362 372 38424 386
rect 38454 488 38520 502
rect 38454 454 38470 488
rect 38504 454 38520 488
rect 38454 420 38520 454
rect 38454 386 38470 420
rect 38504 386 38520 420
rect 38454 372 38520 386
rect 38550 488 38612 502
rect 38550 454 38566 488
rect 38600 454 38612 488
rect 38550 420 38612 454
rect 38550 386 38566 420
rect 38600 386 38612 420
rect 38550 372 38612 386
rect 40250 488 40312 502
rect 40250 454 40262 488
rect 40296 454 40312 488
rect 40250 420 40312 454
rect 40250 386 40262 420
rect 40296 386 40312 420
rect 40250 372 40312 386
rect 40342 488 40408 502
rect 40342 454 40358 488
rect 40392 454 40408 488
rect 40342 420 40408 454
rect 40342 386 40358 420
rect 40392 386 40408 420
rect 40342 372 40408 386
rect 40438 488 40500 502
rect 40438 454 40454 488
rect 40488 454 40500 488
rect 40438 420 40500 454
rect 40438 386 40454 420
rect 40488 386 40500 420
rect 40438 372 40500 386
rect 42138 488 42200 502
rect 42138 454 42150 488
rect 42184 454 42200 488
rect 42138 420 42200 454
rect 42138 386 42150 420
rect 42184 386 42200 420
rect 42138 372 42200 386
rect 42230 488 42296 502
rect 42230 454 42246 488
rect 42280 454 42296 488
rect 42230 420 42296 454
rect 42230 386 42246 420
rect 42280 386 42296 420
rect 42230 372 42296 386
rect 42326 488 42388 502
rect 42326 454 42342 488
rect 42376 454 42388 488
rect 42326 420 42388 454
rect 42326 386 42342 420
rect 42376 386 42388 420
rect 42326 372 42388 386
rect 44026 488 44088 502
rect 44026 454 44038 488
rect 44072 454 44088 488
rect 44026 420 44088 454
rect 44026 386 44038 420
rect 44072 386 44088 420
rect 44026 372 44088 386
rect 44118 488 44184 502
rect 44118 454 44134 488
rect 44168 454 44184 488
rect 44118 420 44184 454
rect 44118 386 44134 420
rect 44168 386 44184 420
rect 44118 372 44184 386
rect 44214 488 44276 502
rect 44214 454 44230 488
rect 44264 454 44276 488
rect 44214 420 44276 454
rect 44214 386 44230 420
rect 44264 386 44276 420
rect 44214 372 44276 386
rect 45908 488 45970 502
rect 45908 454 45920 488
rect 45954 454 45970 488
rect 45908 420 45970 454
rect 45908 386 45920 420
rect 45954 386 45970 420
rect 45908 372 45970 386
rect 46000 488 46066 502
rect 46000 454 46016 488
rect 46050 454 46066 488
rect 46000 420 46066 454
rect 46000 386 46016 420
rect 46050 386 46066 420
rect 46000 372 46066 386
rect 46096 488 46158 502
rect 46096 454 46112 488
rect 46146 454 46158 488
rect 46096 420 46158 454
rect 46096 386 46112 420
rect 46146 386 46158 420
rect 46096 372 46158 386
rect 47796 488 47858 502
rect 47796 454 47808 488
rect 47842 454 47858 488
rect 47796 420 47858 454
rect 47796 386 47808 420
rect 47842 386 47858 420
rect 47796 372 47858 386
rect 47888 488 47954 502
rect 47888 454 47904 488
rect 47938 454 47954 488
rect 47888 420 47954 454
rect 47888 386 47904 420
rect 47938 386 47954 420
rect 47888 372 47954 386
rect 47984 488 48046 502
rect 47984 454 48000 488
rect 48034 454 48046 488
rect 47984 420 48046 454
rect 47984 386 48000 420
rect 48034 386 48046 420
rect 47984 372 48046 386
rect 49684 488 49746 502
rect 49684 454 49696 488
rect 49730 454 49746 488
rect 49684 420 49746 454
rect 49684 386 49696 420
rect 49730 386 49746 420
rect 49684 372 49746 386
rect 49776 488 49842 502
rect 49776 454 49792 488
rect 49826 454 49842 488
rect 49776 420 49842 454
rect 49776 386 49792 420
rect 49826 386 49842 420
rect 49776 372 49842 386
rect 49872 488 49934 502
rect 49872 454 49888 488
rect 49922 454 49934 488
rect 49872 420 49934 454
rect 49872 386 49888 420
rect 49922 386 49934 420
rect 49872 372 49934 386
rect 51572 488 51634 502
rect 51572 454 51584 488
rect 51618 454 51634 488
rect 51572 420 51634 454
rect 51572 386 51584 420
rect 51618 386 51634 420
rect 51572 372 51634 386
rect 51664 488 51730 502
rect 51664 454 51680 488
rect 51714 454 51730 488
rect 51664 420 51730 454
rect 51664 386 51680 420
rect 51714 386 51730 420
rect 51664 372 51730 386
rect 51760 488 51822 502
rect 51760 454 51776 488
rect 51810 454 51822 488
rect 51760 420 51822 454
rect 51760 386 51776 420
rect 51810 386 51822 420
rect 51760 372 51822 386
rect 53460 488 53522 502
rect 53460 454 53472 488
rect 53506 454 53522 488
rect 53460 420 53522 454
rect 53460 386 53472 420
rect 53506 386 53522 420
rect 53460 372 53522 386
rect 53552 488 53618 502
rect 53552 454 53568 488
rect 53602 454 53618 488
rect 53552 420 53618 454
rect 53552 386 53568 420
rect 53602 386 53618 420
rect 53552 372 53618 386
rect 53648 488 53710 502
rect 53648 454 53664 488
rect 53698 454 53710 488
rect 53648 420 53710 454
rect 53648 386 53664 420
rect 53698 386 53710 420
rect 53648 372 53710 386
rect 55348 488 55410 502
rect 55348 454 55360 488
rect 55394 454 55410 488
rect 55348 420 55410 454
rect 55348 386 55360 420
rect 55394 386 55410 420
rect 55348 372 55410 386
rect 55440 488 55506 502
rect 55440 454 55456 488
rect 55490 454 55506 488
rect 55440 420 55506 454
rect 55440 386 55456 420
rect 55490 386 55506 420
rect 55440 372 55506 386
rect 55536 488 55598 502
rect 55536 454 55552 488
rect 55586 454 55598 488
rect 55536 420 55598 454
rect 55536 386 55552 420
rect 55586 386 55598 420
rect 55536 372 55598 386
rect 57236 488 57298 502
rect 57236 454 57248 488
rect 57282 454 57298 488
rect 57236 420 57298 454
rect 57236 386 57248 420
rect 57282 386 57298 420
rect 57236 372 57298 386
rect 57328 488 57394 502
rect 57328 454 57344 488
rect 57378 454 57394 488
rect 57328 420 57394 454
rect 57328 386 57344 420
rect 57378 386 57394 420
rect 57328 372 57394 386
rect 57424 488 57486 502
rect 57424 454 57440 488
rect 57474 454 57486 488
rect 57424 420 57486 454
rect 57424 386 57440 420
rect 57474 386 57486 420
rect 57424 372 57486 386
rect 59124 488 59186 502
rect 59124 454 59136 488
rect 59170 454 59186 488
rect 59124 420 59186 454
rect 59124 386 59136 420
rect 59170 386 59186 420
rect 59124 372 59186 386
rect 59216 488 59282 502
rect 59216 454 59232 488
rect 59266 454 59282 488
rect 59216 420 59282 454
rect 59216 386 59232 420
rect 59266 386 59282 420
rect 59216 372 59282 386
rect 59312 488 59374 502
rect 59312 454 59328 488
rect 59362 454 59374 488
rect 59312 420 59374 454
rect 59312 386 59328 420
rect 59362 386 59374 420
rect 59312 372 59374 386
<< pdiff >>
rect 624 6723 686 6738
rect 624 6689 636 6723
rect 670 6689 686 6723
rect 624 6655 686 6689
rect 624 6621 636 6655
rect 670 6621 686 6655
rect 624 6587 686 6621
rect 298 6563 356 6578
rect 28 6545 80 6563
rect -365 6500 -313 6523
rect -365 6466 -357 6500
rect -323 6466 -313 6500
rect -365 6419 -313 6466
rect -365 6385 -357 6419
rect -323 6385 -313 6419
rect -365 6365 -313 6385
rect -283 6487 -225 6523
rect -283 6453 -271 6487
rect -237 6453 -225 6487
rect -283 6419 -225 6453
rect -283 6385 -271 6419
rect -237 6385 -225 6419
rect -283 6365 -225 6385
rect -195 6487 -143 6523
rect -195 6453 -185 6487
rect -151 6453 -143 6487
rect -195 6419 -143 6453
rect -195 6385 -185 6419
rect -151 6385 -143 6419
rect -195 6365 -143 6385
rect 28 6511 36 6545
rect 70 6511 80 6545
rect 28 6477 80 6511
rect 28 6443 36 6477
rect 70 6443 80 6477
rect 28 6409 80 6443
rect 28 6375 36 6409
rect 70 6375 80 6409
rect 28 6363 80 6375
rect 110 6545 162 6563
rect 110 6511 120 6545
rect 154 6511 162 6545
rect 110 6477 162 6511
rect 110 6443 120 6477
rect 154 6443 162 6477
rect 110 6409 162 6443
rect 110 6375 120 6409
rect 154 6375 162 6409
rect 298 6529 310 6563
rect 344 6529 356 6563
rect 298 6495 356 6529
rect 298 6461 310 6495
rect 344 6461 356 6495
rect 298 6427 356 6461
rect 298 6393 310 6427
rect 344 6393 356 6427
rect 298 6378 356 6393
rect 386 6563 444 6578
rect 386 6529 398 6563
rect 432 6529 444 6563
rect 624 6553 636 6587
rect 670 6553 686 6587
rect 624 6538 686 6553
rect 716 6723 782 6738
rect 716 6689 732 6723
rect 766 6689 782 6723
rect 716 6655 782 6689
rect 716 6621 732 6655
rect 766 6621 782 6655
rect 716 6587 782 6621
rect 716 6553 732 6587
rect 766 6553 782 6587
rect 716 6538 782 6553
rect 812 6723 874 6738
rect 812 6689 828 6723
rect 862 6689 874 6723
rect 812 6655 874 6689
rect 812 6621 828 6655
rect 862 6621 874 6655
rect 812 6587 874 6621
rect 2512 6723 2574 6738
rect 2512 6689 2524 6723
rect 2558 6689 2574 6723
rect 812 6553 828 6587
rect 862 6553 874 6587
rect 812 6538 874 6553
rect 944 6563 1002 6578
rect 386 6495 444 6529
rect 386 6461 398 6495
rect 432 6461 444 6495
rect 386 6427 444 6461
rect 944 6529 956 6563
rect 990 6529 1002 6563
rect 944 6495 1002 6529
rect 944 6461 956 6495
rect 990 6461 1002 6495
rect 386 6393 398 6427
rect 432 6393 444 6427
rect 386 6378 444 6393
rect 110 6363 162 6375
rect 944 6427 1002 6461
rect 944 6393 956 6427
rect 990 6393 1002 6427
rect 944 6378 1002 6393
rect 1032 6563 1090 6578
rect 1032 6529 1044 6563
rect 1078 6529 1090 6563
rect 1032 6495 1090 6529
rect 1032 6461 1044 6495
rect 1078 6461 1090 6495
rect 1032 6427 1090 6461
rect 1032 6393 1044 6427
rect 1078 6393 1090 6427
rect 1032 6378 1090 6393
rect 1224 6553 1276 6571
rect 1224 6519 1232 6553
rect 1266 6519 1276 6553
rect 1224 6485 1276 6519
rect 1224 6451 1232 6485
rect 1266 6451 1276 6485
rect 1224 6417 1276 6451
rect 1224 6383 1232 6417
rect 1266 6383 1276 6417
rect 1224 6371 1276 6383
rect 1306 6553 1358 6571
rect 1306 6519 1316 6553
rect 1350 6519 1358 6553
rect 2512 6655 2574 6689
rect 2512 6621 2524 6655
rect 2558 6621 2574 6655
rect 2512 6587 2574 6621
rect 2186 6563 2244 6578
rect 1916 6545 1968 6563
rect 1306 6485 1358 6519
rect 1306 6451 1316 6485
rect 1350 6451 1358 6485
rect 1306 6417 1358 6451
rect 1306 6383 1316 6417
rect 1350 6383 1358 6417
rect 1306 6371 1358 6383
rect 1523 6500 1575 6523
rect 1523 6466 1531 6500
rect 1565 6466 1575 6500
rect 1523 6419 1575 6466
rect 1523 6385 1531 6419
rect 1565 6385 1575 6419
rect 1523 6365 1575 6385
rect 1605 6487 1663 6523
rect 1605 6453 1617 6487
rect 1651 6453 1663 6487
rect 1605 6419 1663 6453
rect 1605 6385 1617 6419
rect 1651 6385 1663 6419
rect 1605 6365 1663 6385
rect 1693 6487 1745 6523
rect 1693 6453 1703 6487
rect 1737 6453 1745 6487
rect 1693 6419 1745 6453
rect 1693 6385 1703 6419
rect 1737 6385 1745 6419
rect 1693 6365 1745 6385
rect 1916 6511 1924 6545
rect 1958 6511 1968 6545
rect 1916 6477 1968 6511
rect 1916 6443 1924 6477
rect 1958 6443 1968 6477
rect 1916 6409 1968 6443
rect 1916 6375 1924 6409
rect 1958 6375 1968 6409
rect 1916 6363 1968 6375
rect 1998 6545 2050 6563
rect 1998 6511 2008 6545
rect 2042 6511 2050 6545
rect 1998 6477 2050 6511
rect 1998 6443 2008 6477
rect 2042 6443 2050 6477
rect 1998 6409 2050 6443
rect 1998 6375 2008 6409
rect 2042 6375 2050 6409
rect 2186 6529 2198 6563
rect 2232 6529 2244 6563
rect 2186 6495 2244 6529
rect 2186 6461 2198 6495
rect 2232 6461 2244 6495
rect 2186 6427 2244 6461
rect 2186 6393 2198 6427
rect 2232 6393 2244 6427
rect 2186 6378 2244 6393
rect 2274 6563 2332 6578
rect 2274 6529 2286 6563
rect 2320 6529 2332 6563
rect 2512 6553 2524 6587
rect 2558 6553 2574 6587
rect 2512 6538 2574 6553
rect 2604 6723 2670 6738
rect 2604 6689 2620 6723
rect 2654 6689 2670 6723
rect 2604 6655 2670 6689
rect 2604 6621 2620 6655
rect 2654 6621 2670 6655
rect 2604 6587 2670 6621
rect 2604 6553 2620 6587
rect 2654 6553 2670 6587
rect 2604 6538 2670 6553
rect 2700 6723 2762 6738
rect 2700 6689 2716 6723
rect 2750 6689 2762 6723
rect 2700 6655 2762 6689
rect 2700 6621 2716 6655
rect 2750 6621 2762 6655
rect 2700 6587 2762 6621
rect 4400 6723 4462 6738
rect 4400 6689 4412 6723
rect 4446 6689 4462 6723
rect 2700 6553 2716 6587
rect 2750 6553 2762 6587
rect 2700 6538 2762 6553
rect 2832 6563 2890 6578
rect 2274 6495 2332 6529
rect 2274 6461 2286 6495
rect 2320 6461 2332 6495
rect 2274 6427 2332 6461
rect 2832 6529 2844 6563
rect 2878 6529 2890 6563
rect 2832 6495 2890 6529
rect 2832 6461 2844 6495
rect 2878 6461 2890 6495
rect 2274 6393 2286 6427
rect 2320 6393 2332 6427
rect 2274 6378 2332 6393
rect 1998 6363 2050 6375
rect 2832 6427 2890 6461
rect 2832 6393 2844 6427
rect 2878 6393 2890 6427
rect 2832 6378 2890 6393
rect 2920 6563 2978 6578
rect 2920 6529 2932 6563
rect 2966 6529 2978 6563
rect 2920 6495 2978 6529
rect 2920 6461 2932 6495
rect 2966 6461 2978 6495
rect 2920 6427 2978 6461
rect 2920 6393 2932 6427
rect 2966 6393 2978 6427
rect 2920 6378 2978 6393
rect 3112 6553 3164 6571
rect 3112 6519 3120 6553
rect 3154 6519 3164 6553
rect 3112 6485 3164 6519
rect 3112 6451 3120 6485
rect 3154 6451 3164 6485
rect 3112 6417 3164 6451
rect 3112 6383 3120 6417
rect 3154 6383 3164 6417
rect 3112 6371 3164 6383
rect 3194 6553 3246 6571
rect 3194 6519 3204 6553
rect 3238 6519 3246 6553
rect 4400 6655 4462 6689
rect 4400 6621 4412 6655
rect 4446 6621 4462 6655
rect 4400 6587 4462 6621
rect 4074 6563 4132 6578
rect 3804 6545 3856 6563
rect 3194 6485 3246 6519
rect 3194 6451 3204 6485
rect 3238 6451 3246 6485
rect 3194 6417 3246 6451
rect 3194 6383 3204 6417
rect 3238 6383 3246 6417
rect 3194 6371 3246 6383
rect 3411 6500 3463 6523
rect 3411 6466 3419 6500
rect 3453 6466 3463 6500
rect 3411 6419 3463 6466
rect 3411 6385 3419 6419
rect 3453 6385 3463 6419
rect 3411 6365 3463 6385
rect 3493 6487 3551 6523
rect 3493 6453 3505 6487
rect 3539 6453 3551 6487
rect 3493 6419 3551 6453
rect 3493 6385 3505 6419
rect 3539 6385 3551 6419
rect 3493 6365 3551 6385
rect 3581 6487 3633 6523
rect 3581 6453 3591 6487
rect 3625 6453 3633 6487
rect 3581 6419 3633 6453
rect 3581 6385 3591 6419
rect 3625 6385 3633 6419
rect 3581 6365 3633 6385
rect 3804 6511 3812 6545
rect 3846 6511 3856 6545
rect 3804 6477 3856 6511
rect 3804 6443 3812 6477
rect 3846 6443 3856 6477
rect 3804 6409 3856 6443
rect 3804 6375 3812 6409
rect 3846 6375 3856 6409
rect 3804 6363 3856 6375
rect 3886 6545 3938 6563
rect 3886 6511 3896 6545
rect 3930 6511 3938 6545
rect 3886 6477 3938 6511
rect 3886 6443 3896 6477
rect 3930 6443 3938 6477
rect 3886 6409 3938 6443
rect 3886 6375 3896 6409
rect 3930 6375 3938 6409
rect 4074 6529 4086 6563
rect 4120 6529 4132 6563
rect 4074 6495 4132 6529
rect 4074 6461 4086 6495
rect 4120 6461 4132 6495
rect 4074 6427 4132 6461
rect 4074 6393 4086 6427
rect 4120 6393 4132 6427
rect 4074 6378 4132 6393
rect 4162 6563 4220 6578
rect 4162 6529 4174 6563
rect 4208 6529 4220 6563
rect 4400 6553 4412 6587
rect 4446 6553 4462 6587
rect 4400 6538 4462 6553
rect 4492 6723 4558 6738
rect 4492 6689 4508 6723
rect 4542 6689 4558 6723
rect 4492 6655 4558 6689
rect 4492 6621 4508 6655
rect 4542 6621 4558 6655
rect 4492 6587 4558 6621
rect 4492 6553 4508 6587
rect 4542 6553 4558 6587
rect 4492 6538 4558 6553
rect 4588 6723 4650 6738
rect 4588 6689 4604 6723
rect 4638 6689 4650 6723
rect 4588 6655 4650 6689
rect 4588 6621 4604 6655
rect 4638 6621 4650 6655
rect 4588 6587 4650 6621
rect 6288 6723 6350 6738
rect 6288 6689 6300 6723
rect 6334 6689 6350 6723
rect 4588 6553 4604 6587
rect 4638 6553 4650 6587
rect 4588 6538 4650 6553
rect 4720 6563 4778 6578
rect 4162 6495 4220 6529
rect 4162 6461 4174 6495
rect 4208 6461 4220 6495
rect 4162 6427 4220 6461
rect 4720 6529 4732 6563
rect 4766 6529 4778 6563
rect 4720 6495 4778 6529
rect 4720 6461 4732 6495
rect 4766 6461 4778 6495
rect 4162 6393 4174 6427
rect 4208 6393 4220 6427
rect 4162 6378 4220 6393
rect 3886 6363 3938 6375
rect 4720 6427 4778 6461
rect 4720 6393 4732 6427
rect 4766 6393 4778 6427
rect 4720 6378 4778 6393
rect 4808 6563 4866 6578
rect 4808 6529 4820 6563
rect 4854 6529 4866 6563
rect 4808 6495 4866 6529
rect 4808 6461 4820 6495
rect 4854 6461 4866 6495
rect 4808 6427 4866 6461
rect 4808 6393 4820 6427
rect 4854 6393 4866 6427
rect 4808 6378 4866 6393
rect 5000 6553 5052 6571
rect 5000 6519 5008 6553
rect 5042 6519 5052 6553
rect 5000 6485 5052 6519
rect 5000 6451 5008 6485
rect 5042 6451 5052 6485
rect 5000 6417 5052 6451
rect 5000 6383 5008 6417
rect 5042 6383 5052 6417
rect 5000 6371 5052 6383
rect 5082 6553 5134 6571
rect 5082 6519 5092 6553
rect 5126 6519 5134 6553
rect 6288 6655 6350 6689
rect 6288 6621 6300 6655
rect 6334 6621 6350 6655
rect 6288 6587 6350 6621
rect 5962 6563 6020 6578
rect 5692 6545 5744 6563
rect 5082 6485 5134 6519
rect 5082 6451 5092 6485
rect 5126 6451 5134 6485
rect 5082 6417 5134 6451
rect 5082 6383 5092 6417
rect 5126 6383 5134 6417
rect 5082 6371 5134 6383
rect 5299 6500 5351 6523
rect 5299 6466 5307 6500
rect 5341 6466 5351 6500
rect 5299 6419 5351 6466
rect 5299 6385 5307 6419
rect 5341 6385 5351 6419
rect 5299 6365 5351 6385
rect 5381 6487 5439 6523
rect 5381 6453 5393 6487
rect 5427 6453 5439 6487
rect 5381 6419 5439 6453
rect 5381 6385 5393 6419
rect 5427 6385 5439 6419
rect 5381 6365 5439 6385
rect 5469 6487 5521 6523
rect 5469 6453 5479 6487
rect 5513 6453 5521 6487
rect 5469 6419 5521 6453
rect 5469 6385 5479 6419
rect 5513 6385 5521 6419
rect 5469 6365 5521 6385
rect 5692 6511 5700 6545
rect 5734 6511 5744 6545
rect 5692 6477 5744 6511
rect 5692 6443 5700 6477
rect 5734 6443 5744 6477
rect 5692 6409 5744 6443
rect 5692 6375 5700 6409
rect 5734 6375 5744 6409
rect 5692 6363 5744 6375
rect 5774 6545 5826 6563
rect 5774 6511 5784 6545
rect 5818 6511 5826 6545
rect 5774 6477 5826 6511
rect 5774 6443 5784 6477
rect 5818 6443 5826 6477
rect 5774 6409 5826 6443
rect 5774 6375 5784 6409
rect 5818 6375 5826 6409
rect 5962 6529 5974 6563
rect 6008 6529 6020 6563
rect 5962 6495 6020 6529
rect 5962 6461 5974 6495
rect 6008 6461 6020 6495
rect 5962 6427 6020 6461
rect 5962 6393 5974 6427
rect 6008 6393 6020 6427
rect 5962 6378 6020 6393
rect 6050 6563 6108 6578
rect 6050 6529 6062 6563
rect 6096 6529 6108 6563
rect 6288 6553 6300 6587
rect 6334 6553 6350 6587
rect 6288 6538 6350 6553
rect 6380 6723 6446 6738
rect 6380 6689 6396 6723
rect 6430 6689 6446 6723
rect 6380 6655 6446 6689
rect 6380 6621 6396 6655
rect 6430 6621 6446 6655
rect 6380 6587 6446 6621
rect 6380 6553 6396 6587
rect 6430 6553 6446 6587
rect 6380 6538 6446 6553
rect 6476 6723 6538 6738
rect 6476 6689 6492 6723
rect 6526 6689 6538 6723
rect 6476 6655 6538 6689
rect 6476 6621 6492 6655
rect 6526 6621 6538 6655
rect 6476 6587 6538 6621
rect 8176 6723 8238 6738
rect 8176 6689 8188 6723
rect 8222 6689 8238 6723
rect 6476 6553 6492 6587
rect 6526 6553 6538 6587
rect 6476 6538 6538 6553
rect 6608 6563 6666 6578
rect 6050 6495 6108 6529
rect 6050 6461 6062 6495
rect 6096 6461 6108 6495
rect 6050 6427 6108 6461
rect 6608 6529 6620 6563
rect 6654 6529 6666 6563
rect 6608 6495 6666 6529
rect 6608 6461 6620 6495
rect 6654 6461 6666 6495
rect 6050 6393 6062 6427
rect 6096 6393 6108 6427
rect 6050 6378 6108 6393
rect 5774 6363 5826 6375
rect 6608 6427 6666 6461
rect 6608 6393 6620 6427
rect 6654 6393 6666 6427
rect 6608 6378 6666 6393
rect 6696 6563 6754 6578
rect 6696 6529 6708 6563
rect 6742 6529 6754 6563
rect 6696 6495 6754 6529
rect 6696 6461 6708 6495
rect 6742 6461 6754 6495
rect 6696 6427 6754 6461
rect 6696 6393 6708 6427
rect 6742 6393 6754 6427
rect 6696 6378 6754 6393
rect 6888 6553 6940 6571
rect 6888 6519 6896 6553
rect 6930 6519 6940 6553
rect 6888 6485 6940 6519
rect 6888 6451 6896 6485
rect 6930 6451 6940 6485
rect 6888 6417 6940 6451
rect 6888 6383 6896 6417
rect 6930 6383 6940 6417
rect 6888 6371 6940 6383
rect 6970 6553 7022 6571
rect 6970 6519 6980 6553
rect 7014 6519 7022 6553
rect 8176 6655 8238 6689
rect 8176 6621 8188 6655
rect 8222 6621 8238 6655
rect 8176 6587 8238 6621
rect 7850 6563 7908 6578
rect 7580 6545 7632 6563
rect 6970 6485 7022 6519
rect 6970 6451 6980 6485
rect 7014 6451 7022 6485
rect 6970 6417 7022 6451
rect 6970 6383 6980 6417
rect 7014 6383 7022 6417
rect 6970 6371 7022 6383
rect 7187 6500 7239 6523
rect 7187 6466 7195 6500
rect 7229 6466 7239 6500
rect 7187 6419 7239 6466
rect 7187 6385 7195 6419
rect 7229 6385 7239 6419
rect 7187 6365 7239 6385
rect 7269 6487 7327 6523
rect 7269 6453 7281 6487
rect 7315 6453 7327 6487
rect 7269 6419 7327 6453
rect 7269 6385 7281 6419
rect 7315 6385 7327 6419
rect 7269 6365 7327 6385
rect 7357 6487 7409 6523
rect 7357 6453 7367 6487
rect 7401 6453 7409 6487
rect 7357 6419 7409 6453
rect 7357 6385 7367 6419
rect 7401 6385 7409 6419
rect 7357 6365 7409 6385
rect 7580 6511 7588 6545
rect 7622 6511 7632 6545
rect 7580 6477 7632 6511
rect 7580 6443 7588 6477
rect 7622 6443 7632 6477
rect 7580 6409 7632 6443
rect 7580 6375 7588 6409
rect 7622 6375 7632 6409
rect 7580 6363 7632 6375
rect 7662 6545 7714 6563
rect 7662 6511 7672 6545
rect 7706 6511 7714 6545
rect 7662 6477 7714 6511
rect 7662 6443 7672 6477
rect 7706 6443 7714 6477
rect 7662 6409 7714 6443
rect 7662 6375 7672 6409
rect 7706 6375 7714 6409
rect 7850 6529 7862 6563
rect 7896 6529 7908 6563
rect 7850 6495 7908 6529
rect 7850 6461 7862 6495
rect 7896 6461 7908 6495
rect 7850 6427 7908 6461
rect 7850 6393 7862 6427
rect 7896 6393 7908 6427
rect 7850 6378 7908 6393
rect 7938 6563 7996 6578
rect 7938 6529 7950 6563
rect 7984 6529 7996 6563
rect 8176 6553 8188 6587
rect 8222 6553 8238 6587
rect 8176 6538 8238 6553
rect 8268 6723 8334 6738
rect 8268 6689 8284 6723
rect 8318 6689 8334 6723
rect 8268 6655 8334 6689
rect 8268 6621 8284 6655
rect 8318 6621 8334 6655
rect 8268 6587 8334 6621
rect 8268 6553 8284 6587
rect 8318 6553 8334 6587
rect 8268 6538 8334 6553
rect 8364 6723 8426 6738
rect 8364 6689 8380 6723
rect 8414 6689 8426 6723
rect 8364 6655 8426 6689
rect 8364 6621 8380 6655
rect 8414 6621 8426 6655
rect 8364 6587 8426 6621
rect 10064 6723 10126 6738
rect 10064 6689 10076 6723
rect 10110 6689 10126 6723
rect 8364 6553 8380 6587
rect 8414 6553 8426 6587
rect 8364 6538 8426 6553
rect 8496 6563 8554 6578
rect 7938 6495 7996 6529
rect 7938 6461 7950 6495
rect 7984 6461 7996 6495
rect 7938 6427 7996 6461
rect 8496 6529 8508 6563
rect 8542 6529 8554 6563
rect 8496 6495 8554 6529
rect 8496 6461 8508 6495
rect 8542 6461 8554 6495
rect 7938 6393 7950 6427
rect 7984 6393 7996 6427
rect 7938 6378 7996 6393
rect 7662 6363 7714 6375
rect 8496 6427 8554 6461
rect 8496 6393 8508 6427
rect 8542 6393 8554 6427
rect 8496 6378 8554 6393
rect 8584 6563 8642 6578
rect 8584 6529 8596 6563
rect 8630 6529 8642 6563
rect 8584 6495 8642 6529
rect 8584 6461 8596 6495
rect 8630 6461 8642 6495
rect 8584 6427 8642 6461
rect 8584 6393 8596 6427
rect 8630 6393 8642 6427
rect 8584 6378 8642 6393
rect 8776 6553 8828 6571
rect 8776 6519 8784 6553
rect 8818 6519 8828 6553
rect 8776 6485 8828 6519
rect 8776 6451 8784 6485
rect 8818 6451 8828 6485
rect 8776 6417 8828 6451
rect 8776 6383 8784 6417
rect 8818 6383 8828 6417
rect 8776 6371 8828 6383
rect 8858 6553 8910 6571
rect 8858 6519 8868 6553
rect 8902 6519 8910 6553
rect 10064 6655 10126 6689
rect 10064 6621 10076 6655
rect 10110 6621 10126 6655
rect 10064 6587 10126 6621
rect 9738 6563 9796 6578
rect 9468 6545 9520 6563
rect 8858 6485 8910 6519
rect 8858 6451 8868 6485
rect 8902 6451 8910 6485
rect 8858 6417 8910 6451
rect 8858 6383 8868 6417
rect 8902 6383 8910 6417
rect 8858 6371 8910 6383
rect 9075 6500 9127 6523
rect 9075 6466 9083 6500
rect 9117 6466 9127 6500
rect 9075 6419 9127 6466
rect 9075 6385 9083 6419
rect 9117 6385 9127 6419
rect 9075 6365 9127 6385
rect 9157 6487 9215 6523
rect 9157 6453 9169 6487
rect 9203 6453 9215 6487
rect 9157 6419 9215 6453
rect 9157 6385 9169 6419
rect 9203 6385 9215 6419
rect 9157 6365 9215 6385
rect 9245 6487 9297 6523
rect 9245 6453 9255 6487
rect 9289 6453 9297 6487
rect 9245 6419 9297 6453
rect 9245 6385 9255 6419
rect 9289 6385 9297 6419
rect 9245 6365 9297 6385
rect 9468 6511 9476 6545
rect 9510 6511 9520 6545
rect 9468 6477 9520 6511
rect 9468 6443 9476 6477
rect 9510 6443 9520 6477
rect 9468 6409 9520 6443
rect 9468 6375 9476 6409
rect 9510 6375 9520 6409
rect 9468 6363 9520 6375
rect 9550 6545 9602 6563
rect 9550 6511 9560 6545
rect 9594 6511 9602 6545
rect 9550 6477 9602 6511
rect 9550 6443 9560 6477
rect 9594 6443 9602 6477
rect 9550 6409 9602 6443
rect 9550 6375 9560 6409
rect 9594 6375 9602 6409
rect 9738 6529 9750 6563
rect 9784 6529 9796 6563
rect 9738 6495 9796 6529
rect 9738 6461 9750 6495
rect 9784 6461 9796 6495
rect 9738 6427 9796 6461
rect 9738 6393 9750 6427
rect 9784 6393 9796 6427
rect 9738 6378 9796 6393
rect 9826 6563 9884 6578
rect 9826 6529 9838 6563
rect 9872 6529 9884 6563
rect 10064 6553 10076 6587
rect 10110 6553 10126 6587
rect 10064 6538 10126 6553
rect 10156 6723 10222 6738
rect 10156 6689 10172 6723
rect 10206 6689 10222 6723
rect 10156 6655 10222 6689
rect 10156 6621 10172 6655
rect 10206 6621 10222 6655
rect 10156 6587 10222 6621
rect 10156 6553 10172 6587
rect 10206 6553 10222 6587
rect 10156 6538 10222 6553
rect 10252 6723 10314 6738
rect 10252 6689 10268 6723
rect 10302 6689 10314 6723
rect 10252 6655 10314 6689
rect 10252 6621 10268 6655
rect 10302 6621 10314 6655
rect 10252 6587 10314 6621
rect 11952 6723 12014 6738
rect 11952 6689 11964 6723
rect 11998 6689 12014 6723
rect 10252 6553 10268 6587
rect 10302 6553 10314 6587
rect 10252 6538 10314 6553
rect 10384 6563 10442 6578
rect 9826 6495 9884 6529
rect 9826 6461 9838 6495
rect 9872 6461 9884 6495
rect 9826 6427 9884 6461
rect 10384 6529 10396 6563
rect 10430 6529 10442 6563
rect 10384 6495 10442 6529
rect 10384 6461 10396 6495
rect 10430 6461 10442 6495
rect 9826 6393 9838 6427
rect 9872 6393 9884 6427
rect 9826 6378 9884 6393
rect 9550 6363 9602 6375
rect 10384 6427 10442 6461
rect 10384 6393 10396 6427
rect 10430 6393 10442 6427
rect 10384 6378 10442 6393
rect 10472 6563 10530 6578
rect 10472 6529 10484 6563
rect 10518 6529 10530 6563
rect 10472 6495 10530 6529
rect 10472 6461 10484 6495
rect 10518 6461 10530 6495
rect 10472 6427 10530 6461
rect 10472 6393 10484 6427
rect 10518 6393 10530 6427
rect 10472 6378 10530 6393
rect 10664 6553 10716 6571
rect 10664 6519 10672 6553
rect 10706 6519 10716 6553
rect 10664 6485 10716 6519
rect 10664 6451 10672 6485
rect 10706 6451 10716 6485
rect 10664 6417 10716 6451
rect 10664 6383 10672 6417
rect 10706 6383 10716 6417
rect 10664 6371 10716 6383
rect 10746 6553 10798 6571
rect 10746 6519 10756 6553
rect 10790 6519 10798 6553
rect 11952 6655 12014 6689
rect 11952 6621 11964 6655
rect 11998 6621 12014 6655
rect 11952 6587 12014 6621
rect 11626 6563 11684 6578
rect 11356 6545 11408 6563
rect 10746 6485 10798 6519
rect 10746 6451 10756 6485
rect 10790 6451 10798 6485
rect 10746 6417 10798 6451
rect 10746 6383 10756 6417
rect 10790 6383 10798 6417
rect 10746 6371 10798 6383
rect 10963 6500 11015 6523
rect 10963 6466 10971 6500
rect 11005 6466 11015 6500
rect 10963 6419 11015 6466
rect 10963 6385 10971 6419
rect 11005 6385 11015 6419
rect 10963 6365 11015 6385
rect 11045 6487 11103 6523
rect 11045 6453 11057 6487
rect 11091 6453 11103 6487
rect 11045 6419 11103 6453
rect 11045 6385 11057 6419
rect 11091 6385 11103 6419
rect 11045 6365 11103 6385
rect 11133 6487 11185 6523
rect 11133 6453 11143 6487
rect 11177 6453 11185 6487
rect 11133 6419 11185 6453
rect 11133 6385 11143 6419
rect 11177 6385 11185 6419
rect 11133 6365 11185 6385
rect 11356 6511 11364 6545
rect 11398 6511 11408 6545
rect 11356 6477 11408 6511
rect 11356 6443 11364 6477
rect 11398 6443 11408 6477
rect 11356 6409 11408 6443
rect 11356 6375 11364 6409
rect 11398 6375 11408 6409
rect 11356 6363 11408 6375
rect 11438 6545 11490 6563
rect 11438 6511 11448 6545
rect 11482 6511 11490 6545
rect 11438 6477 11490 6511
rect 11438 6443 11448 6477
rect 11482 6443 11490 6477
rect 11438 6409 11490 6443
rect 11438 6375 11448 6409
rect 11482 6375 11490 6409
rect 11626 6529 11638 6563
rect 11672 6529 11684 6563
rect 11626 6495 11684 6529
rect 11626 6461 11638 6495
rect 11672 6461 11684 6495
rect 11626 6427 11684 6461
rect 11626 6393 11638 6427
rect 11672 6393 11684 6427
rect 11626 6378 11684 6393
rect 11714 6563 11772 6578
rect 11714 6529 11726 6563
rect 11760 6529 11772 6563
rect 11952 6553 11964 6587
rect 11998 6553 12014 6587
rect 11952 6538 12014 6553
rect 12044 6723 12110 6738
rect 12044 6689 12060 6723
rect 12094 6689 12110 6723
rect 12044 6655 12110 6689
rect 12044 6621 12060 6655
rect 12094 6621 12110 6655
rect 12044 6587 12110 6621
rect 12044 6553 12060 6587
rect 12094 6553 12110 6587
rect 12044 6538 12110 6553
rect 12140 6723 12202 6738
rect 12140 6689 12156 6723
rect 12190 6689 12202 6723
rect 12140 6655 12202 6689
rect 12140 6621 12156 6655
rect 12190 6621 12202 6655
rect 12140 6587 12202 6621
rect 13840 6723 13902 6738
rect 13840 6689 13852 6723
rect 13886 6689 13902 6723
rect 12140 6553 12156 6587
rect 12190 6553 12202 6587
rect 12140 6538 12202 6553
rect 12272 6563 12330 6578
rect 11714 6495 11772 6529
rect 11714 6461 11726 6495
rect 11760 6461 11772 6495
rect 11714 6427 11772 6461
rect 12272 6529 12284 6563
rect 12318 6529 12330 6563
rect 12272 6495 12330 6529
rect 12272 6461 12284 6495
rect 12318 6461 12330 6495
rect 11714 6393 11726 6427
rect 11760 6393 11772 6427
rect 11714 6378 11772 6393
rect 11438 6363 11490 6375
rect 12272 6427 12330 6461
rect 12272 6393 12284 6427
rect 12318 6393 12330 6427
rect 12272 6378 12330 6393
rect 12360 6563 12418 6578
rect 12360 6529 12372 6563
rect 12406 6529 12418 6563
rect 12360 6495 12418 6529
rect 12360 6461 12372 6495
rect 12406 6461 12418 6495
rect 12360 6427 12418 6461
rect 12360 6393 12372 6427
rect 12406 6393 12418 6427
rect 12360 6378 12418 6393
rect 12552 6553 12604 6571
rect 12552 6519 12560 6553
rect 12594 6519 12604 6553
rect 12552 6485 12604 6519
rect 12552 6451 12560 6485
rect 12594 6451 12604 6485
rect 12552 6417 12604 6451
rect 12552 6383 12560 6417
rect 12594 6383 12604 6417
rect 12552 6371 12604 6383
rect 12634 6553 12686 6571
rect 12634 6519 12644 6553
rect 12678 6519 12686 6553
rect 13840 6655 13902 6689
rect 13840 6621 13852 6655
rect 13886 6621 13902 6655
rect 13840 6587 13902 6621
rect 13514 6563 13572 6578
rect 13244 6545 13296 6563
rect 12634 6485 12686 6519
rect 12634 6451 12644 6485
rect 12678 6451 12686 6485
rect 12634 6417 12686 6451
rect 12634 6383 12644 6417
rect 12678 6383 12686 6417
rect 12634 6371 12686 6383
rect 12851 6500 12903 6523
rect 12851 6466 12859 6500
rect 12893 6466 12903 6500
rect 12851 6419 12903 6466
rect 12851 6385 12859 6419
rect 12893 6385 12903 6419
rect 12851 6365 12903 6385
rect 12933 6487 12991 6523
rect 12933 6453 12945 6487
rect 12979 6453 12991 6487
rect 12933 6419 12991 6453
rect 12933 6385 12945 6419
rect 12979 6385 12991 6419
rect 12933 6365 12991 6385
rect 13021 6487 13073 6523
rect 13021 6453 13031 6487
rect 13065 6453 13073 6487
rect 13021 6419 13073 6453
rect 13021 6385 13031 6419
rect 13065 6385 13073 6419
rect 13021 6365 13073 6385
rect 13244 6511 13252 6545
rect 13286 6511 13296 6545
rect 13244 6477 13296 6511
rect 13244 6443 13252 6477
rect 13286 6443 13296 6477
rect 13244 6409 13296 6443
rect 13244 6375 13252 6409
rect 13286 6375 13296 6409
rect 13244 6363 13296 6375
rect 13326 6545 13378 6563
rect 13326 6511 13336 6545
rect 13370 6511 13378 6545
rect 13326 6477 13378 6511
rect 13326 6443 13336 6477
rect 13370 6443 13378 6477
rect 13326 6409 13378 6443
rect 13326 6375 13336 6409
rect 13370 6375 13378 6409
rect 13514 6529 13526 6563
rect 13560 6529 13572 6563
rect 13514 6495 13572 6529
rect 13514 6461 13526 6495
rect 13560 6461 13572 6495
rect 13514 6427 13572 6461
rect 13514 6393 13526 6427
rect 13560 6393 13572 6427
rect 13514 6378 13572 6393
rect 13602 6563 13660 6578
rect 13602 6529 13614 6563
rect 13648 6529 13660 6563
rect 13840 6553 13852 6587
rect 13886 6553 13902 6587
rect 13840 6538 13902 6553
rect 13932 6723 13998 6738
rect 13932 6689 13948 6723
rect 13982 6689 13998 6723
rect 13932 6655 13998 6689
rect 13932 6621 13948 6655
rect 13982 6621 13998 6655
rect 13932 6587 13998 6621
rect 13932 6553 13948 6587
rect 13982 6553 13998 6587
rect 13932 6538 13998 6553
rect 14028 6723 14090 6738
rect 14028 6689 14044 6723
rect 14078 6689 14090 6723
rect 14028 6655 14090 6689
rect 14028 6621 14044 6655
rect 14078 6621 14090 6655
rect 14028 6587 14090 6621
rect 15722 6723 15784 6738
rect 15722 6689 15734 6723
rect 15768 6689 15784 6723
rect 14028 6553 14044 6587
rect 14078 6553 14090 6587
rect 14028 6538 14090 6553
rect 14160 6563 14218 6578
rect 13602 6495 13660 6529
rect 13602 6461 13614 6495
rect 13648 6461 13660 6495
rect 13602 6427 13660 6461
rect 14160 6529 14172 6563
rect 14206 6529 14218 6563
rect 14160 6495 14218 6529
rect 14160 6461 14172 6495
rect 14206 6461 14218 6495
rect 13602 6393 13614 6427
rect 13648 6393 13660 6427
rect 13602 6378 13660 6393
rect 13326 6363 13378 6375
rect 14160 6427 14218 6461
rect 14160 6393 14172 6427
rect 14206 6393 14218 6427
rect 14160 6378 14218 6393
rect 14248 6563 14306 6578
rect 14248 6529 14260 6563
rect 14294 6529 14306 6563
rect 14248 6495 14306 6529
rect 14248 6461 14260 6495
rect 14294 6461 14306 6495
rect 14248 6427 14306 6461
rect 14248 6393 14260 6427
rect 14294 6393 14306 6427
rect 14248 6378 14306 6393
rect 14440 6553 14492 6571
rect 14440 6519 14448 6553
rect 14482 6519 14492 6553
rect 14440 6485 14492 6519
rect 14440 6451 14448 6485
rect 14482 6451 14492 6485
rect 14440 6417 14492 6451
rect 14440 6383 14448 6417
rect 14482 6383 14492 6417
rect 14440 6371 14492 6383
rect 14522 6553 14574 6571
rect 14522 6519 14532 6553
rect 14566 6519 14574 6553
rect 15722 6655 15784 6689
rect 15722 6621 15734 6655
rect 15768 6621 15784 6655
rect 15722 6587 15784 6621
rect 15396 6563 15454 6578
rect 15126 6545 15178 6563
rect 14522 6485 14574 6519
rect 14522 6451 14532 6485
rect 14566 6451 14574 6485
rect 14522 6417 14574 6451
rect 14522 6383 14532 6417
rect 14566 6383 14574 6417
rect 14522 6371 14574 6383
rect 14733 6500 14785 6523
rect 14733 6466 14741 6500
rect 14775 6466 14785 6500
rect 14733 6419 14785 6466
rect 14733 6385 14741 6419
rect 14775 6385 14785 6419
rect 14733 6365 14785 6385
rect 14815 6487 14873 6523
rect 14815 6453 14827 6487
rect 14861 6453 14873 6487
rect 14815 6419 14873 6453
rect 14815 6385 14827 6419
rect 14861 6385 14873 6419
rect 14815 6365 14873 6385
rect 14903 6487 14955 6523
rect 14903 6453 14913 6487
rect 14947 6453 14955 6487
rect 14903 6419 14955 6453
rect 14903 6385 14913 6419
rect 14947 6385 14955 6419
rect 14903 6365 14955 6385
rect 15126 6511 15134 6545
rect 15168 6511 15178 6545
rect 15126 6477 15178 6511
rect 15126 6443 15134 6477
rect 15168 6443 15178 6477
rect 15126 6409 15178 6443
rect 15126 6375 15134 6409
rect 15168 6375 15178 6409
rect 15126 6363 15178 6375
rect 15208 6545 15260 6563
rect 15208 6511 15218 6545
rect 15252 6511 15260 6545
rect 15208 6477 15260 6511
rect 15208 6443 15218 6477
rect 15252 6443 15260 6477
rect 15208 6409 15260 6443
rect 15208 6375 15218 6409
rect 15252 6375 15260 6409
rect 15396 6529 15408 6563
rect 15442 6529 15454 6563
rect 15396 6495 15454 6529
rect 15396 6461 15408 6495
rect 15442 6461 15454 6495
rect 15396 6427 15454 6461
rect 15396 6393 15408 6427
rect 15442 6393 15454 6427
rect 15396 6378 15454 6393
rect 15484 6563 15542 6578
rect 15484 6529 15496 6563
rect 15530 6529 15542 6563
rect 15722 6553 15734 6587
rect 15768 6553 15784 6587
rect 15722 6538 15784 6553
rect 15814 6723 15880 6738
rect 15814 6689 15830 6723
rect 15864 6689 15880 6723
rect 15814 6655 15880 6689
rect 15814 6621 15830 6655
rect 15864 6621 15880 6655
rect 15814 6587 15880 6621
rect 15814 6553 15830 6587
rect 15864 6553 15880 6587
rect 15814 6538 15880 6553
rect 15910 6723 15972 6738
rect 15910 6689 15926 6723
rect 15960 6689 15972 6723
rect 15910 6655 15972 6689
rect 15910 6621 15926 6655
rect 15960 6621 15972 6655
rect 15910 6587 15972 6621
rect 17610 6723 17672 6738
rect 17610 6689 17622 6723
rect 17656 6689 17672 6723
rect 15910 6553 15926 6587
rect 15960 6553 15972 6587
rect 15910 6538 15972 6553
rect 16042 6563 16100 6578
rect 15484 6495 15542 6529
rect 15484 6461 15496 6495
rect 15530 6461 15542 6495
rect 15484 6427 15542 6461
rect 16042 6529 16054 6563
rect 16088 6529 16100 6563
rect 16042 6495 16100 6529
rect 16042 6461 16054 6495
rect 16088 6461 16100 6495
rect 15484 6393 15496 6427
rect 15530 6393 15542 6427
rect 15484 6378 15542 6393
rect 15208 6363 15260 6375
rect 16042 6427 16100 6461
rect 16042 6393 16054 6427
rect 16088 6393 16100 6427
rect 16042 6378 16100 6393
rect 16130 6563 16188 6578
rect 16130 6529 16142 6563
rect 16176 6529 16188 6563
rect 16130 6495 16188 6529
rect 16130 6461 16142 6495
rect 16176 6461 16188 6495
rect 16130 6427 16188 6461
rect 16130 6393 16142 6427
rect 16176 6393 16188 6427
rect 16130 6378 16188 6393
rect 16322 6553 16374 6571
rect 16322 6519 16330 6553
rect 16364 6519 16374 6553
rect 16322 6485 16374 6519
rect 16322 6451 16330 6485
rect 16364 6451 16374 6485
rect 16322 6417 16374 6451
rect 16322 6383 16330 6417
rect 16364 6383 16374 6417
rect 16322 6371 16374 6383
rect 16404 6553 16456 6571
rect 16404 6519 16414 6553
rect 16448 6519 16456 6553
rect 17610 6655 17672 6689
rect 17610 6621 17622 6655
rect 17656 6621 17672 6655
rect 17610 6587 17672 6621
rect 17284 6563 17342 6578
rect 17014 6545 17066 6563
rect 16404 6485 16456 6519
rect 16404 6451 16414 6485
rect 16448 6451 16456 6485
rect 16404 6417 16456 6451
rect 16404 6383 16414 6417
rect 16448 6383 16456 6417
rect 16404 6371 16456 6383
rect 16621 6500 16673 6523
rect 16621 6466 16629 6500
rect 16663 6466 16673 6500
rect 16621 6419 16673 6466
rect 16621 6385 16629 6419
rect 16663 6385 16673 6419
rect 16621 6365 16673 6385
rect 16703 6487 16761 6523
rect 16703 6453 16715 6487
rect 16749 6453 16761 6487
rect 16703 6419 16761 6453
rect 16703 6385 16715 6419
rect 16749 6385 16761 6419
rect 16703 6365 16761 6385
rect 16791 6487 16843 6523
rect 16791 6453 16801 6487
rect 16835 6453 16843 6487
rect 16791 6419 16843 6453
rect 16791 6385 16801 6419
rect 16835 6385 16843 6419
rect 16791 6365 16843 6385
rect 17014 6511 17022 6545
rect 17056 6511 17066 6545
rect 17014 6477 17066 6511
rect 17014 6443 17022 6477
rect 17056 6443 17066 6477
rect 17014 6409 17066 6443
rect 17014 6375 17022 6409
rect 17056 6375 17066 6409
rect 17014 6363 17066 6375
rect 17096 6545 17148 6563
rect 17096 6511 17106 6545
rect 17140 6511 17148 6545
rect 17096 6477 17148 6511
rect 17096 6443 17106 6477
rect 17140 6443 17148 6477
rect 17096 6409 17148 6443
rect 17096 6375 17106 6409
rect 17140 6375 17148 6409
rect 17284 6529 17296 6563
rect 17330 6529 17342 6563
rect 17284 6495 17342 6529
rect 17284 6461 17296 6495
rect 17330 6461 17342 6495
rect 17284 6427 17342 6461
rect 17284 6393 17296 6427
rect 17330 6393 17342 6427
rect 17284 6378 17342 6393
rect 17372 6563 17430 6578
rect 17372 6529 17384 6563
rect 17418 6529 17430 6563
rect 17610 6553 17622 6587
rect 17656 6553 17672 6587
rect 17610 6538 17672 6553
rect 17702 6723 17768 6738
rect 17702 6689 17718 6723
rect 17752 6689 17768 6723
rect 17702 6655 17768 6689
rect 17702 6621 17718 6655
rect 17752 6621 17768 6655
rect 17702 6587 17768 6621
rect 17702 6553 17718 6587
rect 17752 6553 17768 6587
rect 17702 6538 17768 6553
rect 17798 6723 17860 6738
rect 17798 6689 17814 6723
rect 17848 6689 17860 6723
rect 17798 6655 17860 6689
rect 17798 6621 17814 6655
rect 17848 6621 17860 6655
rect 17798 6587 17860 6621
rect 19498 6723 19560 6738
rect 19498 6689 19510 6723
rect 19544 6689 19560 6723
rect 17798 6553 17814 6587
rect 17848 6553 17860 6587
rect 17798 6538 17860 6553
rect 17930 6563 17988 6578
rect 17372 6495 17430 6529
rect 17372 6461 17384 6495
rect 17418 6461 17430 6495
rect 17372 6427 17430 6461
rect 17930 6529 17942 6563
rect 17976 6529 17988 6563
rect 17930 6495 17988 6529
rect 17930 6461 17942 6495
rect 17976 6461 17988 6495
rect 17372 6393 17384 6427
rect 17418 6393 17430 6427
rect 17372 6378 17430 6393
rect 17096 6363 17148 6375
rect 17930 6427 17988 6461
rect 17930 6393 17942 6427
rect 17976 6393 17988 6427
rect 17930 6378 17988 6393
rect 18018 6563 18076 6578
rect 18018 6529 18030 6563
rect 18064 6529 18076 6563
rect 18018 6495 18076 6529
rect 18018 6461 18030 6495
rect 18064 6461 18076 6495
rect 18018 6427 18076 6461
rect 18018 6393 18030 6427
rect 18064 6393 18076 6427
rect 18018 6378 18076 6393
rect 18210 6553 18262 6571
rect 18210 6519 18218 6553
rect 18252 6519 18262 6553
rect 18210 6485 18262 6519
rect 18210 6451 18218 6485
rect 18252 6451 18262 6485
rect 18210 6417 18262 6451
rect 18210 6383 18218 6417
rect 18252 6383 18262 6417
rect 18210 6371 18262 6383
rect 18292 6553 18344 6571
rect 18292 6519 18302 6553
rect 18336 6519 18344 6553
rect 19498 6655 19560 6689
rect 19498 6621 19510 6655
rect 19544 6621 19560 6655
rect 19498 6587 19560 6621
rect 19172 6563 19230 6578
rect 18902 6545 18954 6563
rect 18292 6485 18344 6519
rect 18292 6451 18302 6485
rect 18336 6451 18344 6485
rect 18292 6417 18344 6451
rect 18292 6383 18302 6417
rect 18336 6383 18344 6417
rect 18292 6371 18344 6383
rect 18509 6500 18561 6523
rect 18509 6466 18517 6500
rect 18551 6466 18561 6500
rect 18509 6419 18561 6466
rect 18509 6385 18517 6419
rect 18551 6385 18561 6419
rect 18509 6365 18561 6385
rect 18591 6487 18649 6523
rect 18591 6453 18603 6487
rect 18637 6453 18649 6487
rect 18591 6419 18649 6453
rect 18591 6385 18603 6419
rect 18637 6385 18649 6419
rect 18591 6365 18649 6385
rect 18679 6487 18731 6523
rect 18679 6453 18689 6487
rect 18723 6453 18731 6487
rect 18679 6419 18731 6453
rect 18679 6385 18689 6419
rect 18723 6385 18731 6419
rect 18679 6365 18731 6385
rect 18902 6511 18910 6545
rect 18944 6511 18954 6545
rect 18902 6477 18954 6511
rect 18902 6443 18910 6477
rect 18944 6443 18954 6477
rect 18902 6409 18954 6443
rect 18902 6375 18910 6409
rect 18944 6375 18954 6409
rect 18902 6363 18954 6375
rect 18984 6545 19036 6563
rect 18984 6511 18994 6545
rect 19028 6511 19036 6545
rect 18984 6477 19036 6511
rect 18984 6443 18994 6477
rect 19028 6443 19036 6477
rect 18984 6409 19036 6443
rect 18984 6375 18994 6409
rect 19028 6375 19036 6409
rect 19172 6529 19184 6563
rect 19218 6529 19230 6563
rect 19172 6495 19230 6529
rect 19172 6461 19184 6495
rect 19218 6461 19230 6495
rect 19172 6427 19230 6461
rect 19172 6393 19184 6427
rect 19218 6393 19230 6427
rect 19172 6378 19230 6393
rect 19260 6563 19318 6578
rect 19260 6529 19272 6563
rect 19306 6529 19318 6563
rect 19498 6553 19510 6587
rect 19544 6553 19560 6587
rect 19498 6538 19560 6553
rect 19590 6723 19656 6738
rect 19590 6689 19606 6723
rect 19640 6689 19656 6723
rect 19590 6655 19656 6689
rect 19590 6621 19606 6655
rect 19640 6621 19656 6655
rect 19590 6587 19656 6621
rect 19590 6553 19606 6587
rect 19640 6553 19656 6587
rect 19590 6538 19656 6553
rect 19686 6723 19748 6738
rect 19686 6689 19702 6723
rect 19736 6689 19748 6723
rect 19686 6655 19748 6689
rect 19686 6621 19702 6655
rect 19736 6621 19748 6655
rect 19686 6587 19748 6621
rect 21386 6723 21448 6738
rect 21386 6689 21398 6723
rect 21432 6689 21448 6723
rect 19686 6553 19702 6587
rect 19736 6553 19748 6587
rect 19686 6538 19748 6553
rect 19818 6563 19876 6578
rect 19260 6495 19318 6529
rect 19260 6461 19272 6495
rect 19306 6461 19318 6495
rect 19260 6427 19318 6461
rect 19818 6529 19830 6563
rect 19864 6529 19876 6563
rect 19818 6495 19876 6529
rect 19818 6461 19830 6495
rect 19864 6461 19876 6495
rect 19260 6393 19272 6427
rect 19306 6393 19318 6427
rect 19260 6378 19318 6393
rect 18984 6363 19036 6375
rect 19818 6427 19876 6461
rect 19818 6393 19830 6427
rect 19864 6393 19876 6427
rect 19818 6378 19876 6393
rect 19906 6563 19964 6578
rect 19906 6529 19918 6563
rect 19952 6529 19964 6563
rect 19906 6495 19964 6529
rect 19906 6461 19918 6495
rect 19952 6461 19964 6495
rect 19906 6427 19964 6461
rect 19906 6393 19918 6427
rect 19952 6393 19964 6427
rect 19906 6378 19964 6393
rect 20098 6553 20150 6571
rect 20098 6519 20106 6553
rect 20140 6519 20150 6553
rect 20098 6485 20150 6519
rect 20098 6451 20106 6485
rect 20140 6451 20150 6485
rect 20098 6417 20150 6451
rect 20098 6383 20106 6417
rect 20140 6383 20150 6417
rect 20098 6371 20150 6383
rect 20180 6553 20232 6571
rect 20180 6519 20190 6553
rect 20224 6519 20232 6553
rect 21386 6655 21448 6689
rect 21386 6621 21398 6655
rect 21432 6621 21448 6655
rect 21386 6587 21448 6621
rect 21060 6563 21118 6578
rect 20790 6545 20842 6563
rect 20180 6485 20232 6519
rect 20180 6451 20190 6485
rect 20224 6451 20232 6485
rect 20180 6417 20232 6451
rect 20180 6383 20190 6417
rect 20224 6383 20232 6417
rect 20180 6371 20232 6383
rect 20397 6500 20449 6523
rect 20397 6466 20405 6500
rect 20439 6466 20449 6500
rect 20397 6419 20449 6466
rect 20397 6385 20405 6419
rect 20439 6385 20449 6419
rect 20397 6365 20449 6385
rect 20479 6487 20537 6523
rect 20479 6453 20491 6487
rect 20525 6453 20537 6487
rect 20479 6419 20537 6453
rect 20479 6385 20491 6419
rect 20525 6385 20537 6419
rect 20479 6365 20537 6385
rect 20567 6487 20619 6523
rect 20567 6453 20577 6487
rect 20611 6453 20619 6487
rect 20567 6419 20619 6453
rect 20567 6385 20577 6419
rect 20611 6385 20619 6419
rect 20567 6365 20619 6385
rect 20790 6511 20798 6545
rect 20832 6511 20842 6545
rect 20790 6477 20842 6511
rect 20790 6443 20798 6477
rect 20832 6443 20842 6477
rect 20790 6409 20842 6443
rect 20790 6375 20798 6409
rect 20832 6375 20842 6409
rect 20790 6363 20842 6375
rect 20872 6545 20924 6563
rect 20872 6511 20882 6545
rect 20916 6511 20924 6545
rect 20872 6477 20924 6511
rect 20872 6443 20882 6477
rect 20916 6443 20924 6477
rect 20872 6409 20924 6443
rect 20872 6375 20882 6409
rect 20916 6375 20924 6409
rect 21060 6529 21072 6563
rect 21106 6529 21118 6563
rect 21060 6495 21118 6529
rect 21060 6461 21072 6495
rect 21106 6461 21118 6495
rect 21060 6427 21118 6461
rect 21060 6393 21072 6427
rect 21106 6393 21118 6427
rect 21060 6378 21118 6393
rect 21148 6563 21206 6578
rect 21148 6529 21160 6563
rect 21194 6529 21206 6563
rect 21386 6553 21398 6587
rect 21432 6553 21448 6587
rect 21386 6538 21448 6553
rect 21478 6723 21544 6738
rect 21478 6689 21494 6723
rect 21528 6689 21544 6723
rect 21478 6655 21544 6689
rect 21478 6621 21494 6655
rect 21528 6621 21544 6655
rect 21478 6587 21544 6621
rect 21478 6553 21494 6587
rect 21528 6553 21544 6587
rect 21478 6538 21544 6553
rect 21574 6723 21636 6738
rect 21574 6689 21590 6723
rect 21624 6689 21636 6723
rect 21574 6655 21636 6689
rect 21574 6621 21590 6655
rect 21624 6621 21636 6655
rect 21574 6587 21636 6621
rect 23274 6723 23336 6738
rect 23274 6689 23286 6723
rect 23320 6689 23336 6723
rect 21574 6553 21590 6587
rect 21624 6553 21636 6587
rect 21574 6538 21636 6553
rect 21706 6563 21764 6578
rect 21148 6495 21206 6529
rect 21148 6461 21160 6495
rect 21194 6461 21206 6495
rect 21148 6427 21206 6461
rect 21706 6529 21718 6563
rect 21752 6529 21764 6563
rect 21706 6495 21764 6529
rect 21706 6461 21718 6495
rect 21752 6461 21764 6495
rect 21148 6393 21160 6427
rect 21194 6393 21206 6427
rect 21148 6378 21206 6393
rect 20872 6363 20924 6375
rect 21706 6427 21764 6461
rect 21706 6393 21718 6427
rect 21752 6393 21764 6427
rect 21706 6378 21764 6393
rect 21794 6563 21852 6578
rect 21794 6529 21806 6563
rect 21840 6529 21852 6563
rect 21794 6495 21852 6529
rect 21794 6461 21806 6495
rect 21840 6461 21852 6495
rect 21794 6427 21852 6461
rect 21794 6393 21806 6427
rect 21840 6393 21852 6427
rect 21794 6378 21852 6393
rect 21986 6553 22038 6571
rect 21986 6519 21994 6553
rect 22028 6519 22038 6553
rect 21986 6485 22038 6519
rect 21986 6451 21994 6485
rect 22028 6451 22038 6485
rect 21986 6417 22038 6451
rect 21986 6383 21994 6417
rect 22028 6383 22038 6417
rect 21986 6371 22038 6383
rect 22068 6553 22120 6571
rect 22068 6519 22078 6553
rect 22112 6519 22120 6553
rect 23274 6655 23336 6689
rect 23274 6621 23286 6655
rect 23320 6621 23336 6655
rect 23274 6587 23336 6621
rect 22948 6563 23006 6578
rect 22678 6545 22730 6563
rect 22068 6485 22120 6519
rect 22068 6451 22078 6485
rect 22112 6451 22120 6485
rect 22068 6417 22120 6451
rect 22068 6383 22078 6417
rect 22112 6383 22120 6417
rect 22068 6371 22120 6383
rect 22285 6500 22337 6523
rect 22285 6466 22293 6500
rect 22327 6466 22337 6500
rect 22285 6419 22337 6466
rect 22285 6385 22293 6419
rect 22327 6385 22337 6419
rect 22285 6365 22337 6385
rect 22367 6487 22425 6523
rect 22367 6453 22379 6487
rect 22413 6453 22425 6487
rect 22367 6419 22425 6453
rect 22367 6385 22379 6419
rect 22413 6385 22425 6419
rect 22367 6365 22425 6385
rect 22455 6487 22507 6523
rect 22455 6453 22465 6487
rect 22499 6453 22507 6487
rect 22455 6419 22507 6453
rect 22455 6385 22465 6419
rect 22499 6385 22507 6419
rect 22455 6365 22507 6385
rect 22678 6511 22686 6545
rect 22720 6511 22730 6545
rect 22678 6477 22730 6511
rect 22678 6443 22686 6477
rect 22720 6443 22730 6477
rect 22678 6409 22730 6443
rect 22678 6375 22686 6409
rect 22720 6375 22730 6409
rect 22678 6363 22730 6375
rect 22760 6545 22812 6563
rect 22760 6511 22770 6545
rect 22804 6511 22812 6545
rect 22760 6477 22812 6511
rect 22760 6443 22770 6477
rect 22804 6443 22812 6477
rect 22760 6409 22812 6443
rect 22760 6375 22770 6409
rect 22804 6375 22812 6409
rect 22948 6529 22960 6563
rect 22994 6529 23006 6563
rect 22948 6495 23006 6529
rect 22948 6461 22960 6495
rect 22994 6461 23006 6495
rect 22948 6427 23006 6461
rect 22948 6393 22960 6427
rect 22994 6393 23006 6427
rect 22948 6378 23006 6393
rect 23036 6563 23094 6578
rect 23036 6529 23048 6563
rect 23082 6529 23094 6563
rect 23274 6553 23286 6587
rect 23320 6553 23336 6587
rect 23274 6538 23336 6553
rect 23366 6723 23432 6738
rect 23366 6689 23382 6723
rect 23416 6689 23432 6723
rect 23366 6655 23432 6689
rect 23366 6621 23382 6655
rect 23416 6621 23432 6655
rect 23366 6587 23432 6621
rect 23366 6553 23382 6587
rect 23416 6553 23432 6587
rect 23366 6538 23432 6553
rect 23462 6723 23524 6738
rect 23462 6689 23478 6723
rect 23512 6689 23524 6723
rect 23462 6655 23524 6689
rect 23462 6621 23478 6655
rect 23512 6621 23524 6655
rect 23462 6587 23524 6621
rect 25162 6723 25224 6738
rect 25162 6689 25174 6723
rect 25208 6689 25224 6723
rect 23462 6553 23478 6587
rect 23512 6553 23524 6587
rect 23462 6538 23524 6553
rect 23594 6563 23652 6578
rect 23036 6495 23094 6529
rect 23036 6461 23048 6495
rect 23082 6461 23094 6495
rect 23036 6427 23094 6461
rect 23594 6529 23606 6563
rect 23640 6529 23652 6563
rect 23594 6495 23652 6529
rect 23594 6461 23606 6495
rect 23640 6461 23652 6495
rect 23036 6393 23048 6427
rect 23082 6393 23094 6427
rect 23036 6378 23094 6393
rect 22760 6363 22812 6375
rect 23594 6427 23652 6461
rect 23594 6393 23606 6427
rect 23640 6393 23652 6427
rect 23594 6378 23652 6393
rect 23682 6563 23740 6578
rect 23682 6529 23694 6563
rect 23728 6529 23740 6563
rect 23682 6495 23740 6529
rect 23682 6461 23694 6495
rect 23728 6461 23740 6495
rect 23682 6427 23740 6461
rect 23682 6393 23694 6427
rect 23728 6393 23740 6427
rect 23682 6378 23740 6393
rect 23874 6553 23926 6571
rect 23874 6519 23882 6553
rect 23916 6519 23926 6553
rect 23874 6485 23926 6519
rect 23874 6451 23882 6485
rect 23916 6451 23926 6485
rect 23874 6417 23926 6451
rect 23874 6383 23882 6417
rect 23916 6383 23926 6417
rect 23874 6371 23926 6383
rect 23956 6553 24008 6571
rect 23956 6519 23966 6553
rect 24000 6519 24008 6553
rect 25162 6655 25224 6689
rect 25162 6621 25174 6655
rect 25208 6621 25224 6655
rect 25162 6587 25224 6621
rect 24836 6563 24894 6578
rect 24566 6545 24618 6563
rect 23956 6485 24008 6519
rect 23956 6451 23966 6485
rect 24000 6451 24008 6485
rect 23956 6417 24008 6451
rect 23956 6383 23966 6417
rect 24000 6383 24008 6417
rect 23956 6371 24008 6383
rect 24173 6500 24225 6523
rect 24173 6466 24181 6500
rect 24215 6466 24225 6500
rect 24173 6419 24225 6466
rect 24173 6385 24181 6419
rect 24215 6385 24225 6419
rect 24173 6365 24225 6385
rect 24255 6487 24313 6523
rect 24255 6453 24267 6487
rect 24301 6453 24313 6487
rect 24255 6419 24313 6453
rect 24255 6385 24267 6419
rect 24301 6385 24313 6419
rect 24255 6365 24313 6385
rect 24343 6487 24395 6523
rect 24343 6453 24353 6487
rect 24387 6453 24395 6487
rect 24343 6419 24395 6453
rect 24343 6385 24353 6419
rect 24387 6385 24395 6419
rect 24343 6365 24395 6385
rect 24566 6511 24574 6545
rect 24608 6511 24618 6545
rect 24566 6477 24618 6511
rect 24566 6443 24574 6477
rect 24608 6443 24618 6477
rect 24566 6409 24618 6443
rect 24566 6375 24574 6409
rect 24608 6375 24618 6409
rect 24566 6363 24618 6375
rect 24648 6545 24700 6563
rect 24648 6511 24658 6545
rect 24692 6511 24700 6545
rect 24648 6477 24700 6511
rect 24648 6443 24658 6477
rect 24692 6443 24700 6477
rect 24648 6409 24700 6443
rect 24648 6375 24658 6409
rect 24692 6375 24700 6409
rect 24836 6529 24848 6563
rect 24882 6529 24894 6563
rect 24836 6495 24894 6529
rect 24836 6461 24848 6495
rect 24882 6461 24894 6495
rect 24836 6427 24894 6461
rect 24836 6393 24848 6427
rect 24882 6393 24894 6427
rect 24836 6378 24894 6393
rect 24924 6563 24982 6578
rect 24924 6529 24936 6563
rect 24970 6529 24982 6563
rect 25162 6553 25174 6587
rect 25208 6553 25224 6587
rect 25162 6538 25224 6553
rect 25254 6723 25320 6738
rect 25254 6689 25270 6723
rect 25304 6689 25320 6723
rect 25254 6655 25320 6689
rect 25254 6621 25270 6655
rect 25304 6621 25320 6655
rect 25254 6587 25320 6621
rect 25254 6553 25270 6587
rect 25304 6553 25320 6587
rect 25254 6538 25320 6553
rect 25350 6723 25412 6738
rect 25350 6689 25366 6723
rect 25400 6689 25412 6723
rect 25350 6655 25412 6689
rect 25350 6621 25366 6655
rect 25400 6621 25412 6655
rect 25350 6587 25412 6621
rect 27050 6723 27112 6738
rect 27050 6689 27062 6723
rect 27096 6689 27112 6723
rect 25350 6553 25366 6587
rect 25400 6553 25412 6587
rect 25350 6538 25412 6553
rect 25482 6563 25540 6578
rect 24924 6495 24982 6529
rect 24924 6461 24936 6495
rect 24970 6461 24982 6495
rect 24924 6427 24982 6461
rect 25482 6529 25494 6563
rect 25528 6529 25540 6563
rect 25482 6495 25540 6529
rect 25482 6461 25494 6495
rect 25528 6461 25540 6495
rect 24924 6393 24936 6427
rect 24970 6393 24982 6427
rect 24924 6378 24982 6393
rect 24648 6363 24700 6375
rect 25482 6427 25540 6461
rect 25482 6393 25494 6427
rect 25528 6393 25540 6427
rect 25482 6378 25540 6393
rect 25570 6563 25628 6578
rect 25570 6529 25582 6563
rect 25616 6529 25628 6563
rect 25570 6495 25628 6529
rect 25570 6461 25582 6495
rect 25616 6461 25628 6495
rect 25570 6427 25628 6461
rect 25570 6393 25582 6427
rect 25616 6393 25628 6427
rect 25570 6378 25628 6393
rect 25762 6553 25814 6571
rect 25762 6519 25770 6553
rect 25804 6519 25814 6553
rect 25762 6485 25814 6519
rect 25762 6451 25770 6485
rect 25804 6451 25814 6485
rect 25762 6417 25814 6451
rect 25762 6383 25770 6417
rect 25804 6383 25814 6417
rect 25762 6371 25814 6383
rect 25844 6553 25896 6571
rect 25844 6519 25854 6553
rect 25888 6519 25896 6553
rect 27050 6655 27112 6689
rect 27050 6621 27062 6655
rect 27096 6621 27112 6655
rect 27050 6587 27112 6621
rect 26724 6563 26782 6578
rect 26454 6545 26506 6563
rect 25844 6485 25896 6519
rect 25844 6451 25854 6485
rect 25888 6451 25896 6485
rect 25844 6417 25896 6451
rect 25844 6383 25854 6417
rect 25888 6383 25896 6417
rect 25844 6371 25896 6383
rect 26061 6500 26113 6523
rect 26061 6466 26069 6500
rect 26103 6466 26113 6500
rect 26061 6419 26113 6466
rect 26061 6385 26069 6419
rect 26103 6385 26113 6419
rect 26061 6365 26113 6385
rect 26143 6487 26201 6523
rect 26143 6453 26155 6487
rect 26189 6453 26201 6487
rect 26143 6419 26201 6453
rect 26143 6385 26155 6419
rect 26189 6385 26201 6419
rect 26143 6365 26201 6385
rect 26231 6487 26283 6523
rect 26231 6453 26241 6487
rect 26275 6453 26283 6487
rect 26231 6419 26283 6453
rect 26231 6385 26241 6419
rect 26275 6385 26283 6419
rect 26231 6365 26283 6385
rect 26454 6511 26462 6545
rect 26496 6511 26506 6545
rect 26454 6477 26506 6511
rect 26454 6443 26462 6477
rect 26496 6443 26506 6477
rect 26454 6409 26506 6443
rect 26454 6375 26462 6409
rect 26496 6375 26506 6409
rect 26454 6363 26506 6375
rect 26536 6545 26588 6563
rect 26536 6511 26546 6545
rect 26580 6511 26588 6545
rect 26536 6477 26588 6511
rect 26536 6443 26546 6477
rect 26580 6443 26588 6477
rect 26536 6409 26588 6443
rect 26536 6375 26546 6409
rect 26580 6375 26588 6409
rect 26724 6529 26736 6563
rect 26770 6529 26782 6563
rect 26724 6495 26782 6529
rect 26724 6461 26736 6495
rect 26770 6461 26782 6495
rect 26724 6427 26782 6461
rect 26724 6393 26736 6427
rect 26770 6393 26782 6427
rect 26724 6378 26782 6393
rect 26812 6563 26870 6578
rect 26812 6529 26824 6563
rect 26858 6529 26870 6563
rect 27050 6553 27062 6587
rect 27096 6553 27112 6587
rect 27050 6538 27112 6553
rect 27142 6723 27208 6738
rect 27142 6689 27158 6723
rect 27192 6689 27208 6723
rect 27142 6655 27208 6689
rect 27142 6621 27158 6655
rect 27192 6621 27208 6655
rect 27142 6587 27208 6621
rect 27142 6553 27158 6587
rect 27192 6553 27208 6587
rect 27142 6538 27208 6553
rect 27238 6723 27300 6738
rect 27238 6689 27254 6723
rect 27288 6689 27300 6723
rect 27238 6655 27300 6689
rect 27238 6621 27254 6655
rect 27288 6621 27300 6655
rect 27238 6587 27300 6621
rect 28938 6723 29000 6738
rect 28938 6689 28950 6723
rect 28984 6689 29000 6723
rect 27238 6553 27254 6587
rect 27288 6553 27300 6587
rect 27238 6538 27300 6553
rect 27370 6563 27428 6578
rect 26812 6495 26870 6529
rect 26812 6461 26824 6495
rect 26858 6461 26870 6495
rect 26812 6427 26870 6461
rect 27370 6529 27382 6563
rect 27416 6529 27428 6563
rect 27370 6495 27428 6529
rect 27370 6461 27382 6495
rect 27416 6461 27428 6495
rect 26812 6393 26824 6427
rect 26858 6393 26870 6427
rect 26812 6378 26870 6393
rect 26536 6363 26588 6375
rect 27370 6427 27428 6461
rect 27370 6393 27382 6427
rect 27416 6393 27428 6427
rect 27370 6378 27428 6393
rect 27458 6563 27516 6578
rect 27458 6529 27470 6563
rect 27504 6529 27516 6563
rect 27458 6495 27516 6529
rect 27458 6461 27470 6495
rect 27504 6461 27516 6495
rect 27458 6427 27516 6461
rect 27458 6393 27470 6427
rect 27504 6393 27516 6427
rect 27458 6378 27516 6393
rect 27650 6553 27702 6571
rect 27650 6519 27658 6553
rect 27692 6519 27702 6553
rect 27650 6485 27702 6519
rect 27650 6451 27658 6485
rect 27692 6451 27702 6485
rect 27650 6417 27702 6451
rect 27650 6383 27658 6417
rect 27692 6383 27702 6417
rect 27650 6371 27702 6383
rect 27732 6553 27784 6571
rect 27732 6519 27742 6553
rect 27776 6519 27784 6553
rect 28938 6655 29000 6689
rect 28938 6621 28950 6655
rect 28984 6621 29000 6655
rect 28938 6587 29000 6621
rect 28612 6563 28670 6578
rect 28342 6545 28394 6563
rect 27732 6485 27784 6519
rect 27732 6451 27742 6485
rect 27776 6451 27784 6485
rect 27732 6417 27784 6451
rect 27732 6383 27742 6417
rect 27776 6383 27784 6417
rect 27732 6371 27784 6383
rect 27949 6500 28001 6523
rect 27949 6466 27957 6500
rect 27991 6466 28001 6500
rect 27949 6419 28001 6466
rect 27949 6385 27957 6419
rect 27991 6385 28001 6419
rect 27949 6365 28001 6385
rect 28031 6487 28089 6523
rect 28031 6453 28043 6487
rect 28077 6453 28089 6487
rect 28031 6419 28089 6453
rect 28031 6385 28043 6419
rect 28077 6385 28089 6419
rect 28031 6365 28089 6385
rect 28119 6487 28171 6523
rect 28119 6453 28129 6487
rect 28163 6453 28171 6487
rect 28119 6419 28171 6453
rect 28119 6385 28129 6419
rect 28163 6385 28171 6419
rect 28119 6365 28171 6385
rect 28342 6511 28350 6545
rect 28384 6511 28394 6545
rect 28342 6477 28394 6511
rect 28342 6443 28350 6477
rect 28384 6443 28394 6477
rect 28342 6409 28394 6443
rect 28342 6375 28350 6409
rect 28384 6375 28394 6409
rect 28342 6363 28394 6375
rect 28424 6545 28476 6563
rect 28424 6511 28434 6545
rect 28468 6511 28476 6545
rect 28424 6477 28476 6511
rect 28424 6443 28434 6477
rect 28468 6443 28476 6477
rect 28424 6409 28476 6443
rect 28424 6375 28434 6409
rect 28468 6375 28476 6409
rect 28612 6529 28624 6563
rect 28658 6529 28670 6563
rect 28612 6495 28670 6529
rect 28612 6461 28624 6495
rect 28658 6461 28670 6495
rect 28612 6427 28670 6461
rect 28612 6393 28624 6427
rect 28658 6393 28670 6427
rect 28612 6378 28670 6393
rect 28700 6563 28758 6578
rect 28700 6529 28712 6563
rect 28746 6529 28758 6563
rect 28938 6553 28950 6587
rect 28984 6553 29000 6587
rect 28938 6538 29000 6553
rect 29030 6723 29096 6738
rect 29030 6689 29046 6723
rect 29080 6689 29096 6723
rect 29030 6655 29096 6689
rect 29030 6621 29046 6655
rect 29080 6621 29096 6655
rect 29030 6587 29096 6621
rect 29030 6553 29046 6587
rect 29080 6553 29096 6587
rect 29030 6538 29096 6553
rect 29126 6723 29188 6738
rect 29126 6689 29142 6723
rect 29176 6689 29188 6723
rect 29126 6655 29188 6689
rect 29126 6621 29142 6655
rect 29176 6621 29188 6655
rect 29126 6587 29188 6621
rect 30826 6723 30888 6738
rect 30826 6689 30838 6723
rect 30872 6689 30888 6723
rect 29126 6553 29142 6587
rect 29176 6553 29188 6587
rect 29126 6538 29188 6553
rect 29258 6563 29316 6578
rect 28700 6495 28758 6529
rect 28700 6461 28712 6495
rect 28746 6461 28758 6495
rect 28700 6427 28758 6461
rect 29258 6529 29270 6563
rect 29304 6529 29316 6563
rect 29258 6495 29316 6529
rect 29258 6461 29270 6495
rect 29304 6461 29316 6495
rect 28700 6393 28712 6427
rect 28746 6393 28758 6427
rect 28700 6378 28758 6393
rect 28424 6363 28476 6375
rect 29258 6427 29316 6461
rect 29258 6393 29270 6427
rect 29304 6393 29316 6427
rect 29258 6378 29316 6393
rect 29346 6563 29404 6578
rect 29346 6529 29358 6563
rect 29392 6529 29404 6563
rect 29346 6495 29404 6529
rect 29346 6461 29358 6495
rect 29392 6461 29404 6495
rect 29346 6427 29404 6461
rect 29346 6393 29358 6427
rect 29392 6393 29404 6427
rect 29346 6378 29404 6393
rect 29538 6553 29590 6571
rect 29538 6519 29546 6553
rect 29580 6519 29590 6553
rect 29538 6485 29590 6519
rect 29538 6451 29546 6485
rect 29580 6451 29590 6485
rect 29538 6417 29590 6451
rect 29538 6383 29546 6417
rect 29580 6383 29590 6417
rect 29538 6371 29590 6383
rect 29620 6553 29672 6571
rect 29620 6519 29630 6553
rect 29664 6519 29672 6553
rect 30826 6655 30888 6689
rect 30826 6621 30838 6655
rect 30872 6621 30888 6655
rect 30826 6587 30888 6621
rect 30500 6563 30558 6578
rect 30230 6545 30282 6563
rect 29620 6485 29672 6519
rect 29620 6451 29630 6485
rect 29664 6451 29672 6485
rect 29620 6417 29672 6451
rect 29620 6383 29630 6417
rect 29664 6383 29672 6417
rect 29620 6371 29672 6383
rect 29837 6500 29889 6523
rect 29837 6466 29845 6500
rect 29879 6466 29889 6500
rect 29837 6419 29889 6466
rect 29837 6385 29845 6419
rect 29879 6385 29889 6419
rect 29837 6365 29889 6385
rect 29919 6487 29977 6523
rect 29919 6453 29931 6487
rect 29965 6453 29977 6487
rect 29919 6419 29977 6453
rect 29919 6385 29931 6419
rect 29965 6385 29977 6419
rect 29919 6365 29977 6385
rect 30007 6487 30059 6523
rect 30007 6453 30017 6487
rect 30051 6453 30059 6487
rect 30007 6419 30059 6453
rect 30007 6385 30017 6419
rect 30051 6385 30059 6419
rect 30007 6365 30059 6385
rect 30230 6511 30238 6545
rect 30272 6511 30282 6545
rect 30230 6477 30282 6511
rect 30230 6443 30238 6477
rect 30272 6443 30282 6477
rect 30230 6409 30282 6443
rect 30230 6375 30238 6409
rect 30272 6375 30282 6409
rect 30230 6363 30282 6375
rect 30312 6545 30364 6563
rect 30312 6511 30322 6545
rect 30356 6511 30364 6545
rect 30312 6477 30364 6511
rect 30312 6443 30322 6477
rect 30356 6443 30364 6477
rect 30312 6409 30364 6443
rect 30312 6375 30322 6409
rect 30356 6375 30364 6409
rect 30500 6529 30512 6563
rect 30546 6529 30558 6563
rect 30500 6495 30558 6529
rect 30500 6461 30512 6495
rect 30546 6461 30558 6495
rect 30500 6427 30558 6461
rect 30500 6393 30512 6427
rect 30546 6393 30558 6427
rect 30500 6378 30558 6393
rect 30588 6563 30646 6578
rect 30588 6529 30600 6563
rect 30634 6529 30646 6563
rect 30826 6553 30838 6587
rect 30872 6553 30888 6587
rect 30826 6538 30888 6553
rect 30918 6723 30984 6738
rect 30918 6689 30934 6723
rect 30968 6689 30984 6723
rect 30918 6655 30984 6689
rect 30918 6621 30934 6655
rect 30968 6621 30984 6655
rect 30918 6587 30984 6621
rect 30918 6553 30934 6587
rect 30968 6553 30984 6587
rect 30918 6538 30984 6553
rect 31014 6723 31076 6738
rect 31014 6689 31030 6723
rect 31064 6689 31076 6723
rect 31014 6655 31076 6689
rect 31014 6621 31030 6655
rect 31064 6621 31076 6655
rect 31014 6587 31076 6621
rect 32714 6723 32776 6738
rect 32714 6689 32726 6723
rect 32760 6689 32776 6723
rect 31014 6553 31030 6587
rect 31064 6553 31076 6587
rect 31014 6538 31076 6553
rect 31146 6563 31204 6578
rect 30588 6495 30646 6529
rect 30588 6461 30600 6495
rect 30634 6461 30646 6495
rect 30588 6427 30646 6461
rect 31146 6529 31158 6563
rect 31192 6529 31204 6563
rect 31146 6495 31204 6529
rect 31146 6461 31158 6495
rect 31192 6461 31204 6495
rect 30588 6393 30600 6427
rect 30634 6393 30646 6427
rect 30588 6378 30646 6393
rect 30312 6363 30364 6375
rect 31146 6427 31204 6461
rect 31146 6393 31158 6427
rect 31192 6393 31204 6427
rect 31146 6378 31204 6393
rect 31234 6563 31292 6578
rect 31234 6529 31246 6563
rect 31280 6529 31292 6563
rect 31234 6495 31292 6529
rect 31234 6461 31246 6495
rect 31280 6461 31292 6495
rect 31234 6427 31292 6461
rect 31234 6393 31246 6427
rect 31280 6393 31292 6427
rect 31234 6378 31292 6393
rect 31426 6553 31478 6571
rect 31426 6519 31434 6553
rect 31468 6519 31478 6553
rect 31426 6485 31478 6519
rect 31426 6451 31434 6485
rect 31468 6451 31478 6485
rect 31426 6417 31478 6451
rect 31426 6383 31434 6417
rect 31468 6383 31478 6417
rect 31426 6371 31478 6383
rect 31508 6553 31560 6571
rect 31508 6519 31518 6553
rect 31552 6519 31560 6553
rect 32714 6655 32776 6689
rect 32714 6621 32726 6655
rect 32760 6621 32776 6655
rect 32714 6587 32776 6621
rect 32388 6563 32446 6578
rect 32118 6545 32170 6563
rect 31508 6485 31560 6519
rect 31508 6451 31518 6485
rect 31552 6451 31560 6485
rect 31508 6417 31560 6451
rect 31508 6383 31518 6417
rect 31552 6383 31560 6417
rect 31508 6371 31560 6383
rect 31725 6500 31777 6523
rect 31725 6466 31733 6500
rect 31767 6466 31777 6500
rect 31725 6419 31777 6466
rect 31725 6385 31733 6419
rect 31767 6385 31777 6419
rect 31725 6365 31777 6385
rect 31807 6487 31865 6523
rect 31807 6453 31819 6487
rect 31853 6453 31865 6487
rect 31807 6419 31865 6453
rect 31807 6385 31819 6419
rect 31853 6385 31865 6419
rect 31807 6365 31865 6385
rect 31895 6487 31947 6523
rect 31895 6453 31905 6487
rect 31939 6453 31947 6487
rect 31895 6419 31947 6453
rect 31895 6385 31905 6419
rect 31939 6385 31947 6419
rect 31895 6365 31947 6385
rect 32118 6511 32126 6545
rect 32160 6511 32170 6545
rect 32118 6477 32170 6511
rect 32118 6443 32126 6477
rect 32160 6443 32170 6477
rect 32118 6409 32170 6443
rect 32118 6375 32126 6409
rect 32160 6375 32170 6409
rect 32118 6363 32170 6375
rect 32200 6545 32252 6563
rect 32200 6511 32210 6545
rect 32244 6511 32252 6545
rect 32200 6477 32252 6511
rect 32200 6443 32210 6477
rect 32244 6443 32252 6477
rect 32200 6409 32252 6443
rect 32200 6375 32210 6409
rect 32244 6375 32252 6409
rect 32388 6529 32400 6563
rect 32434 6529 32446 6563
rect 32388 6495 32446 6529
rect 32388 6461 32400 6495
rect 32434 6461 32446 6495
rect 32388 6427 32446 6461
rect 32388 6393 32400 6427
rect 32434 6393 32446 6427
rect 32388 6378 32446 6393
rect 32476 6563 32534 6578
rect 32476 6529 32488 6563
rect 32522 6529 32534 6563
rect 32714 6553 32726 6587
rect 32760 6553 32776 6587
rect 32714 6538 32776 6553
rect 32806 6723 32872 6738
rect 32806 6689 32822 6723
rect 32856 6689 32872 6723
rect 32806 6655 32872 6689
rect 32806 6621 32822 6655
rect 32856 6621 32872 6655
rect 32806 6587 32872 6621
rect 32806 6553 32822 6587
rect 32856 6553 32872 6587
rect 32806 6538 32872 6553
rect 32902 6723 32964 6738
rect 32902 6689 32918 6723
rect 32952 6689 32964 6723
rect 32902 6655 32964 6689
rect 32902 6621 32918 6655
rect 32952 6621 32964 6655
rect 32902 6587 32964 6621
rect 34602 6723 34664 6738
rect 34602 6689 34614 6723
rect 34648 6689 34664 6723
rect 32902 6553 32918 6587
rect 32952 6553 32964 6587
rect 32902 6538 32964 6553
rect 33034 6563 33092 6578
rect 32476 6495 32534 6529
rect 32476 6461 32488 6495
rect 32522 6461 32534 6495
rect 32476 6427 32534 6461
rect 33034 6529 33046 6563
rect 33080 6529 33092 6563
rect 33034 6495 33092 6529
rect 33034 6461 33046 6495
rect 33080 6461 33092 6495
rect 32476 6393 32488 6427
rect 32522 6393 32534 6427
rect 32476 6378 32534 6393
rect 32200 6363 32252 6375
rect 33034 6427 33092 6461
rect 33034 6393 33046 6427
rect 33080 6393 33092 6427
rect 33034 6378 33092 6393
rect 33122 6563 33180 6578
rect 33122 6529 33134 6563
rect 33168 6529 33180 6563
rect 33122 6495 33180 6529
rect 33122 6461 33134 6495
rect 33168 6461 33180 6495
rect 33122 6427 33180 6461
rect 33122 6393 33134 6427
rect 33168 6393 33180 6427
rect 33122 6378 33180 6393
rect 33314 6553 33366 6571
rect 33314 6519 33322 6553
rect 33356 6519 33366 6553
rect 33314 6485 33366 6519
rect 33314 6451 33322 6485
rect 33356 6451 33366 6485
rect 33314 6417 33366 6451
rect 33314 6383 33322 6417
rect 33356 6383 33366 6417
rect 33314 6371 33366 6383
rect 33396 6553 33448 6571
rect 33396 6519 33406 6553
rect 33440 6519 33448 6553
rect 34602 6655 34664 6689
rect 34602 6621 34614 6655
rect 34648 6621 34664 6655
rect 34602 6587 34664 6621
rect 34276 6563 34334 6578
rect 34006 6545 34058 6563
rect 33396 6485 33448 6519
rect 33396 6451 33406 6485
rect 33440 6451 33448 6485
rect 33396 6417 33448 6451
rect 33396 6383 33406 6417
rect 33440 6383 33448 6417
rect 33396 6371 33448 6383
rect 33613 6500 33665 6523
rect 33613 6466 33621 6500
rect 33655 6466 33665 6500
rect 33613 6419 33665 6466
rect 33613 6385 33621 6419
rect 33655 6385 33665 6419
rect 33613 6365 33665 6385
rect 33695 6487 33753 6523
rect 33695 6453 33707 6487
rect 33741 6453 33753 6487
rect 33695 6419 33753 6453
rect 33695 6385 33707 6419
rect 33741 6385 33753 6419
rect 33695 6365 33753 6385
rect 33783 6487 33835 6523
rect 33783 6453 33793 6487
rect 33827 6453 33835 6487
rect 33783 6419 33835 6453
rect 33783 6385 33793 6419
rect 33827 6385 33835 6419
rect 33783 6365 33835 6385
rect 34006 6511 34014 6545
rect 34048 6511 34058 6545
rect 34006 6477 34058 6511
rect 34006 6443 34014 6477
rect 34048 6443 34058 6477
rect 34006 6409 34058 6443
rect 34006 6375 34014 6409
rect 34048 6375 34058 6409
rect 34006 6363 34058 6375
rect 34088 6545 34140 6563
rect 34088 6511 34098 6545
rect 34132 6511 34140 6545
rect 34088 6477 34140 6511
rect 34088 6443 34098 6477
rect 34132 6443 34140 6477
rect 34088 6409 34140 6443
rect 34088 6375 34098 6409
rect 34132 6375 34140 6409
rect 34276 6529 34288 6563
rect 34322 6529 34334 6563
rect 34276 6495 34334 6529
rect 34276 6461 34288 6495
rect 34322 6461 34334 6495
rect 34276 6427 34334 6461
rect 34276 6393 34288 6427
rect 34322 6393 34334 6427
rect 34276 6378 34334 6393
rect 34364 6563 34422 6578
rect 34364 6529 34376 6563
rect 34410 6529 34422 6563
rect 34602 6553 34614 6587
rect 34648 6553 34664 6587
rect 34602 6538 34664 6553
rect 34694 6723 34760 6738
rect 34694 6689 34710 6723
rect 34744 6689 34760 6723
rect 34694 6655 34760 6689
rect 34694 6621 34710 6655
rect 34744 6621 34760 6655
rect 34694 6587 34760 6621
rect 34694 6553 34710 6587
rect 34744 6553 34760 6587
rect 34694 6538 34760 6553
rect 34790 6723 34852 6738
rect 34790 6689 34806 6723
rect 34840 6689 34852 6723
rect 34790 6655 34852 6689
rect 34790 6621 34806 6655
rect 34840 6621 34852 6655
rect 34790 6587 34852 6621
rect 36490 6723 36552 6738
rect 36490 6689 36502 6723
rect 36536 6689 36552 6723
rect 34790 6553 34806 6587
rect 34840 6553 34852 6587
rect 34790 6538 34852 6553
rect 34922 6563 34980 6578
rect 34364 6495 34422 6529
rect 34364 6461 34376 6495
rect 34410 6461 34422 6495
rect 34364 6427 34422 6461
rect 34922 6529 34934 6563
rect 34968 6529 34980 6563
rect 34922 6495 34980 6529
rect 34922 6461 34934 6495
rect 34968 6461 34980 6495
rect 34364 6393 34376 6427
rect 34410 6393 34422 6427
rect 34364 6378 34422 6393
rect 34088 6363 34140 6375
rect 34922 6427 34980 6461
rect 34922 6393 34934 6427
rect 34968 6393 34980 6427
rect 34922 6378 34980 6393
rect 35010 6563 35068 6578
rect 35010 6529 35022 6563
rect 35056 6529 35068 6563
rect 35010 6495 35068 6529
rect 35010 6461 35022 6495
rect 35056 6461 35068 6495
rect 35010 6427 35068 6461
rect 35010 6393 35022 6427
rect 35056 6393 35068 6427
rect 35010 6378 35068 6393
rect 35202 6553 35254 6571
rect 35202 6519 35210 6553
rect 35244 6519 35254 6553
rect 35202 6485 35254 6519
rect 35202 6451 35210 6485
rect 35244 6451 35254 6485
rect 35202 6417 35254 6451
rect 35202 6383 35210 6417
rect 35244 6383 35254 6417
rect 35202 6371 35254 6383
rect 35284 6553 35336 6571
rect 35284 6519 35294 6553
rect 35328 6519 35336 6553
rect 36490 6655 36552 6689
rect 36490 6621 36502 6655
rect 36536 6621 36552 6655
rect 36490 6587 36552 6621
rect 36164 6563 36222 6578
rect 35894 6545 35946 6563
rect 35284 6485 35336 6519
rect 35284 6451 35294 6485
rect 35328 6451 35336 6485
rect 35284 6417 35336 6451
rect 35284 6383 35294 6417
rect 35328 6383 35336 6417
rect 35284 6371 35336 6383
rect 35501 6500 35553 6523
rect 35501 6466 35509 6500
rect 35543 6466 35553 6500
rect 35501 6419 35553 6466
rect 35501 6385 35509 6419
rect 35543 6385 35553 6419
rect 35501 6365 35553 6385
rect 35583 6487 35641 6523
rect 35583 6453 35595 6487
rect 35629 6453 35641 6487
rect 35583 6419 35641 6453
rect 35583 6385 35595 6419
rect 35629 6385 35641 6419
rect 35583 6365 35641 6385
rect 35671 6487 35723 6523
rect 35671 6453 35681 6487
rect 35715 6453 35723 6487
rect 35671 6419 35723 6453
rect 35671 6385 35681 6419
rect 35715 6385 35723 6419
rect 35671 6365 35723 6385
rect 35894 6511 35902 6545
rect 35936 6511 35946 6545
rect 35894 6477 35946 6511
rect 35894 6443 35902 6477
rect 35936 6443 35946 6477
rect 35894 6409 35946 6443
rect 35894 6375 35902 6409
rect 35936 6375 35946 6409
rect 35894 6363 35946 6375
rect 35976 6545 36028 6563
rect 35976 6511 35986 6545
rect 36020 6511 36028 6545
rect 35976 6477 36028 6511
rect 35976 6443 35986 6477
rect 36020 6443 36028 6477
rect 35976 6409 36028 6443
rect 35976 6375 35986 6409
rect 36020 6375 36028 6409
rect 36164 6529 36176 6563
rect 36210 6529 36222 6563
rect 36164 6495 36222 6529
rect 36164 6461 36176 6495
rect 36210 6461 36222 6495
rect 36164 6427 36222 6461
rect 36164 6393 36176 6427
rect 36210 6393 36222 6427
rect 36164 6378 36222 6393
rect 36252 6563 36310 6578
rect 36252 6529 36264 6563
rect 36298 6529 36310 6563
rect 36490 6553 36502 6587
rect 36536 6553 36552 6587
rect 36490 6538 36552 6553
rect 36582 6723 36648 6738
rect 36582 6689 36598 6723
rect 36632 6689 36648 6723
rect 36582 6655 36648 6689
rect 36582 6621 36598 6655
rect 36632 6621 36648 6655
rect 36582 6587 36648 6621
rect 36582 6553 36598 6587
rect 36632 6553 36648 6587
rect 36582 6538 36648 6553
rect 36678 6723 36740 6738
rect 36678 6689 36694 6723
rect 36728 6689 36740 6723
rect 36678 6655 36740 6689
rect 36678 6621 36694 6655
rect 36728 6621 36740 6655
rect 36678 6587 36740 6621
rect 38378 6723 38440 6738
rect 38378 6689 38390 6723
rect 38424 6689 38440 6723
rect 36678 6553 36694 6587
rect 36728 6553 36740 6587
rect 36678 6538 36740 6553
rect 36810 6563 36868 6578
rect 36252 6495 36310 6529
rect 36252 6461 36264 6495
rect 36298 6461 36310 6495
rect 36252 6427 36310 6461
rect 36810 6529 36822 6563
rect 36856 6529 36868 6563
rect 36810 6495 36868 6529
rect 36810 6461 36822 6495
rect 36856 6461 36868 6495
rect 36252 6393 36264 6427
rect 36298 6393 36310 6427
rect 36252 6378 36310 6393
rect 35976 6363 36028 6375
rect 36810 6427 36868 6461
rect 36810 6393 36822 6427
rect 36856 6393 36868 6427
rect 36810 6378 36868 6393
rect 36898 6563 36956 6578
rect 36898 6529 36910 6563
rect 36944 6529 36956 6563
rect 36898 6495 36956 6529
rect 36898 6461 36910 6495
rect 36944 6461 36956 6495
rect 36898 6427 36956 6461
rect 36898 6393 36910 6427
rect 36944 6393 36956 6427
rect 36898 6378 36956 6393
rect 37090 6553 37142 6571
rect 37090 6519 37098 6553
rect 37132 6519 37142 6553
rect 37090 6485 37142 6519
rect 37090 6451 37098 6485
rect 37132 6451 37142 6485
rect 37090 6417 37142 6451
rect 37090 6383 37098 6417
rect 37132 6383 37142 6417
rect 37090 6371 37142 6383
rect 37172 6553 37224 6571
rect 37172 6519 37182 6553
rect 37216 6519 37224 6553
rect 38378 6655 38440 6689
rect 38378 6621 38390 6655
rect 38424 6621 38440 6655
rect 38378 6587 38440 6621
rect 38052 6563 38110 6578
rect 37782 6545 37834 6563
rect 37172 6485 37224 6519
rect 37172 6451 37182 6485
rect 37216 6451 37224 6485
rect 37172 6417 37224 6451
rect 37172 6383 37182 6417
rect 37216 6383 37224 6417
rect 37172 6371 37224 6383
rect 37389 6500 37441 6523
rect 37389 6466 37397 6500
rect 37431 6466 37441 6500
rect 37389 6419 37441 6466
rect 37389 6385 37397 6419
rect 37431 6385 37441 6419
rect 37389 6365 37441 6385
rect 37471 6487 37529 6523
rect 37471 6453 37483 6487
rect 37517 6453 37529 6487
rect 37471 6419 37529 6453
rect 37471 6385 37483 6419
rect 37517 6385 37529 6419
rect 37471 6365 37529 6385
rect 37559 6487 37611 6523
rect 37559 6453 37569 6487
rect 37603 6453 37611 6487
rect 37559 6419 37611 6453
rect 37559 6385 37569 6419
rect 37603 6385 37611 6419
rect 37559 6365 37611 6385
rect 37782 6511 37790 6545
rect 37824 6511 37834 6545
rect 37782 6477 37834 6511
rect 37782 6443 37790 6477
rect 37824 6443 37834 6477
rect 37782 6409 37834 6443
rect 37782 6375 37790 6409
rect 37824 6375 37834 6409
rect 37782 6363 37834 6375
rect 37864 6545 37916 6563
rect 37864 6511 37874 6545
rect 37908 6511 37916 6545
rect 37864 6477 37916 6511
rect 37864 6443 37874 6477
rect 37908 6443 37916 6477
rect 37864 6409 37916 6443
rect 37864 6375 37874 6409
rect 37908 6375 37916 6409
rect 38052 6529 38064 6563
rect 38098 6529 38110 6563
rect 38052 6495 38110 6529
rect 38052 6461 38064 6495
rect 38098 6461 38110 6495
rect 38052 6427 38110 6461
rect 38052 6393 38064 6427
rect 38098 6393 38110 6427
rect 38052 6378 38110 6393
rect 38140 6563 38198 6578
rect 38140 6529 38152 6563
rect 38186 6529 38198 6563
rect 38378 6553 38390 6587
rect 38424 6553 38440 6587
rect 38378 6538 38440 6553
rect 38470 6723 38536 6738
rect 38470 6689 38486 6723
rect 38520 6689 38536 6723
rect 38470 6655 38536 6689
rect 38470 6621 38486 6655
rect 38520 6621 38536 6655
rect 38470 6587 38536 6621
rect 38470 6553 38486 6587
rect 38520 6553 38536 6587
rect 38470 6538 38536 6553
rect 38566 6723 38628 6738
rect 38566 6689 38582 6723
rect 38616 6689 38628 6723
rect 38566 6655 38628 6689
rect 38566 6621 38582 6655
rect 38616 6621 38628 6655
rect 38566 6587 38628 6621
rect 40266 6723 40328 6738
rect 40266 6689 40278 6723
rect 40312 6689 40328 6723
rect 38566 6553 38582 6587
rect 38616 6553 38628 6587
rect 38566 6538 38628 6553
rect 38698 6563 38756 6578
rect 38140 6495 38198 6529
rect 38140 6461 38152 6495
rect 38186 6461 38198 6495
rect 38140 6427 38198 6461
rect 38698 6529 38710 6563
rect 38744 6529 38756 6563
rect 38698 6495 38756 6529
rect 38698 6461 38710 6495
rect 38744 6461 38756 6495
rect 38140 6393 38152 6427
rect 38186 6393 38198 6427
rect 38140 6378 38198 6393
rect 37864 6363 37916 6375
rect 38698 6427 38756 6461
rect 38698 6393 38710 6427
rect 38744 6393 38756 6427
rect 38698 6378 38756 6393
rect 38786 6563 38844 6578
rect 38786 6529 38798 6563
rect 38832 6529 38844 6563
rect 38786 6495 38844 6529
rect 38786 6461 38798 6495
rect 38832 6461 38844 6495
rect 38786 6427 38844 6461
rect 38786 6393 38798 6427
rect 38832 6393 38844 6427
rect 38786 6378 38844 6393
rect 38978 6553 39030 6571
rect 38978 6519 38986 6553
rect 39020 6519 39030 6553
rect 38978 6485 39030 6519
rect 38978 6451 38986 6485
rect 39020 6451 39030 6485
rect 38978 6417 39030 6451
rect 38978 6383 38986 6417
rect 39020 6383 39030 6417
rect 38978 6371 39030 6383
rect 39060 6553 39112 6571
rect 39060 6519 39070 6553
rect 39104 6519 39112 6553
rect 40266 6655 40328 6689
rect 40266 6621 40278 6655
rect 40312 6621 40328 6655
rect 40266 6587 40328 6621
rect 39940 6563 39998 6578
rect 39670 6545 39722 6563
rect 39060 6485 39112 6519
rect 39060 6451 39070 6485
rect 39104 6451 39112 6485
rect 39060 6417 39112 6451
rect 39060 6383 39070 6417
rect 39104 6383 39112 6417
rect 39060 6371 39112 6383
rect 39277 6500 39329 6523
rect 39277 6466 39285 6500
rect 39319 6466 39329 6500
rect 39277 6419 39329 6466
rect 39277 6385 39285 6419
rect 39319 6385 39329 6419
rect 39277 6365 39329 6385
rect 39359 6487 39417 6523
rect 39359 6453 39371 6487
rect 39405 6453 39417 6487
rect 39359 6419 39417 6453
rect 39359 6385 39371 6419
rect 39405 6385 39417 6419
rect 39359 6365 39417 6385
rect 39447 6487 39499 6523
rect 39447 6453 39457 6487
rect 39491 6453 39499 6487
rect 39447 6419 39499 6453
rect 39447 6385 39457 6419
rect 39491 6385 39499 6419
rect 39447 6365 39499 6385
rect 39670 6511 39678 6545
rect 39712 6511 39722 6545
rect 39670 6477 39722 6511
rect 39670 6443 39678 6477
rect 39712 6443 39722 6477
rect 39670 6409 39722 6443
rect 39670 6375 39678 6409
rect 39712 6375 39722 6409
rect 39670 6363 39722 6375
rect 39752 6545 39804 6563
rect 39752 6511 39762 6545
rect 39796 6511 39804 6545
rect 39752 6477 39804 6511
rect 39752 6443 39762 6477
rect 39796 6443 39804 6477
rect 39752 6409 39804 6443
rect 39752 6375 39762 6409
rect 39796 6375 39804 6409
rect 39940 6529 39952 6563
rect 39986 6529 39998 6563
rect 39940 6495 39998 6529
rect 39940 6461 39952 6495
rect 39986 6461 39998 6495
rect 39940 6427 39998 6461
rect 39940 6393 39952 6427
rect 39986 6393 39998 6427
rect 39940 6378 39998 6393
rect 40028 6563 40086 6578
rect 40028 6529 40040 6563
rect 40074 6529 40086 6563
rect 40266 6553 40278 6587
rect 40312 6553 40328 6587
rect 40266 6538 40328 6553
rect 40358 6723 40424 6738
rect 40358 6689 40374 6723
rect 40408 6689 40424 6723
rect 40358 6655 40424 6689
rect 40358 6621 40374 6655
rect 40408 6621 40424 6655
rect 40358 6587 40424 6621
rect 40358 6553 40374 6587
rect 40408 6553 40424 6587
rect 40358 6538 40424 6553
rect 40454 6723 40516 6738
rect 40454 6689 40470 6723
rect 40504 6689 40516 6723
rect 40454 6655 40516 6689
rect 40454 6621 40470 6655
rect 40504 6621 40516 6655
rect 40454 6587 40516 6621
rect 42154 6723 42216 6738
rect 42154 6689 42166 6723
rect 42200 6689 42216 6723
rect 40454 6553 40470 6587
rect 40504 6553 40516 6587
rect 40454 6538 40516 6553
rect 40586 6563 40644 6578
rect 40028 6495 40086 6529
rect 40028 6461 40040 6495
rect 40074 6461 40086 6495
rect 40028 6427 40086 6461
rect 40586 6529 40598 6563
rect 40632 6529 40644 6563
rect 40586 6495 40644 6529
rect 40586 6461 40598 6495
rect 40632 6461 40644 6495
rect 40028 6393 40040 6427
rect 40074 6393 40086 6427
rect 40028 6378 40086 6393
rect 39752 6363 39804 6375
rect 40586 6427 40644 6461
rect 40586 6393 40598 6427
rect 40632 6393 40644 6427
rect 40586 6378 40644 6393
rect 40674 6563 40732 6578
rect 40674 6529 40686 6563
rect 40720 6529 40732 6563
rect 40674 6495 40732 6529
rect 40674 6461 40686 6495
rect 40720 6461 40732 6495
rect 40674 6427 40732 6461
rect 40674 6393 40686 6427
rect 40720 6393 40732 6427
rect 40674 6378 40732 6393
rect 40866 6553 40918 6571
rect 40866 6519 40874 6553
rect 40908 6519 40918 6553
rect 40866 6485 40918 6519
rect 40866 6451 40874 6485
rect 40908 6451 40918 6485
rect 40866 6417 40918 6451
rect 40866 6383 40874 6417
rect 40908 6383 40918 6417
rect 40866 6371 40918 6383
rect 40948 6553 41000 6571
rect 40948 6519 40958 6553
rect 40992 6519 41000 6553
rect 42154 6655 42216 6689
rect 42154 6621 42166 6655
rect 42200 6621 42216 6655
rect 42154 6587 42216 6621
rect 41828 6563 41886 6578
rect 41558 6545 41610 6563
rect 40948 6485 41000 6519
rect 40948 6451 40958 6485
rect 40992 6451 41000 6485
rect 40948 6417 41000 6451
rect 40948 6383 40958 6417
rect 40992 6383 41000 6417
rect 40948 6371 41000 6383
rect 41165 6500 41217 6523
rect 41165 6466 41173 6500
rect 41207 6466 41217 6500
rect 41165 6419 41217 6466
rect 41165 6385 41173 6419
rect 41207 6385 41217 6419
rect 41165 6365 41217 6385
rect 41247 6487 41305 6523
rect 41247 6453 41259 6487
rect 41293 6453 41305 6487
rect 41247 6419 41305 6453
rect 41247 6385 41259 6419
rect 41293 6385 41305 6419
rect 41247 6365 41305 6385
rect 41335 6487 41387 6523
rect 41335 6453 41345 6487
rect 41379 6453 41387 6487
rect 41335 6419 41387 6453
rect 41335 6385 41345 6419
rect 41379 6385 41387 6419
rect 41335 6365 41387 6385
rect 41558 6511 41566 6545
rect 41600 6511 41610 6545
rect 41558 6477 41610 6511
rect 41558 6443 41566 6477
rect 41600 6443 41610 6477
rect 41558 6409 41610 6443
rect 41558 6375 41566 6409
rect 41600 6375 41610 6409
rect 41558 6363 41610 6375
rect 41640 6545 41692 6563
rect 41640 6511 41650 6545
rect 41684 6511 41692 6545
rect 41640 6477 41692 6511
rect 41640 6443 41650 6477
rect 41684 6443 41692 6477
rect 41640 6409 41692 6443
rect 41640 6375 41650 6409
rect 41684 6375 41692 6409
rect 41828 6529 41840 6563
rect 41874 6529 41886 6563
rect 41828 6495 41886 6529
rect 41828 6461 41840 6495
rect 41874 6461 41886 6495
rect 41828 6427 41886 6461
rect 41828 6393 41840 6427
rect 41874 6393 41886 6427
rect 41828 6378 41886 6393
rect 41916 6563 41974 6578
rect 41916 6529 41928 6563
rect 41962 6529 41974 6563
rect 42154 6553 42166 6587
rect 42200 6553 42216 6587
rect 42154 6538 42216 6553
rect 42246 6723 42312 6738
rect 42246 6689 42262 6723
rect 42296 6689 42312 6723
rect 42246 6655 42312 6689
rect 42246 6621 42262 6655
rect 42296 6621 42312 6655
rect 42246 6587 42312 6621
rect 42246 6553 42262 6587
rect 42296 6553 42312 6587
rect 42246 6538 42312 6553
rect 42342 6723 42404 6738
rect 42342 6689 42358 6723
rect 42392 6689 42404 6723
rect 42342 6655 42404 6689
rect 42342 6621 42358 6655
rect 42392 6621 42404 6655
rect 42342 6587 42404 6621
rect 44042 6723 44104 6738
rect 44042 6689 44054 6723
rect 44088 6689 44104 6723
rect 42342 6553 42358 6587
rect 42392 6553 42404 6587
rect 42342 6538 42404 6553
rect 42474 6563 42532 6578
rect 41916 6495 41974 6529
rect 41916 6461 41928 6495
rect 41962 6461 41974 6495
rect 41916 6427 41974 6461
rect 42474 6529 42486 6563
rect 42520 6529 42532 6563
rect 42474 6495 42532 6529
rect 42474 6461 42486 6495
rect 42520 6461 42532 6495
rect 41916 6393 41928 6427
rect 41962 6393 41974 6427
rect 41916 6378 41974 6393
rect 41640 6363 41692 6375
rect 42474 6427 42532 6461
rect 42474 6393 42486 6427
rect 42520 6393 42532 6427
rect 42474 6378 42532 6393
rect 42562 6563 42620 6578
rect 42562 6529 42574 6563
rect 42608 6529 42620 6563
rect 42562 6495 42620 6529
rect 42562 6461 42574 6495
rect 42608 6461 42620 6495
rect 42562 6427 42620 6461
rect 42562 6393 42574 6427
rect 42608 6393 42620 6427
rect 42562 6378 42620 6393
rect 42754 6553 42806 6571
rect 42754 6519 42762 6553
rect 42796 6519 42806 6553
rect 42754 6485 42806 6519
rect 42754 6451 42762 6485
rect 42796 6451 42806 6485
rect 42754 6417 42806 6451
rect 42754 6383 42762 6417
rect 42796 6383 42806 6417
rect 42754 6371 42806 6383
rect 42836 6553 42888 6571
rect 42836 6519 42846 6553
rect 42880 6519 42888 6553
rect 44042 6655 44104 6689
rect 44042 6621 44054 6655
rect 44088 6621 44104 6655
rect 44042 6587 44104 6621
rect 43716 6563 43774 6578
rect 43446 6545 43498 6563
rect 42836 6485 42888 6519
rect 42836 6451 42846 6485
rect 42880 6451 42888 6485
rect 42836 6417 42888 6451
rect 42836 6383 42846 6417
rect 42880 6383 42888 6417
rect 42836 6371 42888 6383
rect 43053 6500 43105 6523
rect 43053 6466 43061 6500
rect 43095 6466 43105 6500
rect 43053 6419 43105 6466
rect 43053 6385 43061 6419
rect 43095 6385 43105 6419
rect 43053 6365 43105 6385
rect 43135 6487 43193 6523
rect 43135 6453 43147 6487
rect 43181 6453 43193 6487
rect 43135 6419 43193 6453
rect 43135 6385 43147 6419
rect 43181 6385 43193 6419
rect 43135 6365 43193 6385
rect 43223 6487 43275 6523
rect 43223 6453 43233 6487
rect 43267 6453 43275 6487
rect 43223 6419 43275 6453
rect 43223 6385 43233 6419
rect 43267 6385 43275 6419
rect 43223 6365 43275 6385
rect 43446 6511 43454 6545
rect 43488 6511 43498 6545
rect 43446 6477 43498 6511
rect 43446 6443 43454 6477
rect 43488 6443 43498 6477
rect 43446 6409 43498 6443
rect 43446 6375 43454 6409
rect 43488 6375 43498 6409
rect 43446 6363 43498 6375
rect 43528 6545 43580 6563
rect 43528 6511 43538 6545
rect 43572 6511 43580 6545
rect 43528 6477 43580 6511
rect 43528 6443 43538 6477
rect 43572 6443 43580 6477
rect 43528 6409 43580 6443
rect 43528 6375 43538 6409
rect 43572 6375 43580 6409
rect 43716 6529 43728 6563
rect 43762 6529 43774 6563
rect 43716 6495 43774 6529
rect 43716 6461 43728 6495
rect 43762 6461 43774 6495
rect 43716 6427 43774 6461
rect 43716 6393 43728 6427
rect 43762 6393 43774 6427
rect 43716 6378 43774 6393
rect 43804 6563 43862 6578
rect 43804 6529 43816 6563
rect 43850 6529 43862 6563
rect 44042 6553 44054 6587
rect 44088 6553 44104 6587
rect 44042 6538 44104 6553
rect 44134 6723 44200 6738
rect 44134 6689 44150 6723
rect 44184 6689 44200 6723
rect 44134 6655 44200 6689
rect 44134 6621 44150 6655
rect 44184 6621 44200 6655
rect 44134 6587 44200 6621
rect 44134 6553 44150 6587
rect 44184 6553 44200 6587
rect 44134 6538 44200 6553
rect 44230 6723 44292 6738
rect 44230 6689 44246 6723
rect 44280 6689 44292 6723
rect 44230 6655 44292 6689
rect 44230 6621 44246 6655
rect 44280 6621 44292 6655
rect 44230 6587 44292 6621
rect 45924 6723 45986 6738
rect 45924 6689 45936 6723
rect 45970 6689 45986 6723
rect 44230 6553 44246 6587
rect 44280 6553 44292 6587
rect 44230 6538 44292 6553
rect 44362 6563 44420 6578
rect 43804 6495 43862 6529
rect 43804 6461 43816 6495
rect 43850 6461 43862 6495
rect 43804 6427 43862 6461
rect 44362 6529 44374 6563
rect 44408 6529 44420 6563
rect 44362 6495 44420 6529
rect 44362 6461 44374 6495
rect 44408 6461 44420 6495
rect 43804 6393 43816 6427
rect 43850 6393 43862 6427
rect 43804 6378 43862 6393
rect 43528 6363 43580 6375
rect 44362 6427 44420 6461
rect 44362 6393 44374 6427
rect 44408 6393 44420 6427
rect 44362 6378 44420 6393
rect 44450 6563 44508 6578
rect 44450 6529 44462 6563
rect 44496 6529 44508 6563
rect 44450 6495 44508 6529
rect 44450 6461 44462 6495
rect 44496 6461 44508 6495
rect 44450 6427 44508 6461
rect 44450 6393 44462 6427
rect 44496 6393 44508 6427
rect 44450 6378 44508 6393
rect 44642 6553 44694 6571
rect 44642 6519 44650 6553
rect 44684 6519 44694 6553
rect 44642 6485 44694 6519
rect 44642 6451 44650 6485
rect 44684 6451 44694 6485
rect 44642 6417 44694 6451
rect 44642 6383 44650 6417
rect 44684 6383 44694 6417
rect 44642 6371 44694 6383
rect 44724 6553 44776 6571
rect 44724 6519 44734 6553
rect 44768 6519 44776 6553
rect 45924 6655 45986 6689
rect 45924 6621 45936 6655
rect 45970 6621 45986 6655
rect 45924 6587 45986 6621
rect 45598 6563 45656 6578
rect 45328 6545 45380 6563
rect 44724 6485 44776 6519
rect 44724 6451 44734 6485
rect 44768 6451 44776 6485
rect 44724 6417 44776 6451
rect 44724 6383 44734 6417
rect 44768 6383 44776 6417
rect 44724 6371 44776 6383
rect 44935 6500 44987 6523
rect 44935 6466 44943 6500
rect 44977 6466 44987 6500
rect 44935 6419 44987 6466
rect 44935 6385 44943 6419
rect 44977 6385 44987 6419
rect 44935 6365 44987 6385
rect 45017 6487 45075 6523
rect 45017 6453 45029 6487
rect 45063 6453 45075 6487
rect 45017 6419 45075 6453
rect 45017 6385 45029 6419
rect 45063 6385 45075 6419
rect 45017 6365 45075 6385
rect 45105 6487 45157 6523
rect 45105 6453 45115 6487
rect 45149 6453 45157 6487
rect 45105 6419 45157 6453
rect 45105 6385 45115 6419
rect 45149 6385 45157 6419
rect 45105 6365 45157 6385
rect 45328 6511 45336 6545
rect 45370 6511 45380 6545
rect 45328 6477 45380 6511
rect 45328 6443 45336 6477
rect 45370 6443 45380 6477
rect 45328 6409 45380 6443
rect 45328 6375 45336 6409
rect 45370 6375 45380 6409
rect 45328 6363 45380 6375
rect 45410 6545 45462 6563
rect 45410 6511 45420 6545
rect 45454 6511 45462 6545
rect 45410 6477 45462 6511
rect 45410 6443 45420 6477
rect 45454 6443 45462 6477
rect 45410 6409 45462 6443
rect 45410 6375 45420 6409
rect 45454 6375 45462 6409
rect 45598 6529 45610 6563
rect 45644 6529 45656 6563
rect 45598 6495 45656 6529
rect 45598 6461 45610 6495
rect 45644 6461 45656 6495
rect 45598 6427 45656 6461
rect 45598 6393 45610 6427
rect 45644 6393 45656 6427
rect 45598 6378 45656 6393
rect 45686 6563 45744 6578
rect 45686 6529 45698 6563
rect 45732 6529 45744 6563
rect 45924 6553 45936 6587
rect 45970 6553 45986 6587
rect 45924 6538 45986 6553
rect 46016 6723 46082 6738
rect 46016 6689 46032 6723
rect 46066 6689 46082 6723
rect 46016 6655 46082 6689
rect 46016 6621 46032 6655
rect 46066 6621 46082 6655
rect 46016 6587 46082 6621
rect 46016 6553 46032 6587
rect 46066 6553 46082 6587
rect 46016 6538 46082 6553
rect 46112 6723 46174 6738
rect 46112 6689 46128 6723
rect 46162 6689 46174 6723
rect 46112 6655 46174 6689
rect 46112 6621 46128 6655
rect 46162 6621 46174 6655
rect 46112 6587 46174 6621
rect 47812 6723 47874 6738
rect 47812 6689 47824 6723
rect 47858 6689 47874 6723
rect 46112 6553 46128 6587
rect 46162 6553 46174 6587
rect 46112 6538 46174 6553
rect 46244 6563 46302 6578
rect 45686 6495 45744 6529
rect 45686 6461 45698 6495
rect 45732 6461 45744 6495
rect 45686 6427 45744 6461
rect 46244 6529 46256 6563
rect 46290 6529 46302 6563
rect 46244 6495 46302 6529
rect 46244 6461 46256 6495
rect 46290 6461 46302 6495
rect 45686 6393 45698 6427
rect 45732 6393 45744 6427
rect 45686 6378 45744 6393
rect 45410 6363 45462 6375
rect 46244 6427 46302 6461
rect 46244 6393 46256 6427
rect 46290 6393 46302 6427
rect 46244 6378 46302 6393
rect 46332 6563 46390 6578
rect 46332 6529 46344 6563
rect 46378 6529 46390 6563
rect 46332 6495 46390 6529
rect 46332 6461 46344 6495
rect 46378 6461 46390 6495
rect 46332 6427 46390 6461
rect 46332 6393 46344 6427
rect 46378 6393 46390 6427
rect 46332 6378 46390 6393
rect 46524 6553 46576 6571
rect 46524 6519 46532 6553
rect 46566 6519 46576 6553
rect 46524 6485 46576 6519
rect 46524 6451 46532 6485
rect 46566 6451 46576 6485
rect 46524 6417 46576 6451
rect 46524 6383 46532 6417
rect 46566 6383 46576 6417
rect 46524 6371 46576 6383
rect 46606 6553 46658 6571
rect 46606 6519 46616 6553
rect 46650 6519 46658 6553
rect 47812 6655 47874 6689
rect 47812 6621 47824 6655
rect 47858 6621 47874 6655
rect 47812 6587 47874 6621
rect 47486 6563 47544 6578
rect 47216 6545 47268 6563
rect 46606 6485 46658 6519
rect 46606 6451 46616 6485
rect 46650 6451 46658 6485
rect 46606 6417 46658 6451
rect 46606 6383 46616 6417
rect 46650 6383 46658 6417
rect 46606 6371 46658 6383
rect 46823 6500 46875 6523
rect 46823 6466 46831 6500
rect 46865 6466 46875 6500
rect 46823 6419 46875 6466
rect 46823 6385 46831 6419
rect 46865 6385 46875 6419
rect 46823 6365 46875 6385
rect 46905 6487 46963 6523
rect 46905 6453 46917 6487
rect 46951 6453 46963 6487
rect 46905 6419 46963 6453
rect 46905 6385 46917 6419
rect 46951 6385 46963 6419
rect 46905 6365 46963 6385
rect 46993 6487 47045 6523
rect 46993 6453 47003 6487
rect 47037 6453 47045 6487
rect 46993 6419 47045 6453
rect 46993 6385 47003 6419
rect 47037 6385 47045 6419
rect 46993 6365 47045 6385
rect 47216 6511 47224 6545
rect 47258 6511 47268 6545
rect 47216 6477 47268 6511
rect 47216 6443 47224 6477
rect 47258 6443 47268 6477
rect 47216 6409 47268 6443
rect 47216 6375 47224 6409
rect 47258 6375 47268 6409
rect 47216 6363 47268 6375
rect 47298 6545 47350 6563
rect 47298 6511 47308 6545
rect 47342 6511 47350 6545
rect 47298 6477 47350 6511
rect 47298 6443 47308 6477
rect 47342 6443 47350 6477
rect 47298 6409 47350 6443
rect 47298 6375 47308 6409
rect 47342 6375 47350 6409
rect 47486 6529 47498 6563
rect 47532 6529 47544 6563
rect 47486 6495 47544 6529
rect 47486 6461 47498 6495
rect 47532 6461 47544 6495
rect 47486 6427 47544 6461
rect 47486 6393 47498 6427
rect 47532 6393 47544 6427
rect 47486 6378 47544 6393
rect 47574 6563 47632 6578
rect 47574 6529 47586 6563
rect 47620 6529 47632 6563
rect 47812 6553 47824 6587
rect 47858 6553 47874 6587
rect 47812 6538 47874 6553
rect 47904 6723 47970 6738
rect 47904 6689 47920 6723
rect 47954 6689 47970 6723
rect 47904 6655 47970 6689
rect 47904 6621 47920 6655
rect 47954 6621 47970 6655
rect 47904 6587 47970 6621
rect 47904 6553 47920 6587
rect 47954 6553 47970 6587
rect 47904 6538 47970 6553
rect 48000 6723 48062 6738
rect 48000 6689 48016 6723
rect 48050 6689 48062 6723
rect 48000 6655 48062 6689
rect 48000 6621 48016 6655
rect 48050 6621 48062 6655
rect 48000 6587 48062 6621
rect 49700 6723 49762 6738
rect 49700 6689 49712 6723
rect 49746 6689 49762 6723
rect 48000 6553 48016 6587
rect 48050 6553 48062 6587
rect 48000 6538 48062 6553
rect 48132 6563 48190 6578
rect 47574 6495 47632 6529
rect 47574 6461 47586 6495
rect 47620 6461 47632 6495
rect 47574 6427 47632 6461
rect 48132 6529 48144 6563
rect 48178 6529 48190 6563
rect 48132 6495 48190 6529
rect 48132 6461 48144 6495
rect 48178 6461 48190 6495
rect 47574 6393 47586 6427
rect 47620 6393 47632 6427
rect 47574 6378 47632 6393
rect 47298 6363 47350 6375
rect 48132 6427 48190 6461
rect 48132 6393 48144 6427
rect 48178 6393 48190 6427
rect 48132 6378 48190 6393
rect 48220 6563 48278 6578
rect 48220 6529 48232 6563
rect 48266 6529 48278 6563
rect 48220 6495 48278 6529
rect 48220 6461 48232 6495
rect 48266 6461 48278 6495
rect 48220 6427 48278 6461
rect 48220 6393 48232 6427
rect 48266 6393 48278 6427
rect 48220 6378 48278 6393
rect 48412 6553 48464 6571
rect 48412 6519 48420 6553
rect 48454 6519 48464 6553
rect 48412 6485 48464 6519
rect 48412 6451 48420 6485
rect 48454 6451 48464 6485
rect 48412 6417 48464 6451
rect 48412 6383 48420 6417
rect 48454 6383 48464 6417
rect 48412 6371 48464 6383
rect 48494 6553 48546 6571
rect 48494 6519 48504 6553
rect 48538 6519 48546 6553
rect 49700 6655 49762 6689
rect 49700 6621 49712 6655
rect 49746 6621 49762 6655
rect 49700 6587 49762 6621
rect 49374 6563 49432 6578
rect 49104 6545 49156 6563
rect 48494 6485 48546 6519
rect 48494 6451 48504 6485
rect 48538 6451 48546 6485
rect 48494 6417 48546 6451
rect 48494 6383 48504 6417
rect 48538 6383 48546 6417
rect 48494 6371 48546 6383
rect 48711 6500 48763 6523
rect 48711 6466 48719 6500
rect 48753 6466 48763 6500
rect 48711 6419 48763 6466
rect 48711 6385 48719 6419
rect 48753 6385 48763 6419
rect 48711 6365 48763 6385
rect 48793 6487 48851 6523
rect 48793 6453 48805 6487
rect 48839 6453 48851 6487
rect 48793 6419 48851 6453
rect 48793 6385 48805 6419
rect 48839 6385 48851 6419
rect 48793 6365 48851 6385
rect 48881 6487 48933 6523
rect 48881 6453 48891 6487
rect 48925 6453 48933 6487
rect 48881 6419 48933 6453
rect 48881 6385 48891 6419
rect 48925 6385 48933 6419
rect 48881 6365 48933 6385
rect 49104 6511 49112 6545
rect 49146 6511 49156 6545
rect 49104 6477 49156 6511
rect 49104 6443 49112 6477
rect 49146 6443 49156 6477
rect 49104 6409 49156 6443
rect 49104 6375 49112 6409
rect 49146 6375 49156 6409
rect 49104 6363 49156 6375
rect 49186 6545 49238 6563
rect 49186 6511 49196 6545
rect 49230 6511 49238 6545
rect 49186 6477 49238 6511
rect 49186 6443 49196 6477
rect 49230 6443 49238 6477
rect 49186 6409 49238 6443
rect 49186 6375 49196 6409
rect 49230 6375 49238 6409
rect 49374 6529 49386 6563
rect 49420 6529 49432 6563
rect 49374 6495 49432 6529
rect 49374 6461 49386 6495
rect 49420 6461 49432 6495
rect 49374 6427 49432 6461
rect 49374 6393 49386 6427
rect 49420 6393 49432 6427
rect 49374 6378 49432 6393
rect 49462 6563 49520 6578
rect 49462 6529 49474 6563
rect 49508 6529 49520 6563
rect 49700 6553 49712 6587
rect 49746 6553 49762 6587
rect 49700 6538 49762 6553
rect 49792 6723 49858 6738
rect 49792 6689 49808 6723
rect 49842 6689 49858 6723
rect 49792 6655 49858 6689
rect 49792 6621 49808 6655
rect 49842 6621 49858 6655
rect 49792 6587 49858 6621
rect 49792 6553 49808 6587
rect 49842 6553 49858 6587
rect 49792 6538 49858 6553
rect 49888 6723 49950 6738
rect 49888 6689 49904 6723
rect 49938 6689 49950 6723
rect 49888 6655 49950 6689
rect 49888 6621 49904 6655
rect 49938 6621 49950 6655
rect 49888 6587 49950 6621
rect 51588 6723 51650 6738
rect 51588 6689 51600 6723
rect 51634 6689 51650 6723
rect 49888 6553 49904 6587
rect 49938 6553 49950 6587
rect 49888 6538 49950 6553
rect 50020 6563 50078 6578
rect 49462 6495 49520 6529
rect 49462 6461 49474 6495
rect 49508 6461 49520 6495
rect 49462 6427 49520 6461
rect 50020 6529 50032 6563
rect 50066 6529 50078 6563
rect 50020 6495 50078 6529
rect 50020 6461 50032 6495
rect 50066 6461 50078 6495
rect 49462 6393 49474 6427
rect 49508 6393 49520 6427
rect 49462 6378 49520 6393
rect 49186 6363 49238 6375
rect 50020 6427 50078 6461
rect 50020 6393 50032 6427
rect 50066 6393 50078 6427
rect 50020 6378 50078 6393
rect 50108 6563 50166 6578
rect 50108 6529 50120 6563
rect 50154 6529 50166 6563
rect 50108 6495 50166 6529
rect 50108 6461 50120 6495
rect 50154 6461 50166 6495
rect 50108 6427 50166 6461
rect 50108 6393 50120 6427
rect 50154 6393 50166 6427
rect 50108 6378 50166 6393
rect 50300 6553 50352 6571
rect 50300 6519 50308 6553
rect 50342 6519 50352 6553
rect 50300 6485 50352 6519
rect 50300 6451 50308 6485
rect 50342 6451 50352 6485
rect 50300 6417 50352 6451
rect 50300 6383 50308 6417
rect 50342 6383 50352 6417
rect 50300 6371 50352 6383
rect 50382 6553 50434 6571
rect 50382 6519 50392 6553
rect 50426 6519 50434 6553
rect 51588 6655 51650 6689
rect 51588 6621 51600 6655
rect 51634 6621 51650 6655
rect 51588 6587 51650 6621
rect 51262 6563 51320 6578
rect 50992 6545 51044 6563
rect 50382 6485 50434 6519
rect 50382 6451 50392 6485
rect 50426 6451 50434 6485
rect 50382 6417 50434 6451
rect 50382 6383 50392 6417
rect 50426 6383 50434 6417
rect 50382 6371 50434 6383
rect 50599 6500 50651 6523
rect 50599 6466 50607 6500
rect 50641 6466 50651 6500
rect 50599 6419 50651 6466
rect 50599 6385 50607 6419
rect 50641 6385 50651 6419
rect 50599 6365 50651 6385
rect 50681 6487 50739 6523
rect 50681 6453 50693 6487
rect 50727 6453 50739 6487
rect 50681 6419 50739 6453
rect 50681 6385 50693 6419
rect 50727 6385 50739 6419
rect 50681 6365 50739 6385
rect 50769 6487 50821 6523
rect 50769 6453 50779 6487
rect 50813 6453 50821 6487
rect 50769 6419 50821 6453
rect 50769 6385 50779 6419
rect 50813 6385 50821 6419
rect 50769 6365 50821 6385
rect 50992 6511 51000 6545
rect 51034 6511 51044 6545
rect 50992 6477 51044 6511
rect 50992 6443 51000 6477
rect 51034 6443 51044 6477
rect 50992 6409 51044 6443
rect 50992 6375 51000 6409
rect 51034 6375 51044 6409
rect 50992 6363 51044 6375
rect 51074 6545 51126 6563
rect 51074 6511 51084 6545
rect 51118 6511 51126 6545
rect 51074 6477 51126 6511
rect 51074 6443 51084 6477
rect 51118 6443 51126 6477
rect 51074 6409 51126 6443
rect 51074 6375 51084 6409
rect 51118 6375 51126 6409
rect 51262 6529 51274 6563
rect 51308 6529 51320 6563
rect 51262 6495 51320 6529
rect 51262 6461 51274 6495
rect 51308 6461 51320 6495
rect 51262 6427 51320 6461
rect 51262 6393 51274 6427
rect 51308 6393 51320 6427
rect 51262 6378 51320 6393
rect 51350 6563 51408 6578
rect 51350 6529 51362 6563
rect 51396 6529 51408 6563
rect 51588 6553 51600 6587
rect 51634 6553 51650 6587
rect 51588 6538 51650 6553
rect 51680 6723 51746 6738
rect 51680 6689 51696 6723
rect 51730 6689 51746 6723
rect 51680 6655 51746 6689
rect 51680 6621 51696 6655
rect 51730 6621 51746 6655
rect 51680 6587 51746 6621
rect 51680 6553 51696 6587
rect 51730 6553 51746 6587
rect 51680 6538 51746 6553
rect 51776 6723 51838 6738
rect 51776 6689 51792 6723
rect 51826 6689 51838 6723
rect 51776 6655 51838 6689
rect 51776 6621 51792 6655
rect 51826 6621 51838 6655
rect 51776 6587 51838 6621
rect 53476 6723 53538 6738
rect 53476 6689 53488 6723
rect 53522 6689 53538 6723
rect 51776 6553 51792 6587
rect 51826 6553 51838 6587
rect 51776 6538 51838 6553
rect 51908 6563 51966 6578
rect 51350 6495 51408 6529
rect 51350 6461 51362 6495
rect 51396 6461 51408 6495
rect 51350 6427 51408 6461
rect 51908 6529 51920 6563
rect 51954 6529 51966 6563
rect 51908 6495 51966 6529
rect 51908 6461 51920 6495
rect 51954 6461 51966 6495
rect 51350 6393 51362 6427
rect 51396 6393 51408 6427
rect 51350 6378 51408 6393
rect 51074 6363 51126 6375
rect 51908 6427 51966 6461
rect 51908 6393 51920 6427
rect 51954 6393 51966 6427
rect 51908 6378 51966 6393
rect 51996 6563 52054 6578
rect 51996 6529 52008 6563
rect 52042 6529 52054 6563
rect 51996 6495 52054 6529
rect 51996 6461 52008 6495
rect 52042 6461 52054 6495
rect 51996 6427 52054 6461
rect 51996 6393 52008 6427
rect 52042 6393 52054 6427
rect 51996 6378 52054 6393
rect 52188 6553 52240 6571
rect 52188 6519 52196 6553
rect 52230 6519 52240 6553
rect 52188 6485 52240 6519
rect 52188 6451 52196 6485
rect 52230 6451 52240 6485
rect 52188 6417 52240 6451
rect 52188 6383 52196 6417
rect 52230 6383 52240 6417
rect 52188 6371 52240 6383
rect 52270 6553 52322 6571
rect 52270 6519 52280 6553
rect 52314 6519 52322 6553
rect 53476 6655 53538 6689
rect 53476 6621 53488 6655
rect 53522 6621 53538 6655
rect 53476 6587 53538 6621
rect 53150 6563 53208 6578
rect 52880 6545 52932 6563
rect 52270 6485 52322 6519
rect 52270 6451 52280 6485
rect 52314 6451 52322 6485
rect 52270 6417 52322 6451
rect 52270 6383 52280 6417
rect 52314 6383 52322 6417
rect 52270 6371 52322 6383
rect 52487 6500 52539 6523
rect 52487 6466 52495 6500
rect 52529 6466 52539 6500
rect 52487 6419 52539 6466
rect 52487 6385 52495 6419
rect 52529 6385 52539 6419
rect 52487 6365 52539 6385
rect 52569 6487 52627 6523
rect 52569 6453 52581 6487
rect 52615 6453 52627 6487
rect 52569 6419 52627 6453
rect 52569 6385 52581 6419
rect 52615 6385 52627 6419
rect 52569 6365 52627 6385
rect 52657 6487 52709 6523
rect 52657 6453 52667 6487
rect 52701 6453 52709 6487
rect 52657 6419 52709 6453
rect 52657 6385 52667 6419
rect 52701 6385 52709 6419
rect 52657 6365 52709 6385
rect 52880 6511 52888 6545
rect 52922 6511 52932 6545
rect 52880 6477 52932 6511
rect 52880 6443 52888 6477
rect 52922 6443 52932 6477
rect 52880 6409 52932 6443
rect 52880 6375 52888 6409
rect 52922 6375 52932 6409
rect 52880 6363 52932 6375
rect 52962 6545 53014 6563
rect 52962 6511 52972 6545
rect 53006 6511 53014 6545
rect 52962 6477 53014 6511
rect 52962 6443 52972 6477
rect 53006 6443 53014 6477
rect 52962 6409 53014 6443
rect 52962 6375 52972 6409
rect 53006 6375 53014 6409
rect 53150 6529 53162 6563
rect 53196 6529 53208 6563
rect 53150 6495 53208 6529
rect 53150 6461 53162 6495
rect 53196 6461 53208 6495
rect 53150 6427 53208 6461
rect 53150 6393 53162 6427
rect 53196 6393 53208 6427
rect 53150 6378 53208 6393
rect 53238 6563 53296 6578
rect 53238 6529 53250 6563
rect 53284 6529 53296 6563
rect 53476 6553 53488 6587
rect 53522 6553 53538 6587
rect 53476 6538 53538 6553
rect 53568 6723 53634 6738
rect 53568 6689 53584 6723
rect 53618 6689 53634 6723
rect 53568 6655 53634 6689
rect 53568 6621 53584 6655
rect 53618 6621 53634 6655
rect 53568 6587 53634 6621
rect 53568 6553 53584 6587
rect 53618 6553 53634 6587
rect 53568 6538 53634 6553
rect 53664 6723 53726 6738
rect 53664 6689 53680 6723
rect 53714 6689 53726 6723
rect 53664 6655 53726 6689
rect 53664 6621 53680 6655
rect 53714 6621 53726 6655
rect 53664 6587 53726 6621
rect 55364 6723 55426 6738
rect 55364 6689 55376 6723
rect 55410 6689 55426 6723
rect 53664 6553 53680 6587
rect 53714 6553 53726 6587
rect 53664 6538 53726 6553
rect 53796 6563 53854 6578
rect 53238 6495 53296 6529
rect 53238 6461 53250 6495
rect 53284 6461 53296 6495
rect 53238 6427 53296 6461
rect 53796 6529 53808 6563
rect 53842 6529 53854 6563
rect 53796 6495 53854 6529
rect 53796 6461 53808 6495
rect 53842 6461 53854 6495
rect 53238 6393 53250 6427
rect 53284 6393 53296 6427
rect 53238 6378 53296 6393
rect 52962 6363 53014 6375
rect 53796 6427 53854 6461
rect 53796 6393 53808 6427
rect 53842 6393 53854 6427
rect 53796 6378 53854 6393
rect 53884 6563 53942 6578
rect 53884 6529 53896 6563
rect 53930 6529 53942 6563
rect 53884 6495 53942 6529
rect 53884 6461 53896 6495
rect 53930 6461 53942 6495
rect 53884 6427 53942 6461
rect 53884 6393 53896 6427
rect 53930 6393 53942 6427
rect 53884 6378 53942 6393
rect 54076 6553 54128 6571
rect 54076 6519 54084 6553
rect 54118 6519 54128 6553
rect 54076 6485 54128 6519
rect 54076 6451 54084 6485
rect 54118 6451 54128 6485
rect 54076 6417 54128 6451
rect 54076 6383 54084 6417
rect 54118 6383 54128 6417
rect 54076 6371 54128 6383
rect 54158 6553 54210 6571
rect 54158 6519 54168 6553
rect 54202 6519 54210 6553
rect 55364 6655 55426 6689
rect 55364 6621 55376 6655
rect 55410 6621 55426 6655
rect 55364 6587 55426 6621
rect 55038 6563 55096 6578
rect 54768 6545 54820 6563
rect 54158 6485 54210 6519
rect 54158 6451 54168 6485
rect 54202 6451 54210 6485
rect 54158 6417 54210 6451
rect 54158 6383 54168 6417
rect 54202 6383 54210 6417
rect 54158 6371 54210 6383
rect 54375 6500 54427 6523
rect 54375 6466 54383 6500
rect 54417 6466 54427 6500
rect 54375 6419 54427 6466
rect 54375 6385 54383 6419
rect 54417 6385 54427 6419
rect 54375 6365 54427 6385
rect 54457 6487 54515 6523
rect 54457 6453 54469 6487
rect 54503 6453 54515 6487
rect 54457 6419 54515 6453
rect 54457 6385 54469 6419
rect 54503 6385 54515 6419
rect 54457 6365 54515 6385
rect 54545 6487 54597 6523
rect 54545 6453 54555 6487
rect 54589 6453 54597 6487
rect 54545 6419 54597 6453
rect 54545 6385 54555 6419
rect 54589 6385 54597 6419
rect 54545 6365 54597 6385
rect 54768 6511 54776 6545
rect 54810 6511 54820 6545
rect 54768 6477 54820 6511
rect 54768 6443 54776 6477
rect 54810 6443 54820 6477
rect 54768 6409 54820 6443
rect 54768 6375 54776 6409
rect 54810 6375 54820 6409
rect 54768 6363 54820 6375
rect 54850 6545 54902 6563
rect 54850 6511 54860 6545
rect 54894 6511 54902 6545
rect 54850 6477 54902 6511
rect 54850 6443 54860 6477
rect 54894 6443 54902 6477
rect 54850 6409 54902 6443
rect 54850 6375 54860 6409
rect 54894 6375 54902 6409
rect 55038 6529 55050 6563
rect 55084 6529 55096 6563
rect 55038 6495 55096 6529
rect 55038 6461 55050 6495
rect 55084 6461 55096 6495
rect 55038 6427 55096 6461
rect 55038 6393 55050 6427
rect 55084 6393 55096 6427
rect 55038 6378 55096 6393
rect 55126 6563 55184 6578
rect 55126 6529 55138 6563
rect 55172 6529 55184 6563
rect 55364 6553 55376 6587
rect 55410 6553 55426 6587
rect 55364 6538 55426 6553
rect 55456 6723 55522 6738
rect 55456 6689 55472 6723
rect 55506 6689 55522 6723
rect 55456 6655 55522 6689
rect 55456 6621 55472 6655
rect 55506 6621 55522 6655
rect 55456 6587 55522 6621
rect 55456 6553 55472 6587
rect 55506 6553 55522 6587
rect 55456 6538 55522 6553
rect 55552 6723 55614 6738
rect 55552 6689 55568 6723
rect 55602 6689 55614 6723
rect 55552 6655 55614 6689
rect 55552 6621 55568 6655
rect 55602 6621 55614 6655
rect 55552 6587 55614 6621
rect 57252 6723 57314 6738
rect 57252 6689 57264 6723
rect 57298 6689 57314 6723
rect 55552 6553 55568 6587
rect 55602 6553 55614 6587
rect 55552 6538 55614 6553
rect 55684 6563 55742 6578
rect 55126 6495 55184 6529
rect 55126 6461 55138 6495
rect 55172 6461 55184 6495
rect 55126 6427 55184 6461
rect 55684 6529 55696 6563
rect 55730 6529 55742 6563
rect 55684 6495 55742 6529
rect 55684 6461 55696 6495
rect 55730 6461 55742 6495
rect 55126 6393 55138 6427
rect 55172 6393 55184 6427
rect 55126 6378 55184 6393
rect 54850 6363 54902 6375
rect 55684 6427 55742 6461
rect 55684 6393 55696 6427
rect 55730 6393 55742 6427
rect 55684 6378 55742 6393
rect 55772 6563 55830 6578
rect 55772 6529 55784 6563
rect 55818 6529 55830 6563
rect 55772 6495 55830 6529
rect 55772 6461 55784 6495
rect 55818 6461 55830 6495
rect 55772 6427 55830 6461
rect 55772 6393 55784 6427
rect 55818 6393 55830 6427
rect 55772 6378 55830 6393
rect 55964 6553 56016 6571
rect 55964 6519 55972 6553
rect 56006 6519 56016 6553
rect 55964 6485 56016 6519
rect 55964 6451 55972 6485
rect 56006 6451 56016 6485
rect 55964 6417 56016 6451
rect 55964 6383 55972 6417
rect 56006 6383 56016 6417
rect 55964 6371 56016 6383
rect 56046 6553 56098 6571
rect 56046 6519 56056 6553
rect 56090 6519 56098 6553
rect 57252 6655 57314 6689
rect 57252 6621 57264 6655
rect 57298 6621 57314 6655
rect 57252 6587 57314 6621
rect 56926 6563 56984 6578
rect 56656 6545 56708 6563
rect 56046 6485 56098 6519
rect 56046 6451 56056 6485
rect 56090 6451 56098 6485
rect 56046 6417 56098 6451
rect 56046 6383 56056 6417
rect 56090 6383 56098 6417
rect 56046 6371 56098 6383
rect 56263 6500 56315 6523
rect 56263 6466 56271 6500
rect 56305 6466 56315 6500
rect 56263 6419 56315 6466
rect 56263 6385 56271 6419
rect 56305 6385 56315 6419
rect 56263 6365 56315 6385
rect 56345 6487 56403 6523
rect 56345 6453 56357 6487
rect 56391 6453 56403 6487
rect 56345 6419 56403 6453
rect 56345 6385 56357 6419
rect 56391 6385 56403 6419
rect 56345 6365 56403 6385
rect 56433 6487 56485 6523
rect 56433 6453 56443 6487
rect 56477 6453 56485 6487
rect 56433 6419 56485 6453
rect 56433 6385 56443 6419
rect 56477 6385 56485 6419
rect 56433 6365 56485 6385
rect 56656 6511 56664 6545
rect 56698 6511 56708 6545
rect 56656 6477 56708 6511
rect 56656 6443 56664 6477
rect 56698 6443 56708 6477
rect 56656 6409 56708 6443
rect 56656 6375 56664 6409
rect 56698 6375 56708 6409
rect 56656 6363 56708 6375
rect 56738 6545 56790 6563
rect 56738 6511 56748 6545
rect 56782 6511 56790 6545
rect 56738 6477 56790 6511
rect 56738 6443 56748 6477
rect 56782 6443 56790 6477
rect 56738 6409 56790 6443
rect 56738 6375 56748 6409
rect 56782 6375 56790 6409
rect 56926 6529 56938 6563
rect 56972 6529 56984 6563
rect 56926 6495 56984 6529
rect 56926 6461 56938 6495
rect 56972 6461 56984 6495
rect 56926 6427 56984 6461
rect 56926 6393 56938 6427
rect 56972 6393 56984 6427
rect 56926 6378 56984 6393
rect 57014 6563 57072 6578
rect 57014 6529 57026 6563
rect 57060 6529 57072 6563
rect 57252 6553 57264 6587
rect 57298 6553 57314 6587
rect 57252 6538 57314 6553
rect 57344 6723 57410 6738
rect 57344 6689 57360 6723
rect 57394 6689 57410 6723
rect 57344 6655 57410 6689
rect 57344 6621 57360 6655
rect 57394 6621 57410 6655
rect 57344 6587 57410 6621
rect 57344 6553 57360 6587
rect 57394 6553 57410 6587
rect 57344 6538 57410 6553
rect 57440 6723 57502 6738
rect 57440 6689 57456 6723
rect 57490 6689 57502 6723
rect 57440 6655 57502 6689
rect 57440 6621 57456 6655
rect 57490 6621 57502 6655
rect 57440 6587 57502 6621
rect 59140 6723 59202 6738
rect 59140 6689 59152 6723
rect 59186 6689 59202 6723
rect 57440 6553 57456 6587
rect 57490 6553 57502 6587
rect 57440 6538 57502 6553
rect 57572 6563 57630 6578
rect 57014 6495 57072 6529
rect 57014 6461 57026 6495
rect 57060 6461 57072 6495
rect 57014 6427 57072 6461
rect 57572 6529 57584 6563
rect 57618 6529 57630 6563
rect 57572 6495 57630 6529
rect 57572 6461 57584 6495
rect 57618 6461 57630 6495
rect 57014 6393 57026 6427
rect 57060 6393 57072 6427
rect 57014 6378 57072 6393
rect 56738 6363 56790 6375
rect 57572 6427 57630 6461
rect 57572 6393 57584 6427
rect 57618 6393 57630 6427
rect 57572 6378 57630 6393
rect 57660 6563 57718 6578
rect 57660 6529 57672 6563
rect 57706 6529 57718 6563
rect 57660 6495 57718 6529
rect 57660 6461 57672 6495
rect 57706 6461 57718 6495
rect 57660 6427 57718 6461
rect 57660 6393 57672 6427
rect 57706 6393 57718 6427
rect 57660 6378 57718 6393
rect 57852 6553 57904 6571
rect 57852 6519 57860 6553
rect 57894 6519 57904 6553
rect 57852 6485 57904 6519
rect 57852 6451 57860 6485
rect 57894 6451 57904 6485
rect 57852 6417 57904 6451
rect 57852 6383 57860 6417
rect 57894 6383 57904 6417
rect 57852 6371 57904 6383
rect 57934 6553 57986 6571
rect 57934 6519 57944 6553
rect 57978 6519 57986 6553
rect 59140 6655 59202 6689
rect 59140 6621 59152 6655
rect 59186 6621 59202 6655
rect 59140 6587 59202 6621
rect 58814 6563 58872 6578
rect 58544 6545 58596 6563
rect 57934 6485 57986 6519
rect 57934 6451 57944 6485
rect 57978 6451 57986 6485
rect 57934 6417 57986 6451
rect 57934 6383 57944 6417
rect 57978 6383 57986 6417
rect 57934 6371 57986 6383
rect 58151 6500 58203 6523
rect 58151 6466 58159 6500
rect 58193 6466 58203 6500
rect 58151 6419 58203 6466
rect 58151 6385 58159 6419
rect 58193 6385 58203 6419
rect 58151 6365 58203 6385
rect 58233 6487 58291 6523
rect 58233 6453 58245 6487
rect 58279 6453 58291 6487
rect 58233 6419 58291 6453
rect 58233 6385 58245 6419
rect 58279 6385 58291 6419
rect 58233 6365 58291 6385
rect 58321 6487 58373 6523
rect 58321 6453 58331 6487
rect 58365 6453 58373 6487
rect 58321 6419 58373 6453
rect 58321 6385 58331 6419
rect 58365 6385 58373 6419
rect 58321 6365 58373 6385
rect 58544 6511 58552 6545
rect 58586 6511 58596 6545
rect 58544 6477 58596 6511
rect 58544 6443 58552 6477
rect 58586 6443 58596 6477
rect 58544 6409 58596 6443
rect 58544 6375 58552 6409
rect 58586 6375 58596 6409
rect 58544 6363 58596 6375
rect 58626 6545 58678 6563
rect 58626 6511 58636 6545
rect 58670 6511 58678 6545
rect 58626 6477 58678 6511
rect 58626 6443 58636 6477
rect 58670 6443 58678 6477
rect 58626 6409 58678 6443
rect 58626 6375 58636 6409
rect 58670 6375 58678 6409
rect 58814 6529 58826 6563
rect 58860 6529 58872 6563
rect 58814 6495 58872 6529
rect 58814 6461 58826 6495
rect 58860 6461 58872 6495
rect 58814 6427 58872 6461
rect 58814 6393 58826 6427
rect 58860 6393 58872 6427
rect 58814 6378 58872 6393
rect 58902 6563 58960 6578
rect 58902 6529 58914 6563
rect 58948 6529 58960 6563
rect 59140 6553 59152 6587
rect 59186 6553 59202 6587
rect 59140 6538 59202 6553
rect 59232 6723 59298 6738
rect 59232 6689 59248 6723
rect 59282 6689 59298 6723
rect 59232 6655 59298 6689
rect 59232 6621 59248 6655
rect 59282 6621 59298 6655
rect 59232 6587 59298 6621
rect 59232 6553 59248 6587
rect 59282 6553 59298 6587
rect 59232 6538 59298 6553
rect 59328 6723 59390 6738
rect 59328 6689 59344 6723
rect 59378 6689 59390 6723
rect 59328 6655 59390 6689
rect 59328 6621 59344 6655
rect 59378 6621 59390 6655
rect 59328 6587 59390 6621
rect 59328 6553 59344 6587
rect 59378 6553 59390 6587
rect 59328 6538 59390 6553
rect 59460 6563 59518 6578
rect 58902 6495 58960 6529
rect 58902 6461 58914 6495
rect 58948 6461 58960 6495
rect 58902 6427 58960 6461
rect 59460 6529 59472 6563
rect 59506 6529 59518 6563
rect 59460 6495 59518 6529
rect 59460 6461 59472 6495
rect 59506 6461 59518 6495
rect 58902 6393 58914 6427
rect 58948 6393 58960 6427
rect 58902 6378 58960 6393
rect 58626 6363 58678 6375
rect 59460 6427 59518 6461
rect 59460 6393 59472 6427
rect 59506 6393 59518 6427
rect 59460 6378 59518 6393
rect 59548 6563 59606 6578
rect 59548 6529 59560 6563
rect 59594 6529 59606 6563
rect 59548 6495 59606 6529
rect 59548 6461 59560 6495
rect 59594 6461 59606 6495
rect 59548 6427 59606 6461
rect 59548 6393 59560 6427
rect 59594 6393 59606 6427
rect 59548 6378 59606 6393
rect 59740 6553 59792 6571
rect 59740 6519 59748 6553
rect 59782 6519 59792 6553
rect 59740 6485 59792 6519
rect 59740 6451 59748 6485
rect 59782 6451 59792 6485
rect 59740 6417 59792 6451
rect 59740 6383 59748 6417
rect 59782 6383 59792 6417
rect 59740 6371 59792 6383
rect 59822 6553 59874 6571
rect 59822 6519 59832 6553
rect 59866 6519 59874 6553
rect 59822 6485 59874 6519
rect 59822 6451 59832 6485
rect 59866 6451 59874 6485
rect 59822 6417 59874 6451
rect 59822 6383 59832 6417
rect 59866 6383 59874 6417
rect 59822 6371 59874 6383
rect 622 5667 684 5682
rect 622 5633 634 5667
rect 668 5633 684 5667
rect 622 5599 684 5633
rect 622 5565 634 5599
rect 668 5565 684 5599
rect 622 5531 684 5565
rect 201 5499 253 5517
rect 201 5465 209 5499
rect 243 5465 253 5499
rect 201 5431 253 5465
rect 201 5397 209 5431
rect 243 5397 253 5431
rect 201 5363 253 5397
rect 201 5329 209 5363
rect 243 5329 253 5363
rect 201 5317 253 5329
rect 283 5317 325 5517
rect 355 5499 407 5517
rect 355 5465 365 5499
rect 399 5465 407 5499
rect 622 5497 634 5531
rect 668 5497 684 5531
rect 622 5482 684 5497
rect 714 5667 780 5682
rect 714 5633 730 5667
rect 764 5633 780 5667
rect 714 5599 780 5633
rect 714 5565 730 5599
rect 764 5565 780 5599
rect 714 5531 780 5565
rect 714 5497 730 5531
rect 764 5497 780 5531
rect 714 5482 780 5497
rect 810 5667 872 5682
rect 810 5633 826 5667
rect 860 5633 872 5667
rect 2510 5667 2572 5682
rect 810 5599 872 5633
rect 810 5565 826 5599
rect 860 5565 872 5599
rect 810 5531 872 5565
rect 810 5497 826 5531
rect 860 5497 872 5531
rect 2510 5633 2522 5667
rect 2556 5633 2572 5667
rect 2510 5599 2572 5633
rect 2510 5565 2522 5599
rect 2556 5565 2572 5599
rect 2510 5531 2572 5565
rect 810 5482 872 5497
rect 1015 5499 1067 5517
rect 355 5431 407 5465
rect 1015 5465 1023 5499
rect 1057 5465 1067 5499
rect 355 5397 365 5431
rect 399 5397 407 5431
rect 355 5363 407 5397
rect 1015 5431 1067 5465
rect 1015 5397 1023 5431
rect 1057 5397 1067 5431
rect 355 5329 365 5363
rect 399 5329 407 5363
rect 1015 5363 1067 5397
rect 355 5317 407 5329
rect 1015 5329 1023 5363
rect 1057 5329 1067 5363
rect 1015 5317 1067 5329
rect 1097 5317 1139 5517
rect 1169 5499 1221 5517
rect 1169 5465 1179 5499
rect 1213 5465 1221 5499
rect 1169 5431 1221 5465
rect 1169 5397 1179 5431
rect 1213 5397 1221 5431
rect 1169 5363 1221 5397
rect 1169 5329 1179 5363
rect 1213 5329 1221 5363
rect 1169 5317 1221 5329
rect 2089 5499 2141 5517
rect 2089 5465 2097 5499
rect 2131 5465 2141 5499
rect 2089 5431 2141 5465
rect 2089 5397 2097 5431
rect 2131 5397 2141 5431
rect 2089 5363 2141 5397
rect 2089 5329 2097 5363
rect 2131 5329 2141 5363
rect 2089 5317 2141 5329
rect 2171 5317 2213 5517
rect 2243 5499 2295 5517
rect 2243 5465 2253 5499
rect 2287 5465 2295 5499
rect 2510 5497 2522 5531
rect 2556 5497 2572 5531
rect 2510 5482 2572 5497
rect 2602 5667 2668 5682
rect 2602 5633 2618 5667
rect 2652 5633 2668 5667
rect 2602 5599 2668 5633
rect 2602 5565 2618 5599
rect 2652 5565 2668 5599
rect 2602 5531 2668 5565
rect 2602 5497 2618 5531
rect 2652 5497 2668 5531
rect 2602 5482 2668 5497
rect 2698 5667 2760 5682
rect 2698 5633 2714 5667
rect 2748 5633 2760 5667
rect 4398 5667 4460 5682
rect 2698 5599 2760 5633
rect 2698 5565 2714 5599
rect 2748 5565 2760 5599
rect 2698 5531 2760 5565
rect 2698 5497 2714 5531
rect 2748 5497 2760 5531
rect 4398 5633 4410 5667
rect 4444 5633 4460 5667
rect 4398 5599 4460 5633
rect 4398 5565 4410 5599
rect 4444 5565 4460 5599
rect 4398 5531 4460 5565
rect 2698 5482 2760 5497
rect 2903 5499 2955 5517
rect 2243 5431 2295 5465
rect 2903 5465 2911 5499
rect 2945 5465 2955 5499
rect 2243 5397 2253 5431
rect 2287 5397 2295 5431
rect 2243 5363 2295 5397
rect 2903 5431 2955 5465
rect 2903 5397 2911 5431
rect 2945 5397 2955 5431
rect 2243 5329 2253 5363
rect 2287 5329 2295 5363
rect 2903 5363 2955 5397
rect 2243 5317 2295 5329
rect 2903 5329 2911 5363
rect 2945 5329 2955 5363
rect 2903 5317 2955 5329
rect 2985 5317 3027 5517
rect 3057 5499 3109 5517
rect 3057 5465 3067 5499
rect 3101 5465 3109 5499
rect 3057 5431 3109 5465
rect 3057 5397 3067 5431
rect 3101 5397 3109 5431
rect 3057 5363 3109 5397
rect 3057 5329 3067 5363
rect 3101 5329 3109 5363
rect 3057 5317 3109 5329
rect 3977 5499 4029 5517
rect 3977 5465 3985 5499
rect 4019 5465 4029 5499
rect 3977 5431 4029 5465
rect 3977 5397 3985 5431
rect 4019 5397 4029 5431
rect 3977 5363 4029 5397
rect 3977 5329 3985 5363
rect 4019 5329 4029 5363
rect 3977 5317 4029 5329
rect 4059 5317 4101 5517
rect 4131 5499 4183 5517
rect 4131 5465 4141 5499
rect 4175 5465 4183 5499
rect 4398 5497 4410 5531
rect 4444 5497 4460 5531
rect 4398 5482 4460 5497
rect 4490 5667 4556 5682
rect 4490 5633 4506 5667
rect 4540 5633 4556 5667
rect 4490 5599 4556 5633
rect 4490 5565 4506 5599
rect 4540 5565 4556 5599
rect 4490 5531 4556 5565
rect 4490 5497 4506 5531
rect 4540 5497 4556 5531
rect 4490 5482 4556 5497
rect 4586 5667 4648 5682
rect 4586 5633 4602 5667
rect 4636 5633 4648 5667
rect 6286 5667 6348 5682
rect 4586 5599 4648 5633
rect 4586 5565 4602 5599
rect 4636 5565 4648 5599
rect 4586 5531 4648 5565
rect 4586 5497 4602 5531
rect 4636 5497 4648 5531
rect 6286 5633 6298 5667
rect 6332 5633 6348 5667
rect 6286 5599 6348 5633
rect 6286 5565 6298 5599
rect 6332 5565 6348 5599
rect 6286 5531 6348 5565
rect 4586 5482 4648 5497
rect 4791 5499 4843 5517
rect 4131 5431 4183 5465
rect 4791 5465 4799 5499
rect 4833 5465 4843 5499
rect 4131 5397 4141 5431
rect 4175 5397 4183 5431
rect 4131 5363 4183 5397
rect 4791 5431 4843 5465
rect 4791 5397 4799 5431
rect 4833 5397 4843 5431
rect 4131 5329 4141 5363
rect 4175 5329 4183 5363
rect 4791 5363 4843 5397
rect 4131 5317 4183 5329
rect 4791 5329 4799 5363
rect 4833 5329 4843 5363
rect 4791 5317 4843 5329
rect 4873 5317 4915 5517
rect 4945 5499 4997 5517
rect 4945 5465 4955 5499
rect 4989 5465 4997 5499
rect 4945 5431 4997 5465
rect 4945 5397 4955 5431
rect 4989 5397 4997 5431
rect 4945 5363 4997 5397
rect 4945 5329 4955 5363
rect 4989 5329 4997 5363
rect 4945 5317 4997 5329
rect 5865 5499 5917 5517
rect 5865 5465 5873 5499
rect 5907 5465 5917 5499
rect 5865 5431 5917 5465
rect 5865 5397 5873 5431
rect 5907 5397 5917 5431
rect 5865 5363 5917 5397
rect 5865 5329 5873 5363
rect 5907 5329 5917 5363
rect 5865 5317 5917 5329
rect 5947 5317 5989 5517
rect 6019 5499 6071 5517
rect 6019 5465 6029 5499
rect 6063 5465 6071 5499
rect 6286 5497 6298 5531
rect 6332 5497 6348 5531
rect 6286 5482 6348 5497
rect 6378 5667 6444 5682
rect 6378 5633 6394 5667
rect 6428 5633 6444 5667
rect 6378 5599 6444 5633
rect 6378 5565 6394 5599
rect 6428 5565 6444 5599
rect 6378 5531 6444 5565
rect 6378 5497 6394 5531
rect 6428 5497 6444 5531
rect 6378 5482 6444 5497
rect 6474 5667 6536 5682
rect 6474 5633 6490 5667
rect 6524 5633 6536 5667
rect 8174 5667 8236 5682
rect 6474 5599 6536 5633
rect 6474 5565 6490 5599
rect 6524 5565 6536 5599
rect 6474 5531 6536 5565
rect 6474 5497 6490 5531
rect 6524 5497 6536 5531
rect 8174 5633 8186 5667
rect 8220 5633 8236 5667
rect 8174 5599 8236 5633
rect 8174 5565 8186 5599
rect 8220 5565 8236 5599
rect 8174 5531 8236 5565
rect 6474 5482 6536 5497
rect 6679 5499 6731 5517
rect 6019 5431 6071 5465
rect 6679 5465 6687 5499
rect 6721 5465 6731 5499
rect 6019 5397 6029 5431
rect 6063 5397 6071 5431
rect 6019 5363 6071 5397
rect 6679 5431 6731 5465
rect 6679 5397 6687 5431
rect 6721 5397 6731 5431
rect 6019 5329 6029 5363
rect 6063 5329 6071 5363
rect 6679 5363 6731 5397
rect 6019 5317 6071 5329
rect 6679 5329 6687 5363
rect 6721 5329 6731 5363
rect 6679 5317 6731 5329
rect 6761 5317 6803 5517
rect 6833 5499 6885 5517
rect 6833 5465 6843 5499
rect 6877 5465 6885 5499
rect 6833 5431 6885 5465
rect 6833 5397 6843 5431
rect 6877 5397 6885 5431
rect 6833 5363 6885 5397
rect 6833 5329 6843 5363
rect 6877 5329 6885 5363
rect 6833 5317 6885 5329
rect 7753 5499 7805 5517
rect 7753 5465 7761 5499
rect 7795 5465 7805 5499
rect 7753 5431 7805 5465
rect 7753 5397 7761 5431
rect 7795 5397 7805 5431
rect 7753 5363 7805 5397
rect 7753 5329 7761 5363
rect 7795 5329 7805 5363
rect 7753 5317 7805 5329
rect 7835 5317 7877 5517
rect 7907 5499 7959 5517
rect 7907 5465 7917 5499
rect 7951 5465 7959 5499
rect 8174 5497 8186 5531
rect 8220 5497 8236 5531
rect 8174 5482 8236 5497
rect 8266 5667 8332 5682
rect 8266 5633 8282 5667
rect 8316 5633 8332 5667
rect 8266 5599 8332 5633
rect 8266 5565 8282 5599
rect 8316 5565 8332 5599
rect 8266 5531 8332 5565
rect 8266 5497 8282 5531
rect 8316 5497 8332 5531
rect 8266 5482 8332 5497
rect 8362 5667 8424 5682
rect 8362 5633 8378 5667
rect 8412 5633 8424 5667
rect 10062 5667 10124 5682
rect 8362 5599 8424 5633
rect 8362 5565 8378 5599
rect 8412 5565 8424 5599
rect 8362 5531 8424 5565
rect 8362 5497 8378 5531
rect 8412 5497 8424 5531
rect 10062 5633 10074 5667
rect 10108 5633 10124 5667
rect 10062 5599 10124 5633
rect 10062 5565 10074 5599
rect 10108 5565 10124 5599
rect 10062 5531 10124 5565
rect 8362 5482 8424 5497
rect 8567 5499 8619 5517
rect 7907 5431 7959 5465
rect 8567 5465 8575 5499
rect 8609 5465 8619 5499
rect 7907 5397 7917 5431
rect 7951 5397 7959 5431
rect 7907 5363 7959 5397
rect 8567 5431 8619 5465
rect 8567 5397 8575 5431
rect 8609 5397 8619 5431
rect 7907 5329 7917 5363
rect 7951 5329 7959 5363
rect 8567 5363 8619 5397
rect 7907 5317 7959 5329
rect 8567 5329 8575 5363
rect 8609 5329 8619 5363
rect 8567 5317 8619 5329
rect 8649 5317 8691 5517
rect 8721 5499 8773 5517
rect 8721 5465 8731 5499
rect 8765 5465 8773 5499
rect 8721 5431 8773 5465
rect 8721 5397 8731 5431
rect 8765 5397 8773 5431
rect 8721 5363 8773 5397
rect 8721 5329 8731 5363
rect 8765 5329 8773 5363
rect 8721 5317 8773 5329
rect 9641 5499 9693 5517
rect 9641 5465 9649 5499
rect 9683 5465 9693 5499
rect 9641 5431 9693 5465
rect 9641 5397 9649 5431
rect 9683 5397 9693 5431
rect 9641 5363 9693 5397
rect 9641 5329 9649 5363
rect 9683 5329 9693 5363
rect 9641 5317 9693 5329
rect 9723 5317 9765 5517
rect 9795 5499 9847 5517
rect 9795 5465 9805 5499
rect 9839 5465 9847 5499
rect 10062 5497 10074 5531
rect 10108 5497 10124 5531
rect 10062 5482 10124 5497
rect 10154 5667 10220 5682
rect 10154 5633 10170 5667
rect 10204 5633 10220 5667
rect 10154 5599 10220 5633
rect 10154 5565 10170 5599
rect 10204 5565 10220 5599
rect 10154 5531 10220 5565
rect 10154 5497 10170 5531
rect 10204 5497 10220 5531
rect 10154 5482 10220 5497
rect 10250 5667 10312 5682
rect 10250 5633 10266 5667
rect 10300 5633 10312 5667
rect 11950 5667 12012 5682
rect 10250 5599 10312 5633
rect 10250 5565 10266 5599
rect 10300 5565 10312 5599
rect 10250 5531 10312 5565
rect 10250 5497 10266 5531
rect 10300 5497 10312 5531
rect 11950 5633 11962 5667
rect 11996 5633 12012 5667
rect 11950 5599 12012 5633
rect 11950 5565 11962 5599
rect 11996 5565 12012 5599
rect 11950 5531 12012 5565
rect 10250 5482 10312 5497
rect 10455 5499 10507 5517
rect 9795 5431 9847 5465
rect 10455 5465 10463 5499
rect 10497 5465 10507 5499
rect 9795 5397 9805 5431
rect 9839 5397 9847 5431
rect 9795 5363 9847 5397
rect 10455 5431 10507 5465
rect 10455 5397 10463 5431
rect 10497 5397 10507 5431
rect 9795 5329 9805 5363
rect 9839 5329 9847 5363
rect 10455 5363 10507 5397
rect 9795 5317 9847 5329
rect 10455 5329 10463 5363
rect 10497 5329 10507 5363
rect 10455 5317 10507 5329
rect 10537 5317 10579 5517
rect 10609 5499 10661 5517
rect 10609 5465 10619 5499
rect 10653 5465 10661 5499
rect 10609 5431 10661 5465
rect 10609 5397 10619 5431
rect 10653 5397 10661 5431
rect 10609 5363 10661 5397
rect 10609 5329 10619 5363
rect 10653 5329 10661 5363
rect 10609 5317 10661 5329
rect 11529 5499 11581 5517
rect 11529 5465 11537 5499
rect 11571 5465 11581 5499
rect 11529 5431 11581 5465
rect 11529 5397 11537 5431
rect 11571 5397 11581 5431
rect 11529 5363 11581 5397
rect 11529 5329 11537 5363
rect 11571 5329 11581 5363
rect 11529 5317 11581 5329
rect 11611 5317 11653 5517
rect 11683 5499 11735 5517
rect 11683 5465 11693 5499
rect 11727 5465 11735 5499
rect 11950 5497 11962 5531
rect 11996 5497 12012 5531
rect 11950 5482 12012 5497
rect 12042 5667 12108 5682
rect 12042 5633 12058 5667
rect 12092 5633 12108 5667
rect 12042 5599 12108 5633
rect 12042 5565 12058 5599
rect 12092 5565 12108 5599
rect 12042 5531 12108 5565
rect 12042 5497 12058 5531
rect 12092 5497 12108 5531
rect 12042 5482 12108 5497
rect 12138 5667 12200 5682
rect 12138 5633 12154 5667
rect 12188 5633 12200 5667
rect 13838 5667 13900 5682
rect 12138 5599 12200 5633
rect 12138 5565 12154 5599
rect 12188 5565 12200 5599
rect 12138 5531 12200 5565
rect 12138 5497 12154 5531
rect 12188 5497 12200 5531
rect 13838 5633 13850 5667
rect 13884 5633 13900 5667
rect 13838 5599 13900 5633
rect 13838 5565 13850 5599
rect 13884 5565 13900 5599
rect 13838 5531 13900 5565
rect 12138 5482 12200 5497
rect 12343 5499 12395 5517
rect 11683 5431 11735 5465
rect 12343 5465 12351 5499
rect 12385 5465 12395 5499
rect 11683 5397 11693 5431
rect 11727 5397 11735 5431
rect 11683 5363 11735 5397
rect 12343 5431 12395 5465
rect 12343 5397 12351 5431
rect 12385 5397 12395 5431
rect 11683 5329 11693 5363
rect 11727 5329 11735 5363
rect 12343 5363 12395 5397
rect 11683 5317 11735 5329
rect 12343 5329 12351 5363
rect 12385 5329 12395 5363
rect 12343 5317 12395 5329
rect 12425 5317 12467 5517
rect 12497 5499 12549 5517
rect 12497 5465 12507 5499
rect 12541 5465 12549 5499
rect 12497 5431 12549 5465
rect 12497 5397 12507 5431
rect 12541 5397 12549 5431
rect 12497 5363 12549 5397
rect 12497 5329 12507 5363
rect 12541 5329 12549 5363
rect 12497 5317 12549 5329
rect 13417 5499 13469 5517
rect 13417 5465 13425 5499
rect 13459 5465 13469 5499
rect 13417 5431 13469 5465
rect 13417 5397 13425 5431
rect 13459 5397 13469 5431
rect 13417 5363 13469 5397
rect 13417 5329 13425 5363
rect 13459 5329 13469 5363
rect 13417 5317 13469 5329
rect 13499 5317 13541 5517
rect 13571 5499 13623 5517
rect 13571 5465 13581 5499
rect 13615 5465 13623 5499
rect 13838 5497 13850 5531
rect 13884 5497 13900 5531
rect 13838 5482 13900 5497
rect 13930 5667 13996 5682
rect 13930 5633 13946 5667
rect 13980 5633 13996 5667
rect 13930 5599 13996 5633
rect 13930 5565 13946 5599
rect 13980 5565 13996 5599
rect 13930 5531 13996 5565
rect 13930 5497 13946 5531
rect 13980 5497 13996 5531
rect 13930 5482 13996 5497
rect 14026 5667 14088 5682
rect 14026 5633 14042 5667
rect 14076 5633 14088 5667
rect 15720 5667 15782 5682
rect 14026 5599 14088 5633
rect 14026 5565 14042 5599
rect 14076 5565 14088 5599
rect 14026 5531 14088 5565
rect 14026 5497 14042 5531
rect 14076 5497 14088 5531
rect 15720 5633 15732 5667
rect 15766 5633 15782 5667
rect 15720 5599 15782 5633
rect 15720 5565 15732 5599
rect 15766 5565 15782 5599
rect 15720 5531 15782 5565
rect 14026 5482 14088 5497
rect 14231 5499 14283 5517
rect 13571 5431 13623 5465
rect 14231 5465 14239 5499
rect 14273 5465 14283 5499
rect 13571 5397 13581 5431
rect 13615 5397 13623 5431
rect 13571 5363 13623 5397
rect 14231 5431 14283 5465
rect 14231 5397 14239 5431
rect 14273 5397 14283 5431
rect 13571 5329 13581 5363
rect 13615 5329 13623 5363
rect 14231 5363 14283 5397
rect 13571 5317 13623 5329
rect 14231 5329 14239 5363
rect 14273 5329 14283 5363
rect 14231 5317 14283 5329
rect 14313 5317 14355 5517
rect 14385 5499 14437 5517
rect 14385 5465 14395 5499
rect 14429 5465 14437 5499
rect 14385 5431 14437 5465
rect 14385 5397 14395 5431
rect 14429 5397 14437 5431
rect 14385 5363 14437 5397
rect 14385 5329 14395 5363
rect 14429 5329 14437 5363
rect 14385 5317 14437 5329
rect 15299 5499 15351 5517
rect 15299 5465 15307 5499
rect 15341 5465 15351 5499
rect 15299 5431 15351 5465
rect 15299 5397 15307 5431
rect 15341 5397 15351 5431
rect 15299 5363 15351 5397
rect 15299 5329 15307 5363
rect 15341 5329 15351 5363
rect 15299 5317 15351 5329
rect 15381 5317 15423 5517
rect 15453 5499 15505 5517
rect 15453 5465 15463 5499
rect 15497 5465 15505 5499
rect 15720 5497 15732 5531
rect 15766 5497 15782 5531
rect 15720 5482 15782 5497
rect 15812 5667 15878 5682
rect 15812 5633 15828 5667
rect 15862 5633 15878 5667
rect 15812 5599 15878 5633
rect 15812 5565 15828 5599
rect 15862 5565 15878 5599
rect 15812 5531 15878 5565
rect 15812 5497 15828 5531
rect 15862 5497 15878 5531
rect 15812 5482 15878 5497
rect 15908 5667 15970 5682
rect 15908 5633 15924 5667
rect 15958 5633 15970 5667
rect 17608 5667 17670 5682
rect 15908 5599 15970 5633
rect 15908 5565 15924 5599
rect 15958 5565 15970 5599
rect 15908 5531 15970 5565
rect 15908 5497 15924 5531
rect 15958 5497 15970 5531
rect 17608 5633 17620 5667
rect 17654 5633 17670 5667
rect 17608 5599 17670 5633
rect 17608 5565 17620 5599
rect 17654 5565 17670 5599
rect 17608 5531 17670 5565
rect 15908 5482 15970 5497
rect 16113 5499 16165 5517
rect 15453 5431 15505 5465
rect 16113 5465 16121 5499
rect 16155 5465 16165 5499
rect 15453 5397 15463 5431
rect 15497 5397 15505 5431
rect 15453 5363 15505 5397
rect 16113 5431 16165 5465
rect 16113 5397 16121 5431
rect 16155 5397 16165 5431
rect 15453 5329 15463 5363
rect 15497 5329 15505 5363
rect 16113 5363 16165 5397
rect 15453 5317 15505 5329
rect 16113 5329 16121 5363
rect 16155 5329 16165 5363
rect 16113 5317 16165 5329
rect 16195 5317 16237 5517
rect 16267 5499 16319 5517
rect 16267 5465 16277 5499
rect 16311 5465 16319 5499
rect 16267 5431 16319 5465
rect 16267 5397 16277 5431
rect 16311 5397 16319 5431
rect 16267 5363 16319 5397
rect 16267 5329 16277 5363
rect 16311 5329 16319 5363
rect 16267 5317 16319 5329
rect 17187 5499 17239 5517
rect 17187 5465 17195 5499
rect 17229 5465 17239 5499
rect 17187 5431 17239 5465
rect 17187 5397 17195 5431
rect 17229 5397 17239 5431
rect 17187 5363 17239 5397
rect 17187 5329 17195 5363
rect 17229 5329 17239 5363
rect 17187 5317 17239 5329
rect 17269 5317 17311 5517
rect 17341 5499 17393 5517
rect 17341 5465 17351 5499
rect 17385 5465 17393 5499
rect 17608 5497 17620 5531
rect 17654 5497 17670 5531
rect 17608 5482 17670 5497
rect 17700 5667 17766 5682
rect 17700 5633 17716 5667
rect 17750 5633 17766 5667
rect 17700 5599 17766 5633
rect 17700 5565 17716 5599
rect 17750 5565 17766 5599
rect 17700 5531 17766 5565
rect 17700 5497 17716 5531
rect 17750 5497 17766 5531
rect 17700 5482 17766 5497
rect 17796 5667 17858 5682
rect 17796 5633 17812 5667
rect 17846 5633 17858 5667
rect 19496 5667 19558 5682
rect 17796 5599 17858 5633
rect 17796 5565 17812 5599
rect 17846 5565 17858 5599
rect 17796 5531 17858 5565
rect 17796 5497 17812 5531
rect 17846 5497 17858 5531
rect 19496 5633 19508 5667
rect 19542 5633 19558 5667
rect 19496 5599 19558 5633
rect 19496 5565 19508 5599
rect 19542 5565 19558 5599
rect 19496 5531 19558 5565
rect 17796 5482 17858 5497
rect 18001 5499 18053 5517
rect 17341 5431 17393 5465
rect 18001 5465 18009 5499
rect 18043 5465 18053 5499
rect 17341 5397 17351 5431
rect 17385 5397 17393 5431
rect 17341 5363 17393 5397
rect 18001 5431 18053 5465
rect 18001 5397 18009 5431
rect 18043 5397 18053 5431
rect 17341 5329 17351 5363
rect 17385 5329 17393 5363
rect 18001 5363 18053 5397
rect 17341 5317 17393 5329
rect 18001 5329 18009 5363
rect 18043 5329 18053 5363
rect 18001 5317 18053 5329
rect 18083 5317 18125 5517
rect 18155 5499 18207 5517
rect 18155 5465 18165 5499
rect 18199 5465 18207 5499
rect 18155 5431 18207 5465
rect 18155 5397 18165 5431
rect 18199 5397 18207 5431
rect 18155 5363 18207 5397
rect 18155 5329 18165 5363
rect 18199 5329 18207 5363
rect 18155 5317 18207 5329
rect 19075 5499 19127 5517
rect 19075 5465 19083 5499
rect 19117 5465 19127 5499
rect 19075 5431 19127 5465
rect 19075 5397 19083 5431
rect 19117 5397 19127 5431
rect 19075 5363 19127 5397
rect 19075 5329 19083 5363
rect 19117 5329 19127 5363
rect 19075 5317 19127 5329
rect 19157 5317 19199 5517
rect 19229 5499 19281 5517
rect 19229 5465 19239 5499
rect 19273 5465 19281 5499
rect 19496 5497 19508 5531
rect 19542 5497 19558 5531
rect 19496 5482 19558 5497
rect 19588 5667 19654 5682
rect 19588 5633 19604 5667
rect 19638 5633 19654 5667
rect 19588 5599 19654 5633
rect 19588 5565 19604 5599
rect 19638 5565 19654 5599
rect 19588 5531 19654 5565
rect 19588 5497 19604 5531
rect 19638 5497 19654 5531
rect 19588 5482 19654 5497
rect 19684 5667 19746 5682
rect 19684 5633 19700 5667
rect 19734 5633 19746 5667
rect 21384 5667 21446 5682
rect 19684 5599 19746 5633
rect 19684 5565 19700 5599
rect 19734 5565 19746 5599
rect 19684 5531 19746 5565
rect 19684 5497 19700 5531
rect 19734 5497 19746 5531
rect 21384 5633 21396 5667
rect 21430 5633 21446 5667
rect 21384 5599 21446 5633
rect 21384 5565 21396 5599
rect 21430 5565 21446 5599
rect 21384 5531 21446 5565
rect 19684 5482 19746 5497
rect 19889 5499 19941 5517
rect 19229 5431 19281 5465
rect 19889 5465 19897 5499
rect 19931 5465 19941 5499
rect 19229 5397 19239 5431
rect 19273 5397 19281 5431
rect 19229 5363 19281 5397
rect 19889 5431 19941 5465
rect 19889 5397 19897 5431
rect 19931 5397 19941 5431
rect 19229 5329 19239 5363
rect 19273 5329 19281 5363
rect 19889 5363 19941 5397
rect 19229 5317 19281 5329
rect 19889 5329 19897 5363
rect 19931 5329 19941 5363
rect 19889 5317 19941 5329
rect 19971 5317 20013 5517
rect 20043 5499 20095 5517
rect 20043 5465 20053 5499
rect 20087 5465 20095 5499
rect 20043 5431 20095 5465
rect 20043 5397 20053 5431
rect 20087 5397 20095 5431
rect 20043 5363 20095 5397
rect 20043 5329 20053 5363
rect 20087 5329 20095 5363
rect 20043 5317 20095 5329
rect 20963 5499 21015 5517
rect 20963 5465 20971 5499
rect 21005 5465 21015 5499
rect 20963 5431 21015 5465
rect 20963 5397 20971 5431
rect 21005 5397 21015 5431
rect 20963 5363 21015 5397
rect 20963 5329 20971 5363
rect 21005 5329 21015 5363
rect 20963 5317 21015 5329
rect 21045 5317 21087 5517
rect 21117 5499 21169 5517
rect 21117 5465 21127 5499
rect 21161 5465 21169 5499
rect 21384 5497 21396 5531
rect 21430 5497 21446 5531
rect 21384 5482 21446 5497
rect 21476 5667 21542 5682
rect 21476 5633 21492 5667
rect 21526 5633 21542 5667
rect 21476 5599 21542 5633
rect 21476 5565 21492 5599
rect 21526 5565 21542 5599
rect 21476 5531 21542 5565
rect 21476 5497 21492 5531
rect 21526 5497 21542 5531
rect 21476 5482 21542 5497
rect 21572 5667 21634 5682
rect 21572 5633 21588 5667
rect 21622 5633 21634 5667
rect 23272 5667 23334 5682
rect 21572 5599 21634 5633
rect 21572 5565 21588 5599
rect 21622 5565 21634 5599
rect 21572 5531 21634 5565
rect 21572 5497 21588 5531
rect 21622 5497 21634 5531
rect 23272 5633 23284 5667
rect 23318 5633 23334 5667
rect 23272 5599 23334 5633
rect 23272 5565 23284 5599
rect 23318 5565 23334 5599
rect 23272 5531 23334 5565
rect 21572 5482 21634 5497
rect 21777 5499 21829 5517
rect 21117 5431 21169 5465
rect 21777 5465 21785 5499
rect 21819 5465 21829 5499
rect 21117 5397 21127 5431
rect 21161 5397 21169 5431
rect 21117 5363 21169 5397
rect 21777 5431 21829 5465
rect 21777 5397 21785 5431
rect 21819 5397 21829 5431
rect 21117 5329 21127 5363
rect 21161 5329 21169 5363
rect 21777 5363 21829 5397
rect 21117 5317 21169 5329
rect 21777 5329 21785 5363
rect 21819 5329 21829 5363
rect 21777 5317 21829 5329
rect 21859 5317 21901 5517
rect 21931 5499 21983 5517
rect 21931 5465 21941 5499
rect 21975 5465 21983 5499
rect 21931 5431 21983 5465
rect 21931 5397 21941 5431
rect 21975 5397 21983 5431
rect 21931 5363 21983 5397
rect 21931 5329 21941 5363
rect 21975 5329 21983 5363
rect 21931 5317 21983 5329
rect 22851 5499 22903 5517
rect 22851 5465 22859 5499
rect 22893 5465 22903 5499
rect 22851 5431 22903 5465
rect 22851 5397 22859 5431
rect 22893 5397 22903 5431
rect 22851 5363 22903 5397
rect 22851 5329 22859 5363
rect 22893 5329 22903 5363
rect 22851 5317 22903 5329
rect 22933 5317 22975 5517
rect 23005 5499 23057 5517
rect 23005 5465 23015 5499
rect 23049 5465 23057 5499
rect 23272 5497 23284 5531
rect 23318 5497 23334 5531
rect 23272 5482 23334 5497
rect 23364 5667 23430 5682
rect 23364 5633 23380 5667
rect 23414 5633 23430 5667
rect 23364 5599 23430 5633
rect 23364 5565 23380 5599
rect 23414 5565 23430 5599
rect 23364 5531 23430 5565
rect 23364 5497 23380 5531
rect 23414 5497 23430 5531
rect 23364 5482 23430 5497
rect 23460 5667 23522 5682
rect 23460 5633 23476 5667
rect 23510 5633 23522 5667
rect 25160 5667 25222 5682
rect 23460 5599 23522 5633
rect 23460 5565 23476 5599
rect 23510 5565 23522 5599
rect 23460 5531 23522 5565
rect 23460 5497 23476 5531
rect 23510 5497 23522 5531
rect 25160 5633 25172 5667
rect 25206 5633 25222 5667
rect 25160 5599 25222 5633
rect 25160 5565 25172 5599
rect 25206 5565 25222 5599
rect 25160 5531 25222 5565
rect 23460 5482 23522 5497
rect 23665 5499 23717 5517
rect 23005 5431 23057 5465
rect 23665 5465 23673 5499
rect 23707 5465 23717 5499
rect 23005 5397 23015 5431
rect 23049 5397 23057 5431
rect 23005 5363 23057 5397
rect 23665 5431 23717 5465
rect 23665 5397 23673 5431
rect 23707 5397 23717 5431
rect 23005 5329 23015 5363
rect 23049 5329 23057 5363
rect 23665 5363 23717 5397
rect 23005 5317 23057 5329
rect 23665 5329 23673 5363
rect 23707 5329 23717 5363
rect 23665 5317 23717 5329
rect 23747 5317 23789 5517
rect 23819 5499 23871 5517
rect 23819 5465 23829 5499
rect 23863 5465 23871 5499
rect 23819 5431 23871 5465
rect 23819 5397 23829 5431
rect 23863 5397 23871 5431
rect 23819 5363 23871 5397
rect 23819 5329 23829 5363
rect 23863 5329 23871 5363
rect 23819 5317 23871 5329
rect 24739 5499 24791 5517
rect 24739 5465 24747 5499
rect 24781 5465 24791 5499
rect 24739 5431 24791 5465
rect 24739 5397 24747 5431
rect 24781 5397 24791 5431
rect 24739 5363 24791 5397
rect 24739 5329 24747 5363
rect 24781 5329 24791 5363
rect 24739 5317 24791 5329
rect 24821 5317 24863 5517
rect 24893 5499 24945 5517
rect 24893 5465 24903 5499
rect 24937 5465 24945 5499
rect 25160 5497 25172 5531
rect 25206 5497 25222 5531
rect 25160 5482 25222 5497
rect 25252 5667 25318 5682
rect 25252 5633 25268 5667
rect 25302 5633 25318 5667
rect 25252 5599 25318 5633
rect 25252 5565 25268 5599
rect 25302 5565 25318 5599
rect 25252 5531 25318 5565
rect 25252 5497 25268 5531
rect 25302 5497 25318 5531
rect 25252 5482 25318 5497
rect 25348 5667 25410 5682
rect 25348 5633 25364 5667
rect 25398 5633 25410 5667
rect 27048 5667 27110 5682
rect 25348 5599 25410 5633
rect 25348 5565 25364 5599
rect 25398 5565 25410 5599
rect 25348 5531 25410 5565
rect 25348 5497 25364 5531
rect 25398 5497 25410 5531
rect 27048 5633 27060 5667
rect 27094 5633 27110 5667
rect 27048 5599 27110 5633
rect 27048 5565 27060 5599
rect 27094 5565 27110 5599
rect 27048 5531 27110 5565
rect 25348 5482 25410 5497
rect 25553 5499 25605 5517
rect 24893 5431 24945 5465
rect 25553 5465 25561 5499
rect 25595 5465 25605 5499
rect 24893 5397 24903 5431
rect 24937 5397 24945 5431
rect 24893 5363 24945 5397
rect 25553 5431 25605 5465
rect 25553 5397 25561 5431
rect 25595 5397 25605 5431
rect 24893 5329 24903 5363
rect 24937 5329 24945 5363
rect 25553 5363 25605 5397
rect 24893 5317 24945 5329
rect 25553 5329 25561 5363
rect 25595 5329 25605 5363
rect 25553 5317 25605 5329
rect 25635 5317 25677 5517
rect 25707 5499 25759 5517
rect 25707 5465 25717 5499
rect 25751 5465 25759 5499
rect 25707 5431 25759 5465
rect 25707 5397 25717 5431
rect 25751 5397 25759 5431
rect 25707 5363 25759 5397
rect 25707 5329 25717 5363
rect 25751 5329 25759 5363
rect 25707 5317 25759 5329
rect 26627 5499 26679 5517
rect 26627 5465 26635 5499
rect 26669 5465 26679 5499
rect 26627 5431 26679 5465
rect 26627 5397 26635 5431
rect 26669 5397 26679 5431
rect 26627 5363 26679 5397
rect 26627 5329 26635 5363
rect 26669 5329 26679 5363
rect 26627 5317 26679 5329
rect 26709 5317 26751 5517
rect 26781 5499 26833 5517
rect 26781 5465 26791 5499
rect 26825 5465 26833 5499
rect 27048 5497 27060 5531
rect 27094 5497 27110 5531
rect 27048 5482 27110 5497
rect 27140 5667 27206 5682
rect 27140 5633 27156 5667
rect 27190 5633 27206 5667
rect 27140 5599 27206 5633
rect 27140 5565 27156 5599
rect 27190 5565 27206 5599
rect 27140 5531 27206 5565
rect 27140 5497 27156 5531
rect 27190 5497 27206 5531
rect 27140 5482 27206 5497
rect 27236 5667 27298 5682
rect 27236 5633 27252 5667
rect 27286 5633 27298 5667
rect 28936 5667 28998 5682
rect 27236 5599 27298 5633
rect 27236 5565 27252 5599
rect 27286 5565 27298 5599
rect 27236 5531 27298 5565
rect 27236 5497 27252 5531
rect 27286 5497 27298 5531
rect 28936 5633 28948 5667
rect 28982 5633 28998 5667
rect 28936 5599 28998 5633
rect 28936 5565 28948 5599
rect 28982 5565 28998 5599
rect 28936 5531 28998 5565
rect 27236 5482 27298 5497
rect 27441 5499 27493 5517
rect 26781 5431 26833 5465
rect 27441 5465 27449 5499
rect 27483 5465 27493 5499
rect 26781 5397 26791 5431
rect 26825 5397 26833 5431
rect 26781 5363 26833 5397
rect 27441 5431 27493 5465
rect 27441 5397 27449 5431
rect 27483 5397 27493 5431
rect 26781 5329 26791 5363
rect 26825 5329 26833 5363
rect 27441 5363 27493 5397
rect 26781 5317 26833 5329
rect 27441 5329 27449 5363
rect 27483 5329 27493 5363
rect 27441 5317 27493 5329
rect 27523 5317 27565 5517
rect 27595 5499 27647 5517
rect 27595 5465 27605 5499
rect 27639 5465 27647 5499
rect 27595 5431 27647 5465
rect 27595 5397 27605 5431
rect 27639 5397 27647 5431
rect 27595 5363 27647 5397
rect 27595 5329 27605 5363
rect 27639 5329 27647 5363
rect 27595 5317 27647 5329
rect 28515 5499 28567 5517
rect 28515 5465 28523 5499
rect 28557 5465 28567 5499
rect 28515 5431 28567 5465
rect 28515 5397 28523 5431
rect 28557 5397 28567 5431
rect 28515 5363 28567 5397
rect 28515 5329 28523 5363
rect 28557 5329 28567 5363
rect 28515 5317 28567 5329
rect 28597 5317 28639 5517
rect 28669 5499 28721 5517
rect 28669 5465 28679 5499
rect 28713 5465 28721 5499
rect 28936 5497 28948 5531
rect 28982 5497 28998 5531
rect 28936 5482 28998 5497
rect 29028 5667 29094 5682
rect 29028 5633 29044 5667
rect 29078 5633 29094 5667
rect 29028 5599 29094 5633
rect 29028 5565 29044 5599
rect 29078 5565 29094 5599
rect 29028 5531 29094 5565
rect 29028 5497 29044 5531
rect 29078 5497 29094 5531
rect 29028 5482 29094 5497
rect 29124 5667 29186 5682
rect 29124 5633 29140 5667
rect 29174 5633 29186 5667
rect 30824 5667 30886 5682
rect 29124 5599 29186 5633
rect 29124 5565 29140 5599
rect 29174 5565 29186 5599
rect 29124 5531 29186 5565
rect 29124 5497 29140 5531
rect 29174 5497 29186 5531
rect 30824 5633 30836 5667
rect 30870 5633 30886 5667
rect 30824 5599 30886 5633
rect 30824 5565 30836 5599
rect 30870 5565 30886 5599
rect 30824 5531 30886 5565
rect 29124 5482 29186 5497
rect 29329 5499 29381 5517
rect 28669 5431 28721 5465
rect 29329 5465 29337 5499
rect 29371 5465 29381 5499
rect 28669 5397 28679 5431
rect 28713 5397 28721 5431
rect 28669 5363 28721 5397
rect 29329 5431 29381 5465
rect 29329 5397 29337 5431
rect 29371 5397 29381 5431
rect 28669 5329 28679 5363
rect 28713 5329 28721 5363
rect 29329 5363 29381 5397
rect 28669 5317 28721 5329
rect 29329 5329 29337 5363
rect 29371 5329 29381 5363
rect 29329 5317 29381 5329
rect 29411 5317 29453 5517
rect 29483 5499 29535 5517
rect 29483 5465 29493 5499
rect 29527 5465 29535 5499
rect 29483 5431 29535 5465
rect 29483 5397 29493 5431
rect 29527 5397 29535 5431
rect 29483 5363 29535 5397
rect 29483 5329 29493 5363
rect 29527 5329 29535 5363
rect 29483 5317 29535 5329
rect 30403 5499 30455 5517
rect 30403 5465 30411 5499
rect 30445 5465 30455 5499
rect 30403 5431 30455 5465
rect 30403 5397 30411 5431
rect 30445 5397 30455 5431
rect 30403 5363 30455 5397
rect 30403 5329 30411 5363
rect 30445 5329 30455 5363
rect 30403 5317 30455 5329
rect 30485 5317 30527 5517
rect 30557 5499 30609 5517
rect 30557 5465 30567 5499
rect 30601 5465 30609 5499
rect 30824 5497 30836 5531
rect 30870 5497 30886 5531
rect 30824 5482 30886 5497
rect 30916 5667 30982 5682
rect 30916 5633 30932 5667
rect 30966 5633 30982 5667
rect 30916 5599 30982 5633
rect 30916 5565 30932 5599
rect 30966 5565 30982 5599
rect 30916 5531 30982 5565
rect 30916 5497 30932 5531
rect 30966 5497 30982 5531
rect 30916 5482 30982 5497
rect 31012 5667 31074 5682
rect 31012 5633 31028 5667
rect 31062 5633 31074 5667
rect 32712 5667 32774 5682
rect 31012 5599 31074 5633
rect 31012 5565 31028 5599
rect 31062 5565 31074 5599
rect 31012 5531 31074 5565
rect 31012 5497 31028 5531
rect 31062 5497 31074 5531
rect 32712 5633 32724 5667
rect 32758 5633 32774 5667
rect 32712 5599 32774 5633
rect 32712 5565 32724 5599
rect 32758 5565 32774 5599
rect 32712 5531 32774 5565
rect 31012 5482 31074 5497
rect 31217 5499 31269 5517
rect 30557 5431 30609 5465
rect 31217 5465 31225 5499
rect 31259 5465 31269 5499
rect 30557 5397 30567 5431
rect 30601 5397 30609 5431
rect 30557 5363 30609 5397
rect 31217 5431 31269 5465
rect 31217 5397 31225 5431
rect 31259 5397 31269 5431
rect 30557 5329 30567 5363
rect 30601 5329 30609 5363
rect 31217 5363 31269 5397
rect 30557 5317 30609 5329
rect 31217 5329 31225 5363
rect 31259 5329 31269 5363
rect 31217 5317 31269 5329
rect 31299 5317 31341 5517
rect 31371 5499 31423 5517
rect 31371 5465 31381 5499
rect 31415 5465 31423 5499
rect 31371 5431 31423 5465
rect 31371 5397 31381 5431
rect 31415 5397 31423 5431
rect 31371 5363 31423 5397
rect 31371 5329 31381 5363
rect 31415 5329 31423 5363
rect 31371 5317 31423 5329
rect 32291 5499 32343 5517
rect 32291 5465 32299 5499
rect 32333 5465 32343 5499
rect 32291 5431 32343 5465
rect 32291 5397 32299 5431
rect 32333 5397 32343 5431
rect 32291 5363 32343 5397
rect 32291 5329 32299 5363
rect 32333 5329 32343 5363
rect 32291 5317 32343 5329
rect 32373 5317 32415 5517
rect 32445 5499 32497 5517
rect 32445 5465 32455 5499
rect 32489 5465 32497 5499
rect 32712 5497 32724 5531
rect 32758 5497 32774 5531
rect 32712 5482 32774 5497
rect 32804 5667 32870 5682
rect 32804 5633 32820 5667
rect 32854 5633 32870 5667
rect 32804 5599 32870 5633
rect 32804 5565 32820 5599
rect 32854 5565 32870 5599
rect 32804 5531 32870 5565
rect 32804 5497 32820 5531
rect 32854 5497 32870 5531
rect 32804 5482 32870 5497
rect 32900 5667 32962 5682
rect 32900 5633 32916 5667
rect 32950 5633 32962 5667
rect 34600 5667 34662 5682
rect 32900 5599 32962 5633
rect 32900 5565 32916 5599
rect 32950 5565 32962 5599
rect 32900 5531 32962 5565
rect 32900 5497 32916 5531
rect 32950 5497 32962 5531
rect 34600 5633 34612 5667
rect 34646 5633 34662 5667
rect 34600 5599 34662 5633
rect 34600 5565 34612 5599
rect 34646 5565 34662 5599
rect 34600 5531 34662 5565
rect 32900 5482 32962 5497
rect 33105 5499 33157 5517
rect 32445 5431 32497 5465
rect 33105 5465 33113 5499
rect 33147 5465 33157 5499
rect 32445 5397 32455 5431
rect 32489 5397 32497 5431
rect 32445 5363 32497 5397
rect 33105 5431 33157 5465
rect 33105 5397 33113 5431
rect 33147 5397 33157 5431
rect 32445 5329 32455 5363
rect 32489 5329 32497 5363
rect 33105 5363 33157 5397
rect 32445 5317 32497 5329
rect 33105 5329 33113 5363
rect 33147 5329 33157 5363
rect 33105 5317 33157 5329
rect 33187 5317 33229 5517
rect 33259 5499 33311 5517
rect 33259 5465 33269 5499
rect 33303 5465 33311 5499
rect 33259 5431 33311 5465
rect 33259 5397 33269 5431
rect 33303 5397 33311 5431
rect 33259 5363 33311 5397
rect 33259 5329 33269 5363
rect 33303 5329 33311 5363
rect 33259 5317 33311 5329
rect 34179 5499 34231 5517
rect 34179 5465 34187 5499
rect 34221 5465 34231 5499
rect 34179 5431 34231 5465
rect 34179 5397 34187 5431
rect 34221 5397 34231 5431
rect 34179 5363 34231 5397
rect 34179 5329 34187 5363
rect 34221 5329 34231 5363
rect 34179 5317 34231 5329
rect 34261 5317 34303 5517
rect 34333 5499 34385 5517
rect 34333 5465 34343 5499
rect 34377 5465 34385 5499
rect 34600 5497 34612 5531
rect 34646 5497 34662 5531
rect 34600 5482 34662 5497
rect 34692 5667 34758 5682
rect 34692 5633 34708 5667
rect 34742 5633 34758 5667
rect 34692 5599 34758 5633
rect 34692 5565 34708 5599
rect 34742 5565 34758 5599
rect 34692 5531 34758 5565
rect 34692 5497 34708 5531
rect 34742 5497 34758 5531
rect 34692 5482 34758 5497
rect 34788 5667 34850 5682
rect 34788 5633 34804 5667
rect 34838 5633 34850 5667
rect 36488 5667 36550 5682
rect 34788 5599 34850 5633
rect 34788 5565 34804 5599
rect 34838 5565 34850 5599
rect 34788 5531 34850 5565
rect 34788 5497 34804 5531
rect 34838 5497 34850 5531
rect 36488 5633 36500 5667
rect 36534 5633 36550 5667
rect 36488 5599 36550 5633
rect 36488 5565 36500 5599
rect 36534 5565 36550 5599
rect 36488 5531 36550 5565
rect 34788 5482 34850 5497
rect 34993 5499 35045 5517
rect 34333 5431 34385 5465
rect 34993 5465 35001 5499
rect 35035 5465 35045 5499
rect 34333 5397 34343 5431
rect 34377 5397 34385 5431
rect 34333 5363 34385 5397
rect 34993 5431 35045 5465
rect 34993 5397 35001 5431
rect 35035 5397 35045 5431
rect 34333 5329 34343 5363
rect 34377 5329 34385 5363
rect 34993 5363 35045 5397
rect 34333 5317 34385 5329
rect 34993 5329 35001 5363
rect 35035 5329 35045 5363
rect 34993 5317 35045 5329
rect 35075 5317 35117 5517
rect 35147 5499 35199 5517
rect 35147 5465 35157 5499
rect 35191 5465 35199 5499
rect 35147 5431 35199 5465
rect 35147 5397 35157 5431
rect 35191 5397 35199 5431
rect 35147 5363 35199 5397
rect 35147 5329 35157 5363
rect 35191 5329 35199 5363
rect 35147 5317 35199 5329
rect 36067 5499 36119 5517
rect 36067 5465 36075 5499
rect 36109 5465 36119 5499
rect 36067 5431 36119 5465
rect 36067 5397 36075 5431
rect 36109 5397 36119 5431
rect 36067 5363 36119 5397
rect 36067 5329 36075 5363
rect 36109 5329 36119 5363
rect 36067 5317 36119 5329
rect 36149 5317 36191 5517
rect 36221 5499 36273 5517
rect 36221 5465 36231 5499
rect 36265 5465 36273 5499
rect 36488 5497 36500 5531
rect 36534 5497 36550 5531
rect 36488 5482 36550 5497
rect 36580 5667 36646 5682
rect 36580 5633 36596 5667
rect 36630 5633 36646 5667
rect 36580 5599 36646 5633
rect 36580 5565 36596 5599
rect 36630 5565 36646 5599
rect 36580 5531 36646 5565
rect 36580 5497 36596 5531
rect 36630 5497 36646 5531
rect 36580 5482 36646 5497
rect 36676 5667 36738 5682
rect 36676 5633 36692 5667
rect 36726 5633 36738 5667
rect 38376 5667 38438 5682
rect 36676 5599 36738 5633
rect 36676 5565 36692 5599
rect 36726 5565 36738 5599
rect 36676 5531 36738 5565
rect 36676 5497 36692 5531
rect 36726 5497 36738 5531
rect 38376 5633 38388 5667
rect 38422 5633 38438 5667
rect 38376 5599 38438 5633
rect 38376 5565 38388 5599
rect 38422 5565 38438 5599
rect 38376 5531 38438 5565
rect 36676 5482 36738 5497
rect 36881 5499 36933 5517
rect 36221 5431 36273 5465
rect 36881 5465 36889 5499
rect 36923 5465 36933 5499
rect 36221 5397 36231 5431
rect 36265 5397 36273 5431
rect 36221 5363 36273 5397
rect 36881 5431 36933 5465
rect 36881 5397 36889 5431
rect 36923 5397 36933 5431
rect 36221 5329 36231 5363
rect 36265 5329 36273 5363
rect 36881 5363 36933 5397
rect 36221 5317 36273 5329
rect 36881 5329 36889 5363
rect 36923 5329 36933 5363
rect 36881 5317 36933 5329
rect 36963 5317 37005 5517
rect 37035 5499 37087 5517
rect 37035 5465 37045 5499
rect 37079 5465 37087 5499
rect 37035 5431 37087 5465
rect 37035 5397 37045 5431
rect 37079 5397 37087 5431
rect 37035 5363 37087 5397
rect 37035 5329 37045 5363
rect 37079 5329 37087 5363
rect 37035 5317 37087 5329
rect 37955 5499 38007 5517
rect 37955 5465 37963 5499
rect 37997 5465 38007 5499
rect 37955 5431 38007 5465
rect 37955 5397 37963 5431
rect 37997 5397 38007 5431
rect 37955 5363 38007 5397
rect 37955 5329 37963 5363
rect 37997 5329 38007 5363
rect 37955 5317 38007 5329
rect 38037 5317 38079 5517
rect 38109 5499 38161 5517
rect 38109 5465 38119 5499
rect 38153 5465 38161 5499
rect 38376 5497 38388 5531
rect 38422 5497 38438 5531
rect 38376 5482 38438 5497
rect 38468 5667 38534 5682
rect 38468 5633 38484 5667
rect 38518 5633 38534 5667
rect 38468 5599 38534 5633
rect 38468 5565 38484 5599
rect 38518 5565 38534 5599
rect 38468 5531 38534 5565
rect 38468 5497 38484 5531
rect 38518 5497 38534 5531
rect 38468 5482 38534 5497
rect 38564 5667 38626 5682
rect 38564 5633 38580 5667
rect 38614 5633 38626 5667
rect 40264 5667 40326 5682
rect 38564 5599 38626 5633
rect 38564 5565 38580 5599
rect 38614 5565 38626 5599
rect 38564 5531 38626 5565
rect 38564 5497 38580 5531
rect 38614 5497 38626 5531
rect 40264 5633 40276 5667
rect 40310 5633 40326 5667
rect 40264 5599 40326 5633
rect 40264 5565 40276 5599
rect 40310 5565 40326 5599
rect 40264 5531 40326 5565
rect 38564 5482 38626 5497
rect 38769 5499 38821 5517
rect 38109 5431 38161 5465
rect 38769 5465 38777 5499
rect 38811 5465 38821 5499
rect 38109 5397 38119 5431
rect 38153 5397 38161 5431
rect 38109 5363 38161 5397
rect 38769 5431 38821 5465
rect 38769 5397 38777 5431
rect 38811 5397 38821 5431
rect 38109 5329 38119 5363
rect 38153 5329 38161 5363
rect 38769 5363 38821 5397
rect 38109 5317 38161 5329
rect 38769 5329 38777 5363
rect 38811 5329 38821 5363
rect 38769 5317 38821 5329
rect 38851 5317 38893 5517
rect 38923 5499 38975 5517
rect 38923 5465 38933 5499
rect 38967 5465 38975 5499
rect 38923 5431 38975 5465
rect 38923 5397 38933 5431
rect 38967 5397 38975 5431
rect 38923 5363 38975 5397
rect 38923 5329 38933 5363
rect 38967 5329 38975 5363
rect 38923 5317 38975 5329
rect 39843 5499 39895 5517
rect 39843 5465 39851 5499
rect 39885 5465 39895 5499
rect 39843 5431 39895 5465
rect 39843 5397 39851 5431
rect 39885 5397 39895 5431
rect 39843 5363 39895 5397
rect 39843 5329 39851 5363
rect 39885 5329 39895 5363
rect 39843 5317 39895 5329
rect 39925 5317 39967 5517
rect 39997 5499 40049 5517
rect 39997 5465 40007 5499
rect 40041 5465 40049 5499
rect 40264 5497 40276 5531
rect 40310 5497 40326 5531
rect 40264 5482 40326 5497
rect 40356 5667 40422 5682
rect 40356 5633 40372 5667
rect 40406 5633 40422 5667
rect 40356 5599 40422 5633
rect 40356 5565 40372 5599
rect 40406 5565 40422 5599
rect 40356 5531 40422 5565
rect 40356 5497 40372 5531
rect 40406 5497 40422 5531
rect 40356 5482 40422 5497
rect 40452 5667 40514 5682
rect 40452 5633 40468 5667
rect 40502 5633 40514 5667
rect 42152 5667 42214 5682
rect 40452 5599 40514 5633
rect 40452 5565 40468 5599
rect 40502 5565 40514 5599
rect 40452 5531 40514 5565
rect 40452 5497 40468 5531
rect 40502 5497 40514 5531
rect 42152 5633 42164 5667
rect 42198 5633 42214 5667
rect 42152 5599 42214 5633
rect 42152 5565 42164 5599
rect 42198 5565 42214 5599
rect 42152 5531 42214 5565
rect 40452 5482 40514 5497
rect 40657 5499 40709 5517
rect 39997 5431 40049 5465
rect 40657 5465 40665 5499
rect 40699 5465 40709 5499
rect 39997 5397 40007 5431
rect 40041 5397 40049 5431
rect 39997 5363 40049 5397
rect 40657 5431 40709 5465
rect 40657 5397 40665 5431
rect 40699 5397 40709 5431
rect 39997 5329 40007 5363
rect 40041 5329 40049 5363
rect 40657 5363 40709 5397
rect 39997 5317 40049 5329
rect 40657 5329 40665 5363
rect 40699 5329 40709 5363
rect 40657 5317 40709 5329
rect 40739 5317 40781 5517
rect 40811 5499 40863 5517
rect 40811 5465 40821 5499
rect 40855 5465 40863 5499
rect 40811 5431 40863 5465
rect 40811 5397 40821 5431
rect 40855 5397 40863 5431
rect 40811 5363 40863 5397
rect 40811 5329 40821 5363
rect 40855 5329 40863 5363
rect 40811 5317 40863 5329
rect 41731 5499 41783 5517
rect 41731 5465 41739 5499
rect 41773 5465 41783 5499
rect 41731 5431 41783 5465
rect 41731 5397 41739 5431
rect 41773 5397 41783 5431
rect 41731 5363 41783 5397
rect 41731 5329 41739 5363
rect 41773 5329 41783 5363
rect 41731 5317 41783 5329
rect 41813 5317 41855 5517
rect 41885 5499 41937 5517
rect 41885 5465 41895 5499
rect 41929 5465 41937 5499
rect 42152 5497 42164 5531
rect 42198 5497 42214 5531
rect 42152 5482 42214 5497
rect 42244 5667 42310 5682
rect 42244 5633 42260 5667
rect 42294 5633 42310 5667
rect 42244 5599 42310 5633
rect 42244 5565 42260 5599
rect 42294 5565 42310 5599
rect 42244 5531 42310 5565
rect 42244 5497 42260 5531
rect 42294 5497 42310 5531
rect 42244 5482 42310 5497
rect 42340 5667 42402 5682
rect 42340 5633 42356 5667
rect 42390 5633 42402 5667
rect 44040 5667 44102 5682
rect 42340 5599 42402 5633
rect 42340 5565 42356 5599
rect 42390 5565 42402 5599
rect 42340 5531 42402 5565
rect 42340 5497 42356 5531
rect 42390 5497 42402 5531
rect 44040 5633 44052 5667
rect 44086 5633 44102 5667
rect 44040 5599 44102 5633
rect 44040 5565 44052 5599
rect 44086 5565 44102 5599
rect 44040 5531 44102 5565
rect 42340 5482 42402 5497
rect 42545 5499 42597 5517
rect 41885 5431 41937 5465
rect 42545 5465 42553 5499
rect 42587 5465 42597 5499
rect 41885 5397 41895 5431
rect 41929 5397 41937 5431
rect 41885 5363 41937 5397
rect 42545 5431 42597 5465
rect 42545 5397 42553 5431
rect 42587 5397 42597 5431
rect 41885 5329 41895 5363
rect 41929 5329 41937 5363
rect 42545 5363 42597 5397
rect 41885 5317 41937 5329
rect 42545 5329 42553 5363
rect 42587 5329 42597 5363
rect 42545 5317 42597 5329
rect 42627 5317 42669 5517
rect 42699 5499 42751 5517
rect 42699 5465 42709 5499
rect 42743 5465 42751 5499
rect 42699 5431 42751 5465
rect 42699 5397 42709 5431
rect 42743 5397 42751 5431
rect 42699 5363 42751 5397
rect 42699 5329 42709 5363
rect 42743 5329 42751 5363
rect 42699 5317 42751 5329
rect 43619 5499 43671 5517
rect 43619 5465 43627 5499
rect 43661 5465 43671 5499
rect 43619 5431 43671 5465
rect 43619 5397 43627 5431
rect 43661 5397 43671 5431
rect 43619 5363 43671 5397
rect 43619 5329 43627 5363
rect 43661 5329 43671 5363
rect 43619 5317 43671 5329
rect 43701 5317 43743 5517
rect 43773 5499 43825 5517
rect 43773 5465 43783 5499
rect 43817 5465 43825 5499
rect 44040 5497 44052 5531
rect 44086 5497 44102 5531
rect 44040 5482 44102 5497
rect 44132 5667 44198 5682
rect 44132 5633 44148 5667
rect 44182 5633 44198 5667
rect 44132 5599 44198 5633
rect 44132 5565 44148 5599
rect 44182 5565 44198 5599
rect 44132 5531 44198 5565
rect 44132 5497 44148 5531
rect 44182 5497 44198 5531
rect 44132 5482 44198 5497
rect 44228 5667 44290 5682
rect 44228 5633 44244 5667
rect 44278 5633 44290 5667
rect 45922 5667 45984 5682
rect 44228 5599 44290 5633
rect 44228 5565 44244 5599
rect 44278 5565 44290 5599
rect 44228 5531 44290 5565
rect 44228 5497 44244 5531
rect 44278 5497 44290 5531
rect 45922 5633 45934 5667
rect 45968 5633 45984 5667
rect 45922 5599 45984 5633
rect 45922 5565 45934 5599
rect 45968 5565 45984 5599
rect 45922 5531 45984 5565
rect 44228 5482 44290 5497
rect 44433 5499 44485 5517
rect 43773 5431 43825 5465
rect 44433 5465 44441 5499
rect 44475 5465 44485 5499
rect 43773 5397 43783 5431
rect 43817 5397 43825 5431
rect 43773 5363 43825 5397
rect 44433 5431 44485 5465
rect 44433 5397 44441 5431
rect 44475 5397 44485 5431
rect 43773 5329 43783 5363
rect 43817 5329 43825 5363
rect 44433 5363 44485 5397
rect 43773 5317 43825 5329
rect 44433 5329 44441 5363
rect 44475 5329 44485 5363
rect 44433 5317 44485 5329
rect 44515 5317 44557 5517
rect 44587 5499 44639 5517
rect 44587 5465 44597 5499
rect 44631 5465 44639 5499
rect 44587 5431 44639 5465
rect 44587 5397 44597 5431
rect 44631 5397 44639 5431
rect 44587 5363 44639 5397
rect 44587 5329 44597 5363
rect 44631 5329 44639 5363
rect 44587 5317 44639 5329
rect 45501 5499 45553 5517
rect 45501 5465 45509 5499
rect 45543 5465 45553 5499
rect 45501 5431 45553 5465
rect 45501 5397 45509 5431
rect 45543 5397 45553 5431
rect 45501 5363 45553 5397
rect 45501 5329 45509 5363
rect 45543 5329 45553 5363
rect 45501 5317 45553 5329
rect 45583 5317 45625 5517
rect 45655 5499 45707 5517
rect 45655 5465 45665 5499
rect 45699 5465 45707 5499
rect 45922 5497 45934 5531
rect 45968 5497 45984 5531
rect 45922 5482 45984 5497
rect 46014 5667 46080 5682
rect 46014 5633 46030 5667
rect 46064 5633 46080 5667
rect 46014 5599 46080 5633
rect 46014 5565 46030 5599
rect 46064 5565 46080 5599
rect 46014 5531 46080 5565
rect 46014 5497 46030 5531
rect 46064 5497 46080 5531
rect 46014 5482 46080 5497
rect 46110 5667 46172 5682
rect 46110 5633 46126 5667
rect 46160 5633 46172 5667
rect 47810 5667 47872 5682
rect 46110 5599 46172 5633
rect 46110 5565 46126 5599
rect 46160 5565 46172 5599
rect 46110 5531 46172 5565
rect 46110 5497 46126 5531
rect 46160 5497 46172 5531
rect 47810 5633 47822 5667
rect 47856 5633 47872 5667
rect 47810 5599 47872 5633
rect 47810 5565 47822 5599
rect 47856 5565 47872 5599
rect 47810 5531 47872 5565
rect 46110 5482 46172 5497
rect 46315 5499 46367 5517
rect 45655 5431 45707 5465
rect 46315 5465 46323 5499
rect 46357 5465 46367 5499
rect 45655 5397 45665 5431
rect 45699 5397 45707 5431
rect 45655 5363 45707 5397
rect 46315 5431 46367 5465
rect 46315 5397 46323 5431
rect 46357 5397 46367 5431
rect 45655 5329 45665 5363
rect 45699 5329 45707 5363
rect 46315 5363 46367 5397
rect 45655 5317 45707 5329
rect 46315 5329 46323 5363
rect 46357 5329 46367 5363
rect 46315 5317 46367 5329
rect 46397 5317 46439 5517
rect 46469 5499 46521 5517
rect 46469 5465 46479 5499
rect 46513 5465 46521 5499
rect 46469 5431 46521 5465
rect 46469 5397 46479 5431
rect 46513 5397 46521 5431
rect 46469 5363 46521 5397
rect 46469 5329 46479 5363
rect 46513 5329 46521 5363
rect 46469 5317 46521 5329
rect 47389 5499 47441 5517
rect 47389 5465 47397 5499
rect 47431 5465 47441 5499
rect 47389 5431 47441 5465
rect 47389 5397 47397 5431
rect 47431 5397 47441 5431
rect 47389 5363 47441 5397
rect 47389 5329 47397 5363
rect 47431 5329 47441 5363
rect 47389 5317 47441 5329
rect 47471 5317 47513 5517
rect 47543 5499 47595 5517
rect 47543 5465 47553 5499
rect 47587 5465 47595 5499
rect 47810 5497 47822 5531
rect 47856 5497 47872 5531
rect 47810 5482 47872 5497
rect 47902 5667 47968 5682
rect 47902 5633 47918 5667
rect 47952 5633 47968 5667
rect 47902 5599 47968 5633
rect 47902 5565 47918 5599
rect 47952 5565 47968 5599
rect 47902 5531 47968 5565
rect 47902 5497 47918 5531
rect 47952 5497 47968 5531
rect 47902 5482 47968 5497
rect 47998 5667 48060 5682
rect 47998 5633 48014 5667
rect 48048 5633 48060 5667
rect 49698 5667 49760 5682
rect 47998 5599 48060 5633
rect 47998 5565 48014 5599
rect 48048 5565 48060 5599
rect 47998 5531 48060 5565
rect 47998 5497 48014 5531
rect 48048 5497 48060 5531
rect 49698 5633 49710 5667
rect 49744 5633 49760 5667
rect 49698 5599 49760 5633
rect 49698 5565 49710 5599
rect 49744 5565 49760 5599
rect 49698 5531 49760 5565
rect 47998 5482 48060 5497
rect 48203 5499 48255 5517
rect 47543 5431 47595 5465
rect 48203 5465 48211 5499
rect 48245 5465 48255 5499
rect 47543 5397 47553 5431
rect 47587 5397 47595 5431
rect 47543 5363 47595 5397
rect 48203 5431 48255 5465
rect 48203 5397 48211 5431
rect 48245 5397 48255 5431
rect 47543 5329 47553 5363
rect 47587 5329 47595 5363
rect 48203 5363 48255 5397
rect 47543 5317 47595 5329
rect 48203 5329 48211 5363
rect 48245 5329 48255 5363
rect 48203 5317 48255 5329
rect 48285 5317 48327 5517
rect 48357 5499 48409 5517
rect 48357 5465 48367 5499
rect 48401 5465 48409 5499
rect 48357 5431 48409 5465
rect 48357 5397 48367 5431
rect 48401 5397 48409 5431
rect 48357 5363 48409 5397
rect 48357 5329 48367 5363
rect 48401 5329 48409 5363
rect 48357 5317 48409 5329
rect 49277 5499 49329 5517
rect 49277 5465 49285 5499
rect 49319 5465 49329 5499
rect 49277 5431 49329 5465
rect 49277 5397 49285 5431
rect 49319 5397 49329 5431
rect 49277 5363 49329 5397
rect 49277 5329 49285 5363
rect 49319 5329 49329 5363
rect 49277 5317 49329 5329
rect 49359 5317 49401 5517
rect 49431 5499 49483 5517
rect 49431 5465 49441 5499
rect 49475 5465 49483 5499
rect 49698 5497 49710 5531
rect 49744 5497 49760 5531
rect 49698 5482 49760 5497
rect 49790 5667 49856 5682
rect 49790 5633 49806 5667
rect 49840 5633 49856 5667
rect 49790 5599 49856 5633
rect 49790 5565 49806 5599
rect 49840 5565 49856 5599
rect 49790 5531 49856 5565
rect 49790 5497 49806 5531
rect 49840 5497 49856 5531
rect 49790 5482 49856 5497
rect 49886 5667 49948 5682
rect 49886 5633 49902 5667
rect 49936 5633 49948 5667
rect 51586 5667 51648 5682
rect 49886 5599 49948 5633
rect 49886 5565 49902 5599
rect 49936 5565 49948 5599
rect 49886 5531 49948 5565
rect 49886 5497 49902 5531
rect 49936 5497 49948 5531
rect 51586 5633 51598 5667
rect 51632 5633 51648 5667
rect 51586 5599 51648 5633
rect 51586 5565 51598 5599
rect 51632 5565 51648 5599
rect 51586 5531 51648 5565
rect 49886 5482 49948 5497
rect 50091 5499 50143 5517
rect 49431 5431 49483 5465
rect 50091 5465 50099 5499
rect 50133 5465 50143 5499
rect 49431 5397 49441 5431
rect 49475 5397 49483 5431
rect 49431 5363 49483 5397
rect 50091 5431 50143 5465
rect 50091 5397 50099 5431
rect 50133 5397 50143 5431
rect 49431 5329 49441 5363
rect 49475 5329 49483 5363
rect 50091 5363 50143 5397
rect 49431 5317 49483 5329
rect 50091 5329 50099 5363
rect 50133 5329 50143 5363
rect 50091 5317 50143 5329
rect 50173 5317 50215 5517
rect 50245 5499 50297 5517
rect 50245 5465 50255 5499
rect 50289 5465 50297 5499
rect 50245 5431 50297 5465
rect 50245 5397 50255 5431
rect 50289 5397 50297 5431
rect 50245 5363 50297 5397
rect 50245 5329 50255 5363
rect 50289 5329 50297 5363
rect 50245 5317 50297 5329
rect 51165 5499 51217 5517
rect 51165 5465 51173 5499
rect 51207 5465 51217 5499
rect 51165 5431 51217 5465
rect 51165 5397 51173 5431
rect 51207 5397 51217 5431
rect 51165 5363 51217 5397
rect 51165 5329 51173 5363
rect 51207 5329 51217 5363
rect 51165 5317 51217 5329
rect 51247 5317 51289 5517
rect 51319 5499 51371 5517
rect 51319 5465 51329 5499
rect 51363 5465 51371 5499
rect 51586 5497 51598 5531
rect 51632 5497 51648 5531
rect 51586 5482 51648 5497
rect 51678 5667 51744 5682
rect 51678 5633 51694 5667
rect 51728 5633 51744 5667
rect 51678 5599 51744 5633
rect 51678 5565 51694 5599
rect 51728 5565 51744 5599
rect 51678 5531 51744 5565
rect 51678 5497 51694 5531
rect 51728 5497 51744 5531
rect 51678 5482 51744 5497
rect 51774 5667 51836 5682
rect 51774 5633 51790 5667
rect 51824 5633 51836 5667
rect 53474 5667 53536 5682
rect 51774 5599 51836 5633
rect 51774 5565 51790 5599
rect 51824 5565 51836 5599
rect 51774 5531 51836 5565
rect 51774 5497 51790 5531
rect 51824 5497 51836 5531
rect 53474 5633 53486 5667
rect 53520 5633 53536 5667
rect 53474 5599 53536 5633
rect 53474 5565 53486 5599
rect 53520 5565 53536 5599
rect 53474 5531 53536 5565
rect 51774 5482 51836 5497
rect 51979 5499 52031 5517
rect 51319 5431 51371 5465
rect 51979 5465 51987 5499
rect 52021 5465 52031 5499
rect 51319 5397 51329 5431
rect 51363 5397 51371 5431
rect 51319 5363 51371 5397
rect 51979 5431 52031 5465
rect 51979 5397 51987 5431
rect 52021 5397 52031 5431
rect 51319 5329 51329 5363
rect 51363 5329 51371 5363
rect 51979 5363 52031 5397
rect 51319 5317 51371 5329
rect 51979 5329 51987 5363
rect 52021 5329 52031 5363
rect 51979 5317 52031 5329
rect 52061 5317 52103 5517
rect 52133 5499 52185 5517
rect 52133 5465 52143 5499
rect 52177 5465 52185 5499
rect 52133 5431 52185 5465
rect 52133 5397 52143 5431
rect 52177 5397 52185 5431
rect 52133 5363 52185 5397
rect 52133 5329 52143 5363
rect 52177 5329 52185 5363
rect 52133 5317 52185 5329
rect 53053 5499 53105 5517
rect 53053 5465 53061 5499
rect 53095 5465 53105 5499
rect 53053 5431 53105 5465
rect 53053 5397 53061 5431
rect 53095 5397 53105 5431
rect 53053 5363 53105 5397
rect 53053 5329 53061 5363
rect 53095 5329 53105 5363
rect 53053 5317 53105 5329
rect 53135 5317 53177 5517
rect 53207 5499 53259 5517
rect 53207 5465 53217 5499
rect 53251 5465 53259 5499
rect 53474 5497 53486 5531
rect 53520 5497 53536 5531
rect 53474 5482 53536 5497
rect 53566 5667 53632 5682
rect 53566 5633 53582 5667
rect 53616 5633 53632 5667
rect 53566 5599 53632 5633
rect 53566 5565 53582 5599
rect 53616 5565 53632 5599
rect 53566 5531 53632 5565
rect 53566 5497 53582 5531
rect 53616 5497 53632 5531
rect 53566 5482 53632 5497
rect 53662 5667 53724 5682
rect 53662 5633 53678 5667
rect 53712 5633 53724 5667
rect 55362 5667 55424 5682
rect 53662 5599 53724 5633
rect 53662 5565 53678 5599
rect 53712 5565 53724 5599
rect 53662 5531 53724 5565
rect 53662 5497 53678 5531
rect 53712 5497 53724 5531
rect 55362 5633 55374 5667
rect 55408 5633 55424 5667
rect 55362 5599 55424 5633
rect 55362 5565 55374 5599
rect 55408 5565 55424 5599
rect 55362 5531 55424 5565
rect 53662 5482 53724 5497
rect 53867 5499 53919 5517
rect 53207 5431 53259 5465
rect 53867 5465 53875 5499
rect 53909 5465 53919 5499
rect 53207 5397 53217 5431
rect 53251 5397 53259 5431
rect 53207 5363 53259 5397
rect 53867 5431 53919 5465
rect 53867 5397 53875 5431
rect 53909 5397 53919 5431
rect 53207 5329 53217 5363
rect 53251 5329 53259 5363
rect 53867 5363 53919 5397
rect 53207 5317 53259 5329
rect 53867 5329 53875 5363
rect 53909 5329 53919 5363
rect 53867 5317 53919 5329
rect 53949 5317 53991 5517
rect 54021 5499 54073 5517
rect 54021 5465 54031 5499
rect 54065 5465 54073 5499
rect 54021 5431 54073 5465
rect 54021 5397 54031 5431
rect 54065 5397 54073 5431
rect 54021 5363 54073 5397
rect 54021 5329 54031 5363
rect 54065 5329 54073 5363
rect 54021 5317 54073 5329
rect 54941 5499 54993 5517
rect 54941 5465 54949 5499
rect 54983 5465 54993 5499
rect 54941 5431 54993 5465
rect 54941 5397 54949 5431
rect 54983 5397 54993 5431
rect 54941 5363 54993 5397
rect 54941 5329 54949 5363
rect 54983 5329 54993 5363
rect 54941 5317 54993 5329
rect 55023 5317 55065 5517
rect 55095 5499 55147 5517
rect 55095 5465 55105 5499
rect 55139 5465 55147 5499
rect 55362 5497 55374 5531
rect 55408 5497 55424 5531
rect 55362 5482 55424 5497
rect 55454 5667 55520 5682
rect 55454 5633 55470 5667
rect 55504 5633 55520 5667
rect 55454 5599 55520 5633
rect 55454 5565 55470 5599
rect 55504 5565 55520 5599
rect 55454 5531 55520 5565
rect 55454 5497 55470 5531
rect 55504 5497 55520 5531
rect 55454 5482 55520 5497
rect 55550 5667 55612 5682
rect 55550 5633 55566 5667
rect 55600 5633 55612 5667
rect 57250 5667 57312 5682
rect 55550 5599 55612 5633
rect 55550 5565 55566 5599
rect 55600 5565 55612 5599
rect 55550 5531 55612 5565
rect 55550 5497 55566 5531
rect 55600 5497 55612 5531
rect 57250 5633 57262 5667
rect 57296 5633 57312 5667
rect 57250 5599 57312 5633
rect 57250 5565 57262 5599
rect 57296 5565 57312 5599
rect 57250 5531 57312 5565
rect 55550 5482 55612 5497
rect 55755 5499 55807 5517
rect 55095 5431 55147 5465
rect 55755 5465 55763 5499
rect 55797 5465 55807 5499
rect 55095 5397 55105 5431
rect 55139 5397 55147 5431
rect 55095 5363 55147 5397
rect 55755 5431 55807 5465
rect 55755 5397 55763 5431
rect 55797 5397 55807 5431
rect 55095 5329 55105 5363
rect 55139 5329 55147 5363
rect 55755 5363 55807 5397
rect 55095 5317 55147 5329
rect 55755 5329 55763 5363
rect 55797 5329 55807 5363
rect 55755 5317 55807 5329
rect 55837 5317 55879 5517
rect 55909 5499 55961 5517
rect 55909 5465 55919 5499
rect 55953 5465 55961 5499
rect 55909 5431 55961 5465
rect 55909 5397 55919 5431
rect 55953 5397 55961 5431
rect 55909 5363 55961 5397
rect 55909 5329 55919 5363
rect 55953 5329 55961 5363
rect 55909 5317 55961 5329
rect 56829 5499 56881 5517
rect 56829 5465 56837 5499
rect 56871 5465 56881 5499
rect 56829 5431 56881 5465
rect 56829 5397 56837 5431
rect 56871 5397 56881 5431
rect 56829 5363 56881 5397
rect 56829 5329 56837 5363
rect 56871 5329 56881 5363
rect 56829 5317 56881 5329
rect 56911 5317 56953 5517
rect 56983 5499 57035 5517
rect 56983 5465 56993 5499
rect 57027 5465 57035 5499
rect 57250 5497 57262 5531
rect 57296 5497 57312 5531
rect 57250 5482 57312 5497
rect 57342 5667 57408 5682
rect 57342 5633 57358 5667
rect 57392 5633 57408 5667
rect 57342 5599 57408 5633
rect 57342 5565 57358 5599
rect 57392 5565 57408 5599
rect 57342 5531 57408 5565
rect 57342 5497 57358 5531
rect 57392 5497 57408 5531
rect 57342 5482 57408 5497
rect 57438 5667 57500 5682
rect 57438 5633 57454 5667
rect 57488 5633 57500 5667
rect 59138 5667 59200 5682
rect 57438 5599 57500 5633
rect 57438 5565 57454 5599
rect 57488 5565 57500 5599
rect 57438 5531 57500 5565
rect 57438 5497 57454 5531
rect 57488 5497 57500 5531
rect 59138 5633 59150 5667
rect 59184 5633 59200 5667
rect 59138 5599 59200 5633
rect 59138 5565 59150 5599
rect 59184 5565 59200 5599
rect 59138 5531 59200 5565
rect 57438 5482 57500 5497
rect 57643 5499 57695 5517
rect 56983 5431 57035 5465
rect 57643 5465 57651 5499
rect 57685 5465 57695 5499
rect 56983 5397 56993 5431
rect 57027 5397 57035 5431
rect 56983 5363 57035 5397
rect 57643 5431 57695 5465
rect 57643 5397 57651 5431
rect 57685 5397 57695 5431
rect 56983 5329 56993 5363
rect 57027 5329 57035 5363
rect 57643 5363 57695 5397
rect 56983 5317 57035 5329
rect 57643 5329 57651 5363
rect 57685 5329 57695 5363
rect 57643 5317 57695 5329
rect 57725 5317 57767 5517
rect 57797 5499 57849 5517
rect 57797 5465 57807 5499
rect 57841 5465 57849 5499
rect 57797 5431 57849 5465
rect 57797 5397 57807 5431
rect 57841 5397 57849 5431
rect 57797 5363 57849 5397
rect 57797 5329 57807 5363
rect 57841 5329 57849 5363
rect 57797 5317 57849 5329
rect 58717 5499 58769 5517
rect 58717 5465 58725 5499
rect 58759 5465 58769 5499
rect 58717 5431 58769 5465
rect 58717 5397 58725 5431
rect 58759 5397 58769 5431
rect 58717 5363 58769 5397
rect 58717 5329 58725 5363
rect 58759 5329 58769 5363
rect 58717 5317 58769 5329
rect 58799 5317 58841 5517
rect 58871 5499 58923 5517
rect 58871 5465 58881 5499
rect 58915 5465 58923 5499
rect 59138 5497 59150 5531
rect 59184 5497 59200 5531
rect 59138 5482 59200 5497
rect 59230 5667 59296 5682
rect 59230 5633 59246 5667
rect 59280 5633 59296 5667
rect 59230 5599 59296 5633
rect 59230 5565 59246 5599
rect 59280 5565 59296 5599
rect 59230 5531 59296 5565
rect 59230 5497 59246 5531
rect 59280 5497 59296 5531
rect 59230 5482 59296 5497
rect 59326 5667 59388 5682
rect 59326 5633 59342 5667
rect 59376 5633 59388 5667
rect 59326 5599 59388 5633
rect 59326 5565 59342 5599
rect 59376 5565 59388 5599
rect 59326 5531 59388 5565
rect 59326 5497 59342 5531
rect 59376 5497 59388 5531
rect 59326 5482 59388 5497
rect 59531 5499 59583 5517
rect 58871 5431 58923 5465
rect 59531 5465 59539 5499
rect 59573 5465 59583 5499
rect 58871 5397 58881 5431
rect 58915 5397 58923 5431
rect 58871 5363 58923 5397
rect 59531 5431 59583 5465
rect 59531 5397 59539 5431
rect 59573 5397 59583 5431
rect 58871 5329 58881 5363
rect 58915 5329 58923 5363
rect 59531 5363 59583 5397
rect 58871 5317 58923 5329
rect 59531 5329 59539 5363
rect 59573 5329 59583 5363
rect 59531 5317 59583 5329
rect 59613 5317 59655 5517
rect 59685 5499 59737 5517
rect 59685 5465 59695 5499
rect 59729 5465 59737 5499
rect 59685 5431 59737 5465
rect 59685 5397 59695 5431
rect 59729 5397 59737 5431
rect 59685 5363 59737 5397
rect 59685 5329 59695 5363
rect 59729 5329 59737 5363
rect 59685 5317 59737 5329
rect 5702 5133 5754 5145
rect 5702 5099 5710 5133
rect 5744 5099 5754 5133
rect 5702 5065 5754 5099
rect 5702 5031 5710 5065
rect 5744 5031 5754 5065
rect 5702 4945 5754 5031
rect 5784 5133 5838 5145
rect 5784 5099 5794 5133
rect 5828 5099 5838 5133
rect 5784 5065 5838 5099
rect 5784 5031 5794 5065
rect 5828 5031 5838 5065
rect 5784 4995 5838 5031
rect 5784 4961 5794 4995
rect 5828 4961 5838 4995
rect 5784 4945 5838 4961
rect 5868 5133 5922 5145
rect 5868 5099 5878 5133
rect 5912 5099 5922 5133
rect 5868 5065 5922 5099
rect 5868 5031 5878 5065
rect 5912 5031 5922 5065
rect 5868 4945 5922 5031
rect 5952 5133 6006 5145
rect 5952 5099 5962 5133
rect 5996 5099 6006 5133
rect 5952 5065 6006 5099
rect 5952 5031 5962 5065
rect 5996 5031 6006 5065
rect 5952 4995 6006 5031
rect 5952 4961 5962 4995
rect 5996 4961 6006 4995
rect 5952 4945 6006 4961
rect 6036 5133 6090 5145
rect 6036 5099 6046 5133
rect 6080 5099 6090 5133
rect 6036 5065 6090 5099
rect 6036 5031 6046 5065
rect 6080 5031 6090 5065
rect 6036 4945 6090 5031
rect 6120 5133 6174 5145
rect 6120 5099 6130 5133
rect 6164 5099 6174 5133
rect 6120 5065 6174 5099
rect 6120 5031 6130 5065
rect 6164 5031 6174 5065
rect 6120 4995 6174 5031
rect 6120 4961 6130 4995
rect 6164 4961 6174 4995
rect 6120 4945 6174 4961
rect 6204 5133 6258 5145
rect 6204 5099 6214 5133
rect 6248 5099 6258 5133
rect 6204 5065 6258 5099
rect 6204 5031 6214 5065
rect 6248 5031 6258 5065
rect 6204 4945 6258 5031
rect 6288 5133 6342 5145
rect 6288 5099 6298 5133
rect 6332 5099 6342 5133
rect 6288 5065 6342 5099
rect 6288 5031 6298 5065
rect 6332 5031 6342 5065
rect 6288 4995 6342 5031
rect 6288 4961 6298 4995
rect 6332 4961 6342 4995
rect 6288 4945 6342 4961
rect 6372 5133 6426 5145
rect 6372 5099 6382 5133
rect 6416 5099 6426 5133
rect 6372 5065 6426 5099
rect 6372 5031 6382 5065
rect 6416 5031 6426 5065
rect 6372 4945 6426 5031
rect 6456 5133 6510 5145
rect 6456 5099 6466 5133
rect 6500 5099 6510 5133
rect 6456 5065 6510 5099
rect 6456 5031 6466 5065
rect 6500 5031 6510 5065
rect 6456 4995 6510 5031
rect 6456 4961 6466 4995
rect 6500 4961 6510 4995
rect 6456 4945 6510 4961
rect 6540 5133 6594 5145
rect 6540 5099 6550 5133
rect 6584 5099 6594 5133
rect 6540 5065 6594 5099
rect 6540 5031 6550 5065
rect 6584 5031 6594 5065
rect 6540 4945 6594 5031
rect 6624 5133 6678 5145
rect 6624 5099 6634 5133
rect 6668 5099 6678 5133
rect 6624 5065 6678 5099
rect 6624 5031 6634 5065
rect 6668 5031 6678 5065
rect 6624 4995 6678 5031
rect 6624 4961 6634 4995
rect 6668 4961 6678 4995
rect 6624 4945 6678 4961
rect 6708 5133 6762 5145
rect 6708 5099 6718 5133
rect 6752 5099 6762 5133
rect 6708 5065 6762 5099
rect 6708 5031 6718 5065
rect 6752 5031 6762 5065
rect 6708 4945 6762 5031
rect 6792 5133 6846 5145
rect 6792 5099 6802 5133
rect 6836 5099 6846 5133
rect 6792 5065 6846 5099
rect 6792 5031 6802 5065
rect 6836 5031 6846 5065
rect 6792 4995 6846 5031
rect 6792 4961 6802 4995
rect 6836 4961 6846 4995
rect 6792 4945 6846 4961
rect 6876 5133 6930 5145
rect 6876 5099 6886 5133
rect 6920 5099 6930 5133
rect 6876 5065 6930 5099
rect 6876 5031 6886 5065
rect 6920 5031 6930 5065
rect 6876 4945 6930 5031
rect 6960 5133 7014 5145
rect 6960 5099 6970 5133
rect 7004 5099 7014 5133
rect 6960 5065 7014 5099
rect 6960 5031 6970 5065
rect 7004 5031 7014 5065
rect 6960 4995 7014 5031
rect 6960 4961 6970 4995
rect 7004 4961 7014 4995
rect 6960 4945 7014 4961
rect 7044 5133 7096 5145
rect 7044 5099 7054 5133
rect 7088 5099 7096 5133
rect 7044 5065 7096 5099
rect 7044 5031 7054 5065
rect 7088 5031 7096 5065
rect 7044 4995 7096 5031
rect 7044 4961 7054 4995
rect 7088 4961 7096 4995
rect 7044 4945 7096 4961
rect 7584 5131 7636 5143
rect 7584 5097 7592 5131
rect 7626 5097 7636 5131
rect 7584 5063 7636 5097
rect 7584 5029 7592 5063
rect 7626 5029 7636 5063
rect 7584 4943 7636 5029
rect 7666 5131 7720 5143
rect 7666 5097 7676 5131
rect 7710 5097 7720 5131
rect 7666 5063 7720 5097
rect 7666 5029 7676 5063
rect 7710 5029 7720 5063
rect 7666 4993 7720 5029
rect 7666 4959 7676 4993
rect 7710 4959 7720 4993
rect 7666 4943 7720 4959
rect 7750 5131 7804 5143
rect 7750 5097 7760 5131
rect 7794 5097 7804 5131
rect 7750 5063 7804 5097
rect 7750 5029 7760 5063
rect 7794 5029 7804 5063
rect 7750 4943 7804 5029
rect 7834 5131 7888 5143
rect 7834 5097 7844 5131
rect 7878 5097 7888 5131
rect 7834 5063 7888 5097
rect 7834 5029 7844 5063
rect 7878 5029 7888 5063
rect 7834 4993 7888 5029
rect 7834 4959 7844 4993
rect 7878 4959 7888 4993
rect 7834 4943 7888 4959
rect 7918 5131 7972 5143
rect 7918 5097 7928 5131
rect 7962 5097 7972 5131
rect 7918 5063 7972 5097
rect 7918 5029 7928 5063
rect 7962 5029 7972 5063
rect 7918 4943 7972 5029
rect 8002 5131 8056 5143
rect 8002 5097 8012 5131
rect 8046 5097 8056 5131
rect 8002 5063 8056 5097
rect 8002 5029 8012 5063
rect 8046 5029 8056 5063
rect 8002 4993 8056 5029
rect 8002 4959 8012 4993
rect 8046 4959 8056 4993
rect 8002 4943 8056 4959
rect 8086 5131 8140 5143
rect 8086 5097 8096 5131
rect 8130 5097 8140 5131
rect 8086 5063 8140 5097
rect 8086 5029 8096 5063
rect 8130 5029 8140 5063
rect 8086 4943 8140 5029
rect 8170 5131 8224 5143
rect 8170 5097 8180 5131
rect 8214 5097 8224 5131
rect 8170 5063 8224 5097
rect 8170 5029 8180 5063
rect 8214 5029 8224 5063
rect 8170 4993 8224 5029
rect 8170 4959 8180 4993
rect 8214 4959 8224 4993
rect 8170 4943 8224 4959
rect 8254 5131 8308 5143
rect 8254 5097 8264 5131
rect 8298 5097 8308 5131
rect 8254 5063 8308 5097
rect 8254 5029 8264 5063
rect 8298 5029 8308 5063
rect 8254 4943 8308 5029
rect 8338 5131 8392 5143
rect 8338 5097 8348 5131
rect 8382 5097 8392 5131
rect 8338 5063 8392 5097
rect 8338 5029 8348 5063
rect 8382 5029 8392 5063
rect 8338 4993 8392 5029
rect 8338 4959 8348 4993
rect 8382 4959 8392 4993
rect 8338 4943 8392 4959
rect 8422 5131 8476 5143
rect 8422 5097 8432 5131
rect 8466 5097 8476 5131
rect 8422 5063 8476 5097
rect 8422 5029 8432 5063
rect 8466 5029 8476 5063
rect 8422 4943 8476 5029
rect 8506 5131 8560 5143
rect 8506 5097 8516 5131
rect 8550 5097 8560 5131
rect 8506 5063 8560 5097
rect 8506 5029 8516 5063
rect 8550 5029 8560 5063
rect 8506 4993 8560 5029
rect 8506 4959 8516 4993
rect 8550 4959 8560 4993
rect 8506 4943 8560 4959
rect 8590 5131 8644 5143
rect 8590 5097 8600 5131
rect 8634 5097 8644 5131
rect 8590 5063 8644 5097
rect 8590 5029 8600 5063
rect 8634 5029 8644 5063
rect 8590 4943 8644 5029
rect 8674 5131 8728 5143
rect 8674 5097 8684 5131
rect 8718 5097 8728 5131
rect 8674 5063 8728 5097
rect 8674 5029 8684 5063
rect 8718 5029 8728 5063
rect 8674 4993 8728 5029
rect 8674 4959 8684 4993
rect 8718 4959 8728 4993
rect 8674 4943 8728 4959
rect 8758 5131 8812 5143
rect 8758 5097 8768 5131
rect 8802 5097 8812 5131
rect 8758 5063 8812 5097
rect 8758 5029 8768 5063
rect 8802 5029 8812 5063
rect 8758 4943 8812 5029
rect 8842 5131 8896 5143
rect 8842 5097 8852 5131
rect 8886 5097 8896 5131
rect 8842 5063 8896 5097
rect 8842 5029 8852 5063
rect 8886 5029 8896 5063
rect 8842 4993 8896 5029
rect 8842 4959 8852 4993
rect 8886 4959 8896 4993
rect 8842 4943 8896 4959
rect 8926 5131 8978 5143
rect 8926 5097 8936 5131
rect 8970 5097 8978 5131
rect 8926 5063 8978 5097
rect 8926 5029 8936 5063
rect 8970 5029 8978 5063
rect 8926 4993 8978 5029
rect 8926 4959 8936 4993
rect 8970 4959 8978 4993
rect 8926 4943 8978 4959
rect 20800 5133 20852 5145
rect 20800 5099 20808 5133
rect 20842 5099 20852 5133
rect 20800 5065 20852 5099
rect 20800 5031 20808 5065
rect 20842 5031 20852 5065
rect 20800 4945 20852 5031
rect 20882 5133 20936 5145
rect 20882 5099 20892 5133
rect 20926 5099 20936 5133
rect 20882 5065 20936 5099
rect 20882 5031 20892 5065
rect 20926 5031 20936 5065
rect 20882 4995 20936 5031
rect 20882 4961 20892 4995
rect 20926 4961 20936 4995
rect 20882 4945 20936 4961
rect 20966 5133 21020 5145
rect 20966 5099 20976 5133
rect 21010 5099 21020 5133
rect 20966 5065 21020 5099
rect 20966 5031 20976 5065
rect 21010 5031 21020 5065
rect 20966 4945 21020 5031
rect 21050 5133 21104 5145
rect 21050 5099 21060 5133
rect 21094 5099 21104 5133
rect 21050 5065 21104 5099
rect 21050 5031 21060 5065
rect 21094 5031 21104 5065
rect 21050 4995 21104 5031
rect 21050 4961 21060 4995
rect 21094 4961 21104 4995
rect 21050 4945 21104 4961
rect 21134 5133 21188 5145
rect 21134 5099 21144 5133
rect 21178 5099 21188 5133
rect 21134 5065 21188 5099
rect 21134 5031 21144 5065
rect 21178 5031 21188 5065
rect 21134 4945 21188 5031
rect 21218 5133 21272 5145
rect 21218 5099 21228 5133
rect 21262 5099 21272 5133
rect 21218 5065 21272 5099
rect 21218 5031 21228 5065
rect 21262 5031 21272 5065
rect 21218 4995 21272 5031
rect 21218 4961 21228 4995
rect 21262 4961 21272 4995
rect 21218 4945 21272 4961
rect 21302 5133 21356 5145
rect 21302 5099 21312 5133
rect 21346 5099 21356 5133
rect 21302 5065 21356 5099
rect 21302 5031 21312 5065
rect 21346 5031 21356 5065
rect 21302 4945 21356 5031
rect 21386 5133 21440 5145
rect 21386 5099 21396 5133
rect 21430 5099 21440 5133
rect 21386 5065 21440 5099
rect 21386 5031 21396 5065
rect 21430 5031 21440 5065
rect 21386 4995 21440 5031
rect 21386 4961 21396 4995
rect 21430 4961 21440 4995
rect 21386 4945 21440 4961
rect 21470 5133 21524 5145
rect 21470 5099 21480 5133
rect 21514 5099 21524 5133
rect 21470 5065 21524 5099
rect 21470 5031 21480 5065
rect 21514 5031 21524 5065
rect 21470 4945 21524 5031
rect 21554 5133 21608 5145
rect 21554 5099 21564 5133
rect 21598 5099 21608 5133
rect 21554 5065 21608 5099
rect 21554 5031 21564 5065
rect 21598 5031 21608 5065
rect 21554 4995 21608 5031
rect 21554 4961 21564 4995
rect 21598 4961 21608 4995
rect 21554 4945 21608 4961
rect 21638 5133 21692 5145
rect 21638 5099 21648 5133
rect 21682 5099 21692 5133
rect 21638 5065 21692 5099
rect 21638 5031 21648 5065
rect 21682 5031 21692 5065
rect 21638 4945 21692 5031
rect 21722 5133 21776 5145
rect 21722 5099 21732 5133
rect 21766 5099 21776 5133
rect 21722 5065 21776 5099
rect 21722 5031 21732 5065
rect 21766 5031 21776 5065
rect 21722 4995 21776 5031
rect 21722 4961 21732 4995
rect 21766 4961 21776 4995
rect 21722 4945 21776 4961
rect 21806 5133 21860 5145
rect 21806 5099 21816 5133
rect 21850 5099 21860 5133
rect 21806 5065 21860 5099
rect 21806 5031 21816 5065
rect 21850 5031 21860 5065
rect 21806 4945 21860 5031
rect 21890 5133 21944 5145
rect 21890 5099 21900 5133
rect 21934 5099 21944 5133
rect 21890 5065 21944 5099
rect 21890 5031 21900 5065
rect 21934 5031 21944 5065
rect 21890 4995 21944 5031
rect 21890 4961 21900 4995
rect 21934 4961 21944 4995
rect 21890 4945 21944 4961
rect 21974 5133 22028 5145
rect 21974 5099 21984 5133
rect 22018 5099 22028 5133
rect 21974 5065 22028 5099
rect 21974 5031 21984 5065
rect 22018 5031 22028 5065
rect 21974 4945 22028 5031
rect 22058 5133 22112 5145
rect 22058 5099 22068 5133
rect 22102 5099 22112 5133
rect 22058 5065 22112 5099
rect 22058 5031 22068 5065
rect 22102 5031 22112 5065
rect 22058 4995 22112 5031
rect 22058 4961 22068 4995
rect 22102 4961 22112 4995
rect 22058 4945 22112 4961
rect 22142 5133 22194 5145
rect 22142 5099 22152 5133
rect 22186 5099 22194 5133
rect 22142 5065 22194 5099
rect 22142 5031 22152 5065
rect 22186 5031 22194 5065
rect 22142 4995 22194 5031
rect 22142 4961 22152 4995
rect 22186 4961 22194 4995
rect 22142 4945 22194 4961
rect 22682 5131 22734 5143
rect 22682 5097 22690 5131
rect 22724 5097 22734 5131
rect 22682 5063 22734 5097
rect 22682 5029 22690 5063
rect 22724 5029 22734 5063
rect 22682 4943 22734 5029
rect 22764 5131 22818 5143
rect 22764 5097 22774 5131
rect 22808 5097 22818 5131
rect 22764 5063 22818 5097
rect 22764 5029 22774 5063
rect 22808 5029 22818 5063
rect 22764 4993 22818 5029
rect 22764 4959 22774 4993
rect 22808 4959 22818 4993
rect 22764 4943 22818 4959
rect 22848 5131 22902 5143
rect 22848 5097 22858 5131
rect 22892 5097 22902 5131
rect 22848 5063 22902 5097
rect 22848 5029 22858 5063
rect 22892 5029 22902 5063
rect 22848 4943 22902 5029
rect 22932 5131 22986 5143
rect 22932 5097 22942 5131
rect 22976 5097 22986 5131
rect 22932 5063 22986 5097
rect 22932 5029 22942 5063
rect 22976 5029 22986 5063
rect 22932 4993 22986 5029
rect 22932 4959 22942 4993
rect 22976 4959 22986 4993
rect 22932 4943 22986 4959
rect 23016 5131 23070 5143
rect 23016 5097 23026 5131
rect 23060 5097 23070 5131
rect 23016 5063 23070 5097
rect 23016 5029 23026 5063
rect 23060 5029 23070 5063
rect 23016 4943 23070 5029
rect 23100 5131 23154 5143
rect 23100 5097 23110 5131
rect 23144 5097 23154 5131
rect 23100 5063 23154 5097
rect 23100 5029 23110 5063
rect 23144 5029 23154 5063
rect 23100 4993 23154 5029
rect 23100 4959 23110 4993
rect 23144 4959 23154 4993
rect 23100 4943 23154 4959
rect 23184 5131 23238 5143
rect 23184 5097 23194 5131
rect 23228 5097 23238 5131
rect 23184 5063 23238 5097
rect 23184 5029 23194 5063
rect 23228 5029 23238 5063
rect 23184 4943 23238 5029
rect 23268 5131 23322 5143
rect 23268 5097 23278 5131
rect 23312 5097 23322 5131
rect 23268 5063 23322 5097
rect 23268 5029 23278 5063
rect 23312 5029 23322 5063
rect 23268 4993 23322 5029
rect 23268 4959 23278 4993
rect 23312 4959 23322 4993
rect 23268 4943 23322 4959
rect 23352 5131 23406 5143
rect 23352 5097 23362 5131
rect 23396 5097 23406 5131
rect 23352 5063 23406 5097
rect 23352 5029 23362 5063
rect 23396 5029 23406 5063
rect 23352 4943 23406 5029
rect 23436 5131 23490 5143
rect 23436 5097 23446 5131
rect 23480 5097 23490 5131
rect 23436 5063 23490 5097
rect 23436 5029 23446 5063
rect 23480 5029 23490 5063
rect 23436 4993 23490 5029
rect 23436 4959 23446 4993
rect 23480 4959 23490 4993
rect 23436 4943 23490 4959
rect 23520 5131 23574 5143
rect 23520 5097 23530 5131
rect 23564 5097 23574 5131
rect 23520 5063 23574 5097
rect 23520 5029 23530 5063
rect 23564 5029 23574 5063
rect 23520 4943 23574 5029
rect 23604 5131 23658 5143
rect 23604 5097 23614 5131
rect 23648 5097 23658 5131
rect 23604 5063 23658 5097
rect 23604 5029 23614 5063
rect 23648 5029 23658 5063
rect 23604 4993 23658 5029
rect 23604 4959 23614 4993
rect 23648 4959 23658 4993
rect 23604 4943 23658 4959
rect 23688 5131 23742 5143
rect 23688 5097 23698 5131
rect 23732 5097 23742 5131
rect 23688 5063 23742 5097
rect 23688 5029 23698 5063
rect 23732 5029 23742 5063
rect 23688 4943 23742 5029
rect 23772 5131 23826 5143
rect 23772 5097 23782 5131
rect 23816 5097 23826 5131
rect 23772 5063 23826 5097
rect 23772 5029 23782 5063
rect 23816 5029 23826 5063
rect 23772 4993 23826 5029
rect 23772 4959 23782 4993
rect 23816 4959 23826 4993
rect 23772 4943 23826 4959
rect 23856 5131 23910 5143
rect 23856 5097 23866 5131
rect 23900 5097 23910 5131
rect 23856 5063 23910 5097
rect 23856 5029 23866 5063
rect 23900 5029 23910 5063
rect 23856 4943 23910 5029
rect 23940 5131 23994 5143
rect 23940 5097 23950 5131
rect 23984 5097 23994 5131
rect 23940 5063 23994 5097
rect 23940 5029 23950 5063
rect 23984 5029 23994 5063
rect 23940 4993 23994 5029
rect 23940 4959 23950 4993
rect 23984 4959 23994 4993
rect 23940 4943 23994 4959
rect 24024 5131 24076 5143
rect 24024 5097 24034 5131
rect 24068 5097 24076 5131
rect 24024 5063 24076 5097
rect 24024 5029 24034 5063
rect 24068 5029 24076 5063
rect 24024 4993 24076 5029
rect 24024 4959 24034 4993
rect 24068 4959 24076 4993
rect 24024 4943 24076 4959
rect 35904 5133 35956 5145
rect 35904 5099 35912 5133
rect 35946 5099 35956 5133
rect 35904 5065 35956 5099
rect 35904 5031 35912 5065
rect 35946 5031 35956 5065
rect 35904 4945 35956 5031
rect 35986 5133 36040 5145
rect 35986 5099 35996 5133
rect 36030 5099 36040 5133
rect 35986 5065 36040 5099
rect 35986 5031 35996 5065
rect 36030 5031 36040 5065
rect 35986 4995 36040 5031
rect 35986 4961 35996 4995
rect 36030 4961 36040 4995
rect 35986 4945 36040 4961
rect 36070 5133 36124 5145
rect 36070 5099 36080 5133
rect 36114 5099 36124 5133
rect 36070 5065 36124 5099
rect 36070 5031 36080 5065
rect 36114 5031 36124 5065
rect 36070 4945 36124 5031
rect 36154 5133 36208 5145
rect 36154 5099 36164 5133
rect 36198 5099 36208 5133
rect 36154 5065 36208 5099
rect 36154 5031 36164 5065
rect 36198 5031 36208 5065
rect 36154 4995 36208 5031
rect 36154 4961 36164 4995
rect 36198 4961 36208 4995
rect 36154 4945 36208 4961
rect 36238 5133 36292 5145
rect 36238 5099 36248 5133
rect 36282 5099 36292 5133
rect 36238 5065 36292 5099
rect 36238 5031 36248 5065
rect 36282 5031 36292 5065
rect 36238 4945 36292 5031
rect 36322 5133 36376 5145
rect 36322 5099 36332 5133
rect 36366 5099 36376 5133
rect 36322 5065 36376 5099
rect 36322 5031 36332 5065
rect 36366 5031 36376 5065
rect 36322 4995 36376 5031
rect 36322 4961 36332 4995
rect 36366 4961 36376 4995
rect 36322 4945 36376 4961
rect 36406 5133 36460 5145
rect 36406 5099 36416 5133
rect 36450 5099 36460 5133
rect 36406 5065 36460 5099
rect 36406 5031 36416 5065
rect 36450 5031 36460 5065
rect 36406 4945 36460 5031
rect 36490 5133 36544 5145
rect 36490 5099 36500 5133
rect 36534 5099 36544 5133
rect 36490 5065 36544 5099
rect 36490 5031 36500 5065
rect 36534 5031 36544 5065
rect 36490 4995 36544 5031
rect 36490 4961 36500 4995
rect 36534 4961 36544 4995
rect 36490 4945 36544 4961
rect 36574 5133 36628 5145
rect 36574 5099 36584 5133
rect 36618 5099 36628 5133
rect 36574 5065 36628 5099
rect 36574 5031 36584 5065
rect 36618 5031 36628 5065
rect 36574 4945 36628 5031
rect 36658 5133 36712 5145
rect 36658 5099 36668 5133
rect 36702 5099 36712 5133
rect 36658 5065 36712 5099
rect 36658 5031 36668 5065
rect 36702 5031 36712 5065
rect 36658 4995 36712 5031
rect 36658 4961 36668 4995
rect 36702 4961 36712 4995
rect 36658 4945 36712 4961
rect 36742 5133 36796 5145
rect 36742 5099 36752 5133
rect 36786 5099 36796 5133
rect 36742 5065 36796 5099
rect 36742 5031 36752 5065
rect 36786 5031 36796 5065
rect 36742 4945 36796 5031
rect 36826 5133 36880 5145
rect 36826 5099 36836 5133
rect 36870 5099 36880 5133
rect 36826 5065 36880 5099
rect 36826 5031 36836 5065
rect 36870 5031 36880 5065
rect 36826 4995 36880 5031
rect 36826 4961 36836 4995
rect 36870 4961 36880 4995
rect 36826 4945 36880 4961
rect 36910 5133 36964 5145
rect 36910 5099 36920 5133
rect 36954 5099 36964 5133
rect 36910 5065 36964 5099
rect 36910 5031 36920 5065
rect 36954 5031 36964 5065
rect 36910 4945 36964 5031
rect 36994 5133 37048 5145
rect 36994 5099 37004 5133
rect 37038 5099 37048 5133
rect 36994 5065 37048 5099
rect 36994 5031 37004 5065
rect 37038 5031 37048 5065
rect 36994 4995 37048 5031
rect 36994 4961 37004 4995
rect 37038 4961 37048 4995
rect 36994 4945 37048 4961
rect 37078 5133 37132 5145
rect 37078 5099 37088 5133
rect 37122 5099 37132 5133
rect 37078 5065 37132 5099
rect 37078 5031 37088 5065
rect 37122 5031 37132 5065
rect 37078 4945 37132 5031
rect 37162 5133 37216 5145
rect 37162 5099 37172 5133
rect 37206 5099 37216 5133
rect 37162 5065 37216 5099
rect 37162 5031 37172 5065
rect 37206 5031 37216 5065
rect 37162 4995 37216 5031
rect 37162 4961 37172 4995
rect 37206 4961 37216 4995
rect 37162 4945 37216 4961
rect 37246 5133 37298 5145
rect 37246 5099 37256 5133
rect 37290 5099 37298 5133
rect 37246 5065 37298 5099
rect 37246 5031 37256 5065
rect 37290 5031 37298 5065
rect 37246 4995 37298 5031
rect 37246 4961 37256 4995
rect 37290 4961 37298 4995
rect 37246 4945 37298 4961
rect 37786 5131 37838 5143
rect 37786 5097 37794 5131
rect 37828 5097 37838 5131
rect 37786 5063 37838 5097
rect 37786 5029 37794 5063
rect 37828 5029 37838 5063
rect 37786 4943 37838 5029
rect 37868 5131 37922 5143
rect 37868 5097 37878 5131
rect 37912 5097 37922 5131
rect 37868 5063 37922 5097
rect 37868 5029 37878 5063
rect 37912 5029 37922 5063
rect 37868 4993 37922 5029
rect 37868 4959 37878 4993
rect 37912 4959 37922 4993
rect 37868 4943 37922 4959
rect 37952 5131 38006 5143
rect 37952 5097 37962 5131
rect 37996 5097 38006 5131
rect 37952 5063 38006 5097
rect 37952 5029 37962 5063
rect 37996 5029 38006 5063
rect 37952 4943 38006 5029
rect 38036 5131 38090 5143
rect 38036 5097 38046 5131
rect 38080 5097 38090 5131
rect 38036 5063 38090 5097
rect 38036 5029 38046 5063
rect 38080 5029 38090 5063
rect 38036 4993 38090 5029
rect 38036 4959 38046 4993
rect 38080 4959 38090 4993
rect 38036 4943 38090 4959
rect 38120 5131 38174 5143
rect 38120 5097 38130 5131
rect 38164 5097 38174 5131
rect 38120 5063 38174 5097
rect 38120 5029 38130 5063
rect 38164 5029 38174 5063
rect 38120 4943 38174 5029
rect 38204 5131 38258 5143
rect 38204 5097 38214 5131
rect 38248 5097 38258 5131
rect 38204 5063 38258 5097
rect 38204 5029 38214 5063
rect 38248 5029 38258 5063
rect 38204 4993 38258 5029
rect 38204 4959 38214 4993
rect 38248 4959 38258 4993
rect 38204 4943 38258 4959
rect 38288 5131 38342 5143
rect 38288 5097 38298 5131
rect 38332 5097 38342 5131
rect 38288 5063 38342 5097
rect 38288 5029 38298 5063
rect 38332 5029 38342 5063
rect 38288 4943 38342 5029
rect 38372 5131 38426 5143
rect 38372 5097 38382 5131
rect 38416 5097 38426 5131
rect 38372 5063 38426 5097
rect 38372 5029 38382 5063
rect 38416 5029 38426 5063
rect 38372 4993 38426 5029
rect 38372 4959 38382 4993
rect 38416 4959 38426 4993
rect 38372 4943 38426 4959
rect 38456 5131 38510 5143
rect 38456 5097 38466 5131
rect 38500 5097 38510 5131
rect 38456 5063 38510 5097
rect 38456 5029 38466 5063
rect 38500 5029 38510 5063
rect 38456 4943 38510 5029
rect 38540 5131 38594 5143
rect 38540 5097 38550 5131
rect 38584 5097 38594 5131
rect 38540 5063 38594 5097
rect 38540 5029 38550 5063
rect 38584 5029 38594 5063
rect 38540 4993 38594 5029
rect 38540 4959 38550 4993
rect 38584 4959 38594 4993
rect 38540 4943 38594 4959
rect 38624 5131 38678 5143
rect 38624 5097 38634 5131
rect 38668 5097 38678 5131
rect 38624 5063 38678 5097
rect 38624 5029 38634 5063
rect 38668 5029 38678 5063
rect 38624 4943 38678 5029
rect 38708 5131 38762 5143
rect 38708 5097 38718 5131
rect 38752 5097 38762 5131
rect 38708 5063 38762 5097
rect 38708 5029 38718 5063
rect 38752 5029 38762 5063
rect 38708 4993 38762 5029
rect 38708 4959 38718 4993
rect 38752 4959 38762 4993
rect 38708 4943 38762 4959
rect 38792 5131 38846 5143
rect 38792 5097 38802 5131
rect 38836 5097 38846 5131
rect 38792 5063 38846 5097
rect 38792 5029 38802 5063
rect 38836 5029 38846 5063
rect 38792 4943 38846 5029
rect 38876 5131 38930 5143
rect 38876 5097 38886 5131
rect 38920 5097 38930 5131
rect 38876 5063 38930 5097
rect 38876 5029 38886 5063
rect 38920 5029 38930 5063
rect 38876 4993 38930 5029
rect 38876 4959 38886 4993
rect 38920 4959 38930 4993
rect 38876 4943 38930 4959
rect 38960 5131 39014 5143
rect 38960 5097 38970 5131
rect 39004 5097 39014 5131
rect 38960 5063 39014 5097
rect 38960 5029 38970 5063
rect 39004 5029 39014 5063
rect 38960 4943 39014 5029
rect 39044 5131 39098 5143
rect 39044 5097 39054 5131
rect 39088 5097 39098 5131
rect 39044 5063 39098 5097
rect 39044 5029 39054 5063
rect 39088 5029 39098 5063
rect 39044 4993 39098 5029
rect 39044 4959 39054 4993
rect 39088 4959 39098 4993
rect 39044 4943 39098 4959
rect 39128 5131 39180 5143
rect 39128 5097 39138 5131
rect 39172 5097 39180 5131
rect 39128 5063 39180 5097
rect 39128 5029 39138 5063
rect 39172 5029 39180 5063
rect 39128 4993 39180 5029
rect 39128 4959 39138 4993
rect 39172 4959 39180 4993
rect 39128 4943 39180 4959
rect 51002 5133 51054 5145
rect 51002 5099 51010 5133
rect 51044 5099 51054 5133
rect 51002 5065 51054 5099
rect 51002 5031 51010 5065
rect 51044 5031 51054 5065
rect 51002 4945 51054 5031
rect 51084 5133 51138 5145
rect 51084 5099 51094 5133
rect 51128 5099 51138 5133
rect 51084 5065 51138 5099
rect 51084 5031 51094 5065
rect 51128 5031 51138 5065
rect 51084 4995 51138 5031
rect 51084 4961 51094 4995
rect 51128 4961 51138 4995
rect 51084 4945 51138 4961
rect 51168 5133 51222 5145
rect 51168 5099 51178 5133
rect 51212 5099 51222 5133
rect 51168 5065 51222 5099
rect 51168 5031 51178 5065
rect 51212 5031 51222 5065
rect 51168 4945 51222 5031
rect 51252 5133 51306 5145
rect 51252 5099 51262 5133
rect 51296 5099 51306 5133
rect 51252 5065 51306 5099
rect 51252 5031 51262 5065
rect 51296 5031 51306 5065
rect 51252 4995 51306 5031
rect 51252 4961 51262 4995
rect 51296 4961 51306 4995
rect 51252 4945 51306 4961
rect 51336 5133 51390 5145
rect 51336 5099 51346 5133
rect 51380 5099 51390 5133
rect 51336 5065 51390 5099
rect 51336 5031 51346 5065
rect 51380 5031 51390 5065
rect 51336 4945 51390 5031
rect 51420 5133 51474 5145
rect 51420 5099 51430 5133
rect 51464 5099 51474 5133
rect 51420 5065 51474 5099
rect 51420 5031 51430 5065
rect 51464 5031 51474 5065
rect 51420 4995 51474 5031
rect 51420 4961 51430 4995
rect 51464 4961 51474 4995
rect 51420 4945 51474 4961
rect 51504 5133 51558 5145
rect 51504 5099 51514 5133
rect 51548 5099 51558 5133
rect 51504 5065 51558 5099
rect 51504 5031 51514 5065
rect 51548 5031 51558 5065
rect 51504 4945 51558 5031
rect 51588 5133 51642 5145
rect 51588 5099 51598 5133
rect 51632 5099 51642 5133
rect 51588 5065 51642 5099
rect 51588 5031 51598 5065
rect 51632 5031 51642 5065
rect 51588 4995 51642 5031
rect 51588 4961 51598 4995
rect 51632 4961 51642 4995
rect 51588 4945 51642 4961
rect 51672 5133 51726 5145
rect 51672 5099 51682 5133
rect 51716 5099 51726 5133
rect 51672 5065 51726 5099
rect 51672 5031 51682 5065
rect 51716 5031 51726 5065
rect 51672 4945 51726 5031
rect 51756 5133 51810 5145
rect 51756 5099 51766 5133
rect 51800 5099 51810 5133
rect 51756 5065 51810 5099
rect 51756 5031 51766 5065
rect 51800 5031 51810 5065
rect 51756 4995 51810 5031
rect 51756 4961 51766 4995
rect 51800 4961 51810 4995
rect 51756 4945 51810 4961
rect 51840 5133 51894 5145
rect 51840 5099 51850 5133
rect 51884 5099 51894 5133
rect 51840 5065 51894 5099
rect 51840 5031 51850 5065
rect 51884 5031 51894 5065
rect 51840 4945 51894 5031
rect 51924 5133 51978 5145
rect 51924 5099 51934 5133
rect 51968 5099 51978 5133
rect 51924 5065 51978 5099
rect 51924 5031 51934 5065
rect 51968 5031 51978 5065
rect 51924 4995 51978 5031
rect 51924 4961 51934 4995
rect 51968 4961 51978 4995
rect 51924 4945 51978 4961
rect 52008 5133 52062 5145
rect 52008 5099 52018 5133
rect 52052 5099 52062 5133
rect 52008 5065 52062 5099
rect 52008 5031 52018 5065
rect 52052 5031 52062 5065
rect 52008 4945 52062 5031
rect 52092 5133 52146 5145
rect 52092 5099 52102 5133
rect 52136 5099 52146 5133
rect 52092 5065 52146 5099
rect 52092 5031 52102 5065
rect 52136 5031 52146 5065
rect 52092 4995 52146 5031
rect 52092 4961 52102 4995
rect 52136 4961 52146 4995
rect 52092 4945 52146 4961
rect 52176 5133 52230 5145
rect 52176 5099 52186 5133
rect 52220 5099 52230 5133
rect 52176 5065 52230 5099
rect 52176 5031 52186 5065
rect 52220 5031 52230 5065
rect 52176 4945 52230 5031
rect 52260 5133 52314 5145
rect 52260 5099 52270 5133
rect 52304 5099 52314 5133
rect 52260 5065 52314 5099
rect 52260 5031 52270 5065
rect 52304 5031 52314 5065
rect 52260 4995 52314 5031
rect 52260 4961 52270 4995
rect 52304 4961 52314 4995
rect 52260 4945 52314 4961
rect 52344 5133 52396 5145
rect 52344 5099 52354 5133
rect 52388 5099 52396 5133
rect 52344 5065 52396 5099
rect 52344 5031 52354 5065
rect 52388 5031 52396 5065
rect 52344 4995 52396 5031
rect 52344 4961 52354 4995
rect 52388 4961 52396 4995
rect 52344 4945 52396 4961
rect 52884 5131 52936 5143
rect 52884 5097 52892 5131
rect 52926 5097 52936 5131
rect 52884 5063 52936 5097
rect 52884 5029 52892 5063
rect 52926 5029 52936 5063
rect 52884 4943 52936 5029
rect 52966 5131 53020 5143
rect 52966 5097 52976 5131
rect 53010 5097 53020 5131
rect 52966 5063 53020 5097
rect 52966 5029 52976 5063
rect 53010 5029 53020 5063
rect 52966 4993 53020 5029
rect 52966 4959 52976 4993
rect 53010 4959 53020 4993
rect 52966 4943 53020 4959
rect 53050 5131 53104 5143
rect 53050 5097 53060 5131
rect 53094 5097 53104 5131
rect 53050 5063 53104 5097
rect 53050 5029 53060 5063
rect 53094 5029 53104 5063
rect 53050 4943 53104 5029
rect 53134 5131 53188 5143
rect 53134 5097 53144 5131
rect 53178 5097 53188 5131
rect 53134 5063 53188 5097
rect 53134 5029 53144 5063
rect 53178 5029 53188 5063
rect 53134 4993 53188 5029
rect 53134 4959 53144 4993
rect 53178 4959 53188 4993
rect 53134 4943 53188 4959
rect 53218 5131 53272 5143
rect 53218 5097 53228 5131
rect 53262 5097 53272 5131
rect 53218 5063 53272 5097
rect 53218 5029 53228 5063
rect 53262 5029 53272 5063
rect 53218 4943 53272 5029
rect 53302 5131 53356 5143
rect 53302 5097 53312 5131
rect 53346 5097 53356 5131
rect 53302 5063 53356 5097
rect 53302 5029 53312 5063
rect 53346 5029 53356 5063
rect 53302 4993 53356 5029
rect 53302 4959 53312 4993
rect 53346 4959 53356 4993
rect 53302 4943 53356 4959
rect 53386 5131 53440 5143
rect 53386 5097 53396 5131
rect 53430 5097 53440 5131
rect 53386 5063 53440 5097
rect 53386 5029 53396 5063
rect 53430 5029 53440 5063
rect 53386 4943 53440 5029
rect 53470 5131 53524 5143
rect 53470 5097 53480 5131
rect 53514 5097 53524 5131
rect 53470 5063 53524 5097
rect 53470 5029 53480 5063
rect 53514 5029 53524 5063
rect 53470 4993 53524 5029
rect 53470 4959 53480 4993
rect 53514 4959 53524 4993
rect 53470 4943 53524 4959
rect 53554 5131 53608 5143
rect 53554 5097 53564 5131
rect 53598 5097 53608 5131
rect 53554 5063 53608 5097
rect 53554 5029 53564 5063
rect 53598 5029 53608 5063
rect 53554 4943 53608 5029
rect 53638 5131 53692 5143
rect 53638 5097 53648 5131
rect 53682 5097 53692 5131
rect 53638 5063 53692 5097
rect 53638 5029 53648 5063
rect 53682 5029 53692 5063
rect 53638 4993 53692 5029
rect 53638 4959 53648 4993
rect 53682 4959 53692 4993
rect 53638 4943 53692 4959
rect 53722 5131 53776 5143
rect 53722 5097 53732 5131
rect 53766 5097 53776 5131
rect 53722 5063 53776 5097
rect 53722 5029 53732 5063
rect 53766 5029 53776 5063
rect 53722 4943 53776 5029
rect 53806 5131 53860 5143
rect 53806 5097 53816 5131
rect 53850 5097 53860 5131
rect 53806 5063 53860 5097
rect 53806 5029 53816 5063
rect 53850 5029 53860 5063
rect 53806 4993 53860 5029
rect 53806 4959 53816 4993
rect 53850 4959 53860 4993
rect 53806 4943 53860 4959
rect 53890 5131 53944 5143
rect 53890 5097 53900 5131
rect 53934 5097 53944 5131
rect 53890 5063 53944 5097
rect 53890 5029 53900 5063
rect 53934 5029 53944 5063
rect 53890 4943 53944 5029
rect 53974 5131 54028 5143
rect 53974 5097 53984 5131
rect 54018 5097 54028 5131
rect 53974 5063 54028 5097
rect 53974 5029 53984 5063
rect 54018 5029 54028 5063
rect 53974 4993 54028 5029
rect 53974 4959 53984 4993
rect 54018 4959 54028 4993
rect 53974 4943 54028 4959
rect 54058 5131 54112 5143
rect 54058 5097 54068 5131
rect 54102 5097 54112 5131
rect 54058 5063 54112 5097
rect 54058 5029 54068 5063
rect 54102 5029 54112 5063
rect 54058 4943 54112 5029
rect 54142 5131 54196 5143
rect 54142 5097 54152 5131
rect 54186 5097 54196 5131
rect 54142 5063 54196 5097
rect 54142 5029 54152 5063
rect 54186 5029 54196 5063
rect 54142 4993 54196 5029
rect 54142 4959 54152 4993
rect 54186 4959 54196 4993
rect 54142 4943 54196 4959
rect 54226 5131 54278 5143
rect 54226 5097 54236 5131
rect 54270 5097 54278 5131
rect 54226 5063 54278 5097
rect 54226 5029 54236 5063
rect 54270 5029 54278 5063
rect 54226 4993 54278 5029
rect 54226 4959 54236 4993
rect 54270 4959 54278 4993
rect 54226 4943 54278 4959
rect 30064 4056 30116 4068
rect 30064 4022 30072 4056
rect 30106 4022 30116 4056
rect 30064 3988 30116 4022
rect 30064 3954 30072 3988
rect 30106 3954 30116 3988
rect 30064 3920 30116 3954
rect 30064 3886 30072 3920
rect 30106 3886 30116 3920
rect 30064 3868 30116 3886
rect 30146 4056 30200 4068
rect 30146 4022 30156 4056
rect 30190 4022 30200 4056
rect 30146 3988 30200 4022
rect 30146 3954 30156 3988
rect 30190 3954 30200 3988
rect 30146 3920 30200 3954
rect 30146 3886 30156 3920
rect 30190 3886 30200 3920
rect 30146 3868 30200 3886
rect 30230 4056 30284 4068
rect 30230 4022 30240 4056
rect 30274 4022 30284 4056
rect 30230 3988 30284 4022
rect 30230 3954 30240 3988
rect 30274 3954 30284 3988
rect 30230 3868 30284 3954
rect 30314 4056 30368 4068
rect 30314 4022 30324 4056
rect 30358 4022 30368 4056
rect 30314 3988 30368 4022
rect 30314 3954 30324 3988
rect 30358 3954 30368 3988
rect 30314 3920 30368 3954
rect 30314 3886 30324 3920
rect 30358 3886 30368 3920
rect 30314 3868 30368 3886
rect 30398 4056 30450 4068
rect 30398 4022 30408 4056
rect 30442 4022 30450 4056
rect 30398 3868 30450 4022
rect 30595 4056 30647 4068
rect 30595 4022 30603 4056
rect 30637 4022 30647 4056
rect 30595 3988 30647 4022
rect 30595 3954 30603 3988
rect 30637 3954 30647 3988
rect 30595 3918 30647 3954
rect 30595 3884 30603 3918
rect 30637 3884 30647 3918
rect 30595 3868 30647 3884
rect 30677 4056 30731 4068
rect 30677 4022 30687 4056
rect 30721 4022 30731 4056
rect 30677 3988 30731 4022
rect 30677 3954 30687 3988
rect 30721 3954 30731 3988
rect 30677 3918 30731 3954
rect 30677 3884 30687 3918
rect 30721 3884 30731 3918
rect 30677 3868 30731 3884
rect 30761 4056 30815 4068
rect 30761 4022 30771 4056
rect 30805 4022 30815 4056
rect 30761 3988 30815 4022
rect 30761 3954 30771 3988
rect 30805 3954 30815 3988
rect 30761 3868 30815 3954
rect 30845 4056 30899 4068
rect 30845 4022 30855 4056
rect 30889 4022 30899 4056
rect 30845 3988 30899 4022
rect 30845 3954 30855 3988
rect 30889 3954 30899 3988
rect 30845 3918 30899 3954
rect 30845 3884 30855 3918
rect 30889 3884 30899 3918
rect 30845 3868 30899 3884
rect 30929 4056 30983 4068
rect 30929 4022 30939 4056
rect 30973 4022 30983 4056
rect 30929 3988 30983 4022
rect 30929 3954 30939 3988
rect 30973 3954 30983 3988
rect 30929 3868 30983 3954
rect 31013 4056 31067 4068
rect 31013 4022 31023 4056
rect 31057 4022 31067 4056
rect 31013 3988 31067 4022
rect 31013 3954 31023 3988
rect 31057 3954 31067 3988
rect 31013 3918 31067 3954
rect 31013 3884 31023 3918
rect 31057 3884 31067 3918
rect 31013 3868 31067 3884
rect 31097 4056 31151 4068
rect 31097 4022 31107 4056
rect 31141 4022 31151 4056
rect 31097 3988 31151 4022
rect 31097 3954 31107 3988
rect 31141 3954 31151 3988
rect 31097 3868 31151 3954
rect 31181 4056 31235 4068
rect 31181 4022 31191 4056
rect 31225 4022 31235 4056
rect 31181 3988 31235 4022
rect 31181 3954 31191 3988
rect 31225 3954 31235 3988
rect 31181 3918 31235 3954
rect 31181 3884 31191 3918
rect 31225 3884 31235 3918
rect 31181 3868 31235 3884
rect 31265 4056 31319 4068
rect 31265 4022 31275 4056
rect 31309 4022 31319 4056
rect 31265 3988 31319 4022
rect 31265 3954 31275 3988
rect 31309 3954 31319 3988
rect 31265 3868 31319 3954
rect 31349 4056 31403 4068
rect 31349 4022 31359 4056
rect 31393 4022 31403 4056
rect 31349 3988 31403 4022
rect 31349 3954 31359 3988
rect 31393 3954 31403 3988
rect 31349 3918 31403 3954
rect 31349 3884 31359 3918
rect 31393 3884 31403 3918
rect 31349 3868 31403 3884
rect 31433 4056 31487 4068
rect 31433 4022 31443 4056
rect 31477 4022 31487 4056
rect 31433 3988 31487 4022
rect 31433 3954 31443 3988
rect 31477 3954 31487 3988
rect 31433 3868 31487 3954
rect 31517 4056 31571 4068
rect 31517 4022 31527 4056
rect 31561 4022 31571 4056
rect 31517 3988 31571 4022
rect 31517 3954 31527 3988
rect 31561 3954 31571 3988
rect 31517 3918 31571 3954
rect 31517 3884 31527 3918
rect 31561 3884 31571 3918
rect 31517 3868 31571 3884
rect 31601 4056 31655 4068
rect 31601 4022 31611 4056
rect 31645 4022 31655 4056
rect 31601 3988 31655 4022
rect 31601 3954 31611 3988
rect 31645 3954 31655 3988
rect 31601 3868 31655 3954
rect 31685 4056 31739 4068
rect 31685 4022 31695 4056
rect 31729 4022 31739 4056
rect 31685 3988 31739 4022
rect 31685 3954 31695 3988
rect 31729 3954 31739 3988
rect 31685 3918 31739 3954
rect 31685 3884 31695 3918
rect 31729 3884 31739 3918
rect 31685 3868 31739 3884
rect 31769 4056 31823 4068
rect 31769 4022 31779 4056
rect 31813 4022 31823 4056
rect 31769 3988 31823 4022
rect 31769 3954 31779 3988
rect 31813 3954 31823 3988
rect 31769 3868 31823 3954
rect 31853 4056 31907 4068
rect 31853 4022 31863 4056
rect 31897 4022 31907 4056
rect 31853 3988 31907 4022
rect 31853 3954 31863 3988
rect 31897 3954 31907 3988
rect 31853 3918 31907 3954
rect 31853 3884 31863 3918
rect 31897 3884 31907 3918
rect 31853 3868 31907 3884
rect 31937 4056 31989 4068
rect 31937 4022 31947 4056
rect 31981 4022 31989 4056
rect 31937 3988 31989 4022
rect 31937 3954 31947 3988
rect 31981 3954 31989 3988
rect 31937 3868 31989 3954
rect 43421 3840 43473 3852
rect 43421 3806 43429 3840
rect 43463 3806 43473 3840
rect 43421 3772 43473 3806
rect 13279 3680 13331 3692
rect 13279 3646 13287 3680
rect 13321 3646 13331 3680
rect 13279 3612 13331 3646
rect 13279 3578 13287 3612
rect 13321 3578 13331 3612
rect 13279 3542 13331 3578
rect 13279 3508 13287 3542
rect 13321 3508 13331 3542
rect 13279 3492 13331 3508
rect 13361 3680 13415 3692
rect 13361 3646 13371 3680
rect 13405 3646 13415 3680
rect 13361 3612 13415 3646
rect 13361 3578 13371 3612
rect 13405 3578 13415 3612
rect 13361 3542 13415 3578
rect 13361 3508 13371 3542
rect 13405 3508 13415 3542
rect 13361 3492 13415 3508
rect 13445 3680 13499 3692
rect 13445 3646 13455 3680
rect 13489 3646 13499 3680
rect 13445 3612 13499 3646
rect 13445 3578 13455 3612
rect 13489 3578 13499 3612
rect 13445 3492 13499 3578
rect 13529 3680 13583 3692
rect 13529 3646 13539 3680
rect 13573 3646 13583 3680
rect 13529 3612 13583 3646
rect 13529 3578 13539 3612
rect 13573 3578 13583 3612
rect 13529 3542 13583 3578
rect 13529 3508 13539 3542
rect 13573 3508 13583 3542
rect 13529 3492 13583 3508
rect 13613 3680 13667 3692
rect 13613 3646 13623 3680
rect 13657 3646 13667 3680
rect 13613 3612 13667 3646
rect 13613 3578 13623 3612
rect 13657 3578 13667 3612
rect 13613 3492 13667 3578
rect 13697 3680 13751 3692
rect 13697 3646 13707 3680
rect 13741 3646 13751 3680
rect 13697 3612 13751 3646
rect 13697 3578 13707 3612
rect 13741 3578 13751 3612
rect 13697 3542 13751 3578
rect 13697 3508 13707 3542
rect 13741 3508 13751 3542
rect 13697 3492 13751 3508
rect 13781 3680 13835 3692
rect 13781 3646 13791 3680
rect 13825 3646 13835 3680
rect 13781 3612 13835 3646
rect 13781 3578 13791 3612
rect 13825 3578 13835 3612
rect 13781 3492 13835 3578
rect 13865 3680 13919 3692
rect 13865 3646 13875 3680
rect 13909 3646 13919 3680
rect 13865 3612 13919 3646
rect 13865 3578 13875 3612
rect 13909 3578 13919 3612
rect 13865 3542 13919 3578
rect 13865 3508 13875 3542
rect 13909 3508 13919 3542
rect 13865 3492 13919 3508
rect 13949 3680 14003 3692
rect 13949 3646 13959 3680
rect 13993 3646 14003 3680
rect 13949 3612 14003 3646
rect 13949 3578 13959 3612
rect 13993 3578 14003 3612
rect 13949 3492 14003 3578
rect 14033 3680 14087 3692
rect 14033 3646 14043 3680
rect 14077 3646 14087 3680
rect 14033 3612 14087 3646
rect 14033 3578 14043 3612
rect 14077 3578 14087 3612
rect 14033 3542 14087 3578
rect 14033 3508 14043 3542
rect 14077 3508 14087 3542
rect 14033 3492 14087 3508
rect 14117 3680 14171 3692
rect 14117 3646 14127 3680
rect 14161 3646 14171 3680
rect 14117 3612 14171 3646
rect 14117 3578 14127 3612
rect 14161 3578 14171 3612
rect 14117 3492 14171 3578
rect 14201 3680 14255 3692
rect 14201 3646 14211 3680
rect 14245 3646 14255 3680
rect 14201 3612 14255 3646
rect 14201 3578 14211 3612
rect 14245 3578 14255 3612
rect 14201 3542 14255 3578
rect 14201 3508 14211 3542
rect 14245 3508 14255 3542
rect 14201 3492 14255 3508
rect 14285 3680 14339 3692
rect 14285 3646 14295 3680
rect 14329 3646 14339 3680
rect 14285 3612 14339 3646
rect 14285 3578 14295 3612
rect 14329 3578 14339 3612
rect 14285 3492 14339 3578
rect 14369 3680 14423 3692
rect 14369 3646 14379 3680
rect 14413 3646 14423 3680
rect 14369 3612 14423 3646
rect 14369 3578 14379 3612
rect 14413 3578 14423 3612
rect 14369 3542 14423 3578
rect 14369 3508 14379 3542
rect 14413 3508 14423 3542
rect 14369 3492 14423 3508
rect 14453 3680 14507 3692
rect 14453 3646 14463 3680
rect 14497 3646 14507 3680
rect 14453 3612 14507 3646
rect 14453 3578 14463 3612
rect 14497 3578 14507 3612
rect 14453 3492 14507 3578
rect 14537 3680 14591 3692
rect 14537 3646 14547 3680
rect 14581 3646 14591 3680
rect 14537 3612 14591 3646
rect 14537 3578 14547 3612
rect 14581 3578 14591 3612
rect 14537 3542 14591 3578
rect 14537 3508 14547 3542
rect 14581 3508 14591 3542
rect 14537 3492 14591 3508
rect 14621 3680 14673 3692
rect 14621 3646 14631 3680
rect 14665 3646 14673 3680
rect 15209 3680 15261 3692
rect 14621 3612 14673 3646
rect 14621 3578 14631 3612
rect 14665 3578 14673 3612
rect 15209 3646 15217 3680
rect 15251 3646 15261 3680
rect 15209 3612 15261 3646
rect 15209 3578 15217 3612
rect 15251 3578 15261 3612
rect 14621 3492 14673 3578
rect 15209 3542 15261 3578
rect 15209 3508 15217 3542
rect 15251 3508 15261 3542
rect 15209 3492 15261 3508
rect 15291 3680 15345 3692
rect 15291 3646 15301 3680
rect 15335 3646 15345 3680
rect 15291 3612 15345 3646
rect 15291 3578 15301 3612
rect 15335 3578 15345 3612
rect 15291 3542 15345 3578
rect 15291 3508 15301 3542
rect 15335 3508 15345 3542
rect 15291 3492 15345 3508
rect 15375 3680 15429 3692
rect 15375 3646 15385 3680
rect 15419 3646 15429 3680
rect 15375 3612 15429 3646
rect 15375 3578 15385 3612
rect 15419 3578 15429 3612
rect 15375 3492 15429 3578
rect 15459 3680 15513 3692
rect 15459 3646 15469 3680
rect 15503 3646 15513 3680
rect 15459 3612 15513 3646
rect 15459 3578 15469 3612
rect 15503 3578 15513 3612
rect 15459 3542 15513 3578
rect 15459 3508 15469 3542
rect 15503 3508 15513 3542
rect 15459 3492 15513 3508
rect 15543 3680 15597 3692
rect 15543 3646 15553 3680
rect 15587 3646 15597 3680
rect 15543 3612 15597 3646
rect 15543 3578 15553 3612
rect 15587 3578 15597 3612
rect 15543 3492 15597 3578
rect 15627 3680 15681 3692
rect 15627 3646 15637 3680
rect 15671 3646 15681 3680
rect 15627 3612 15681 3646
rect 15627 3578 15637 3612
rect 15671 3578 15681 3612
rect 15627 3542 15681 3578
rect 15627 3508 15637 3542
rect 15671 3508 15681 3542
rect 15627 3492 15681 3508
rect 15711 3680 15765 3692
rect 15711 3646 15721 3680
rect 15755 3646 15765 3680
rect 15711 3612 15765 3646
rect 15711 3578 15721 3612
rect 15755 3578 15765 3612
rect 15711 3492 15765 3578
rect 15795 3680 15849 3692
rect 15795 3646 15805 3680
rect 15839 3646 15849 3680
rect 15795 3612 15849 3646
rect 15795 3578 15805 3612
rect 15839 3578 15849 3612
rect 15795 3542 15849 3578
rect 15795 3508 15805 3542
rect 15839 3508 15849 3542
rect 15795 3492 15849 3508
rect 15879 3680 15933 3692
rect 15879 3646 15889 3680
rect 15923 3646 15933 3680
rect 15879 3612 15933 3646
rect 15879 3578 15889 3612
rect 15923 3578 15933 3612
rect 15879 3492 15933 3578
rect 15963 3680 16017 3692
rect 15963 3646 15973 3680
rect 16007 3646 16017 3680
rect 15963 3612 16017 3646
rect 15963 3578 15973 3612
rect 16007 3578 16017 3612
rect 15963 3542 16017 3578
rect 15963 3508 15973 3542
rect 16007 3508 16017 3542
rect 15963 3492 16017 3508
rect 16047 3680 16101 3692
rect 16047 3646 16057 3680
rect 16091 3646 16101 3680
rect 16047 3612 16101 3646
rect 16047 3578 16057 3612
rect 16091 3578 16101 3612
rect 16047 3492 16101 3578
rect 16131 3680 16185 3692
rect 16131 3646 16141 3680
rect 16175 3646 16185 3680
rect 16131 3612 16185 3646
rect 16131 3578 16141 3612
rect 16175 3578 16185 3612
rect 16131 3542 16185 3578
rect 16131 3508 16141 3542
rect 16175 3508 16185 3542
rect 16131 3492 16185 3508
rect 16215 3680 16269 3692
rect 16215 3646 16225 3680
rect 16259 3646 16269 3680
rect 16215 3612 16269 3646
rect 16215 3578 16225 3612
rect 16259 3578 16269 3612
rect 16215 3492 16269 3578
rect 16299 3680 16353 3692
rect 16299 3646 16309 3680
rect 16343 3646 16353 3680
rect 16299 3612 16353 3646
rect 16299 3578 16309 3612
rect 16343 3578 16353 3612
rect 16299 3542 16353 3578
rect 16299 3508 16309 3542
rect 16343 3508 16353 3542
rect 16299 3492 16353 3508
rect 16383 3680 16437 3692
rect 16383 3646 16393 3680
rect 16427 3646 16437 3680
rect 16383 3612 16437 3646
rect 16383 3578 16393 3612
rect 16427 3578 16437 3612
rect 16383 3492 16437 3578
rect 16467 3680 16521 3692
rect 16467 3646 16477 3680
rect 16511 3646 16521 3680
rect 16467 3612 16521 3646
rect 16467 3578 16477 3612
rect 16511 3578 16521 3612
rect 16467 3542 16521 3578
rect 16467 3508 16477 3542
rect 16511 3508 16521 3542
rect 16467 3492 16521 3508
rect 16551 3680 16603 3692
rect 16551 3646 16561 3680
rect 16595 3646 16603 3680
rect 16551 3612 16603 3646
rect 43421 3738 43429 3772
rect 43463 3738 43473 3772
rect 43421 3702 43473 3738
rect 43421 3668 43429 3702
rect 43463 3668 43473 3702
rect 43421 3652 43473 3668
rect 43503 3840 43557 3852
rect 43503 3806 43513 3840
rect 43547 3806 43557 3840
rect 43503 3772 43557 3806
rect 43503 3738 43513 3772
rect 43547 3738 43557 3772
rect 43503 3702 43557 3738
rect 43503 3668 43513 3702
rect 43547 3668 43557 3702
rect 43503 3652 43557 3668
rect 43587 3840 43641 3852
rect 43587 3806 43597 3840
rect 43631 3806 43641 3840
rect 43587 3772 43641 3806
rect 43587 3738 43597 3772
rect 43631 3738 43641 3772
rect 43587 3652 43641 3738
rect 43671 3840 43725 3852
rect 43671 3806 43681 3840
rect 43715 3806 43725 3840
rect 43671 3772 43725 3806
rect 43671 3738 43681 3772
rect 43715 3738 43725 3772
rect 43671 3702 43725 3738
rect 43671 3668 43681 3702
rect 43715 3668 43725 3702
rect 43671 3652 43725 3668
rect 43755 3840 43809 3852
rect 43755 3806 43765 3840
rect 43799 3806 43809 3840
rect 43755 3772 43809 3806
rect 43755 3738 43765 3772
rect 43799 3738 43809 3772
rect 43755 3652 43809 3738
rect 43839 3840 43893 3852
rect 43839 3806 43849 3840
rect 43883 3806 43893 3840
rect 43839 3772 43893 3806
rect 43839 3738 43849 3772
rect 43883 3738 43893 3772
rect 43839 3702 43893 3738
rect 43839 3668 43849 3702
rect 43883 3668 43893 3702
rect 43839 3652 43893 3668
rect 43923 3840 43977 3852
rect 43923 3806 43933 3840
rect 43967 3806 43977 3840
rect 43923 3772 43977 3806
rect 43923 3738 43933 3772
rect 43967 3738 43977 3772
rect 43923 3652 43977 3738
rect 44007 3840 44061 3852
rect 44007 3806 44017 3840
rect 44051 3806 44061 3840
rect 44007 3772 44061 3806
rect 44007 3738 44017 3772
rect 44051 3738 44061 3772
rect 44007 3702 44061 3738
rect 44007 3668 44017 3702
rect 44051 3668 44061 3702
rect 44007 3652 44061 3668
rect 44091 3840 44145 3852
rect 44091 3806 44101 3840
rect 44135 3806 44145 3840
rect 44091 3772 44145 3806
rect 44091 3738 44101 3772
rect 44135 3738 44145 3772
rect 44091 3652 44145 3738
rect 44175 3840 44229 3852
rect 44175 3806 44185 3840
rect 44219 3806 44229 3840
rect 44175 3772 44229 3806
rect 44175 3738 44185 3772
rect 44219 3738 44229 3772
rect 44175 3702 44229 3738
rect 44175 3668 44185 3702
rect 44219 3668 44229 3702
rect 44175 3652 44229 3668
rect 44259 3840 44313 3852
rect 44259 3806 44269 3840
rect 44303 3806 44313 3840
rect 44259 3772 44313 3806
rect 44259 3738 44269 3772
rect 44303 3738 44313 3772
rect 44259 3652 44313 3738
rect 44343 3840 44397 3852
rect 44343 3806 44353 3840
rect 44387 3806 44397 3840
rect 44343 3772 44397 3806
rect 44343 3738 44353 3772
rect 44387 3738 44397 3772
rect 44343 3702 44397 3738
rect 44343 3668 44353 3702
rect 44387 3668 44397 3702
rect 44343 3652 44397 3668
rect 44427 3840 44481 3852
rect 44427 3806 44437 3840
rect 44471 3806 44481 3840
rect 44427 3772 44481 3806
rect 44427 3738 44437 3772
rect 44471 3738 44481 3772
rect 44427 3652 44481 3738
rect 44511 3840 44565 3852
rect 44511 3806 44521 3840
rect 44555 3806 44565 3840
rect 44511 3772 44565 3806
rect 44511 3738 44521 3772
rect 44555 3738 44565 3772
rect 44511 3702 44565 3738
rect 44511 3668 44521 3702
rect 44555 3668 44565 3702
rect 44511 3652 44565 3668
rect 44595 3840 44649 3852
rect 44595 3806 44605 3840
rect 44639 3806 44649 3840
rect 44595 3772 44649 3806
rect 44595 3738 44605 3772
rect 44639 3738 44649 3772
rect 44595 3652 44649 3738
rect 44679 3840 44733 3852
rect 44679 3806 44689 3840
rect 44723 3806 44733 3840
rect 44679 3772 44733 3806
rect 44679 3738 44689 3772
rect 44723 3738 44733 3772
rect 44679 3702 44733 3738
rect 44679 3668 44689 3702
rect 44723 3668 44733 3702
rect 44679 3652 44733 3668
rect 44763 3840 44815 3852
rect 44763 3806 44773 3840
rect 44807 3806 44815 3840
rect 45351 3840 45403 3852
rect 44763 3772 44815 3806
rect 44763 3738 44773 3772
rect 44807 3738 44815 3772
rect 45351 3806 45359 3840
rect 45393 3806 45403 3840
rect 45351 3772 45403 3806
rect 45351 3738 45359 3772
rect 45393 3738 45403 3772
rect 44763 3652 44815 3738
rect 45351 3702 45403 3738
rect 45351 3668 45359 3702
rect 45393 3668 45403 3702
rect 45351 3652 45403 3668
rect 45433 3840 45487 3852
rect 45433 3806 45443 3840
rect 45477 3806 45487 3840
rect 45433 3772 45487 3806
rect 45433 3738 45443 3772
rect 45477 3738 45487 3772
rect 45433 3702 45487 3738
rect 45433 3668 45443 3702
rect 45477 3668 45487 3702
rect 45433 3652 45487 3668
rect 45517 3840 45571 3852
rect 45517 3806 45527 3840
rect 45561 3806 45571 3840
rect 45517 3772 45571 3806
rect 45517 3738 45527 3772
rect 45561 3738 45571 3772
rect 45517 3652 45571 3738
rect 45601 3840 45655 3852
rect 45601 3806 45611 3840
rect 45645 3806 45655 3840
rect 45601 3772 45655 3806
rect 45601 3738 45611 3772
rect 45645 3738 45655 3772
rect 45601 3702 45655 3738
rect 45601 3668 45611 3702
rect 45645 3668 45655 3702
rect 45601 3652 45655 3668
rect 45685 3840 45739 3852
rect 45685 3806 45695 3840
rect 45729 3806 45739 3840
rect 45685 3772 45739 3806
rect 45685 3738 45695 3772
rect 45729 3738 45739 3772
rect 45685 3652 45739 3738
rect 45769 3840 45823 3852
rect 45769 3806 45779 3840
rect 45813 3806 45823 3840
rect 45769 3772 45823 3806
rect 45769 3738 45779 3772
rect 45813 3738 45823 3772
rect 45769 3702 45823 3738
rect 45769 3668 45779 3702
rect 45813 3668 45823 3702
rect 45769 3652 45823 3668
rect 45853 3840 45907 3852
rect 45853 3806 45863 3840
rect 45897 3806 45907 3840
rect 45853 3772 45907 3806
rect 45853 3738 45863 3772
rect 45897 3738 45907 3772
rect 45853 3652 45907 3738
rect 45937 3840 45991 3852
rect 45937 3806 45947 3840
rect 45981 3806 45991 3840
rect 45937 3772 45991 3806
rect 45937 3738 45947 3772
rect 45981 3738 45991 3772
rect 45937 3702 45991 3738
rect 45937 3668 45947 3702
rect 45981 3668 45991 3702
rect 45937 3652 45991 3668
rect 46021 3840 46075 3852
rect 46021 3806 46031 3840
rect 46065 3806 46075 3840
rect 46021 3772 46075 3806
rect 46021 3738 46031 3772
rect 46065 3738 46075 3772
rect 46021 3652 46075 3738
rect 46105 3840 46159 3852
rect 46105 3806 46115 3840
rect 46149 3806 46159 3840
rect 46105 3772 46159 3806
rect 46105 3738 46115 3772
rect 46149 3738 46159 3772
rect 46105 3702 46159 3738
rect 46105 3668 46115 3702
rect 46149 3668 46159 3702
rect 46105 3652 46159 3668
rect 46189 3840 46243 3852
rect 46189 3806 46199 3840
rect 46233 3806 46243 3840
rect 46189 3772 46243 3806
rect 46189 3738 46199 3772
rect 46233 3738 46243 3772
rect 46189 3652 46243 3738
rect 46273 3840 46327 3852
rect 46273 3806 46283 3840
rect 46317 3806 46327 3840
rect 46273 3772 46327 3806
rect 46273 3738 46283 3772
rect 46317 3738 46327 3772
rect 46273 3702 46327 3738
rect 46273 3668 46283 3702
rect 46317 3668 46327 3702
rect 46273 3652 46327 3668
rect 46357 3840 46411 3852
rect 46357 3806 46367 3840
rect 46401 3806 46411 3840
rect 46357 3772 46411 3806
rect 46357 3738 46367 3772
rect 46401 3738 46411 3772
rect 46357 3652 46411 3738
rect 46441 3840 46495 3852
rect 46441 3806 46451 3840
rect 46485 3806 46495 3840
rect 46441 3772 46495 3806
rect 46441 3738 46451 3772
rect 46485 3738 46495 3772
rect 46441 3702 46495 3738
rect 46441 3668 46451 3702
rect 46485 3668 46495 3702
rect 46441 3652 46495 3668
rect 46525 3840 46579 3852
rect 46525 3806 46535 3840
rect 46569 3806 46579 3840
rect 46525 3772 46579 3806
rect 46525 3738 46535 3772
rect 46569 3738 46579 3772
rect 46525 3652 46579 3738
rect 46609 3840 46663 3852
rect 46609 3806 46619 3840
rect 46653 3806 46663 3840
rect 46609 3772 46663 3806
rect 46609 3738 46619 3772
rect 46653 3738 46663 3772
rect 46609 3702 46663 3738
rect 46609 3668 46619 3702
rect 46653 3668 46663 3702
rect 46609 3652 46663 3668
rect 46693 3840 46745 3852
rect 46693 3806 46703 3840
rect 46737 3806 46745 3840
rect 46693 3772 46745 3806
rect 46693 3738 46703 3772
rect 46737 3738 46745 3772
rect 46693 3652 46745 3738
rect 16551 3578 16561 3612
rect 16595 3578 16603 3612
rect 16551 3492 16603 3578
rect 5704 2481 5756 2497
rect 5704 2447 5712 2481
rect 5746 2447 5756 2481
rect 5704 2411 5756 2447
rect 5704 2377 5712 2411
rect 5746 2377 5756 2411
rect 5704 2343 5756 2377
rect 5704 2309 5712 2343
rect 5746 2309 5756 2343
rect 5704 2297 5756 2309
rect 5786 2481 5840 2497
rect 5786 2447 5796 2481
rect 5830 2447 5840 2481
rect 5786 2411 5840 2447
rect 5786 2377 5796 2411
rect 5830 2377 5840 2411
rect 5786 2343 5840 2377
rect 5786 2309 5796 2343
rect 5830 2309 5840 2343
rect 5786 2297 5840 2309
rect 5870 2411 5924 2497
rect 5870 2377 5880 2411
rect 5914 2377 5924 2411
rect 5870 2343 5924 2377
rect 5870 2309 5880 2343
rect 5914 2309 5924 2343
rect 5870 2297 5924 2309
rect 5954 2481 6008 2497
rect 5954 2447 5964 2481
rect 5998 2447 6008 2481
rect 5954 2411 6008 2447
rect 5954 2377 5964 2411
rect 5998 2377 6008 2411
rect 5954 2343 6008 2377
rect 5954 2309 5964 2343
rect 5998 2309 6008 2343
rect 5954 2297 6008 2309
rect 6038 2411 6092 2497
rect 6038 2377 6048 2411
rect 6082 2377 6092 2411
rect 6038 2343 6092 2377
rect 6038 2309 6048 2343
rect 6082 2309 6092 2343
rect 6038 2297 6092 2309
rect 6122 2481 6176 2497
rect 6122 2447 6132 2481
rect 6166 2447 6176 2481
rect 6122 2411 6176 2447
rect 6122 2377 6132 2411
rect 6166 2377 6176 2411
rect 6122 2343 6176 2377
rect 6122 2309 6132 2343
rect 6166 2309 6176 2343
rect 6122 2297 6176 2309
rect 6206 2411 6260 2497
rect 6206 2377 6216 2411
rect 6250 2377 6260 2411
rect 6206 2343 6260 2377
rect 6206 2309 6216 2343
rect 6250 2309 6260 2343
rect 6206 2297 6260 2309
rect 6290 2481 6344 2497
rect 6290 2447 6300 2481
rect 6334 2447 6344 2481
rect 6290 2411 6344 2447
rect 6290 2377 6300 2411
rect 6334 2377 6344 2411
rect 6290 2343 6344 2377
rect 6290 2309 6300 2343
rect 6334 2309 6344 2343
rect 6290 2297 6344 2309
rect 6374 2411 6428 2497
rect 6374 2377 6384 2411
rect 6418 2377 6428 2411
rect 6374 2343 6428 2377
rect 6374 2309 6384 2343
rect 6418 2309 6428 2343
rect 6374 2297 6428 2309
rect 6458 2481 6512 2497
rect 6458 2447 6468 2481
rect 6502 2447 6512 2481
rect 6458 2411 6512 2447
rect 6458 2377 6468 2411
rect 6502 2377 6512 2411
rect 6458 2343 6512 2377
rect 6458 2309 6468 2343
rect 6502 2309 6512 2343
rect 6458 2297 6512 2309
rect 6542 2411 6596 2497
rect 6542 2377 6552 2411
rect 6586 2377 6596 2411
rect 6542 2343 6596 2377
rect 6542 2309 6552 2343
rect 6586 2309 6596 2343
rect 6542 2297 6596 2309
rect 6626 2481 6680 2497
rect 6626 2447 6636 2481
rect 6670 2447 6680 2481
rect 6626 2411 6680 2447
rect 6626 2377 6636 2411
rect 6670 2377 6680 2411
rect 6626 2343 6680 2377
rect 6626 2309 6636 2343
rect 6670 2309 6680 2343
rect 6626 2297 6680 2309
rect 6710 2411 6764 2497
rect 6710 2377 6720 2411
rect 6754 2377 6764 2411
rect 6710 2343 6764 2377
rect 6710 2309 6720 2343
rect 6754 2309 6764 2343
rect 6710 2297 6764 2309
rect 6794 2481 6848 2497
rect 6794 2447 6804 2481
rect 6838 2447 6848 2481
rect 6794 2411 6848 2447
rect 6794 2377 6804 2411
rect 6838 2377 6848 2411
rect 6794 2343 6848 2377
rect 6794 2309 6804 2343
rect 6838 2309 6848 2343
rect 6794 2297 6848 2309
rect 6878 2411 6932 2497
rect 6878 2377 6888 2411
rect 6922 2377 6932 2411
rect 6878 2343 6932 2377
rect 6878 2309 6888 2343
rect 6922 2309 6932 2343
rect 6878 2297 6932 2309
rect 6962 2481 7016 2497
rect 6962 2447 6972 2481
rect 7006 2447 7016 2481
rect 6962 2411 7016 2447
rect 6962 2377 6972 2411
rect 7006 2377 7016 2411
rect 6962 2343 7016 2377
rect 6962 2309 6972 2343
rect 7006 2309 7016 2343
rect 6962 2297 7016 2309
rect 7046 2411 7098 2497
rect 7046 2377 7056 2411
rect 7090 2377 7098 2411
rect 7046 2343 7098 2377
rect 7046 2309 7056 2343
rect 7090 2309 7098 2343
rect 7046 2297 7098 2309
rect 7586 2479 7638 2495
rect 7586 2445 7594 2479
rect 7628 2445 7638 2479
rect 7586 2409 7638 2445
rect 7586 2375 7594 2409
rect 7628 2375 7638 2409
rect 7586 2341 7638 2375
rect 7586 2307 7594 2341
rect 7628 2307 7638 2341
rect 7586 2295 7638 2307
rect 7668 2479 7722 2495
rect 7668 2445 7678 2479
rect 7712 2445 7722 2479
rect 7668 2409 7722 2445
rect 7668 2375 7678 2409
rect 7712 2375 7722 2409
rect 7668 2341 7722 2375
rect 7668 2307 7678 2341
rect 7712 2307 7722 2341
rect 7668 2295 7722 2307
rect 7752 2409 7806 2495
rect 7752 2375 7762 2409
rect 7796 2375 7806 2409
rect 7752 2341 7806 2375
rect 7752 2307 7762 2341
rect 7796 2307 7806 2341
rect 7752 2295 7806 2307
rect 7836 2479 7890 2495
rect 7836 2445 7846 2479
rect 7880 2445 7890 2479
rect 7836 2409 7890 2445
rect 7836 2375 7846 2409
rect 7880 2375 7890 2409
rect 7836 2341 7890 2375
rect 7836 2307 7846 2341
rect 7880 2307 7890 2341
rect 7836 2295 7890 2307
rect 7920 2409 7974 2495
rect 7920 2375 7930 2409
rect 7964 2375 7974 2409
rect 7920 2341 7974 2375
rect 7920 2307 7930 2341
rect 7964 2307 7974 2341
rect 7920 2295 7974 2307
rect 8004 2479 8058 2495
rect 8004 2445 8014 2479
rect 8048 2445 8058 2479
rect 8004 2409 8058 2445
rect 8004 2375 8014 2409
rect 8048 2375 8058 2409
rect 8004 2341 8058 2375
rect 8004 2307 8014 2341
rect 8048 2307 8058 2341
rect 8004 2295 8058 2307
rect 8088 2409 8142 2495
rect 8088 2375 8098 2409
rect 8132 2375 8142 2409
rect 8088 2341 8142 2375
rect 8088 2307 8098 2341
rect 8132 2307 8142 2341
rect 8088 2295 8142 2307
rect 8172 2479 8226 2495
rect 8172 2445 8182 2479
rect 8216 2445 8226 2479
rect 8172 2409 8226 2445
rect 8172 2375 8182 2409
rect 8216 2375 8226 2409
rect 8172 2341 8226 2375
rect 8172 2307 8182 2341
rect 8216 2307 8226 2341
rect 8172 2295 8226 2307
rect 8256 2409 8310 2495
rect 8256 2375 8266 2409
rect 8300 2375 8310 2409
rect 8256 2341 8310 2375
rect 8256 2307 8266 2341
rect 8300 2307 8310 2341
rect 8256 2295 8310 2307
rect 8340 2479 8394 2495
rect 8340 2445 8350 2479
rect 8384 2445 8394 2479
rect 8340 2409 8394 2445
rect 8340 2375 8350 2409
rect 8384 2375 8394 2409
rect 8340 2341 8394 2375
rect 8340 2307 8350 2341
rect 8384 2307 8394 2341
rect 8340 2295 8394 2307
rect 8424 2409 8478 2495
rect 8424 2375 8434 2409
rect 8468 2375 8478 2409
rect 8424 2341 8478 2375
rect 8424 2307 8434 2341
rect 8468 2307 8478 2341
rect 8424 2295 8478 2307
rect 8508 2479 8562 2495
rect 8508 2445 8518 2479
rect 8552 2445 8562 2479
rect 8508 2409 8562 2445
rect 8508 2375 8518 2409
rect 8552 2375 8562 2409
rect 8508 2341 8562 2375
rect 8508 2307 8518 2341
rect 8552 2307 8562 2341
rect 8508 2295 8562 2307
rect 8592 2409 8646 2495
rect 8592 2375 8602 2409
rect 8636 2375 8646 2409
rect 8592 2341 8646 2375
rect 8592 2307 8602 2341
rect 8636 2307 8646 2341
rect 8592 2295 8646 2307
rect 8676 2479 8730 2495
rect 8676 2445 8686 2479
rect 8720 2445 8730 2479
rect 8676 2409 8730 2445
rect 8676 2375 8686 2409
rect 8720 2375 8730 2409
rect 8676 2341 8730 2375
rect 8676 2307 8686 2341
rect 8720 2307 8730 2341
rect 8676 2295 8730 2307
rect 8760 2409 8814 2495
rect 8760 2375 8770 2409
rect 8804 2375 8814 2409
rect 8760 2341 8814 2375
rect 8760 2307 8770 2341
rect 8804 2307 8814 2341
rect 8760 2295 8814 2307
rect 8844 2479 8898 2495
rect 8844 2445 8854 2479
rect 8888 2445 8898 2479
rect 8844 2409 8898 2445
rect 8844 2375 8854 2409
rect 8888 2375 8898 2409
rect 8844 2341 8898 2375
rect 8844 2307 8854 2341
rect 8888 2307 8898 2341
rect 8844 2295 8898 2307
rect 8928 2409 8980 2495
rect 8928 2375 8938 2409
rect 8972 2375 8980 2409
rect 8928 2341 8980 2375
rect 8928 2307 8938 2341
rect 8972 2307 8980 2341
rect 8928 2295 8980 2307
rect 20802 2481 20854 2497
rect 20802 2447 20810 2481
rect 20844 2447 20854 2481
rect 20802 2411 20854 2447
rect 20802 2377 20810 2411
rect 20844 2377 20854 2411
rect 20802 2343 20854 2377
rect 20802 2309 20810 2343
rect 20844 2309 20854 2343
rect 20802 2297 20854 2309
rect 20884 2481 20938 2497
rect 20884 2447 20894 2481
rect 20928 2447 20938 2481
rect 20884 2411 20938 2447
rect 20884 2377 20894 2411
rect 20928 2377 20938 2411
rect 20884 2343 20938 2377
rect 20884 2309 20894 2343
rect 20928 2309 20938 2343
rect 20884 2297 20938 2309
rect 20968 2411 21022 2497
rect 20968 2377 20978 2411
rect 21012 2377 21022 2411
rect 20968 2343 21022 2377
rect 20968 2309 20978 2343
rect 21012 2309 21022 2343
rect 20968 2297 21022 2309
rect 21052 2481 21106 2497
rect 21052 2447 21062 2481
rect 21096 2447 21106 2481
rect 21052 2411 21106 2447
rect 21052 2377 21062 2411
rect 21096 2377 21106 2411
rect 21052 2343 21106 2377
rect 21052 2309 21062 2343
rect 21096 2309 21106 2343
rect 21052 2297 21106 2309
rect 21136 2411 21190 2497
rect 21136 2377 21146 2411
rect 21180 2377 21190 2411
rect 21136 2343 21190 2377
rect 21136 2309 21146 2343
rect 21180 2309 21190 2343
rect 21136 2297 21190 2309
rect 21220 2481 21274 2497
rect 21220 2447 21230 2481
rect 21264 2447 21274 2481
rect 21220 2411 21274 2447
rect 21220 2377 21230 2411
rect 21264 2377 21274 2411
rect 21220 2343 21274 2377
rect 21220 2309 21230 2343
rect 21264 2309 21274 2343
rect 21220 2297 21274 2309
rect 21304 2411 21358 2497
rect 21304 2377 21314 2411
rect 21348 2377 21358 2411
rect 21304 2343 21358 2377
rect 21304 2309 21314 2343
rect 21348 2309 21358 2343
rect 21304 2297 21358 2309
rect 21388 2481 21442 2497
rect 21388 2447 21398 2481
rect 21432 2447 21442 2481
rect 21388 2411 21442 2447
rect 21388 2377 21398 2411
rect 21432 2377 21442 2411
rect 21388 2343 21442 2377
rect 21388 2309 21398 2343
rect 21432 2309 21442 2343
rect 21388 2297 21442 2309
rect 21472 2411 21526 2497
rect 21472 2377 21482 2411
rect 21516 2377 21526 2411
rect 21472 2343 21526 2377
rect 21472 2309 21482 2343
rect 21516 2309 21526 2343
rect 21472 2297 21526 2309
rect 21556 2481 21610 2497
rect 21556 2447 21566 2481
rect 21600 2447 21610 2481
rect 21556 2411 21610 2447
rect 21556 2377 21566 2411
rect 21600 2377 21610 2411
rect 21556 2343 21610 2377
rect 21556 2309 21566 2343
rect 21600 2309 21610 2343
rect 21556 2297 21610 2309
rect 21640 2411 21694 2497
rect 21640 2377 21650 2411
rect 21684 2377 21694 2411
rect 21640 2343 21694 2377
rect 21640 2309 21650 2343
rect 21684 2309 21694 2343
rect 21640 2297 21694 2309
rect 21724 2481 21778 2497
rect 21724 2447 21734 2481
rect 21768 2447 21778 2481
rect 21724 2411 21778 2447
rect 21724 2377 21734 2411
rect 21768 2377 21778 2411
rect 21724 2343 21778 2377
rect 21724 2309 21734 2343
rect 21768 2309 21778 2343
rect 21724 2297 21778 2309
rect 21808 2411 21862 2497
rect 21808 2377 21818 2411
rect 21852 2377 21862 2411
rect 21808 2343 21862 2377
rect 21808 2309 21818 2343
rect 21852 2309 21862 2343
rect 21808 2297 21862 2309
rect 21892 2481 21946 2497
rect 21892 2447 21902 2481
rect 21936 2447 21946 2481
rect 21892 2411 21946 2447
rect 21892 2377 21902 2411
rect 21936 2377 21946 2411
rect 21892 2343 21946 2377
rect 21892 2309 21902 2343
rect 21936 2309 21946 2343
rect 21892 2297 21946 2309
rect 21976 2411 22030 2497
rect 21976 2377 21986 2411
rect 22020 2377 22030 2411
rect 21976 2343 22030 2377
rect 21976 2309 21986 2343
rect 22020 2309 22030 2343
rect 21976 2297 22030 2309
rect 22060 2481 22114 2497
rect 22060 2447 22070 2481
rect 22104 2447 22114 2481
rect 22060 2411 22114 2447
rect 22060 2377 22070 2411
rect 22104 2377 22114 2411
rect 22060 2343 22114 2377
rect 22060 2309 22070 2343
rect 22104 2309 22114 2343
rect 22060 2297 22114 2309
rect 22144 2411 22196 2497
rect 22144 2377 22154 2411
rect 22188 2377 22196 2411
rect 22144 2343 22196 2377
rect 22144 2309 22154 2343
rect 22188 2309 22196 2343
rect 22144 2297 22196 2309
rect 22684 2479 22736 2495
rect 22684 2445 22692 2479
rect 22726 2445 22736 2479
rect 22684 2409 22736 2445
rect 22684 2375 22692 2409
rect 22726 2375 22736 2409
rect 22684 2341 22736 2375
rect 22684 2307 22692 2341
rect 22726 2307 22736 2341
rect 22684 2295 22736 2307
rect 22766 2479 22820 2495
rect 22766 2445 22776 2479
rect 22810 2445 22820 2479
rect 22766 2409 22820 2445
rect 22766 2375 22776 2409
rect 22810 2375 22820 2409
rect 22766 2341 22820 2375
rect 22766 2307 22776 2341
rect 22810 2307 22820 2341
rect 22766 2295 22820 2307
rect 22850 2409 22904 2495
rect 22850 2375 22860 2409
rect 22894 2375 22904 2409
rect 22850 2341 22904 2375
rect 22850 2307 22860 2341
rect 22894 2307 22904 2341
rect 22850 2295 22904 2307
rect 22934 2479 22988 2495
rect 22934 2445 22944 2479
rect 22978 2445 22988 2479
rect 22934 2409 22988 2445
rect 22934 2375 22944 2409
rect 22978 2375 22988 2409
rect 22934 2341 22988 2375
rect 22934 2307 22944 2341
rect 22978 2307 22988 2341
rect 22934 2295 22988 2307
rect 23018 2409 23072 2495
rect 23018 2375 23028 2409
rect 23062 2375 23072 2409
rect 23018 2341 23072 2375
rect 23018 2307 23028 2341
rect 23062 2307 23072 2341
rect 23018 2295 23072 2307
rect 23102 2479 23156 2495
rect 23102 2445 23112 2479
rect 23146 2445 23156 2479
rect 23102 2409 23156 2445
rect 23102 2375 23112 2409
rect 23146 2375 23156 2409
rect 23102 2341 23156 2375
rect 23102 2307 23112 2341
rect 23146 2307 23156 2341
rect 23102 2295 23156 2307
rect 23186 2409 23240 2495
rect 23186 2375 23196 2409
rect 23230 2375 23240 2409
rect 23186 2341 23240 2375
rect 23186 2307 23196 2341
rect 23230 2307 23240 2341
rect 23186 2295 23240 2307
rect 23270 2479 23324 2495
rect 23270 2445 23280 2479
rect 23314 2445 23324 2479
rect 23270 2409 23324 2445
rect 23270 2375 23280 2409
rect 23314 2375 23324 2409
rect 23270 2341 23324 2375
rect 23270 2307 23280 2341
rect 23314 2307 23324 2341
rect 23270 2295 23324 2307
rect 23354 2409 23408 2495
rect 23354 2375 23364 2409
rect 23398 2375 23408 2409
rect 23354 2341 23408 2375
rect 23354 2307 23364 2341
rect 23398 2307 23408 2341
rect 23354 2295 23408 2307
rect 23438 2479 23492 2495
rect 23438 2445 23448 2479
rect 23482 2445 23492 2479
rect 23438 2409 23492 2445
rect 23438 2375 23448 2409
rect 23482 2375 23492 2409
rect 23438 2341 23492 2375
rect 23438 2307 23448 2341
rect 23482 2307 23492 2341
rect 23438 2295 23492 2307
rect 23522 2409 23576 2495
rect 23522 2375 23532 2409
rect 23566 2375 23576 2409
rect 23522 2341 23576 2375
rect 23522 2307 23532 2341
rect 23566 2307 23576 2341
rect 23522 2295 23576 2307
rect 23606 2479 23660 2495
rect 23606 2445 23616 2479
rect 23650 2445 23660 2479
rect 23606 2409 23660 2445
rect 23606 2375 23616 2409
rect 23650 2375 23660 2409
rect 23606 2341 23660 2375
rect 23606 2307 23616 2341
rect 23650 2307 23660 2341
rect 23606 2295 23660 2307
rect 23690 2409 23744 2495
rect 23690 2375 23700 2409
rect 23734 2375 23744 2409
rect 23690 2341 23744 2375
rect 23690 2307 23700 2341
rect 23734 2307 23744 2341
rect 23690 2295 23744 2307
rect 23774 2479 23828 2495
rect 23774 2445 23784 2479
rect 23818 2445 23828 2479
rect 23774 2409 23828 2445
rect 23774 2375 23784 2409
rect 23818 2375 23828 2409
rect 23774 2341 23828 2375
rect 23774 2307 23784 2341
rect 23818 2307 23828 2341
rect 23774 2295 23828 2307
rect 23858 2409 23912 2495
rect 23858 2375 23868 2409
rect 23902 2375 23912 2409
rect 23858 2341 23912 2375
rect 23858 2307 23868 2341
rect 23902 2307 23912 2341
rect 23858 2295 23912 2307
rect 23942 2479 23996 2495
rect 23942 2445 23952 2479
rect 23986 2445 23996 2479
rect 23942 2409 23996 2445
rect 23942 2375 23952 2409
rect 23986 2375 23996 2409
rect 23942 2341 23996 2375
rect 23942 2307 23952 2341
rect 23986 2307 23996 2341
rect 23942 2295 23996 2307
rect 24026 2409 24078 2495
rect 24026 2375 24036 2409
rect 24070 2375 24078 2409
rect 24026 2341 24078 2375
rect 24026 2307 24036 2341
rect 24070 2307 24078 2341
rect 24026 2295 24078 2307
rect 35906 2481 35958 2497
rect 35906 2447 35914 2481
rect 35948 2447 35958 2481
rect 35906 2411 35958 2447
rect 35906 2377 35914 2411
rect 35948 2377 35958 2411
rect 35906 2343 35958 2377
rect 35906 2309 35914 2343
rect 35948 2309 35958 2343
rect 35906 2297 35958 2309
rect 35988 2481 36042 2497
rect 35988 2447 35998 2481
rect 36032 2447 36042 2481
rect 35988 2411 36042 2447
rect 35988 2377 35998 2411
rect 36032 2377 36042 2411
rect 35988 2343 36042 2377
rect 35988 2309 35998 2343
rect 36032 2309 36042 2343
rect 35988 2297 36042 2309
rect 36072 2411 36126 2497
rect 36072 2377 36082 2411
rect 36116 2377 36126 2411
rect 36072 2343 36126 2377
rect 36072 2309 36082 2343
rect 36116 2309 36126 2343
rect 36072 2297 36126 2309
rect 36156 2481 36210 2497
rect 36156 2447 36166 2481
rect 36200 2447 36210 2481
rect 36156 2411 36210 2447
rect 36156 2377 36166 2411
rect 36200 2377 36210 2411
rect 36156 2343 36210 2377
rect 36156 2309 36166 2343
rect 36200 2309 36210 2343
rect 36156 2297 36210 2309
rect 36240 2411 36294 2497
rect 36240 2377 36250 2411
rect 36284 2377 36294 2411
rect 36240 2343 36294 2377
rect 36240 2309 36250 2343
rect 36284 2309 36294 2343
rect 36240 2297 36294 2309
rect 36324 2481 36378 2497
rect 36324 2447 36334 2481
rect 36368 2447 36378 2481
rect 36324 2411 36378 2447
rect 36324 2377 36334 2411
rect 36368 2377 36378 2411
rect 36324 2343 36378 2377
rect 36324 2309 36334 2343
rect 36368 2309 36378 2343
rect 36324 2297 36378 2309
rect 36408 2411 36462 2497
rect 36408 2377 36418 2411
rect 36452 2377 36462 2411
rect 36408 2343 36462 2377
rect 36408 2309 36418 2343
rect 36452 2309 36462 2343
rect 36408 2297 36462 2309
rect 36492 2481 36546 2497
rect 36492 2447 36502 2481
rect 36536 2447 36546 2481
rect 36492 2411 36546 2447
rect 36492 2377 36502 2411
rect 36536 2377 36546 2411
rect 36492 2343 36546 2377
rect 36492 2309 36502 2343
rect 36536 2309 36546 2343
rect 36492 2297 36546 2309
rect 36576 2411 36630 2497
rect 36576 2377 36586 2411
rect 36620 2377 36630 2411
rect 36576 2343 36630 2377
rect 36576 2309 36586 2343
rect 36620 2309 36630 2343
rect 36576 2297 36630 2309
rect 36660 2481 36714 2497
rect 36660 2447 36670 2481
rect 36704 2447 36714 2481
rect 36660 2411 36714 2447
rect 36660 2377 36670 2411
rect 36704 2377 36714 2411
rect 36660 2343 36714 2377
rect 36660 2309 36670 2343
rect 36704 2309 36714 2343
rect 36660 2297 36714 2309
rect 36744 2411 36798 2497
rect 36744 2377 36754 2411
rect 36788 2377 36798 2411
rect 36744 2343 36798 2377
rect 36744 2309 36754 2343
rect 36788 2309 36798 2343
rect 36744 2297 36798 2309
rect 36828 2481 36882 2497
rect 36828 2447 36838 2481
rect 36872 2447 36882 2481
rect 36828 2411 36882 2447
rect 36828 2377 36838 2411
rect 36872 2377 36882 2411
rect 36828 2343 36882 2377
rect 36828 2309 36838 2343
rect 36872 2309 36882 2343
rect 36828 2297 36882 2309
rect 36912 2411 36966 2497
rect 36912 2377 36922 2411
rect 36956 2377 36966 2411
rect 36912 2343 36966 2377
rect 36912 2309 36922 2343
rect 36956 2309 36966 2343
rect 36912 2297 36966 2309
rect 36996 2481 37050 2497
rect 36996 2447 37006 2481
rect 37040 2447 37050 2481
rect 36996 2411 37050 2447
rect 36996 2377 37006 2411
rect 37040 2377 37050 2411
rect 36996 2343 37050 2377
rect 36996 2309 37006 2343
rect 37040 2309 37050 2343
rect 36996 2297 37050 2309
rect 37080 2411 37134 2497
rect 37080 2377 37090 2411
rect 37124 2377 37134 2411
rect 37080 2343 37134 2377
rect 37080 2309 37090 2343
rect 37124 2309 37134 2343
rect 37080 2297 37134 2309
rect 37164 2481 37218 2497
rect 37164 2447 37174 2481
rect 37208 2447 37218 2481
rect 37164 2411 37218 2447
rect 37164 2377 37174 2411
rect 37208 2377 37218 2411
rect 37164 2343 37218 2377
rect 37164 2309 37174 2343
rect 37208 2309 37218 2343
rect 37164 2297 37218 2309
rect 37248 2411 37300 2497
rect 37248 2377 37258 2411
rect 37292 2377 37300 2411
rect 37248 2343 37300 2377
rect 37248 2309 37258 2343
rect 37292 2309 37300 2343
rect 37248 2297 37300 2309
rect 37788 2479 37840 2495
rect 37788 2445 37796 2479
rect 37830 2445 37840 2479
rect 37788 2409 37840 2445
rect 37788 2375 37796 2409
rect 37830 2375 37840 2409
rect 37788 2341 37840 2375
rect 37788 2307 37796 2341
rect 37830 2307 37840 2341
rect 37788 2295 37840 2307
rect 37870 2479 37924 2495
rect 37870 2445 37880 2479
rect 37914 2445 37924 2479
rect 37870 2409 37924 2445
rect 37870 2375 37880 2409
rect 37914 2375 37924 2409
rect 37870 2341 37924 2375
rect 37870 2307 37880 2341
rect 37914 2307 37924 2341
rect 37870 2295 37924 2307
rect 37954 2409 38008 2495
rect 37954 2375 37964 2409
rect 37998 2375 38008 2409
rect 37954 2341 38008 2375
rect 37954 2307 37964 2341
rect 37998 2307 38008 2341
rect 37954 2295 38008 2307
rect 38038 2479 38092 2495
rect 38038 2445 38048 2479
rect 38082 2445 38092 2479
rect 38038 2409 38092 2445
rect 38038 2375 38048 2409
rect 38082 2375 38092 2409
rect 38038 2341 38092 2375
rect 38038 2307 38048 2341
rect 38082 2307 38092 2341
rect 38038 2295 38092 2307
rect 38122 2409 38176 2495
rect 38122 2375 38132 2409
rect 38166 2375 38176 2409
rect 38122 2341 38176 2375
rect 38122 2307 38132 2341
rect 38166 2307 38176 2341
rect 38122 2295 38176 2307
rect 38206 2479 38260 2495
rect 38206 2445 38216 2479
rect 38250 2445 38260 2479
rect 38206 2409 38260 2445
rect 38206 2375 38216 2409
rect 38250 2375 38260 2409
rect 38206 2341 38260 2375
rect 38206 2307 38216 2341
rect 38250 2307 38260 2341
rect 38206 2295 38260 2307
rect 38290 2409 38344 2495
rect 38290 2375 38300 2409
rect 38334 2375 38344 2409
rect 38290 2341 38344 2375
rect 38290 2307 38300 2341
rect 38334 2307 38344 2341
rect 38290 2295 38344 2307
rect 38374 2479 38428 2495
rect 38374 2445 38384 2479
rect 38418 2445 38428 2479
rect 38374 2409 38428 2445
rect 38374 2375 38384 2409
rect 38418 2375 38428 2409
rect 38374 2341 38428 2375
rect 38374 2307 38384 2341
rect 38418 2307 38428 2341
rect 38374 2295 38428 2307
rect 38458 2409 38512 2495
rect 38458 2375 38468 2409
rect 38502 2375 38512 2409
rect 38458 2341 38512 2375
rect 38458 2307 38468 2341
rect 38502 2307 38512 2341
rect 38458 2295 38512 2307
rect 38542 2479 38596 2495
rect 38542 2445 38552 2479
rect 38586 2445 38596 2479
rect 38542 2409 38596 2445
rect 38542 2375 38552 2409
rect 38586 2375 38596 2409
rect 38542 2341 38596 2375
rect 38542 2307 38552 2341
rect 38586 2307 38596 2341
rect 38542 2295 38596 2307
rect 38626 2409 38680 2495
rect 38626 2375 38636 2409
rect 38670 2375 38680 2409
rect 38626 2341 38680 2375
rect 38626 2307 38636 2341
rect 38670 2307 38680 2341
rect 38626 2295 38680 2307
rect 38710 2479 38764 2495
rect 38710 2445 38720 2479
rect 38754 2445 38764 2479
rect 38710 2409 38764 2445
rect 38710 2375 38720 2409
rect 38754 2375 38764 2409
rect 38710 2341 38764 2375
rect 38710 2307 38720 2341
rect 38754 2307 38764 2341
rect 38710 2295 38764 2307
rect 38794 2409 38848 2495
rect 38794 2375 38804 2409
rect 38838 2375 38848 2409
rect 38794 2341 38848 2375
rect 38794 2307 38804 2341
rect 38838 2307 38848 2341
rect 38794 2295 38848 2307
rect 38878 2479 38932 2495
rect 38878 2445 38888 2479
rect 38922 2445 38932 2479
rect 38878 2409 38932 2445
rect 38878 2375 38888 2409
rect 38922 2375 38932 2409
rect 38878 2341 38932 2375
rect 38878 2307 38888 2341
rect 38922 2307 38932 2341
rect 38878 2295 38932 2307
rect 38962 2409 39016 2495
rect 38962 2375 38972 2409
rect 39006 2375 39016 2409
rect 38962 2341 39016 2375
rect 38962 2307 38972 2341
rect 39006 2307 39016 2341
rect 38962 2295 39016 2307
rect 39046 2479 39100 2495
rect 39046 2445 39056 2479
rect 39090 2445 39100 2479
rect 39046 2409 39100 2445
rect 39046 2375 39056 2409
rect 39090 2375 39100 2409
rect 39046 2341 39100 2375
rect 39046 2307 39056 2341
rect 39090 2307 39100 2341
rect 39046 2295 39100 2307
rect 39130 2409 39182 2495
rect 39130 2375 39140 2409
rect 39174 2375 39182 2409
rect 39130 2341 39182 2375
rect 39130 2307 39140 2341
rect 39174 2307 39182 2341
rect 39130 2295 39182 2307
rect 51004 2481 51056 2497
rect 51004 2447 51012 2481
rect 51046 2447 51056 2481
rect 51004 2411 51056 2447
rect 51004 2377 51012 2411
rect 51046 2377 51056 2411
rect 51004 2343 51056 2377
rect 51004 2309 51012 2343
rect 51046 2309 51056 2343
rect 51004 2297 51056 2309
rect 51086 2481 51140 2497
rect 51086 2447 51096 2481
rect 51130 2447 51140 2481
rect 51086 2411 51140 2447
rect 51086 2377 51096 2411
rect 51130 2377 51140 2411
rect 51086 2343 51140 2377
rect 51086 2309 51096 2343
rect 51130 2309 51140 2343
rect 51086 2297 51140 2309
rect 51170 2411 51224 2497
rect 51170 2377 51180 2411
rect 51214 2377 51224 2411
rect 51170 2343 51224 2377
rect 51170 2309 51180 2343
rect 51214 2309 51224 2343
rect 51170 2297 51224 2309
rect 51254 2481 51308 2497
rect 51254 2447 51264 2481
rect 51298 2447 51308 2481
rect 51254 2411 51308 2447
rect 51254 2377 51264 2411
rect 51298 2377 51308 2411
rect 51254 2343 51308 2377
rect 51254 2309 51264 2343
rect 51298 2309 51308 2343
rect 51254 2297 51308 2309
rect 51338 2411 51392 2497
rect 51338 2377 51348 2411
rect 51382 2377 51392 2411
rect 51338 2343 51392 2377
rect 51338 2309 51348 2343
rect 51382 2309 51392 2343
rect 51338 2297 51392 2309
rect 51422 2481 51476 2497
rect 51422 2447 51432 2481
rect 51466 2447 51476 2481
rect 51422 2411 51476 2447
rect 51422 2377 51432 2411
rect 51466 2377 51476 2411
rect 51422 2343 51476 2377
rect 51422 2309 51432 2343
rect 51466 2309 51476 2343
rect 51422 2297 51476 2309
rect 51506 2411 51560 2497
rect 51506 2377 51516 2411
rect 51550 2377 51560 2411
rect 51506 2343 51560 2377
rect 51506 2309 51516 2343
rect 51550 2309 51560 2343
rect 51506 2297 51560 2309
rect 51590 2481 51644 2497
rect 51590 2447 51600 2481
rect 51634 2447 51644 2481
rect 51590 2411 51644 2447
rect 51590 2377 51600 2411
rect 51634 2377 51644 2411
rect 51590 2343 51644 2377
rect 51590 2309 51600 2343
rect 51634 2309 51644 2343
rect 51590 2297 51644 2309
rect 51674 2411 51728 2497
rect 51674 2377 51684 2411
rect 51718 2377 51728 2411
rect 51674 2343 51728 2377
rect 51674 2309 51684 2343
rect 51718 2309 51728 2343
rect 51674 2297 51728 2309
rect 51758 2481 51812 2497
rect 51758 2447 51768 2481
rect 51802 2447 51812 2481
rect 51758 2411 51812 2447
rect 51758 2377 51768 2411
rect 51802 2377 51812 2411
rect 51758 2343 51812 2377
rect 51758 2309 51768 2343
rect 51802 2309 51812 2343
rect 51758 2297 51812 2309
rect 51842 2411 51896 2497
rect 51842 2377 51852 2411
rect 51886 2377 51896 2411
rect 51842 2343 51896 2377
rect 51842 2309 51852 2343
rect 51886 2309 51896 2343
rect 51842 2297 51896 2309
rect 51926 2481 51980 2497
rect 51926 2447 51936 2481
rect 51970 2447 51980 2481
rect 51926 2411 51980 2447
rect 51926 2377 51936 2411
rect 51970 2377 51980 2411
rect 51926 2343 51980 2377
rect 51926 2309 51936 2343
rect 51970 2309 51980 2343
rect 51926 2297 51980 2309
rect 52010 2411 52064 2497
rect 52010 2377 52020 2411
rect 52054 2377 52064 2411
rect 52010 2343 52064 2377
rect 52010 2309 52020 2343
rect 52054 2309 52064 2343
rect 52010 2297 52064 2309
rect 52094 2481 52148 2497
rect 52094 2447 52104 2481
rect 52138 2447 52148 2481
rect 52094 2411 52148 2447
rect 52094 2377 52104 2411
rect 52138 2377 52148 2411
rect 52094 2343 52148 2377
rect 52094 2309 52104 2343
rect 52138 2309 52148 2343
rect 52094 2297 52148 2309
rect 52178 2411 52232 2497
rect 52178 2377 52188 2411
rect 52222 2377 52232 2411
rect 52178 2343 52232 2377
rect 52178 2309 52188 2343
rect 52222 2309 52232 2343
rect 52178 2297 52232 2309
rect 52262 2481 52316 2497
rect 52262 2447 52272 2481
rect 52306 2447 52316 2481
rect 52262 2411 52316 2447
rect 52262 2377 52272 2411
rect 52306 2377 52316 2411
rect 52262 2343 52316 2377
rect 52262 2309 52272 2343
rect 52306 2309 52316 2343
rect 52262 2297 52316 2309
rect 52346 2411 52398 2497
rect 52346 2377 52356 2411
rect 52390 2377 52398 2411
rect 52346 2343 52398 2377
rect 52346 2309 52356 2343
rect 52390 2309 52398 2343
rect 52346 2297 52398 2309
rect 52886 2479 52938 2495
rect 52886 2445 52894 2479
rect 52928 2445 52938 2479
rect 52886 2409 52938 2445
rect 52886 2375 52894 2409
rect 52928 2375 52938 2409
rect 52886 2341 52938 2375
rect 52886 2307 52894 2341
rect 52928 2307 52938 2341
rect 52886 2295 52938 2307
rect 52968 2479 53022 2495
rect 52968 2445 52978 2479
rect 53012 2445 53022 2479
rect 52968 2409 53022 2445
rect 52968 2375 52978 2409
rect 53012 2375 53022 2409
rect 52968 2341 53022 2375
rect 52968 2307 52978 2341
rect 53012 2307 53022 2341
rect 52968 2295 53022 2307
rect 53052 2409 53106 2495
rect 53052 2375 53062 2409
rect 53096 2375 53106 2409
rect 53052 2341 53106 2375
rect 53052 2307 53062 2341
rect 53096 2307 53106 2341
rect 53052 2295 53106 2307
rect 53136 2479 53190 2495
rect 53136 2445 53146 2479
rect 53180 2445 53190 2479
rect 53136 2409 53190 2445
rect 53136 2375 53146 2409
rect 53180 2375 53190 2409
rect 53136 2341 53190 2375
rect 53136 2307 53146 2341
rect 53180 2307 53190 2341
rect 53136 2295 53190 2307
rect 53220 2409 53274 2495
rect 53220 2375 53230 2409
rect 53264 2375 53274 2409
rect 53220 2341 53274 2375
rect 53220 2307 53230 2341
rect 53264 2307 53274 2341
rect 53220 2295 53274 2307
rect 53304 2479 53358 2495
rect 53304 2445 53314 2479
rect 53348 2445 53358 2479
rect 53304 2409 53358 2445
rect 53304 2375 53314 2409
rect 53348 2375 53358 2409
rect 53304 2341 53358 2375
rect 53304 2307 53314 2341
rect 53348 2307 53358 2341
rect 53304 2295 53358 2307
rect 53388 2409 53442 2495
rect 53388 2375 53398 2409
rect 53432 2375 53442 2409
rect 53388 2341 53442 2375
rect 53388 2307 53398 2341
rect 53432 2307 53442 2341
rect 53388 2295 53442 2307
rect 53472 2479 53526 2495
rect 53472 2445 53482 2479
rect 53516 2445 53526 2479
rect 53472 2409 53526 2445
rect 53472 2375 53482 2409
rect 53516 2375 53526 2409
rect 53472 2341 53526 2375
rect 53472 2307 53482 2341
rect 53516 2307 53526 2341
rect 53472 2295 53526 2307
rect 53556 2409 53610 2495
rect 53556 2375 53566 2409
rect 53600 2375 53610 2409
rect 53556 2341 53610 2375
rect 53556 2307 53566 2341
rect 53600 2307 53610 2341
rect 53556 2295 53610 2307
rect 53640 2479 53694 2495
rect 53640 2445 53650 2479
rect 53684 2445 53694 2479
rect 53640 2409 53694 2445
rect 53640 2375 53650 2409
rect 53684 2375 53694 2409
rect 53640 2341 53694 2375
rect 53640 2307 53650 2341
rect 53684 2307 53694 2341
rect 53640 2295 53694 2307
rect 53724 2409 53778 2495
rect 53724 2375 53734 2409
rect 53768 2375 53778 2409
rect 53724 2341 53778 2375
rect 53724 2307 53734 2341
rect 53768 2307 53778 2341
rect 53724 2295 53778 2307
rect 53808 2479 53862 2495
rect 53808 2445 53818 2479
rect 53852 2445 53862 2479
rect 53808 2409 53862 2445
rect 53808 2375 53818 2409
rect 53852 2375 53862 2409
rect 53808 2341 53862 2375
rect 53808 2307 53818 2341
rect 53852 2307 53862 2341
rect 53808 2295 53862 2307
rect 53892 2409 53946 2495
rect 53892 2375 53902 2409
rect 53936 2375 53946 2409
rect 53892 2341 53946 2375
rect 53892 2307 53902 2341
rect 53936 2307 53946 2341
rect 53892 2295 53946 2307
rect 53976 2479 54030 2495
rect 53976 2445 53986 2479
rect 54020 2445 54030 2479
rect 53976 2409 54030 2445
rect 53976 2375 53986 2409
rect 54020 2375 54030 2409
rect 53976 2341 54030 2375
rect 53976 2307 53986 2341
rect 54020 2307 54030 2341
rect 53976 2295 54030 2307
rect 54060 2409 54114 2495
rect 54060 2375 54070 2409
rect 54104 2375 54114 2409
rect 54060 2341 54114 2375
rect 54060 2307 54070 2341
rect 54104 2307 54114 2341
rect 54060 2295 54114 2307
rect 54144 2479 54198 2495
rect 54144 2445 54154 2479
rect 54188 2445 54198 2479
rect 54144 2409 54198 2445
rect 54144 2375 54154 2409
rect 54188 2375 54198 2409
rect 54144 2341 54198 2375
rect 54144 2307 54154 2341
rect 54188 2307 54198 2341
rect 54144 2295 54198 2307
rect 54228 2409 54280 2495
rect 54228 2375 54238 2409
rect 54272 2375 54280 2409
rect 54228 2341 54280 2375
rect 54228 2307 54238 2341
rect 54272 2307 54280 2341
rect 54228 2295 54280 2307
rect 245 2111 297 2123
rect 245 2077 253 2111
rect 287 2077 297 2111
rect 245 2043 297 2077
rect 245 2009 253 2043
rect 287 2009 297 2043
rect 245 1975 297 2009
rect 245 1941 253 1975
rect 287 1941 297 1975
rect 245 1923 297 1941
rect 327 1923 369 2123
rect 399 2111 451 2123
rect 399 2077 409 2111
rect 443 2077 451 2111
rect 1059 2111 1111 2123
rect 399 2043 451 2077
rect 1059 2077 1067 2111
rect 1101 2077 1111 2111
rect 399 2009 409 2043
rect 443 2009 451 2043
rect 399 1975 451 2009
rect 1059 2043 1111 2077
rect 1059 2009 1067 2043
rect 1101 2009 1111 2043
rect 399 1941 409 1975
rect 443 1941 451 1975
rect 1059 1975 1111 2009
rect 399 1923 451 1941
rect 594 1943 656 1958
rect 594 1909 606 1943
rect 640 1909 656 1943
rect 594 1875 656 1909
rect 594 1841 606 1875
rect 640 1841 656 1875
rect 594 1807 656 1841
rect 594 1773 606 1807
rect 640 1773 656 1807
rect 594 1758 656 1773
rect 686 1943 752 1958
rect 686 1909 702 1943
rect 736 1909 752 1943
rect 686 1875 752 1909
rect 686 1841 702 1875
rect 736 1841 752 1875
rect 686 1807 752 1841
rect 686 1773 702 1807
rect 736 1773 752 1807
rect 686 1758 752 1773
rect 782 1943 844 1958
rect 782 1909 798 1943
rect 832 1909 844 1943
rect 1059 1941 1067 1975
rect 1101 1941 1111 1975
rect 1059 1923 1111 1941
rect 1141 1923 1183 2123
rect 1213 2111 1265 2123
rect 1213 2077 1223 2111
rect 1257 2077 1265 2111
rect 1213 2043 1265 2077
rect 1213 2009 1223 2043
rect 1257 2009 1265 2043
rect 1213 1975 1265 2009
rect 1213 1941 1223 1975
rect 1257 1941 1265 1975
rect 1213 1923 1265 1941
rect 2133 2111 2185 2123
rect 2133 2077 2141 2111
rect 2175 2077 2185 2111
rect 2133 2043 2185 2077
rect 2133 2009 2141 2043
rect 2175 2009 2185 2043
rect 2133 1975 2185 2009
rect 2133 1941 2141 1975
rect 2175 1941 2185 1975
rect 2133 1923 2185 1941
rect 2215 1923 2257 2123
rect 2287 2111 2339 2123
rect 2287 2077 2297 2111
rect 2331 2077 2339 2111
rect 2947 2111 2999 2123
rect 2287 2043 2339 2077
rect 2947 2077 2955 2111
rect 2989 2077 2999 2111
rect 2287 2009 2297 2043
rect 2331 2009 2339 2043
rect 2287 1975 2339 2009
rect 2947 2043 2999 2077
rect 2947 2009 2955 2043
rect 2989 2009 2999 2043
rect 2287 1941 2297 1975
rect 2331 1941 2339 1975
rect 2947 1975 2999 2009
rect 2287 1923 2339 1941
rect 2482 1943 2544 1958
rect 782 1875 844 1909
rect 782 1841 798 1875
rect 832 1841 844 1875
rect 782 1807 844 1841
rect 782 1773 798 1807
rect 832 1773 844 1807
rect 2482 1909 2494 1943
rect 2528 1909 2544 1943
rect 2482 1875 2544 1909
rect 2482 1841 2494 1875
rect 2528 1841 2544 1875
rect 2482 1807 2544 1841
rect 782 1758 844 1773
rect 2482 1773 2494 1807
rect 2528 1773 2544 1807
rect 2482 1758 2544 1773
rect 2574 1943 2640 1958
rect 2574 1909 2590 1943
rect 2624 1909 2640 1943
rect 2574 1875 2640 1909
rect 2574 1841 2590 1875
rect 2624 1841 2640 1875
rect 2574 1807 2640 1841
rect 2574 1773 2590 1807
rect 2624 1773 2640 1807
rect 2574 1758 2640 1773
rect 2670 1943 2732 1958
rect 2670 1909 2686 1943
rect 2720 1909 2732 1943
rect 2947 1941 2955 1975
rect 2989 1941 2999 1975
rect 2947 1923 2999 1941
rect 3029 1923 3071 2123
rect 3101 2111 3153 2123
rect 3101 2077 3111 2111
rect 3145 2077 3153 2111
rect 3101 2043 3153 2077
rect 3101 2009 3111 2043
rect 3145 2009 3153 2043
rect 3101 1975 3153 2009
rect 3101 1941 3111 1975
rect 3145 1941 3153 1975
rect 3101 1923 3153 1941
rect 4021 2111 4073 2123
rect 4021 2077 4029 2111
rect 4063 2077 4073 2111
rect 4021 2043 4073 2077
rect 4021 2009 4029 2043
rect 4063 2009 4073 2043
rect 4021 1975 4073 2009
rect 4021 1941 4029 1975
rect 4063 1941 4073 1975
rect 4021 1923 4073 1941
rect 4103 1923 4145 2123
rect 4175 2111 4227 2123
rect 4175 2077 4185 2111
rect 4219 2077 4227 2111
rect 4835 2111 4887 2123
rect 4175 2043 4227 2077
rect 4835 2077 4843 2111
rect 4877 2077 4887 2111
rect 4175 2009 4185 2043
rect 4219 2009 4227 2043
rect 4175 1975 4227 2009
rect 4835 2043 4887 2077
rect 4835 2009 4843 2043
rect 4877 2009 4887 2043
rect 4175 1941 4185 1975
rect 4219 1941 4227 1975
rect 4835 1975 4887 2009
rect 4175 1923 4227 1941
rect 4370 1943 4432 1958
rect 2670 1875 2732 1909
rect 2670 1841 2686 1875
rect 2720 1841 2732 1875
rect 2670 1807 2732 1841
rect 2670 1773 2686 1807
rect 2720 1773 2732 1807
rect 4370 1909 4382 1943
rect 4416 1909 4432 1943
rect 4370 1875 4432 1909
rect 4370 1841 4382 1875
rect 4416 1841 4432 1875
rect 4370 1807 4432 1841
rect 2670 1758 2732 1773
rect 4370 1773 4382 1807
rect 4416 1773 4432 1807
rect 4370 1758 4432 1773
rect 4462 1943 4528 1958
rect 4462 1909 4478 1943
rect 4512 1909 4528 1943
rect 4462 1875 4528 1909
rect 4462 1841 4478 1875
rect 4512 1841 4528 1875
rect 4462 1807 4528 1841
rect 4462 1773 4478 1807
rect 4512 1773 4528 1807
rect 4462 1758 4528 1773
rect 4558 1943 4620 1958
rect 4558 1909 4574 1943
rect 4608 1909 4620 1943
rect 4835 1941 4843 1975
rect 4877 1941 4887 1975
rect 4835 1923 4887 1941
rect 4917 1923 4959 2123
rect 4989 2111 5041 2123
rect 4989 2077 4999 2111
rect 5033 2077 5041 2111
rect 4989 2043 5041 2077
rect 4989 2009 4999 2043
rect 5033 2009 5041 2043
rect 4989 1975 5041 2009
rect 4989 1941 4999 1975
rect 5033 1941 5041 1975
rect 4989 1923 5041 1941
rect 5909 2111 5961 2123
rect 5909 2077 5917 2111
rect 5951 2077 5961 2111
rect 5909 2043 5961 2077
rect 5909 2009 5917 2043
rect 5951 2009 5961 2043
rect 5909 1975 5961 2009
rect 5909 1941 5917 1975
rect 5951 1941 5961 1975
rect 5909 1923 5961 1941
rect 5991 1923 6033 2123
rect 6063 2111 6115 2123
rect 6063 2077 6073 2111
rect 6107 2077 6115 2111
rect 6723 2111 6775 2123
rect 6063 2043 6115 2077
rect 6723 2077 6731 2111
rect 6765 2077 6775 2111
rect 6063 2009 6073 2043
rect 6107 2009 6115 2043
rect 6063 1975 6115 2009
rect 6723 2043 6775 2077
rect 6723 2009 6731 2043
rect 6765 2009 6775 2043
rect 6063 1941 6073 1975
rect 6107 1941 6115 1975
rect 6723 1975 6775 2009
rect 6063 1923 6115 1941
rect 6258 1943 6320 1958
rect 4558 1875 4620 1909
rect 4558 1841 4574 1875
rect 4608 1841 4620 1875
rect 4558 1807 4620 1841
rect 4558 1773 4574 1807
rect 4608 1773 4620 1807
rect 6258 1909 6270 1943
rect 6304 1909 6320 1943
rect 6258 1875 6320 1909
rect 6258 1841 6270 1875
rect 6304 1841 6320 1875
rect 6258 1807 6320 1841
rect 4558 1758 4620 1773
rect 6258 1773 6270 1807
rect 6304 1773 6320 1807
rect 6258 1758 6320 1773
rect 6350 1943 6416 1958
rect 6350 1909 6366 1943
rect 6400 1909 6416 1943
rect 6350 1875 6416 1909
rect 6350 1841 6366 1875
rect 6400 1841 6416 1875
rect 6350 1807 6416 1841
rect 6350 1773 6366 1807
rect 6400 1773 6416 1807
rect 6350 1758 6416 1773
rect 6446 1943 6508 1958
rect 6446 1909 6462 1943
rect 6496 1909 6508 1943
rect 6723 1941 6731 1975
rect 6765 1941 6775 1975
rect 6723 1923 6775 1941
rect 6805 1923 6847 2123
rect 6877 2111 6929 2123
rect 6877 2077 6887 2111
rect 6921 2077 6929 2111
rect 6877 2043 6929 2077
rect 6877 2009 6887 2043
rect 6921 2009 6929 2043
rect 6877 1975 6929 2009
rect 6877 1941 6887 1975
rect 6921 1941 6929 1975
rect 6877 1923 6929 1941
rect 7797 2111 7849 2123
rect 7797 2077 7805 2111
rect 7839 2077 7849 2111
rect 7797 2043 7849 2077
rect 7797 2009 7805 2043
rect 7839 2009 7849 2043
rect 7797 1975 7849 2009
rect 7797 1941 7805 1975
rect 7839 1941 7849 1975
rect 7797 1923 7849 1941
rect 7879 1923 7921 2123
rect 7951 2111 8003 2123
rect 7951 2077 7961 2111
rect 7995 2077 8003 2111
rect 8611 2111 8663 2123
rect 7951 2043 8003 2077
rect 8611 2077 8619 2111
rect 8653 2077 8663 2111
rect 7951 2009 7961 2043
rect 7995 2009 8003 2043
rect 7951 1975 8003 2009
rect 8611 2043 8663 2077
rect 8611 2009 8619 2043
rect 8653 2009 8663 2043
rect 7951 1941 7961 1975
rect 7995 1941 8003 1975
rect 8611 1975 8663 2009
rect 7951 1923 8003 1941
rect 8146 1943 8208 1958
rect 6446 1875 6508 1909
rect 6446 1841 6462 1875
rect 6496 1841 6508 1875
rect 6446 1807 6508 1841
rect 6446 1773 6462 1807
rect 6496 1773 6508 1807
rect 8146 1909 8158 1943
rect 8192 1909 8208 1943
rect 8146 1875 8208 1909
rect 8146 1841 8158 1875
rect 8192 1841 8208 1875
rect 8146 1807 8208 1841
rect 6446 1758 6508 1773
rect 8146 1773 8158 1807
rect 8192 1773 8208 1807
rect 8146 1758 8208 1773
rect 8238 1943 8304 1958
rect 8238 1909 8254 1943
rect 8288 1909 8304 1943
rect 8238 1875 8304 1909
rect 8238 1841 8254 1875
rect 8288 1841 8304 1875
rect 8238 1807 8304 1841
rect 8238 1773 8254 1807
rect 8288 1773 8304 1807
rect 8238 1758 8304 1773
rect 8334 1943 8396 1958
rect 8334 1909 8350 1943
rect 8384 1909 8396 1943
rect 8611 1941 8619 1975
rect 8653 1941 8663 1975
rect 8611 1923 8663 1941
rect 8693 1923 8735 2123
rect 8765 2111 8817 2123
rect 8765 2077 8775 2111
rect 8809 2077 8817 2111
rect 8765 2043 8817 2077
rect 8765 2009 8775 2043
rect 8809 2009 8817 2043
rect 8765 1975 8817 2009
rect 8765 1941 8775 1975
rect 8809 1941 8817 1975
rect 8765 1923 8817 1941
rect 9685 2111 9737 2123
rect 9685 2077 9693 2111
rect 9727 2077 9737 2111
rect 9685 2043 9737 2077
rect 9685 2009 9693 2043
rect 9727 2009 9737 2043
rect 9685 1975 9737 2009
rect 9685 1941 9693 1975
rect 9727 1941 9737 1975
rect 9685 1923 9737 1941
rect 9767 1923 9809 2123
rect 9839 2111 9891 2123
rect 9839 2077 9849 2111
rect 9883 2077 9891 2111
rect 10499 2111 10551 2123
rect 9839 2043 9891 2077
rect 10499 2077 10507 2111
rect 10541 2077 10551 2111
rect 9839 2009 9849 2043
rect 9883 2009 9891 2043
rect 9839 1975 9891 2009
rect 10499 2043 10551 2077
rect 10499 2009 10507 2043
rect 10541 2009 10551 2043
rect 9839 1941 9849 1975
rect 9883 1941 9891 1975
rect 10499 1975 10551 2009
rect 9839 1923 9891 1941
rect 10034 1943 10096 1958
rect 8334 1875 8396 1909
rect 8334 1841 8350 1875
rect 8384 1841 8396 1875
rect 8334 1807 8396 1841
rect 8334 1773 8350 1807
rect 8384 1773 8396 1807
rect 10034 1909 10046 1943
rect 10080 1909 10096 1943
rect 10034 1875 10096 1909
rect 10034 1841 10046 1875
rect 10080 1841 10096 1875
rect 10034 1807 10096 1841
rect 8334 1758 8396 1773
rect 10034 1773 10046 1807
rect 10080 1773 10096 1807
rect 10034 1758 10096 1773
rect 10126 1943 10192 1958
rect 10126 1909 10142 1943
rect 10176 1909 10192 1943
rect 10126 1875 10192 1909
rect 10126 1841 10142 1875
rect 10176 1841 10192 1875
rect 10126 1807 10192 1841
rect 10126 1773 10142 1807
rect 10176 1773 10192 1807
rect 10126 1758 10192 1773
rect 10222 1943 10284 1958
rect 10222 1909 10238 1943
rect 10272 1909 10284 1943
rect 10499 1941 10507 1975
rect 10541 1941 10551 1975
rect 10499 1923 10551 1941
rect 10581 1923 10623 2123
rect 10653 2111 10705 2123
rect 10653 2077 10663 2111
rect 10697 2077 10705 2111
rect 10653 2043 10705 2077
rect 10653 2009 10663 2043
rect 10697 2009 10705 2043
rect 10653 1975 10705 2009
rect 10653 1941 10663 1975
rect 10697 1941 10705 1975
rect 10653 1923 10705 1941
rect 11573 2111 11625 2123
rect 11573 2077 11581 2111
rect 11615 2077 11625 2111
rect 11573 2043 11625 2077
rect 11573 2009 11581 2043
rect 11615 2009 11625 2043
rect 11573 1975 11625 2009
rect 11573 1941 11581 1975
rect 11615 1941 11625 1975
rect 11573 1923 11625 1941
rect 11655 1923 11697 2123
rect 11727 2111 11779 2123
rect 11727 2077 11737 2111
rect 11771 2077 11779 2111
rect 12387 2111 12439 2123
rect 11727 2043 11779 2077
rect 12387 2077 12395 2111
rect 12429 2077 12439 2111
rect 11727 2009 11737 2043
rect 11771 2009 11779 2043
rect 11727 1975 11779 2009
rect 12387 2043 12439 2077
rect 12387 2009 12395 2043
rect 12429 2009 12439 2043
rect 11727 1941 11737 1975
rect 11771 1941 11779 1975
rect 12387 1975 12439 2009
rect 11727 1923 11779 1941
rect 11922 1943 11984 1958
rect 10222 1875 10284 1909
rect 10222 1841 10238 1875
rect 10272 1841 10284 1875
rect 10222 1807 10284 1841
rect 10222 1773 10238 1807
rect 10272 1773 10284 1807
rect 11922 1909 11934 1943
rect 11968 1909 11984 1943
rect 11922 1875 11984 1909
rect 11922 1841 11934 1875
rect 11968 1841 11984 1875
rect 11922 1807 11984 1841
rect 10222 1758 10284 1773
rect 11922 1773 11934 1807
rect 11968 1773 11984 1807
rect 11922 1758 11984 1773
rect 12014 1943 12080 1958
rect 12014 1909 12030 1943
rect 12064 1909 12080 1943
rect 12014 1875 12080 1909
rect 12014 1841 12030 1875
rect 12064 1841 12080 1875
rect 12014 1807 12080 1841
rect 12014 1773 12030 1807
rect 12064 1773 12080 1807
rect 12014 1758 12080 1773
rect 12110 1943 12172 1958
rect 12110 1909 12126 1943
rect 12160 1909 12172 1943
rect 12387 1941 12395 1975
rect 12429 1941 12439 1975
rect 12387 1923 12439 1941
rect 12469 1923 12511 2123
rect 12541 2111 12593 2123
rect 12541 2077 12551 2111
rect 12585 2077 12593 2111
rect 12541 2043 12593 2077
rect 12541 2009 12551 2043
rect 12585 2009 12593 2043
rect 12541 1975 12593 2009
rect 12541 1941 12551 1975
rect 12585 1941 12593 1975
rect 12541 1923 12593 1941
rect 13461 2111 13513 2123
rect 13461 2077 13469 2111
rect 13503 2077 13513 2111
rect 13461 2043 13513 2077
rect 13461 2009 13469 2043
rect 13503 2009 13513 2043
rect 13461 1975 13513 2009
rect 13461 1941 13469 1975
rect 13503 1941 13513 1975
rect 13461 1923 13513 1941
rect 13543 1923 13585 2123
rect 13615 2111 13667 2123
rect 13615 2077 13625 2111
rect 13659 2077 13667 2111
rect 14275 2111 14327 2123
rect 13615 2043 13667 2077
rect 14275 2077 14283 2111
rect 14317 2077 14327 2111
rect 13615 2009 13625 2043
rect 13659 2009 13667 2043
rect 13615 1975 13667 2009
rect 14275 2043 14327 2077
rect 14275 2009 14283 2043
rect 14317 2009 14327 2043
rect 13615 1941 13625 1975
rect 13659 1941 13667 1975
rect 14275 1975 14327 2009
rect 13615 1923 13667 1941
rect 13810 1943 13872 1958
rect 12110 1875 12172 1909
rect 12110 1841 12126 1875
rect 12160 1841 12172 1875
rect 12110 1807 12172 1841
rect 12110 1773 12126 1807
rect 12160 1773 12172 1807
rect 13810 1909 13822 1943
rect 13856 1909 13872 1943
rect 13810 1875 13872 1909
rect 13810 1841 13822 1875
rect 13856 1841 13872 1875
rect 13810 1807 13872 1841
rect 12110 1758 12172 1773
rect 13810 1773 13822 1807
rect 13856 1773 13872 1807
rect 13810 1758 13872 1773
rect 13902 1943 13968 1958
rect 13902 1909 13918 1943
rect 13952 1909 13968 1943
rect 13902 1875 13968 1909
rect 13902 1841 13918 1875
rect 13952 1841 13968 1875
rect 13902 1807 13968 1841
rect 13902 1773 13918 1807
rect 13952 1773 13968 1807
rect 13902 1758 13968 1773
rect 13998 1943 14060 1958
rect 13998 1909 14014 1943
rect 14048 1909 14060 1943
rect 14275 1941 14283 1975
rect 14317 1941 14327 1975
rect 14275 1923 14327 1941
rect 14357 1923 14399 2123
rect 14429 2111 14481 2123
rect 14429 2077 14439 2111
rect 14473 2077 14481 2111
rect 14429 2043 14481 2077
rect 14429 2009 14439 2043
rect 14473 2009 14481 2043
rect 14429 1975 14481 2009
rect 14429 1941 14439 1975
rect 14473 1941 14481 1975
rect 14429 1923 14481 1941
rect 15343 2111 15395 2123
rect 15343 2077 15351 2111
rect 15385 2077 15395 2111
rect 15343 2043 15395 2077
rect 15343 2009 15351 2043
rect 15385 2009 15395 2043
rect 15343 1975 15395 2009
rect 15343 1941 15351 1975
rect 15385 1941 15395 1975
rect 15343 1923 15395 1941
rect 15425 1923 15467 2123
rect 15497 2111 15549 2123
rect 15497 2077 15507 2111
rect 15541 2077 15549 2111
rect 16157 2111 16209 2123
rect 15497 2043 15549 2077
rect 16157 2077 16165 2111
rect 16199 2077 16209 2111
rect 15497 2009 15507 2043
rect 15541 2009 15549 2043
rect 15497 1975 15549 2009
rect 16157 2043 16209 2077
rect 16157 2009 16165 2043
rect 16199 2009 16209 2043
rect 15497 1941 15507 1975
rect 15541 1941 15549 1975
rect 16157 1975 16209 2009
rect 15497 1923 15549 1941
rect 15692 1943 15754 1958
rect 13998 1875 14060 1909
rect 13998 1841 14014 1875
rect 14048 1841 14060 1875
rect 13998 1807 14060 1841
rect 13998 1773 14014 1807
rect 14048 1773 14060 1807
rect 15692 1909 15704 1943
rect 15738 1909 15754 1943
rect 15692 1875 15754 1909
rect 15692 1841 15704 1875
rect 15738 1841 15754 1875
rect 15692 1807 15754 1841
rect 13998 1758 14060 1773
rect 15692 1773 15704 1807
rect 15738 1773 15754 1807
rect 15692 1758 15754 1773
rect 15784 1943 15850 1958
rect 15784 1909 15800 1943
rect 15834 1909 15850 1943
rect 15784 1875 15850 1909
rect 15784 1841 15800 1875
rect 15834 1841 15850 1875
rect 15784 1807 15850 1841
rect 15784 1773 15800 1807
rect 15834 1773 15850 1807
rect 15784 1758 15850 1773
rect 15880 1943 15942 1958
rect 15880 1909 15896 1943
rect 15930 1909 15942 1943
rect 16157 1941 16165 1975
rect 16199 1941 16209 1975
rect 16157 1923 16209 1941
rect 16239 1923 16281 2123
rect 16311 2111 16363 2123
rect 16311 2077 16321 2111
rect 16355 2077 16363 2111
rect 16311 2043 16363 2077
rect 16311 2009 16321 2043
rect 16355 2009 16363 2043
rect 16311 1975 16363 2009
rect 16311 1941 16321 1975
rect 16355 1941 16363 1975
rect 16311 1923 16363 1941
rect 17231 2111 17283 2123
rect 17231 2077 17239 2111
rect 17273 2077 17283 2111
rect 17231 2043 17283 2077
rect 17231 2009 17239 2043
rect 17273 2009 17283 2043
rect 17231 1975 17283 2009
rect 17231 1941 17239 1975
rect 17273 1941 17283 1975
rect 17231 1923 17283 1941
rect 17313 1923 17355 2123
rect 17385 2111 17437 2123
rect 17385 2077 17395 2111
rect 17429 2077 17437 2111
rect 18045 2111 18097 2123
rect 17385 2043 17437 2077
rect 18045 2077 18053 2111
rect 18087 2077 18097 2111
rect 17385 2009 17395 2043
rect 17429 2009 17437 2043
rect 17385 1975 17437 2009
rect 18045 2043 18097 2077
rect 18045 2009 18053 2043
rect 18087 2009 18097 2043
rect 17385 1941 17395 1975
rect 17429 1941 17437 1975
rect 18045 1975 18097 2009
rect 17385 1923 17437 1941
rect 17580 1943 17642 1958
rect 15880 1875 15942 1909
rect 15880 1841 15896 1875
rect 15930 1841 15942 1875
rect 15880 1807 15942 1841
rect 15880 1773 15896 1807
rect 15930 1773 15942 1807
rect 17580 1909 17592 1943
rect 17626 1909 17642 1943
rect 17580 1875 17642 1909
rect 17580 1841 17592 1875
rect 17626 1841 17642 1875
rect 17580 1807 17642 1841
rect 15880 1758 15942 1773
rect 17580 1773 17592 1807
rect 17626 1773 17642 1807
rect 17580 1758 17642 1773
rect 17672 1943 17738 1958
rect 17672 1909 17688 1943
rect 17722 1909 17738 1943
rect 17672 1875 17738 1909
rect 17672 1841 17688 1875
rect 17722 1841 17738 1875
rect 17672 1807 17738 1841
rect 17672 1773 17688 1807
rect 17722 1773 17738 1807
rect 17672 1758 17738 1773
rect 17768 1943 17830 1958
rect 17768 1909 17784 1943
rect 17818 1909 17830 1943
rect 18045 1941 18053 1975
rect 18087 1941 18097 1975
rect 18045 1923 18097 1941
rect 18127 1923 18169 2123
rect 18199 2111 18251 2123
rect 18199 2077 18209 2111
rect 18243 2077 18251 2111
rect 18199 2043 18251 2077
rect 18199 2009 18209 2043
rect 18243 2009 18251 2043
rect 18199 1975 18251 2009
rect 18199 1941 18209 1975
rect 18243 1941 18251 1975
rect 18199 1923 18251 1941
rect 19119 2111 19171 2123
rect 19119 2077 19127 2111
rect 19161 2077 19171 2111
rect 19119 2043 19171 2077
rect 19119 2009 19127 2043
rect 19161 2009 19171 2043
rect 19119 1975 19171 2009
rect 19119 1941 19127 1975
rect 19161 1941 19171 1975
rect 19119 1923 19171 1941
rect 19201 1923 19243 2123
rect 19273 2111 19325 2123
rect 19273 2077 19283 2111
rect 19317 2077 19325 2111
rect 19933 2111 19985 2123
rect 19273 2043 19325 2077
rect 19933 2077 19941 2111
rect 19975 2077 19985 2111
rect 19273 2009 19283 2043
rect 19317 2009 19325 2043
rect 19273 1975 19325 2009
rect 19933 2043 19985 2077
rect 19933 2009 19941 2043
rect 19975 2009 19985 2043
rect 19273 1941 19283 1975
rect 19317 1941 19325 1975
rect 19933 1975 19985 2009
rect 19273 1923 19325 1941
rect 19468 1943 19530 1958
rect 17768 1875 17830 1909
rect 17768 1841 17784 1875
rect 17818 1841 17830 1875
rect 17768 1807 17830 1841
rect 17768 1773 17784 1807
rect 17818 1773 17830 1807
rect 19468 1909 19480 1943
rect 19514 1909 19530 1943
rect 19468 1875 19530 1909
rect 19468 1841 19480 1875
rect 19514 1841 19530 1875
rect 19468 1807 19530 1841
rect 17768 1758 17830 1773
rect 19468 1773 19480 1807
rect 19514 1773 19530 1807
rect 19468 1758 19530 1773
rect 19560 1943 19626 1958
rect 19560 1909 19576 1943
rect 19610 1909 19626 1943
rect 19560 1875 19626 1909
rect 19560 1841 19576 1875
rect 19610 1841 19626 1875
rect 19560 1807 19626 1841
rect 19560 1773 19576 1807
rect 19610 1773 19626 1807
rect 19560 1758 19626 1773
rect 19656 1943 19718 1958
rect 19656 1909 19672 1943
rect 19706 1909 19718 1943
rect 19933 1941 19941 1975
rect 19975 1941 19985 1975
rect 19933 1923 19985 1941
rect 20015 1923 20057 2123
rect 20087 2111 20139 2123
rect 20087 2077 20097 2111
rect 20131 2077 20139 2111
rect 20087 2043 20139 2077
rect 20087 2009 20097 2043
rect 20131 2009 20139 2043
rect 20087 1975 20139 2009
rect 20087 1941 20097 1975
rect 20131 1941 20139 1975
rect 20087 1923 20139 1941
rect 21007 2111 21059 2123
rect 21007 2077 21015 2111
rect 21049 2077 21059 2111
rect 21007 2043 21059 2077
rect 21007 2009 21015 2043
rect 21049 2009 21059 2043
rect 21007 1975 21059 2009
rect 21007 1941 21015 1975
rect 21049 1941 21059 1975
rect 21007 1923 21059 1941
rect 21089 1923 21131 2123
rect 21161 2111 21213 2123
rect 21161 2077 21171 2111
rect 21205 2077 21213 2111
rect 21821 2111 21873 2123
rect 21161 2043 21213 2077
rect 21821 2077 21829 2111
rect 21863 2077 21873 2111
rect 21161 2009 21171 2043
rect 21205 2009 21213 2043
rect 21161 1975 21213 2009
rect 21821 2043 21873 2077
rect 21821 2009 21829 2043
rect 21863 2009 21873 2043
rect 21161 1941 21171 1975
rect 21205 1941 21213 1975
rect 21821 1975 21873 2009
rect 21161 1923 21213 1941
rect 21356 1943 21418 1958
rect 19656 1875 19718 1909
rect 19656 1841 19672 1875
rect 19706 1841 19718 1875
rect 19656 1807 19718 1841
rect 19656 1773 19672 1807
rect 19706 1773 19718 1807
rect 21356 1909 21368 1943
rect 21402 1909 21418 1943
rect 21356 1875 21418 1909
rect 21356 1841 21368 1875
rect 21402 1841 21418 1875
rect 21356 1807 21418 1841
rect 19656 1758 19718 1773
rect 21356 1773 21368 1807
rect 21402 1773 21418 1807
rect 21356 1758 21418 1773
rect 21448 1943 21514 1958
rect 21448 1909 21464 1943
rect 21498 1909 21514 1943
rect 21448 1875 21514 1909
rect 21448 1841 21464 1875
rect 21498 1841 21514 1875
rect 21448 1807 21514 1841
rect 21448 1773 21464 1807
rect 21498 1773 21514 1807
rect 21448 1758 21514 1773
rect 21544 1943 21606 1958
rect 21544 1909 21560 1943
rect 21594 1909 21606 1943
rect 21821 1941 21829 1975
rect 21863 1941 21873 1975
rect 21821 1923 21873 1941
rect 21903 1923 21945 2123
rect 21975 2111 22027 2123
rect 21975 2077 21985 2111
rect 22019 2077 22027 2111
rect 21975 2043 22027 2077
rect 21975 2009 21985 2043
rect 22019 2009 22027 2043
rect 21975 1975 22027 2009
rect 21975 1941 21985 1975
rect 22019 1941 22027 1975
rect 21975 1923 22027 1941
rect 22895 2111 22947 2123
rect 22895 2077 22903 2111
rect 22937 2077 22947 2111
rect 22895 2043 22947 2077
rect 22895 2009 22903 2043
rect 22937 2009 22947 2043
rect 22895 1975 22947 2009
rect 22895 1941 22903 1975
rect 22937 1941 22947 1975
rect 22895 1923 22947 1941
rect 22977 1923 23019 2123
rect 23049 2111 23101 2123
rect 23049 2077 23059 2111
rect 23093 2077 23101 2111
rect 23709 2111 23761 2123
rect 23049 2043 23101 2077
rect 23709 2077 23717 2111
rect 23751 2077 23761 2111
rect 23049 2009 23059 2043
rect 23093 2009 23101 2043
rect 23049 1975 23101 2009
rect 23709 2043 23761 2077
rect 23709 2009 23717 2043
rect 23751 2009 23761 2043
rect 23049 1941 23059 1975
rect 23093 1941 23101 1975
rect 23709 1975 23761 2009
rect 23049 1923 23101 1941
rect 23244 1943 23306 1958
rect 21544 1875 21606 1909
rect 21544 1841 21560 1875
rect 21594 1841 21606 1875
rect 21544 1807 21606 1841
rect 21544 1773 21560 1807
rect 21594 1773 21606 1807
rect 23244 1909 23256 1943
rect 23290 1909 23306 1943
rect 23244 1875 23306 1909
rect 23244 1841 23256 1875
rect 23290 1841 23306 1875
rect 23244 1807 23306 1841
rect 21544 1758 21606 1773
rect 23244 1773 23256 1807
rect 23290 1773 23306 1807
rect 23244 1758 23306 1773
rect 23336 1943 23402 1958
rect 23336 1909 23352 1943
rect 23386 1909 23402 1943
rect 23336 1875 23402 1909
rect 23336 1841 23352 1875
rect 23386 1841 23402 1875
rect 23336 1807 23402 1841
rect 23336 1773 23352 1807
rect 23386 1773 23402 1807
rect 23336 1758 23402 1773
rect 23432 1943 23494 1958
rect 23432 1909 23448 1943
rect 23482 1909 23494 1943
rect 23709 1941 23717 1975
rect 23751 1941 23761 1975
rect 23709 1923 23761 1941
rect 23791 1923 23833 2123
rect 23863 2111 23915 2123
rect 23863 2077 23873 2111
rect 23907 2077 23915 2111
rect 23863 2043 23915 2077
rect 23863 2009 23873 2043
rect 23907 2009 23915 2043
rect 23863 1975 23915 2009
rect 23863 1941 23873 1975
rect 23907 1941 23915 1975
rect 23863 1923 23915 1941
rect 24783 2111 24835 2123
rect 24783 2077 24791 2111
rect 24825 2077 24835 2111
rect 24783 2043 24835 2077
rect 24783 2009 24791 2043
rect 24825 2009 24835 2043
rect 24783 1975 24835 2009
rect 24783 1941 24791 1975
rect 24825 1941 24835 1975
rect 24783 1923 24835 1941
rect 24865 1923 24907 2123
rect 24937 2111 24989 2123
rect 24937 2077 24947 2111
rect 24981 2077 24989 2111
rect 25597 2111 25649 2123
rect 24937 2043 24989 2077
rect 25597 2077 25605 2111
rect 25639 2077 25649 2111
rect 24937 2009 24947 2043
rect 24981 2009 24989 2043
rect 24937 1975 24989 2009
rect 25597 2043 25649 2077
rect 25597 2009 25605 2043
rect 25639 2009 25649 2043
rect 24937 1941 24947 1975
rect 24981 1941 24989 1975
rect 25597 1975 25649 2009
rect 24937 1923 24989 1941
rect 25132 1943 25194 1958
rect 23432 1875 23494 1909
rect 23432 1841 23448 1875
rect 23482 1841 23494 1875
rect 23432 1807 23494 1841
rect 23432 1773 23448 1807
rect 23482 1773 23494 1807
rect 25132 1909 25144 1943
rect 25178 1909 25194 1943
rect 25132 1875 25194 1909
rect 25132 1841 25144 1875
rect 25178 1841 25194 1875
rect 25132 1807 25194 1841
rect 23432 1758 23494 1773
rect 25132 1773 25144 1807
rect 25178 1773 25194 1807
rect 25132 1758 25194 1773
rect 25224 1943 25290 1958
rect 25224 1909 25240 1943
rect 25274 1909 25290 1943
rect 25224 1875 25290 1909
rect 25224 1841 25240 1875
rect 25274 1841 25290 1875
rect 25224 1807 25290 1841
rect 25224 1773 25240 1807
rect 25274 1773 25290 1807
rect 25224 1758 25290 1773
rect 25320 1943 25382 1958
rect 25320 1909 25336 1943
rect 25370 1909 25382 1943
rect 25597 1941 25605 1975
rect 25639 1941 25649 1975
rect 25597 1923 25649 1941
rect 25679 1923 25721 2123
rect 25751 2111 25803 2123
rect 25751 2077 25761 2111
rect 25795 2077 25803 2111
rect 25751 2043 25803 2077
rect 25751 2009 25761 2043
rect 25795 2009 25803 2043
rect 25751 1975 25803 2009
rect 25751 1941 25761 1975
rect 25795 1941 25803 1975
rect 25751 1923 25803 1941
rect 26671 2111 26723 2123
rect 26671 2077 26679 2111
rect 26713 2077 26723 2111
rect 26671 2043 26723 2077
rect 26671 2009 26679 2043
rect 26713 2009 26723 2043
rect 26671 1975 26723 2009
rect 26671 1941 26679 1975
rect 26713 1941 26723 1975
rect 26671 1923 26723 1941
rect 26753 1923 26795 2123
rect 26825 2111 26877 2123
rect 26825 2077 26835 2111
rect 26869 2077 26877 2111
rect 27485 2111 27537 2123
rect 26825 2043 26877 2077
rect 27485 2077 27493 2111
rect 27527 2077 27537 2111
rect 26825 2009 26835 2043
rect 26869 2009 26877 2043
rect 26825 1975 26877 2009
rect 27485 2043 27537 2077
rect 27485 2009 27493 2043
rect 27527 2009 27537 2043
rect 26825 1941 26835 1975
rect 26869 1941 26877 1975
rect 27485 1975 27537 2009
rect 26825 1923 26877 1941
rect 27020 1943 27082 1958
rect 25320 1875 25382 1909
rect 25320 1841 25336 1875
rect 25370 1841 25382 1875
rect 25320 1807 25382 1841
rect 25320 1773 25336 1807
rect 25370 1773 25382 1807
rect 27020 1909 27032 1943
rect 27066 1909 27082 1943
rect 27020 1875 27082 1909
rect 27020 1841 27032 1875
rect 27066 1841 27082 1875
rect 27020 1807 27082 1841
rect 25320 1758 25382 1773
rect 27020 1773 27032 1807
rect 27066 1773 27082 1807
rect 27020 1758 27082 1773
rect 27112 1943 27178 1958
rect 27112 1909 27128 1943
rect 27162 1909 27178 1943
rect 27112 1875 27178 1909
rect 27112 1841 27128 1875
rect 27162 1841 27178 1875
rect 27112 1807 27178 1841
rect 27112 1773 27128 1807
rect 27162 1773 27178 1807
rect 27112 1758 27178 1773
rect 27208 1943 27270 1958
rect 27208 1909 27224 1943
rect 27258 1909 27270 1943
rect 27485 1941 27493 1975
rect 27527 1941 27537 1975
rect 27485 1923 27537 1941
rect 27567 1923 27609 2123
rect 27639 2111 27691 2123
rect 27639 2077 27649 2111
rect 27683 2077 27691 2111
rect 27639 2043 27691 2077
rect 27639 2009 27649 2043
rect 27683 2009 27691 2043
rect 27639 1975 27691 2009
rect 27639 1941 27649 1975
rect 27683 1941 27691 1975
rect 27639 1923 27691 1941
rect 28559 2111 28611 2123
rect 28559 2077 28567 2111
rect 28601 2077 28611 2111
rect 28559 2043 28611 2077
rect 28559 2009 28567 2043
rect 28601 2009 28611 2043
rect 28559 1975 28611 2009
rect 28559 1941 28567 1975
rect 28601 1941 28611 1975
rect 28559 1923 28611 1941
rect 28641 1923 28683 2123
rect 28713 2111 28765 2123
rect 28713 2077 28723 2111
rect 28757 2077 28765 2111
rect 29373 2111 29425 2123
rect 28713 2043 28765 2077
rect 29373 2077 29381 2111
rect 29415 2077 29425 2111
rect 28713 2009 28723 2043
rect 28757 2009 28765 2043
rect 28713 1975 28765 2009
rect 29373 2043 29425 2077
rect 29373 2009 29381 2043
rect 29415 2009 29425 2043
rect 28713 1941 28723 1975
rect 28757 1941 28765 1975
rect 29373 1975 29425 2009
rect 28713 1923 28765 1941
rect 28908 1943 28970 1958
rect 27208 1875 27270 1909
rect 27208 1841 27224 1875
rect 27258 1841 27270 1875
rect 27208 1807 27270 1841
rect 27208 1773 27224 1807
rect 27258 1773 27270 1807
rect 28908 1909 28920 1943
rect 28954 1909 28970 1943
rect 28908 1875 28970 1909
rect 28908 1841 28920 1875
rect 28954 1841 28970 1875
rect 28908 1807 28970 1841
rect 27208 1758 27270 1773
rect 28908 1773 28920 1807
rect 28954 1773 28970 1807
rect 28908 1758 28970 1773
rect 29000 1943 29066 1958
rect 29000 1909 29016 1943
rect 29050 1909 29066 1943
rect 29000 1875 29066 1909
rect 29000 1841 29016 1875
rect 29050 1841 29066 1875
rect 29000 1807 29066 1841
rect 29000 1773 29016 1807
rect 29050 1773 29066 1807
rect 29000 1758 29066 1773
rect 29096 1943 29158 1958
rect 29096 1909 29112 1943
rect 29146 1909 29158 1943
rect 29373 1941 29381 1975
rect 29415 1941 29425 1975
rect 29373 1923 29425 1941
rect 29455 1923 29497 2123
rect 29527 2111 29579 2123
rect 29527 2077 29537 2111
rect 29571 2077 29579 2111
rect 29527 2043 29579 2077
rect 29527 2009 29537 2043
rect 29571 2009 29579 2043
rect 29527 1975 29579 2009
rect 29527 1941 29537 1975
rect 29571 1941 29579 1975
rect 29527 1923 29579 1941
rect 30447 2111 30499 2123
rect 30447 2077 30455 2111
rect 30489 2077 30499 2111
rect 30447 2043 30499 2077
rect 30447 2009 30455 2043
rect 30489 2009 30499 2043
rect 30447 1975 30499 2009
rect 30447 1941 30455 1975
rect 30489 1941 30499 1975
rect 30447 1923 30499 1941
rect 30529 1923 30571 2123
rect 30601 2111 30653 2123
rect 30601 2077 30611 2111
rect 30645 2077 30653 2111
rect 31261 2111 31313 2123
rect 30601 2043 30653 2077
rect 31261 2077 31269 2111
rect 31303 2077 31313 2111
rect 30601 2009 30611 2043
rect 30645 2009 30653 2043
rect 30601 1975 30653 2009
rect 31261 2043 31313 2077
rect 31261 2009 31269 2043
rect 31303 2009 31313 2043
rect 30601 1941 30611 1975
rect 30645 1941 30653 1975
rect 31261 1975 31313 2009
rect 30601 1923 30653 1941
rect 30796 1943 30858 1958
rect 29096 1875 29158 1909
rect 29096 1841 29112 1875
rect 29146 1841 29158 1875
rect 29096 1807 29158 1841
rect 29096 1773 29112 1807
rect 29146 1773 29158 1807
rect 30796 1909 30808 1943
rect 30842 1909 30858 1943
rect 30796 1875 30858 1909
rect 30796 1841 30808 1875
rect 30842 1841 30858 1875
rect 30796 1807 30858 1841
rect 29096 1758 29158 1773
rect 30796 1773 30808 1807
rect 30842 1773 30858 1807
rect 30796 1758 30858 1773
rect 30888 1943 30954 1958
rect 30888 1909 30904 1943
rect 30938 1909 30954 1943
rect 30888 1875 30954 1909
rect 30888 1841 30904 1875
rect 30938 1841 30954 1875
rect 30888 1807 30954 1841
rect 30888 1773 30904 1807
rect 30938 1773 30954 1807
rect 30888 1758 30954 1773
rect 30984 1943 31046 1958
rect 30984 1909 31000 1943
rect 31034 1909 31046 1943
rect 31261 1941 31269 1975
rect 31303 1941 31313 1975
rect 31261 1923 31313 1941
rect 31343 1923 31385 2123
rect 31415 2111 31467 2123
rect 31415 2077 31425 2111
rect 31459 2077 31467 2111
rect 31415 2043 31467 2077
rect 31415 2009 31425 2043
rect 31459 2009 31467 2043
rect 31415 1975 31467 2009
rect 31415 1941 31425 1975
rect 31459 1941 31467 1975
rect 31415 1923 31467 1941
rect 32335 2111 32387 2123
rect 32335 2077 32343 2111
rect 32377 2077 32387 2111
rect 32335 2043 32387 2077
rect 32335 2009 32343 2043
rect 32377 2009 32387 2043
rect 32335 1975 32387 2009
rect 32335 1941 32343 1975
rect 32377 1941 32387 1975
rect 32335 1923 32387 1941
rect 32417 1923 32459 2123
rect 32489 2111 32541 2123
rect 32489 2077 32499 2111
rect 32533 2077 32541 2111
rect 33149 2111 33201 2123
rect 32489 2043 32541 2077
rect 33149 2077 33157 2111
rect 33191 2077 33201 2111
rect 32489 2009 32499 2043
rect 32533 2009 32541 2043
rect 32489 1975 32541 2009
rect 33149 2043 33201 2077
rect 33149 2009 33157 2043
rect 33191 2009 33201 2043
rect 32489 1941 32499 1975
rect 32533 1941 32541 1975
rect 33149 1975 33201 2009
rect 32489 1923 32541 1941
rect 32684 1943 32746 1958
rect 30984 1875 31046 1909
rect 30984 1841 31000 1875
rect 31034 1841 31046 1875
rect 30984 1807 31046 1841
rect 30984 1773 31000 1807
rect 31034 1773 31046 1807
rect 32684 1909 32696 1943
rect 32730 1909 32746 1943
rect 32684 1875 32746 1909
rect 32684 1841 32696 1875
rect 32730 1841 32746 1875
rect 32684 1807 32746 1841
rect 30984 1758 31046 1773
rect 32684 1773 32696 1807
rect 32730 1773 32746 1807
rect 32684 1758 32746 1773
rect 32776 1943 32842 1958
rect 32776 1909 32792 1943
rect 32826 1909 32842 1943
rect 32776 1875 32842 1909
rect 32776 1841 32792 1875
rect 32826 1841 32842 1875
rect 32776 1807 32842 1841
rect 32776 1773 32792 1807
rect 32826 1773 32842 1807
rect 32776 1758 32842 1773
rect 32872 1943 32934 1958
rect 32872 1909 32888 1943
rect 32922 1909 32934 1943
rect 33149 1941 33157 1975
rect 33191 1941 33201 1975
rect 33149 1923 33201 1941
rect 33231 1923 33273 2123
rect 33303 2111 33355 2123
rect 33303 2077 33313 2111
rect 33347 2077 33355 2111
rect 33303 2043 33355 2077
rect 33303 2009 33313 2043
rect 33347 2009 33355 2043
rect 33303 1975 33355 2009
rect 33303 1941 33313 1975
rect 33347 1941 33355 1975
rect 33303 1923 33355 1941
rect 34223 2111 34275 2123
rect 34223 2077 34231 2111
rect 34265 2077 34275 2111
rect 34223 2043 34275 2077
rect 34223 2009 34231 2043
rect 34265 2009 34275 2043
rect 34223 1975 34275 2009
rect 34223 1941 34231 1975
rect 34265 1941 34275 1975
rect 34223 1923 34275 1941
rect 34305 1923 34347 2123
rect 34377 2111 34429 2123
rect 34377 2077 34387 2111
rect 34421 2077 34429 2111
rect 35037 2111 35089 2123
rect 34377 2043 34429 2077
rect 35037 2077 35045 2111
rect 35079 2077 35089 2111
rect 34377 2009 34387 2043
rect 34421 2009 34429 2043
rect 34377 1975 34429 2009
rect 35037 2043 35089 2077
rect 35037 2009 35045 2043
rect 35079 2009 35089 2043
rect 34377 1941 34387 1975
rect 34421 1941 34429 1975
rect 35037 1975 35089 2009
rect 34377 1923 34429 1941
rect 34572 1943 34634 1958
rect 32872 1875 32934 1909
rect 32872 1841 32888 1875
rect 32922 1841 32934 1875
rect 32872 1807 32934 1841
rect 32872 1773 32888 1807
rect 32922 1773 32934 1807
rect 34572 1909 34584 1943
rect 34618 1909 34634 1943
rect 34572 1875 34634 1909
rect 34572 1841 34584 1875
rect 34618 1841 34634 1875
rect 34572 1807 34634 1841
rect 32872 1758 32934 1773
rect 34572 1773 34584 1807
rect 34618 1773 34634 1807
rect 34572 1758 34634 1773
rect 34664 1943 34730 1958
rect 34664 1909 34680 1943
rect 34714 1909 34730 1943
rect 34664 1875 34730 1909
rect 34664 1841 34680 1875
rect 34714 1841 34730 1875
rect 34664 1807 34730 1841
rect 34664 1773 34680 1807
rect 34714 1773 34730 1807
rect 34664 1758 34730 1773
rect 34760 1943 34822 1958
rect 34760 1909 34776 1943
rect 34810 1909 34822 1943
rect 35037 1941 35045 1975
rect 35079 1941 35089 1975
rect 35037 1923 35089 1941
rect 35119 1923 35161 2123
rect 35191 2111 35243 2123
rect 35191 2077 35201 2111
rect 35235 2077 35243 2111
rect 35191 2043 35243 2077
rect 35191 2009 35201 2043
rect 35235 2009 35243 2043
rect 35191 1975 35243 2009
rect 35191 1941 35201 1975
rect 35235 1941 35243 1975
rect 35191 1923 35243 1941
rect 36111 2111 36163 2123
rect 36111 2077 36119 2111
rect 36153 2077 36163 2111
rect 36111 2043 36163 2077
rect 36111 2009 36119 2043
rect 36153 2009 36163 2043
rect 36111 1975 36163 2009
rect 36111 1941 36119 1975
rect 36153 1941 36163 1975
rect 36111 1923 36163 1941
rect 36193 1923 36235 2123
rect 36265 2111 36317 2123
rect 36265 2077 36275 2111
rect 36309 2077 36317 2111
rect 36925 2111 36977 2123
rect 36265 2043 36317 2077
rect 36925 2077 36933 2111
rect 36967 2077 36977 2111
rect 36265 2009 36275 2043
rect 36309 2009 36317 2043
rect 36265 1975 36317 2009
rect 36925 2043 36977 2077
rect 36925 2009 36933 2043
rect 36967 2009 36977 2043
rect 36265 1941 36275 1975
rect 36309 1941 36317 1975
rect 36925 1975 36977 2009
rect 36265 1923 36317 1941
rect 36460 1943 36522 1958
rect 34760 1875 34822 1909
rect 34760 1841 34776 1875
rect 34810 1841 34822 1875
rect 34760 1807 34822 1841
rect 34760 1773 34776 1807
rect 34810 1773 34822 1807
rect 36460 1909 36472 1943
rect 36506 1909 36522 1943
rect 36460 1875 36522 1909
rect 36460 1841 36472 1875
rect 36506 1841 36522 1875
rect 36460 1807 36522 1841
rect 34760 1758 34822 1773
rect 36460 1773 36472 1807
rect 36506 1773 36522 1807
rect 36460 1758 36522 1773
rect 36552 1943 36618 1958
rect 36552 1909 36568 1943
rect 36602 1909 36618 1943
rect 36552 1875 36618 1909
rect 36552 1841 36568 1875
rect 36602 1841 36618 1875
rect 36552 1807 36618 1841
rect 36552 1773 36568 1807
rect 36602 1773 36618 1807
rect 36552 1758 36618 1773
rect 36648 1943 36710 1958
rect 36648 1909 36664 1943
rect 36698 1909 36710 1943
rect 36925 1941 36933 1975
rect 36967 1941 36977 1975
rect 36925 1923 36977 1941
rect 37007 1923 37049 2123
rect 37079 2111 37131 2123
rect 37079 2077 37089 2111
rect 37123 2077 37131 2111
rect 37079 2043 37131 2077
rect 37079 2009 37089 2043
rect 37123 2009 37131 2043
rect 37079 1975 37131 2009
rect 37079 1941 37089 1975
rect 37123 1941 37131 1975
rect 37079 1923 37131 1941
rect 37999 2111 38051 2123
rect 37999 2077 38007 2111
rect 38041 2077 38051 2111
rect 37999 2043 38051 2077
rect 37999 2009 38007 2043
rect 38041 2009 38051 2043
rect 37999 1975 38051 2009
rect 37999 1941 38007 1975
rect 38041 1941 38051 1975
rect 37999 1923 38051 1941
rect 38081 1923 38123 2123
rect 38153 2111 38205 2123
rect 38153 2077 38163 2111
rect 38197 2077 38205 2111
rect 38813 2111 38865 2123
rect 38153 2043 38205 2077
rect 38813 2077 38821 2111
rect 38855 2077 38865 2111
rect 38153 2009 38163 2043
rect 38197 2009 38205 2043
rect 38153 1975 38205 2009
rect 38813 2043 38865 2077
rect 38813 2009 38821 2043
rect 38855 2009 38865 2043
rect 38153 1941 38163 1975
rect 38197 1941 38205 1975
rect 38813 1975 38865 2009
rect 38153 1923 38205 1941
rect 38348 1943 38410 1958
rect 36648 1875 36710 1909
rect 36648 1841 36664 1875
rect 36698 1841 36710 1875
rect 36648 1807 36710 1841
rect 36648 1773 36664 1807
rect 36698 1773 36710 1807
rect 38348 1909 38360 1943
rect 38394 1909 38410 1943
rect 38348 1875 38410 1909
rect 38348 1841 38360 1875
rect 38394 1841 38410 1875
rect 38348 1807 38410 1841
rect 36648 1758 36710 1773
rect 38348 1773 38360 1807
rect 38394 1773 38410 1807
rect 38348 1758 38410 1773
rect 38440 1943 38506 1958
rect 38440 1909 38456 1943
rect 38490 1909 38506 1943
rect 38440 1875 38506 1909
rect 38440 1841 38456 1875
rect 38490 1841 38506 1875
rect 38440 1807 38506 1841
rect 38440 1773 38456 1807
rect 38490 1773 38506 1807
rect 38440 1758 38506 1773
rect 38536 1943 38598 1958
rect 38536 1909 38552 1943
rect 38586 1909 38598 1943
rect 38813 1941 38821 1975
rect 38855 1941 38865 1975
rect 38813 1923 38865 1941
rect 38895 1923 38937 2123
rect 38967 2111 39019 2123
rect 38967 2077 38977 2111
rect 39011 2077 39019 2111
rect 38967 2043 39019 2077
rect 38967 2009 38977 2043
rect 39011 2009 39019 2043
rect 38967 1975 39019 2009
rect 38967 1941 38977 1975
rect 39011 1941 39019 1975
rect 38967 1923 39019 1941
rect 39887 2111 39939 2123
rect 39887 2077 39895 2111
rect 39929 2077 39939 2111
rect 39887 2043 39939 2077
rect 39887 2009 39895 2043
rect 39929 2009 39939 2043
rect 39887 1975 39939 2009
rect 39887 1941 39895 1975
rect 39929 1941 39939 1975
rect 39887 1923 39939 1941
rect 39969 1923 40011 2123
rect 40041 2111 40093 2123
rect 40041 2077 40051 2111
rect 40085 2077 40093 2111
rect 40701 2111 40753 2123
rect 40041 2043 40093 2077
rect 40701 2077 40709 2111
rect 40743 2077 40753 2111
rect 40041 2009 40051 2043
rect 40085 2009 40093 2043
rect 40041 1975 40093 2009
rect 40701 2043 40753 2077
rect 40701 2009 40709 2043
rect 40743 2009 40753 2043
rect 40041 1941 40051 1975
rect 40085 1941 40093 1975
rect 40701 1975 40753 2009
rect 40041 1923 40093 1941
rect 40236 1943 40298 1958
rect 38536 1875 38598 1909
rect 38536 1841 38552 1875
rect 38586 1841 38598 1875
rect 38536 1807 38598 1841
rect 38536 1773 38552 1807
rect 38586 1773 38598 1807
rect 40236 1909 40248 1943
rect 40282 1909 40298 1943
rect 40236 1875 40298 1909
rect 40236 1841 40248 1875
rect 40282 1841 40298 1875
rect 40236 1807 40298 1841
rect 38536 1758 38598 1773
rect 40236 1773 40248 1807
rect 40282 1773 40298 1807
rect 40236 1758 40298 1773
rect 40328 1943 40394 1958
rect 40328 1909 40344 1943
rect 40378 1909 40394 1943
rect 40328 1875 40394 1909
rect 40328 1841 40344 1875
rect 40378 1841 40394 1875
rect 40328 1807 40394 1841
rect 40328 1773 40344 1807
rect 40378 1773 40394 1807
rect 40328 1758 40394 1773
rect 40424 1943 40486 1958
rect 40424 1909 40440 1943
rect 40474 1909 40486 1943
rect 40701 1941 40709 1975
rect 40743 1941 40753 1975
rect 40701 1923 40753 1941
rect 40783 1923 40825 2123
rect 40855 2111 40907 2123
rect 40855 2077 40865 2111
rect 40899 2077 40907 2111
rect 40855 2043 40907 2077
rect 40855 2009 40865 2043
rect 40899 2009 40907 2043
rect 40855 1975 40907 2009
rect 40855 1941 40865 1975
rect 40899 1941 40907 1975
rect 40855 1923 40907 1941
rect 41775 2111 41827 2123
rect 41775 2077 41783 2111
rect 41817 2077 41827 2111
rect 41775 2043 41827 2077
rect 41775 2009 41783 2043
rect 41817 2009 41827 2043
rect 41775 1975 41827 2009
rect 41775 1941 41783 1975
rect 41817 1941 41827 1975
rect 41775 1923 41827 1941
rect 41857 1923 41899 2123
rect 41929 2111 41981 2123
rect 41929 2077 41939 2111
rect 41973 2077 41981 2111
rect 42589 2111 42641 2123
rect 41929 2043 41981 2077
rect 42589 2077 42597 2111
rect 42631 2077 42641 2111
rect 41929 2009 41939 2043
rect 41973 2009 41981 2043
rect 41929 1975 41981 2009
rect 42589 2043 42641 2077
rect 42589 2009 42597 2043
rect 42631 2009 42641 2043
rect 41929 1941 41939 1975
rect 41973 1941 41981 1975
rect 42589 1975 42641 2009
rect 41929 1923 41981 1941
rect 42124 1943 42186 1958
rect 40424 1875 40486 1909
rect 40424 1841 40440 1875
rect 40474 1841 40486 1875
rect 40424 1807 40486 1841
rect 40424 1773 40440 1807
rect 40474 1773 40486 1807
rect 42124 1909 42136 1943
rect 42170 1909 42186 1943
rect 42124 1875 42186 1909
rect 42124 1841 42136 1875
rect 42170 1841 42186 1875
rect 42124 1807 42186 1841
rect 40424 1758 40486 1773
rect 42124 1773 42136 1807
rect 42170 1773 42186 1807
rect 42124 1758 42186 1773
rect 42216 1943 42282 1958
rect 42216 1909 42232 1943
rect 42266 1909 42282 1943
rect 42216 1875 42282 1909
rect 42216 1841 42232 1875
rect 42266 1841 42282 1875
rect 42216 1807 42282 1841
rect 42216 1773 42232 1807
rect 42266 1773 42282 1807
rect 42216 1758 42282 1773
rect 42312 1943 42374 1958
rect 42312 1909 42328 1943
rect 42362 1909 42374 1943
rect 42589 1941 42597 1975
rect 42631 1941 42641 1975
rect 42589 1923 42641 1941
rect 42671 1923 42713 2123
rect 42743 2111 42795 2123
rect 42743 2077 42753 2111
rect 42787 2077 42795 2111
rect 42743 2043 42795 2077
rect 42743 2009 42753 2043
rect 42787 2009 42795 2043
rect 42743 1975 42795 2009
rect 42743 1941 42753 1975
rect 42787 1941 42795 1975
rect 42743 1923 42795 1941
rect 43663 2111 43715 2123
rect 43663 2077 43671 2111
rect 43705 2077 43715 2111
rect 43663 2043 43715 2077
rect 43663 2009 43671 2043
rect 43705 2009 43715 2043
rect 43663 1975 43715 2009
rect 43663 1941 43671 1975
rect 43705 1941 43715 1975
rect 43663 1923 43715 1941
rect 43745 1923 43787 2123
rect 43817 2111 43869 2123
rect 43817 2077 43827 2111
rect 43861 2077 43869 2111
rect 44477 2111 44529 2123
rect 43817 2043 43869 2077
rect 44477 2077 44485 2111
rect 44519 2077 44529 2111
rect 43817 2009 43827 2043
rect 43861 2009 43869 2043
rect 43817 1975 43869 2009
rect 44477 2043 44529 2077
rect 44477 2009 44485 2043
rect 44519 2009 44529 2043
rect 43817 1941 43827 1975
rect 43861 1941 43869 1975
rect 44477 1975 44529 2009
rect 43817 1923 43869 1941
rect 44012 1943 44074 1958
rect 42312 1875 42374 1909
rect 42312 1841 42328 1875
rect 42362 1841 42374 1875
rect 42312 1807 42374 1841
rect 42312 1773 42328 1807
rect 42362 1773 42374 1807
rect 44012 1909 44024 1943
rect 44058 1909 44074 1943
rect 44012 1875 44074 1909
rect 44012 1841 44024 1875
rect 44058 1841 44074 1875
rect 44012 1807 44074 1841
rect 42312 1758 42374 1773
rect 44012 1773 44024 1807
rect 44058 1773 44074 1807
rect 44012 1758 44074 1773
rect 44104 1943 44170 1958
rect 44104 1909 44120 1943
rect 44154 1909 44170 1943
rect 44104 1875 44170 1909
rect 44104 1841 44120 1875
rect 44154 1841 44170 1875
rect 44104 1807 44170 1841
rect 44104 1773 44120 1807
rect 44154 1773 44170 1807
rect 44104 1758 44170 1773
rect 44200 1943 44262 1958
rect 44200 1909 44216 1943
rect 44250 1909 44262 1943
rect 44477 1941 44485 1975
rect 44519 1941 44529 1975
rect 44477 1923 44529 1941
rect 44559 1923 44601 2123
rect 44631 2111 44683 2123
rect 44631 2077 44641 2111
rect 44675 2077 44683 2111
rect 44631 2043 44683 2077
rect 44631 2009 44641 2043
rect 44675 2009 44683 2043
rect 44631 1975 44683 2009
rect 44631 1941 44641 1975
rect 44675 1941 44683 1975
rect 44631 1923 44683 1941
rect 45545 2111 45597 2123
rect 45545 2077 45553 2111
rect 45587 2077 45597 2111
rect 45545 2043 45597 2077
rect 45545 2009 45553 2043
rect 45587 2009 45597 2043
rect 45545 1975 45597 2009
rect 45545 1941 45553 1975
rect 45587 1941 45597 1975
rect 45545 1923 45597 1941
rect 45627 1923 45669 2123
rect 45699 2111 45751 2123
rect 45699 2077 45709 2111
rect 45743 2077 45751 2111
rect 46359 2111 46411 2123
rect 45699 2043 45751 2077
rect 46359 2077 46367 2111
rect 46401 2077 46411 2111
rect 45699 2009 45709 2043
rect 45743 2009 45751 2043
rect 45699 1975 45751 2009
rect 46359 2043 46411 2077
rect 46359 2009 46367 2043
rect 46401 2009 46411 2043
rect 45699 1941 45709 1975
rect 45743 1941 45751 1975
rect 46359 1975 46411 2009
rect 45699 1923 45751 1941
rect 45894 1943 45956 1958
rect 44200 1875 44262 1909
rect 44200 1841 44216 1875
rect 44250 1841 44262 1875
rect 44200 1807 44262 1841
rect 44200 1773 44216 1807
rect 44250 1773 44262 1807
rect 45894 1909 45906 1943
rect 45940 1909 45956 1943
rect 45894 1875 45956 1909
rect 45894 1841 45906 1875
rect 45940 1841 45956 1875
rect 45894 1807 45956 1841
rect 44200 1758 44262 1773
rect 45894 1773 45906 1807
rect 45940 1773 45956 1807
rect 45894 1758 45956 1773
rect 45986 1943 46052 1958
rect 45986 1909 46002 1943
rect 46036 1909 46052 1943
rect 45986 1875 46052 1909
rect 45986 1841 46002 1875
rect 46036 1841 46052 1875
rect 45986 1807 46052 1841
rect 45986 1773 46002 1807
rect 46036 1773 46052 1807
rect 45986 1758 46052 1773
rect 46082 1943 46144 1958
rect 46082 1909 46098 1943
rect 46132 1909 46144 1943
rect 46359 1941 46367 1975
rect 46401 1941 46411 1975
rect 46359 1923 46411 1941
rect 46441 1923 46483 2123
rect 46513 2111 46565 2123
rect 46513 2077 46523 2111
rect 46557 2077 46565 2111
rect 46513 2043 46565 2077
rect 46513 2009 46523 2043
rect 46557 2009 46565 2043
rect 46513 1975 46565 2009
rect 46513 1941 46523 1975
rect 46557 1941 46565 1975
rect 46513 1923 46565 1941
rect 47433 2111 47485 2123
rect 47433 2077 47441 2111
rect 47475 2077 47485 2111
rect 47433 2043 47485 2077
rect 47433 2009 47441 2043
rect 47475 2009 47485 2043
rect 47433 1975 47485 2009
rect 47433 1941 47441 1975
rect 47475 1941 47485 1975
rect 47433 1923 47485 1941
rect 47515 1923 47557 2123
rect 47587 2111 47639 2123
rect 47587 2077 47597 2111
rect 47631 2077 47639 2111
rect 48247 2111 48299 2123
rect 47587 2043 47639 2077
rect 48247 2077 48255 2111
rect 48289 2077 48299 2111
rect 47587 2009 47597 2043
rect 47631 2009 47639 2043
rect 47587 1975 47639 2009
rect 48247 2043 48299 2077
rect 48247 2009 48255 2043
rect 48289 2009 48299 2043
rect 47587 1941 47597 1975
rect 47631 1941 47639 1975
rect 48247 1975 48299 2009
rect 47587 1923 47639 1941
rect 47782 1943 47844 1958
rect 46082 1875 46144 1909
rect 46082 1841 46098 1875
rect 46132 1841 46144 1875
rect 46082 1807 46144 1841
rect 46082 1773 46098 1807
rect 46132 1773 46144 1807
rect 47782 1909 47794 1943
rect 47828 1909 47844 1943
rect 47782 1875 47844 1909
rect 47782 1841 47794 1875
rect 47828 1841 47844 1875
rect 47782 1807 47844 1841
rect 46082 1758 46144 1773
rect 47782 1773 47794 1807
rect 47828 1773 47844 1807
rect 47782 1758 47844 1773
rect 47874 1943 47940 1958
rect 47874 1909 47890 1943
rect 47924 1909 47940 1943
rect 47874 1875 47940 1909
rect 47874 1841 47890 1875
rect 47924 1841 47940 1875
rect 47874 1807 47940 1841
rect 47874 1773 47890 1807
rect 47924 1773 47940 1807
rect 47874 1758 47940 1773
rect 47970 1943 48032 1958
rect 47970 1909 47986 1943
rect 48020 1909 48032 1943
rect 48247 1941 48255 1975
rect 48289 1941 48299 1975
rect 48247 1923 48299 1941
rect 48329 1923 48371 2123
rect 48401 2111 48453 2123
rect 48401 2077 48411 2111
rect 48445 2077 48453 2111
rect 48401 2043 48453 2077
rect 48401 2009 48411 2043
rect 48445 2009 48453 2043
rect 48401 1975 48453 2009
rect 48401 1941 48411 1975
rect 48445 1941 48453 1975
rect 48401 1923 48453 1941
rect 49321 2111 49373 2123
rect 49321 2077 49329 2111
rect 49363 2077 49373 2111
rect 49321 2043 49373 2077
rect 49321 2009 49329 2043
rect 49363 2009 49373 2043
rect 49321 1975 49373 2009
rect 49321 1941 49329 1975
rect 49363 1941 49373 1975
rect 49321 1923 49373 1941
rect 49403 1923 49445 2123
rect 49475 2111 49527 2123
rect 49475 2077 49485 2111
rect 49519 2077 49527 2111
rect 50135 2111 50187 2123
rect 49475 2043 49527 2077
rect 50135 2077 50143 2111
rect 50177 2077 50187 2111
rect 49475 2009 49485 2043
rect 49519 2009 49527 2043
rect 49475 1975 49527 2009
rect 50135 2043 50187 2077
rect 50135 2009 50143 2043
rect 50177 2009 50187 2043
rect 49475 1941 49485 1975
rect 49519 1941 49527 1975
rect 50135 1975 50187 2009
rect 49475 1923 49527 1941
rect 49670 1943 49732 1958
rect 47970 1875 48032 1909
rect 47970 1841 47986 1875
rect 48020 1841 48032 1875
rect 47970 1807 48032 1841
rect 47970 1773 47986 1807
rect 48020 1773 48032 1807
rect 49670 1909 49682 1943
rect 49716 1909 49732 1943
rect 49670 1875 49732 1909
rect 49670 1841 49682 1875
rect 49716 1841 49732 1875
rect 49670 1807 49732 1841
rect 47970 1758 48032 1773
rect 49670 1773 49682 1807
rect 49716 1773 49732 1807
rect 49670 1758 49732 1773
rect 49762 1943 49828 1958
rect 49762 1909 49778 1943
rect 49812 1909 49828 1943
rect 49762 1875 49828 1909
rect 49762 1841 49778 1875
rect 49812 1841 49828 1875
rect 49762 1807 49828 1841
rect 49762 1773 49778 1807
rect 49812 1773 49828 1807
rect 49762 1758 49828 1773
rect 49858 1943 49920 1958
rect 49858 1909 49874 1943
rect 49908 1909 49920 1943
rect 50135 1941 50143 1975
rect 50177 1941 50187 1975
rect 50135 1923 50187 1941
rect 50217 1923 50259 2123
rect 50289 2111 50341 2123
rect 50289 2077 50299 2111
rect 50333 2077 50341 2111
rect 50289 2043 50341 2077
rect 50289 2009 50299 2043
rect 50333 2009 50341 2043
rect 50289 1975 50341 2009
rect 50289 1941 50299 1975
rect 50333 1941 50341 1975
rect 50289 1923 50341 1941
rect 51209 2111 51261 2123
rect 51209 2077 51217 2111
rect 51251 2077 51261 2111
rect 51209 2043 51261 2077
rect 51209 2009 51217 2043
rect 51251 2009 51261 2043
rect 51209 1975 51261 2009
rect 51209 1941 51217 1975
rect 51251 1941 51261 1975
rect 51209 1923 51261 1941
rect 51291 1923 51333 2123
rect 51363 2111 51415 2123
rect 51363 2077 51373 2111
rect 51407 2077 51415 2111
rect 52023 2111 52075 2123
rect 51363 2043 51415 2077
rect 52023 2077 52031 2111
rect 52065 2077 52075 2111
rect 51363 2009 51373 2043
rect 51407 2009 51415 2043
rect 51363 1975 51415 2009
rect 52023 2043 52075 2077
rect 52023 2009 52031 2043
rect 52065 2009 52075 2043
rect 51363 1941 51373 1975
rect 51407 1941 51415 1975
rect 52023 1975 52075 2009
rect 51363 1923 51415 1941
rect 51558 1943 51620 1958
rect 49858 1875 49920 1909
rect 49858 1841 49874 1875
rect 49908 1841 49920 1875
rect 49858 1807 49920 1841
rect 49858 1773 49874 1807
rect 49908 1773 49920 1807
rect 51558 1909 51570 1943
rect 51604 1909 51620 1943
rect 51558 1875 51620 1909
rect 51558 1841 51570 1875
rect 51604 1841 51620 1875
rect 51558 1807 51620 1841
rect 49858 1758 49920 1773
rect 51558 1773 51570 1807
rect 51604 1773 51620 1807
rect 51558 1758 51620 1773
rect 51650 1943 51716 1958
rect 51650 1909 51666 1943
rect 51700 1909 51716 1943
rect 51650 1875 51716 1909
rect 51650 1841 51666 1875
rect 51700 1841 51716 1875
rect 51650 1807 51716 1841
rect 51650 1773 51666 1807
rect 51700 1773 51716 1807
rect 51650 1758 51716 1773
rect 51746 1943 51808 1958
rect 51746 1909 51762 1943
rect 51796 1909 51808 1943
rect 52023 1941 52031 1975
rect 52065 1941 52075 1975
rect 52023 1923 52075 1941
rect 52105 1923 52147 2123
rect 52177 2111 52229 2123
rect 52177 2077 52187 2111
rect 52221 2077 52229 2111
rect 52177 2043 52229 2077
rect 52177 2009 52187 2043
rect 52221 2009 52229 2043
rect 52177 1975 52229 2009
rect 52177 1941 52187 1975
rect 52221 1941 52229 1975
rect 52177 1923 52229 1941
rect 53097 2111 53149 2123
rect 53097 2077 53105 2111
rect 53139 2077 53149 2111
rect 53097 2043 53149 2077
rect 53097 2009 53105 2043
rect 53139 2009 53149 2043
rect 53097 1975 53149 2009
rect 53097 1941 53105 1975
rect 53139 1941 53149 1975
rect 53097 1923 53149 1941
rect 53179 1923 53221 2123
rect 53251 2111 53303 2123
rect 53251 2077 53261 2111
rect 53295 2077 53303 2111
rect 53911 2111 53963 2123
rect 53251 2043 53303 2077
rect 53911 2077 53919 2111
rect 53953 2077 53963 2111
rect 53251 2009 53261 2043
rect 53295 2009 53303 2043
rect 53251 1975 53303 2009
rect 53911 2043 53963 2077
rect 53911 2009 53919 2043
rect 53953 2009 53963 2043
rect 53251 1941 53261 1975
rect 53295 1941 53303 1975
rect 53911 1975 53963 2009
rect 53251 1923 53303 1941
rect 53446 1943 53508 1958
rect 51746 1875 51808 1909
rect 51746 1841 51762 1875
rect 51796 1841 51808 1875
rect 51746 1807 51808 1841
rect 51746 1773 51762 1807
rect 51796 1773 51808 1807
rect 53446 1909 53458 1943
rect 53492 1909 53508 1943
rect 53446 1875 53508 1909
rect 53446 1841 53458 1875
rect 53492 1841 53508 1875
rect 53446 1807 53508 1841
rect 51746 1758 51808 1773
rect 53446 1773 53458 1807
rect 53492 1773 53508 1807
rect 53446 1758 53508 1773
rect 53538 1943 53604 1958
rect 53538 1909 53554 1943
rect 53588 1909 53604 1943
rect 53538 1875 53604 1909
rect 53538 1841 53554 1875
rect 53588 1841 53604 1875
rect 53538 1807 53604 1841
rect 53538 1773 53554 1807
rect 53588 1773 53604 1807
rect 53538 1758 53604 1773
rect 53634 1943 53696 1958
rect 53634 1909 53650 1943
rect 53684 1909 53696 1943
rect 53911 1941 53919 1975
rect 53953 1941 53963 1975
rect 53911 1923 53963 1941
rect 53993 1923 54035 2123
rect 54065 2111 54117 2123
rect 54065 2077 54075 2111
rect 54109 2077 54117 2111
rect 54065 2043 54117 2077
rect 54065 2009 54075 2043
rect 54109 2009 54117 2043
rect 54065 1975 54117 2009
rect 54065 1941 54075 1975
rect 54109 1941 54117 1975
rect 54065 1923 54117 1941
rect 54985 2111 55037 2123
rect 54985 2077 54993 2111
rect 55027 2077 55037 2111
rect 54985 2043 55037 2077
rect 54985 2009 54993 2043
rect 55027 2009 55037 2043
rect 54985 1975 55037 2009
rect 54985 1941 54993 1975
rect 55027 1941 55037 1975
rect 54985 1923 55037 1941
rect 55067 1923 55109 2123
rect 55139 2111 55191 2123
rect 55139 2077 55149 2111
rect 55183 2077 55191 2111
rect 55799 2111 55851 2123
rect 55139 2043 55191 2077
rect 55799 2077 55807 2111
rect 55841 2077 55851 2111
rect 55139 2009 55149 2043
rect 55183 2009 55191 2043
rect 55139 1975 55191 2009
rect 55799 2043 55851 2077
rect 55799 2009 55807 2043
rect 55841 2009 55851 2043
rect 55139 1941 55149 1975
rect 55183 1941 55191 1975
rect 55799 1975 55851 2009
rect 55139 1923 55191 1941
rect 55334 1943 55396 1958
rect 53634 1875 53696 1909
rect 53634 1841 53650 1875
rect 53684 1841 53696 1875
rect 53634 1807 53696 1841
rect 53634 1773 53650 1807
rect 53684 1773 53696 1807
rect 55334 1909 55346 1943
rect 55380 1909 55396 1943
rect 55334 1875 55396 1909
rect 55334 1841 55346 1875
rect 55380 1841 55396 1875
rect 55334 1807 55396 1841
rect 53634 1758 53696 1773
rect 55334 1773 55346 1807
rect 55380 1773 55396 1807
rect 55334 1758 55396 1773
rect 55426 1943 55492 1958
rect 55426 1909 55442 1943
rect 55476 1909 55492 1943
rect 55426 1875 55492 1909
rect 55426 1841 55442 1875
rect 55476 1841 55492 1875
rect 55426 1807 55492 1841
rect 55426 1773 55442 1807
rect 55476 1773 55492 1807
rect 55426 1758 55492 1773
rect 55522 1943 55584 1958
rect 55522 1909 55538 1943
rect 55572 1909 55584 1943
rect 55799 1941 55807 1975
rect 55841 1941 55851 1975
rect 55799 1923 55851 1941
rect 55881 1923 55923 2123
rect 55953 2111 56005 2123
rect 55953 2077 55963 2111
rect 55997 2077 56005 2111
rect 55953 2043 56005 2077
rect 55953 2009 55963 2043
rect 55997 2009 56005 2043
rect 55953 1975 56005 2009
rect 55953 1941 55963 1975
rect 55997 1941 56005 1975
rect 55953 1923 56005 1941
rect 56873 2111 56925 2123
rect 56873 2077 56881 2111
rect 56915 2077 56925 2111
rect 56873 2043 56925 2077
rect 56873 2009 56881 2043
rect 56915 2009 56925 2043
rect 56873 1975 56925 2009
rect 56873 1941 56881 1975
rect 56915 1941 56925 1975
rect 56873 1923 56925 1941
rect 56955 1923 56997 2123
rect 57027 2111 57079 2123
rect 57027 2077 57037 2111
rect 57071 2077 57079 2111
rect 57687 2111 57739 2123
rect 57027 2043 57079 2077
rect 57687 2077 57695 2111
rect 57729 2077 57739 2111
rect 57027 2009 57037 2043
rect 57071 2009 57079 2043
rect 57027 1975 57079 2009
rect 57687 2043 57739 2077
rect 57687 2009 57695 2043
rect 57729 2009 57739 2043
rect 57027 1941 57037 1975
rect 57071 1941 57079 1975
rect 57687 1975 57739 2009
rect 57027 1923 57079 1941
rect 57222 1943 57284 1958
rect 55522 1875 55584 1909
rect 55522 1841 55538 1875
rect 55572 1841 55584 1875
rect 55522 1807 55584 1841
rect 55522 1773 55538 1807
rect 55572 1773 55584 1807
rect 57222 1909 57234 1943
rect 57268 1909 57284 1943
rect 57222 1875 57284 1909
rect 57222 1841 57234 1875
rect 57268 1841 57284 1875
rect 57222 1807 57284 1841
rect 55522 1758 55584 1773
rect 57222 1773 57234 1807
rect 57268 1773 57284 1807
rect 57222 1758 57284 1773
rect 57314 1943 57380 1958
rect 57314 1909 57330 1943
rect 57364 1909 57380 1943
rect 57314 1875 57380 1909
rect 57314 1841 57330 1875
rect 57364 1841 57380 1875
rect 57314 1807 57380 1841
rect 57314 1773 57330 1807
rect 57364 1773 57380 1807
rect 57314 1758 57380 1773
rect 57410 1943 57472 1958
rect 57410 1909 57426 1943
rect 57460 1909 57472 1943
rect 57687 1941 57695 1975
rect 57729 1941 57739 1975
rect 57687 1923 57739 1941
rect 57769 1923 57811 2123
rect 57841 2111 57893 2123
rect 57841 2077 57851 2111
rect 57885 2077 57893 2111
rect 57841 2043 57893 2077
rect 57841 2009 57851 2043
rect 57885 2009 57893 2043
rect 57841 1975 57893 2009
rect 57841 1941 57851 1975
rect 57885 1941 57893 1975
rect 57841 1923 57893 1941
rect 58761 2111 58813 2123
rect 58761 2077 58769 2111
rect 58803 2077 58813 2111
rect 58761 2043 58813 2077
rect 58761 2009 58769 2043
rect 58803 2009 58813 2043
rect 58761 1975 58813 2009
rect 58761 1941 58769 1975
rect 58803 1941 58813 1975
rect 58761 1923 58813 1941
rect 58843 1923 58885 2123
rect 58915 2111 58967 2123
rect 58915 2077 58925 2111
rect 58959 2077 58967 2111
rect 59575 2111 59627 2123
rect 58915 2043 58967 2077
rect 59575 2077 59583 2111
rect 59617 2077 59627 2111
rect 58915 2009 58925 2043
rect 58959 2009 58967 2043
rect 58915 1975 58967 2009
rect 59575 2043 59627 2077
rect 59575 2009 59583 2043
rect 59617 2009 59627 2043
rect 58915 1941 58925 1975
rect 58959 1941 58967 1975
rect 59575 1975 59627 2009
rect 58915 1923 58967 1941
rect 59110 1943 59172 1958
rect 57410 1875 57472 1909
rect 57410 1841 57426 1875
rect 57460 1841 57472 1875
rect 57410 1807 57472 1841
rect 57410 1773 57426 1807
rect 57460 1773 57472 1807
rect 59110 1909 59122 1943
rect 59156 1909 59172 1943
rect 59110 1875 59172 1909
rect 59110 1841 59122 1875
rect 59156 1841 59172 1875
rect 59110 1807 59172 1841
rect 57410 1758 57472 1773
rect 59110 1773 59122 1807
rect 59156 1773 59172 1807
rect 59110 1758 59172 1773
rect 59202 1943 59268 1958
rect 59202 1909 59218 1943
rect 59252 1909 59268 1943
rect 59202 1875 59268 1909
rect 59202 1841 59218 1875
rect 59252 1841 59268 1875
rect 59202 1807 59268 1841
rect 59202 1773 59218 1807
rect 59252 1773 59268 1807
rect 59202 1758 59268 1773
rect 59298 1943 59360 1958
rect 59298 1909 59314 1943
rect 59348 1909 59360 1943
rect 59575 1941 59583 1975
rect 59617 1941 59627 1975
rect 59575 1923 59627 1941
rect 59657 1923 59699 2123
rect 59729 2111 59781 2123
rect 59729 2077 59739 2111
rect 59773 2077 59781 2111
rect 59729 2043 59781 2077
rect 59729 2009 59739 2043
rect 59773 2009 59781 2043
rect 59729 1975 59781 2009
rect 59729 1941 59739 1975
rect 59773 1941 59781 1975
rect 59729 1923 59781 1941
rect 59298 1875 59360 1909
rect 59298 1841 59314 1875
rect 59348 1841 59360 1875
rect 59298 1807 59360 1841
rect 59298 1773 59314 1807
rect 59348 1773 59360 1807
rect 59298 1758 59360 1773
rect 108 1057 160 1069
rect 108 1023 116 1057
rect 150 1023 160 1057
rect 108 989 160 1023
rect 108 955 116 989
rect 150 955 160 989
rect 108 921 160 955
rect 108 887 116 921
rect 150 887 160 921
rect 108 869 160 887
rect 190 1057 242 1069
rect 190 1023 200 1057
rect 234 1023 242 1057
rect 190 989 242 1023
rect 190 955 200 989
rect 234 955 242 989
rect 190 921 242 955
rect 190 887 200 921
rect 234 887 242 921
rect 190 869 242 887
rect 376 1047 434 1062
rect 376 1013 388 1047
rect 422 1013 434 1047
rect 376 979 434 1013
rect 376 945 388 979
rect 422 945 434 979
rect 376 911 434 945
rect 376 877 388 911
rect 422 877 434 911
rect 376 862 434 877
rect 464 1047 522 1062
rect 464 1013 476 1047
rect 510 1013 522 1047
rect 464 979 522 1013
rect 1304 1065 1356 1077
rect 1022 1047 1080 1062
rect 1022 1013 1034 1047
rect 1068 1013 1080 1047
rect 464 945 476 979
rect 510 945 522 979
rect 464 911 522 945
rect 464 877 476 911
rect 510 877 522 911
rect 1022 979 1080 1013
rect 1022 945 1034 979
rect 1068 945 1080 979
rect 1022 911 1080 945
rect 464 862 522 877
rect 592 887 654 902
rect 592 853 604 887
rect 638 853 654 887
rect 592 819 654 853
rect 592 785 604 819
rect 638 785 654 819
rect 592 751 654 785
rect 592 717 604 751
rect 638 717 654 751
rect 592 702 654 717
rect 684 887 750 902
rect 684 853 700 887
rect 734 853 750 887
rect 684 819 750 853
rect 684 785 700 819
rect 734 785 750 819
rect 684 751 750 785
rect 684 717 700 751
rect 734 717 750 751
rect 684 702 750 717
rect 780 887 842 902
rect 780 853 796 887
rect 830 853 842 887
rect 1022 877 1034 911
rect 1068 877 1080 911
rect 1022 862 1080 877
rect 1110 1047 1168 1062
rect 1110 1013 1122 1047
rect 1156 1013 1168 1047
rect 1110 979 1168 1013
rect 1110 945 1122 979
rect 1156 945 1168 979
rect 1110 911 1168 945
rect 1110 877 1122 911
rect 1156 877 1168 911
rect 1304 1031 1312 1065
rect 1346 1031 1356 1065
rect 1304 997 1356 1031
rect 1304 963 1312 997
rect 1346 963 1356 997
rect 1304 929 1356 963
rect 1304 895 1312 929
rect 1346 895 1356 929
rect 1304 877 1356 895
rect 1386 1065 1438 1077
rect 1386 1031 1396 1065
rect 1430 1031 1438 1065
rect 1386 997 1438 1031
rect 1386 963 1396 997
rect 1430 963 1438 997
rect 1386 929 1438 963
rect 1386 895 1396 929
rect 1430 895 1438 929
rect 1609 1055 1661 1075
rect 1609 1021 1617 1055
rect 1651 1021 1661 1055
rect 1609 987 1661 1021
rect 1609 953 1617 987
rect 1651 953 1661 987
rect 1609 917 1661 953
rect 1691 1055 1749 1075
rect 1691 1021 1703 1055
rect 1737 1021 1749 1055
rect 1691 987 1749 1021
rect 1691 953 1703 987
rect 1737 953 1749 987
rect 1691 917 1749 953
rect 1779 1055 1831 1075
rect 1779 1021 1789 1055
rect 1823 1021 1831 1055
rect 1779 974 1831 1021
rect 1779 940 1789 974
rect 1823 940 1831 974
rect 1779 917 1831 940
rect 1996 1057 2048 1069
rect 1996 1023 2004 1057
rect 2038 1023 2048 1057
rect 1996 989 2048 1023
rect 1996 955 2004 989
rect 2038 955 2048 989
rect 1996 921 2048 955
rect 1386 877 1438 895
rect 1110 862 1168 877
rect 780 819 842 853
rect 780 785 796 819
rect 830 785 842 819
rect 780 751 842 785
rect 1996 887 2004 921
rect 2038 887 2048 921
rect 1996 869 2048 887
rect 2078 1057 2130 1069
rect 2078 1023 2088 1057
rect 2122 1023 2130 1057
rect 2078 989 2130 1023
rect 2078 955 2088 989
rect 2122 955 2130 989
rect 2078 921 2130 955
rect 2078 887 2088 921
rect 2122 887 2130 921
rect 2078 869 2130 887
rect 2264 1047 2322 1062
rect 2264 1013 2276 1047
rect 2310 1013 2322 1047
rect 2264 979 2322 1013
rect 2264 945 2276 979
rect 2310 945 2322 979
rect 2264 911 2322 945
rect 2264 877 2276 911
rect 2310 877 2322 911
rect 2264 862 2322 877
rect 2352 1047 2410 1062
rect 2352 1013 2364 1047
rect 2398 1013 2410 1047
rect 2352 979 2410 1013
rect 3192 1065 3244 1077
rect 2910 1047 2968 1062
rect 2910 1013 2922 1047
rect 2956 1013 2968 1047
rect 2352 945 2364 979
rect 2398 945 2410 979
rect 2352 911 2410 945
rect 2352 877 2364 911
rect 2398 877 2410 911
rect 2910 979 2968 1013
rect 2910 945 2922 979
rect 2956 945 2968 979
rect 2910 911 2968 945
rect 2352 862 2410 877
rect 2480 887 2542 902
rect 2480 853 2492 887
rect 2526 853 2542 887
rect 780 717 796 751
rect 830 717 842 751
rect 780 702 842 717
rect 2480 819 2542 853
rect 2480 785 2492 819
rect 2526 785 2542 819
rect 2480 751 2542 785
rect 2480 717 2492 751
rect 2526 717 2542 751
rect 2480 702 2542 717
rect 2572 887 2638 902
rect 2572 853 2588 887
rect 2622 853 2638 887
rect 2572 819 2638 853
rect 2572 785 2588 819
rect 2622 785 2638 819
rect 2572 751 2638 785
rect 2572 717 2588 751
rect 2622 717 2638 751
rect 2572 702 2638 717
rect 2668 887 2730 902
rect 2668 853 2684 887
rect 2718 853 2730 887
rect 2910 877 2922 911
rect 2956 877 2968 911
rect 2910 862 2968 877
rect 2998 1047 3056 1062
rect 2998 1013 3010 1047
rect 3044 1013 3056 1047
rect 2998 979 3056 1013
rect 2998 945 3010 979
rect 3044 945 3056 979
rect 2998 911 3056 945
rect 2998 877 3010 911
rect 3044 877 3056 911
rect 3192 1031 3200 1065
rect 3234 1031 3244 1065
rect 3192 997 3244 1031
rect 3192 963 3200 997
rect 3234 963 3244 997
rect 3192 929 3244 963
rect 3192 895 3200 929
rect 3234 895 3244 929
rect 3192 877 3244 895
rect 3274 1065 3326 1077
rect 3274 1031 3284 1065
rect 3318 1031 3326 1065
rect 3274 997 3326 1031
rect 3274 963 3284 997
rect 3318 963 3326 997
rect 3274 929 3326 963
rect 3274 895 3284 929
rect 3318 895 3326 929
rect 3497 1055 3549 1075
rect 3497 1021 3505 1055
rect 3539 1021 3549 1055
rect 3497 987 3549 1021
rect 3497 953 3505 987
rect 3539 953 3549 987
rect 3497 917 3549 953
rect 3579 1055 3637 1075
rect 3579 1021 3591 1055
rect 3625 1021 3637 1055
rect 3579 987 3637 1021
rect 3579 953 3591 987
rect 3625 953 3637 987
rect 3579 917 3637 953
rect 3667 1055 3719 1075
rect 3667 1021 3677 1055
rect 3711 1021 3719 1055
rect 3667 974 3719 1021
rect 3667 940 3677 974
rect 3711 940 3719 974
rect 3667 917 3719 940
rect 3884 1057 3936 1069
rect 3884 1023 3892 1057
rect 3926 1023 3936 1057
rect 3884 989 3936 1023
rect 3884 955 3892 989
rect 3926 955 3936 989
rect 3884 921 3936 955
rect 3274 877 3326 895
rect 2998 862 3056 877
rect 2668 819 2730 853
rect 2668 785 2684 819
rect 2718 785 2730 819
rect 2668 751 2730 785
rect 3884 887 3892 921
rect 3926 887 3936 921
rect 3884 869 3936 887
rect 3966 1057 4018 1069
rect 3966 1023 3976 1057
rect 4010 1023 4018 1057
rect 3966 989 4018 1023
rect 3966 955 3976 989
rect 4010 955 4018 989
rect 3966 921 4018 955
rect 3966 887 3976 921
rect 4010 887 4018 921
rect 3966 869 4018 887
rect 4152 1047 4210 1062
rect 4152 1013 4164 1047
rect 4198 1013 4210 1047
rect 4152 979 4210 1013
rect 4152 945 4164 979
rect 4198 945 4210 979
rect 4152 911 4210 945
rect 4152 877 4164 911
rect 4198 877 4210 911
rect 4152 862 4210 877
rect 4240 1047 4298 1062
rect 4240 1013 4252 1047
rect 4286 1013 4298 1047
rect 4240 979 4298 1013
rect 5080 1065 5132 1077
rect 4798 1047 4856 1062
rect 4798 1013 4810 1047
rect 4844 1013 4856 1047
rect 4240 945 4252 979
rect 4286 945 4298 979
rect 4240 911 4298 945
rect 4240 877 4252 911
rect 4286 877 4298 911
rect 4798 979 4856 1013
rect 4798 945 4810 979
rect 4844 945 4856 979
rect 4798 911 4856 945
rect 4240 862 4298 877
rect 4368 887 4430 902
rect 4368 853 4380 887
rect 4414 853 4430 887
rect 2668 717 2684 751
rect 2718 717 2730 751
rect 2668 702 2730 717
rect 4368 819 4430 853
rect 4368 785 4380 819
rect 4414 785 4430 819
rect 4368 751 4430 785
rect 4368 717 4380 751
rect 4414 717 4430 751
rect 4368 702 4430 717
rect 4460 887 4526 902
rect 4460 853 4476 887
rect 4510 853 4526 887
rect 4460 819 4526 853
rect 4460 785 4476 819
rect 4510 785 4526 819
rect 4460 751 4526 785
rect 4460 717 4476 751
rect 4510 717 4526 751
rect 4460 702 4526 717
rect 4556 887 4618 902
rect 4556 853 4572 887
rect 4606 853 4618 887
rect 4798 877 4810 911
rect 4844 877 4856 911
rect 4798 862 4856 877
rect 4886 1047 4944 1062
rect 4886 1013 4898 1047
rect 4932 1013 4944 1047
rect 4886 979 4944 1013
rect 4886 945 4898 979
rect 4932 945 4944 979
rect 4886 911 4944 945
rect 4886 877 4898 911
rect 4932 877 4944 911
rect 5080 1031 5088 1065
rect 5122 1031 5132 1065
rect 5080 997 5132 1031
rect 5080 963 5088 997
rect 5122 963 5132 997
rect 5080 929 5132 963
rect 5080 895 5088 929
rect 5122 895 5132 929
rect 5080 877 5132 895
rect 5162 1065 5214 1077
rect 5162 1031 5172 1065
rect 5206 1031 5214 1065
rect 5162 997 5214 1031
rect 5162 963 5172 997
rect 5206 963 5214 997
rect 5162 929 5214 963
rect 5162 895 5172 929
rect 5206 895 5214 929
rect 5385 1055 5437 1075
rect 5385 1021 5393 1055
rect 5427 1021 5437 1055
rect 5385 987 5437 1021
rect 5385 953 5393 987
rect 5427 953 5437 987
rect 5385 917 5437 953
rect 5467 1055 5525 1075
rect 5467 1021 5479 1055
rect 5513 1021 5525 1055
rect 5467 987 5525 1021
rect 5467 953 5479 987
rect 5513 953 5525 987
rect 5467 917 5525 953
rect 5555 1055 5607 1075
rect 5555 1021 5565 1055
rect 5599 1021 5607 1055
rect 5555 974 5607 1021
rect 5555 940 5565 974
rect 5599 940 5607 974
rect 5555 917 5607 940
rect 5772 1057 5824 1069
rect 5772 1023 5780 1057
rect 5814 1023 5824 1057
rect 5772 989 5824 1023
rect 5772 955 5780 989
rect 5814 955 5824 989
rect 5772 921 5824 955
rect 5162 877 5214 895
rect 4886 862 4944 877
rect 4556 819 4618 853
rect 4556 785 4572 819
rect 4606 785 4618 819
rect 4556 751 4618 785
rect 5772 887 5780 921
rect 5814 887 5824 921
rect 5772 869 5824 887
rect 5854 1057 5906 1069
rect 5854 1023 5864 1057
rect 5898 1023 5906 1057
rect 5854 989 5906 1023
rect 5854 955 5864 989
rect 5898 955 5906 989
rect 5854 921 5906 955
rect 5854 887 5864 921
rect 5898 887 5906 921
rect 5854 869 5906 887
rect 6040 1047 6098 1062
rect 6040 1013 6052 1047
rect 6086 1013 6098 1047
rect 6040 979 6098 1013
rect 6040 945 6052 979
rect 6086 945 6098 979
rect 6040 911 6098 945
rect 6040 877 6052 911
rect 6086 877 6098 911
rect 6040 862 6098 877
rect 6128 1047 6186 1062
rect 6128 1013 6140 1047
rect 6174 1013 6186 1047
rect 6128 979 6186 1013
rect 6968 1065 7020 1077
rect 6686 1047 6744 1062
rect 6686 1013 6698 1047
rect 6732 1013 6744 1047
rect 6128 945 6140 979
rect 6174 945 6186 979
rect 6128 911 6186 945
rect 6128 877 6140 911
rect 6174 877 6186 911
rect 6686 979 6744 1013
rect 6686 945 6698 979
rect 6732 945 6744 979
rect 6686 911 6744 945
rect 6128 862 6186 877
rect 6256 887 6318 902
rect 6256 853 6268 887
rect 6302 853 6318 887
rect 4556 717 4572 751
rect 4606 717 4618 751
rect 4556 702 4618 717
rect 6256 819 6318 853
rect 6256 785 6268 819
rect 6302 785 6318 819
rect 6256 751 6318 785
rect 6256 717 6268 751
rect 6302 717 6318 751
rect 6256 702 6318 717
rect 6348 887 6414 902
rect 6348 853 6364 887
rect 6398 853 6414 887
rect 6348 819 6414 853
rect 6348 785 6364 819
rect 6398 785 6414 819
rect 6348 751 6414 785
rect 6348 717 6364 751
rect 6398 717 6414 751
rect 6348 702 6414 717
rect 6444 887 6506 902
rect 6444 853 6460 887
rect 6494 853 6506 887
rect 6686 877 6698 911
rect 6732 877 6744 911
rect 6686 862 6744 877
rect 6774 1047 6832 1062
rect 6774 1013 6786 1047
rect 6820 1013 6832 1047
rect 6774 979 6832 1013
rect 6774 945 6786 979
rect 6820 945 6832 979
rect 6774 911 6832 945
rect 6774 877 6786 911
rect 6820 877 6832 911
rect 6968 1031 6976 1065
rect 7010 1031 7020 1065
rect 6968 997 7020 1031
rect 6968 963 6976 997
rect 7010 963 7020 997
rect 6968 929 7020 963
rect 6968 895 6976 929
rect 7010 895 7020 929
rect 6968 877 7020 895
rect 7050 1065 7102 1077
rect 7050 1031 7060 1065
rect 7094 1031 7102 1065
rect 7050 997 7102 1031
rect 7050 963 7060 997
rect 7094 963 7102 997
rect 7050 929 7102 963
rect 7050 895 7060 929
rect 7094 895 7102 929
rect 7273 1055 7325 1075
rect 7273 1021 7281 1055
rect 7315 1021 7325 1055
rect 7273 987 7325 1021
rect 7273 953 7281 987
rect 7315 953 7325 987
rect 7273 917 7325 953
rect 7355 1055 7413 1075
rect 7355 1021 7367 1055
rect 7401 1021 7413 1055
rect 7355 987 7413 1021
rect 7355 953 7367 987
rect 7401 953 7413 987
rect 7355 917 7413 953
rect 7443 1055 7495 1075
rect 7443 1021 7453 1055
rect 7487 1021 7495 1055
rect 7443 974 7495 1021
rect 7443 940 7453 974
rect 7487 940 7495 974
rect 7443 917 7495 940
rect 7660 1057 7712 1069
rect 7660 1023 7668 1057
rect 7702 1023 7712 1057
rect 7660 989 7712 1023
rect 7660 955 7668 989
rect 7702 955 7712 989
rect 7660 921 7712 955
rect 7050 877 7102 895
rect 6774 862 6832 877
rect 6444 819 6506 853
rect 6444 785 6460 819
rect 6494 785 6506 819
rect 6444 751 6506 785
rect 7660 887 7668 921
rect 7702 887 7712 921
rect 7660 869 7712 887
rect 7742 1057 7794 1069
rect 7742 1023 7752 1057
rect 7786 1023 7794 1057
rect 7742 989 7794 1023
rect 7742 955 7752 989
rect 7786 955 7794 989
rect 7742 921 7794 955
rect 7742 887 7752 921
rect 7786 887 7794 921
rect 7742 869 7794 887
rect 7928 1047 7986 1062
rect 7928 1013 7940 1047
rect 7974 1013 7986 1047
rect 7928 979 7986 1013
rect 7928 945 7940 979
rect 7974 945 7986 979
rect 7928 911 7986 945
rect 7928 877 7940 911
rect 7974 877 7986 911
rect 7928 862 7986 877
rect 8016 1047 8074 1062
rect 8016 1013 8028 1047
rect 8062 1013 8074 1047
rect 8016 979 8074 1013
rect 8856 1065 8908 1077
rect 8574 1047 8632 1062
rect 8574 1013 8586 1047
rect 8620 1013 8632 1047
rect 8016 945 8028 979
rect 8062 945 8074 979
rect 8016 911 8074 945
rect 8016 877 8028 911
rect 8062 877 8074 911
rect 8574 979 8632 1013
rect 8574 945 8586 979
rect 8620 945 8632 979
rect 8574 911 8632 945
rect 8016 862 8074 877
rect 8144 887 8206 902
rect 8144 853 8156 887
rect 8190 853 8206 887
rect 6444 717 6460 751
rect 6494 717 6506 751
rect 6444 702 6506 717
rect 8144 819 8206 853
rect 8144 785 8156 819
rect 8190 785 8206 819
rect 8144 751 8206 785
rect 8144 717 8156 751
rect 8190 717 8206 751
rect 8144 702 8206 717
rect 8236 887 8302 902
rect 8236 853 8252 887
rect 8286 853 8302 887
rect 8236 819 8302 853
rect 8236 785 8252 819
rect 8286 785 8302 819
rect 8236 751 8302 785
rect 8236 717 8252 751
rect 8286 717 8302 751
rect 8236 702 8302 717
rect 8332 887 8394 902
rect 8332 853 8348 887
rect 8382 853 8394 887
rect 8574 877 8586 911
rect 8620 877 8632 911
rect 8574 862 8632 877
rect 8662 1047 8720 1062
rect 8662 1013 8674 1047
rect 8708 1013 8720 1047
rect 8662 979 8720 1013
rect 8662 945 8674 979
rect 8708 945 8720 979
rect 8662 911 8720 945
rect 8662 877 8674 911
rect 8708 877 8720 911
rect 8856 1031 8864 1065
rect 8898 1031 8908 1065
rect 8856 997 8908 1031
rect 8856 963 8864 997
rect 8898 963 8908 997
rect 8856 929 8908 963
rect 8856 895 8864 929
rect 8898 895 8908 929
rect 8856 877 8908 895
rect 8938 1065 8990 1077
rect 8938 1031 8948 1065
rect 8982 1031 8990 1065
rect 8938 997 8990 1031
rect 8938 963 8948 997
rect 8982 963 8990 997
rect 8938 929 8990 963
rect 8938 895 8948 929
rect 8982 895 8990 929
rect 9161 1055 9213 1075
rect 9161 1021 9169 1055
rect 9203 1021 9213 1055
rect 9161 987 9213 1021
rect 9161 953 9169 987
rect 9203 953 9213 987
rect 9161 917 9213 953
rect 9243 1055 9301 1075
rect 9243 1021 9255 1055
rect 9289 1021 9301 1055
rect 9243 987 9301 1021
rect 9243 953 9255 987
rect 9289 953 9301 987
rect 9243 917 9301 953
rect 9331 1055 9383 1075
rect 9331 1021 9341 1055
rect 9375 1021 9383 1055
rect 9331 974 9383 1021
rect 9331 940 9341 974
rect 9375 940 9383 974
rect 9331 917 9383 940
rect 9548 1057 9600 1069
rect 9548 1023 9556 1057
rect 9590 1023 9600 1057
rect 9548 989 9600 1023
rect 9548 955 9556 989
rect 9590 955 9600 989
rect 9548 921 9600 955
rect 8938 877 8990 895
rect 8662 862 8720 877
rect 8332 819 8394 853
rect 8332 785 8348 819
rect 8382 785 8394 819
rect 8332 751 8394 785
rect 9548 887 9556 921
rect 9590 887 9600 921
rect 9548 869 9600 887
rect 9630 1057 9682 1069
rect 9630 1023 9640 1057
rect 9674 1023 9682 1057
rect 9630 989 9682 1023
rect 9630 955 9640 989
rect 9674 955 9682 989
rect 9630 921 9682 955
rect 9630 887 9640 921
rect 9674 887 9682 921
rect 9630 869 9682 887
rect 9816 1047 9874 1062
rect 9816 1013 9828 1047
rect 9862 1013 9874 1047
rect 9816 979 9874 1013
rect 9816 945 9828 979
rect 9862 945 9874 979
rect 9816 911 9874 945
rect 9816 877 9828 911
rect 9862 877 9874 911
rect 9816 862 9874 877
rect 9904 1047 9962 1062
rect 9904 1013 9916 1047
rect 9950 1013 9962 1047
rect 9904 979 9962 1013
rect 10744 1065 10796 1077
rect 10462 1047 10520 1062
rect 10462 1013 10474 1047
rect 10508 1013 10520 1047
rect 9904 945 9916 979
rect 9950 945 9962 979
rect 9904 911 9962 945
rect 9904 877 9916 911
rect 9950 877 9962 911
rect 10462 979 10520 1013
rect 10462 945 10474 979
rect 10508 945 10520 979
rect 10462 911 10520 945
rect 9904 862 9962 877
rect 10032 887 10094 902
rect 10032 853 10044 887
rect 10078 853 10094 887
rect 8332 717 8348 751
rect 8382 717 8394 751
rect 8332 702 8394 717
rect 10032 819 10094 853
rect 10032 785 10044 819
rect 10078 785 10094 819
rect 10032 751 10094 785
rect 10032 717 10044 751
rect 10078 717 10094 751
rect 10032 702 10094 717
rect 10124 887 10190 902
rect 10124 853 10140 887
rect 10174 853 10190 887
rect 10124 819 10190 853
rect 10124 785 10140 819
rect 10174 785 10190 819
rect 10124 751 10190 785
rect 10124 717 10140 751
rect 10174 717 10190 751
rect 10124 702 10190 717
rect 10220 887 10282 902
rect 10220 853 10236 887
rect 10270 853 10282 887
rect 10462 877 10474 911
rect 10508 877 10520 911
rect 10462 862 10520 877
rect 10550 1047 10608 1062
rect 10550 1013 10562 1047
rect 10596 1013 10608 1047
rect 10550 979 10608 1013
rect 10550 945 10562 979
rect 10596 945 10608 979
rect 10550 911 10608 945
rect 10550 877 10562 911
rect 10596 877 10608 911
rect 10744 1031 10752 1065
rect 10786 1031 10796 1065
rect 10744 997 10796 1031
rect 10744 963 10752 997
rect 10786 963 10796 997
rect 10744 929 10796 963
rect 10744 895 10752 929
rect 10786 895 10796 929
rect 10744 877 10796 895
rect 10826 1065 10878 1077
rect 10826 1031 10836 1065
rect 10870 1031 10878 1065
rect 10826 997 10878 1031
rect 10826 963 10836 997
rect 10870 963 10878 997
rect 10826 929 10878 963
rect 10826 895 10836 929
rect 10870 895 10878 929
rect 11049 1055 11101 1075
rect 11049 1021 11057 1055
rect 11091 1021 11101 1055
rect 11049 987 11101 1021
rect 11049 953 11057 987
rect 11091 953 11101 987
rect 11049 917 11101 953
rect 11131 1055 11189 1075
rect 11131 1021 11143 1055
rect 11177 1021 11189 1055
rect 11131 987 11189 1021
rect 11131 953 11143 987
rect 11177 953 11189 987
rect 11131 917 11189 953
rect 11219 1055 11271 1075
rect 11219 1021 11229 1055
rect 11263 1021 11271 1055
rect 11219 974 11271 1021
rect 11219 940 11229 974
rect 11263 940 11271 974
rect 11219 917 11271 940
rect 11436 1057 11488 1069
rect 11436 1023 11444 1057
rect 11478 1023 11488 1057
rect 11436 989 11488 1023
rect 11436 955 11444 989
rect 11478 955 11488 989
rect 11436 921 11488 955
rect 10826 877 10878 895
rect 10550 862 10608 877
rect 10220 819 10282 853
rect 10220 785 10236 819
rect 10270 785 10282 819
rect 10220 751 10282 785
rect 11436 887 11444 921
rect 11478 887 11488 921
rect 11436 869 11488 887
rect 11518 1057 11570 1069
rect 11518 1023 11528 1057
rect 11562 1023 11570 1057
rect 11518 989 11570 1023
rect 11518 955 11528 989
rect 11562 955 11570 989
rect 11518 921 11570 955
rect 11518 887 11528 921
rect 11562 887 11570 921
rect 11518 869 11570 887
rect 11704 1047 11762 1062
rect 11704 1013 11716 1047
rect 11750 1013 11762 1047
rect 11704 979 11762 1013
rect 11704 945 11716 979
rect 11750 945 11762 979
rect 11704 911 11762 945
rect 11704 877 11716 911
rect 11750 877 11762 911
rect 11704 862 11762 877
rect 11792 1047 11850 1062
rect 11792 1013 11804 1047
rect 11838 1013 11850 1047
rect 11792 979 11850 1013
rect 12632 1065 12684 1077
rect 12350 1047 12408 1062
rect 12350 1013 12362 1047
rect 12396 1013 12408 1047
rect 11792 945 11804 979
rect 11838 945 11850 979
rect 11792 911 11850 945
rect 11792 877 11804 911
rect 11838 877 11850 911
rect 12350 979 12408 1013
rect 12350 945 12362 979
rect 12396 945 12408 979
rect 12350 911 12408 945
rect 11792 862 11850 877
rect 11920 887 11982 902
rect 11920 853 11932 887
rect 11966 853 11982 887
rect 10220 717 10236 751
rect 10270 717 10282 751
rect 10220 702 10282 717
rect 11920 819 11982 853
rect 11920 785 11932 819
rect 11966 785 11982 819
rect 11920 751 11982 785
rect 11920 717 11932 751
rect 11966 717 11982 751
rect 11920 702 11982 717
rect 12012 887 12078 902
rect 12012 853 12028 887
rect 12062 853 12078 887
rect 12012 819 12078 853
rect 12012 785 12028 819
rect 12062 785 12078 819
rect 12012 751 12078 785
rect 12012 717 12028 751
rect 12062 717 12078 751
rect 12012 702 12078 717
rect 12108 887 12170 902
rect 12108 853 12124 887
rect 12158 853 12170 887
rect 12350 877 12362 911
rect 12396 877 12408 911
rect 12350 862 12408 877
rect 12438 1047 12496 1062
rect 12438 1013 12450 1047
rect 12484 1013 12496 1047
rect 12438 979 12496 1013
rect 12438 945 12450 979
rect 12484 945 12496 979
rect 12438 911 12496 945
rect 12438 877 12450 911
rect 12484 877 12496 911
rect 12632 1031 12640 1065
rect 12674 1031 12684 1065
rect 12632 997 12684 1031
rect 12632 963 12640 997
rect 12674 963 12684 997
rect 12632 929 12684 963
rect 12632 895 12640 929
rect 12674 895 12684 929
rect 12632 877 12684 895
rect 12714 1065 12766 1077
rect 12714 1031 12724 1065
rect 12758 1031 12766 1065
rect 12714 997 12766 1031
rect 12714 963 12724 997
rect 12758 963 12766 997
rect 12714 929 12766 963
rect 12714 895 12724 929
rect 12758 895 12766 929
rect 12937 1055 12989 1075
rect 12937 1021 12945 1055
rect 12979 1021 12989 1055
rect 12937 987 12989 1021
rect 12937 953 12945 987
rect 12979 953 12989 987
rect 12937 917 12989 953
rect 13019 1055 13077 1075
rect 13019 1021 13031 1055
rect 13065 1021 13077 1055
rect 13019 987 13077 1021
rect 13019 953 13031 987
rect 13065 953 13077 987
rect 13019 917 13077 953
rect 13107 1055 13159 1075
rect 13107 1021 13117 1055
rect 13151 1021 13159 1055
rect 13107 974 13159 1021
rect 13107 940 13117 974
rect 13151 940 13159 974
rect 13107 917 13159 940
rect 13324 1057 13376 1069
rect 13324 1023 13332 1057
rect 13366 1023 13376 1057
rect 13324 989 13376 1023
rect 13324 955 13332 989
rect 13366 955 13376 989
rect 13324 921 13376 955
rect 12714 877 12766 895
rect 12438 862 12496 877
rect 12108 819 12170 853
rect 12108 785 12124 819
rect 12158 785 12170 819
rect 12108 751 12170 785
rect 13324 887 13332 921
rect 13366 887 13376 921
rect 13324 869 13376 887
rect 13406 1057 13458 1069
rect 13406 1023 13416 1057
rect 13450 1023 13458 1057
rect 13406 989 13458 1023
rect 13406 955 13416 989
rect 13450 955 13458 989
rect 13406 921 13458 955
rect 13406 887 13416 921
rect 13450 887 13458 921
rect 13406 869 13458 887
rect 13592 1047 13650 1062
rect 13592 1013 13604 1047
rect 13638 1013 13650 1047
rect 13592 979 13650 1013
rect 13592 945 13604 979
rect 13638 945 13650 979
rect 13592 911 13650 945
rect 13592 877 13604 911
rect 13638 877 13650 911
rect 13592 862 13650 877
rect 13680 1047 13738 1062
rect 13680 1013 13692 1047
rect 13726 1013 13738 1047
rect 13680 979 13738 1013
rect 14520 1065 14572 1077
rect 14238 1047 14296 1062
rect 14238 1013 14250 1047
rect 14284 1013 14296 1047
rect 13680 945 13692 979
rect 13726 945 13738 979
rect 13680 911 13738 945
rect 13680 877 13692 911
rect 13726 877 13738 911
rect 14238 979 14296 1013
rect 14238 945 14250 979
rect 14284 945 14296 979
rect 14238 911 14296 945
rect 13680 862 13738 877
rect 13808 887 13870 902
rect 13808 853 13820 887
rect 13854 853 13870 887
rect 12108 717 12124 751
rect 12158 717 12170 751
rect 12108 702 12170 717
rect 13808 819 13870 853
rect 13808 785 13820 819
rect 13854 785 13870 819
rect 13808 751 13870 785
rect 13808 717 13820 751
rect 13854 717 13870 751
rect 13808 702 13870 717
rect 13900 887 13966 902
rect 13900 853 13916 887
rect 13950 853 13966 887
rect 13900 819 13966 853
rect 13900 785 13916 819
rect 13950 785 13966 819
rect 13900 751 13966 785
rect 13900 717 13916 751
rect 13950 717 13966 751
rect 13900 702 13966 717
rect 13996 887 14058 902
rect 13996 853 14012 887
rect 14046 853 14058 887
rect 14238 877 14250 911
rect 14284 877 14296 911
rect 14238 862 14296 877
rect 14326 1047 14384 1062
rect 14326 1013 14338 1047
rect 14372 1013 14384 1047
rect 14326 979 14384 1013
rect 14326 945 14338 979
rect 14372 945 14384 979
rect 14326 911 14384 945
rect 14326 877 14338 911
rect 14372 877 14384 911
rect 14520 1031 14528 1065
rect 14562 1031 14572 1065
rect 14520 997 14572 1031
rect 14520 963 14528 997
rect 14562 963 14572 997
rect 14520 929 14572 963
rect 14520 895 14528 929
rect 14562 895 14572 929
rect 14520 877 14572 895
rect 14602 1065 14654 1077
rect 14602 1031 14612 1065
rect 14646 1031 14654 1065
rect 14602 997 14654 1031
rect 14602 963 14612 997
rect 14646 963 14654 997
rect 14602 929 14654 963
rect 14602 895 14612 929
rect 14646 895 14654 929
rect 14825 1055 14877 1075
rect 14825 1021 14833 1055
rect 14867 1021 14877 1055
rect 14825 987 14877 1021
rect 14825 953 14833 987
rect 14867 953 14877 987
rect 14825 917 14877 953
rect 14907 1055 14965 1075
rect 14907 1021 14919 1055
rect 14953 1021 14965 1055
rect 14907 987 14965 1021
rect 14907 953 14919 987
rect 14953 953 14965 987
rect 14907 917 14965 953
rect 14995 1055 15047 1075
rect 14995 1021 15005 1055
rect 15039 1021 15047 1055
rect 14995 974 15047 1021
rect 14995 940 15005 974
rect 15039 940 15047 974
rect 14995 917 15047 940
rect 15206 1057 15258 1069
rect 15206 1023 15214 1057
rect 15248 1023 15258 1057
rect 15206 989 15258 1023
rect 15206 955 15214 989
rect 15248 955 15258 989
rect 15206 921 15258 955
rect 14602 877 14654 895
rect 14326 862 14384 877
rect 13996 819 14058 853
rect 13996 785 14012 819
rect 14046 785 14058 819
rect 13996 751 14058 785
rect 15206 887 15214 921
rect 15248 887 15258 921
rect 15206 869 15258 887
rect 15288 1057 15340 1069
rect 15288 1023 15298 1057
rect 15332 1023 15340 1057
rect 15288 989 15340 1023
rect 15288 955 15298 989
rect 15332 955 15340 989
rect 15288 921 15340 955
rect 15288 887 15298 921
rect 15332 887 15340 921
rect 15288 869 15340 887
rect 15474 1047 15532 1062
rect 15474 1013 15486 1047
rect 15520 1013 15532 1047
rect 15474 979 15532 1013
rect 15474 945 15486 979
rect 15520 945 15532 979
rect 15474 911 15532 945
rect 15474 877 15486 911
rect 15520 877 15532 911
rect 15474 862 15532 877
rect 15562 1047 15620 1062
rect 15562 1013 15574 1047
rect 15608 1013 15620 1047
rect 15562 979 15620 1013
rect 16402 1065 16454 1077
rect 16120 1047 16178 1062
rect 16120 1013 16132 1047
rect 16166 1013 16178 1047
rect 15562 945 15574 979
rect 15608 945 15620 979
rect 15562 911 15620 945
rect 15562 877 15574 911
rect 15608 877 15620 911
rect 16120 979 16178 1013
rect 16120 945 16132 979
rect 16166 945 16178 979
rect 16120 911 16178 945
rect 15562 862 15620 877
rect 15690 887 15752 902
rect 15690 853 15702 887
rect 15736 853 15752 887
rect 13996 717 14012 751
rect 14046 717 14058 751
rect 13996 702 14058 717
rect 15690 819 15752 853
rect 15690 785 15702 819
rect 15736 785 15752 819
rect 15690 751 15752 785
rect 15690 717 15702 751
rect 15736 717 15752 751
rect 15690 702 15752 717
rect 15782 887 15848 902
rect 15782 853 15798 887
rect 15832 853 15848 887
rect 15782 819 15848 853
rect 15782 785 15798 819
rect 15832 785 15848 819
rect 15782 751 15848 785
rect 15782 717 15798 751
rect 15832 717 15848 751
rect 15782 702 15848 717
rect 15878 887 15940 902
rect 15878 853 15894 887
rect 15928 853 15940 887
rect 16120 877 16132 911
rect 16166 877 16178 911
rect 16120 862 16178 877
rect 16208 1047 16266 1062
rect 16208 1013 16220 1047
rect 16254 1013 16266 1047
rect 16208 979 16266 1013
rect 16208 945 16220 979
rect 16254 945 16266 979
rect 16208 911 16266 945
rect 16208 877 16220 911
rect 16254 877 16266 911
rect 16402 1031 16410 1065
rect 16444 1031 16454 1065
rect 16402 997 16454 1031
rect 16402 963 16410 997
rect 16444 963 16454 997
rect 16402 929 16454 963
rect 16402 895 16410 929
rect 16444 895 16454 929
rect 16402 877 16454 895
rect 16484 1065 16536 1077
rect 16484 1031 16494 1065
rect 16528 1031 16536 1065
rect 16484 997 16536 1031
rect 16484 963 16494 997
rect 16528 963 16536 997
rect 16484 929 16536 963
rect 16484 895 16494 929
rect 16528 895 16536 929
rect 16707 1055 16759 1075
rect 16707 1021 16715 1055
rect 16749 1021 16759 1055
rect 16707 987 16759 1021
rect 16707 953 16715 987
rect 16749 953 16759 987
rect 16707 917 16759 953
rect 16789 1055 16847 1075
rect 16789 1021 16801 1055
rect 16835 1021 16847 1055
rect 16789 987 16847 1021
rect 16789 953 16801 987
rect 16835 953 16847 987
rect 16789 917 16847 953
rect 16877 1055 16929 1075
rect 16877 1021 16887 1055
rect 16921 1021 16929 1055
rect 16877 974 16929 1021
rect 16877 940 16887 974
rect 16921 940 16929 974
rect 16877 917 16929 940
rect 17094 1057 17146 1069
rect 17094 1023 17102 1057
rect 17136 1023 17146 1057
rect 17094 989 17146 1023
rect 17094 955 17102 989
rect 17136 955 17146 989
rect 17094 921 17146 955
rect 16484 877 16536 895
rect 16208 862 16266 877
rect 15878 819 15940 853
rect 15878 785 15894 819
rect 15928 785 15940 819
rect 15878 751 15940 785
rect 17094 887 17102 921
rect 17136 887 17146 921
rect 17094 869 17146 887
rect 17176 1057 17228 1069
rect 17176 1023 17186 1057
rect 17220 1023 17228 1057
rect 17176 989 17228 1023
rect 17176 955 17186 989
rect 17220 955 17228 989
rect 17176 921 17228 955
rect 17176 887 17186 921
rect 17220 887 17228 921
rect 17176 869 17228 887
rect 17362 1047 17420 1062
rect 17362 1013 17374 1047
rect 17408 1013 17420 1047
rect 17362 979 17420 1013
rect 17362 945 17374 979
rect 17408 945 17420 979
rect 17362 911 17420 945
rect 17362 877 17374 911
rect 17408 877 17420 911
rect 17362 862 17420 877
rect 17450 1047 17508 1062
rect 17450 1013 17462 1047
rect 17496 1013 17508 1047
rect 17450 979 17508 1013
rect 18290 1065 18342 1077
rect 18008 1047 18066 1062
rect 18008 1013 18020 1047
rect 18054 1013 18066 1047
rect 17450 945 17462 979
rect 17496 945 17508 979
rect 17450 911 17508 945
rect 17450 877 17462 911
rect 17496 877 17508 911
rect 18008 979 18066 1013
rect 18008 945 18020 979
rect 18054 945 18066 979
rect 18008 911 18066 945
rect 17450 862 17508 877
rect 17578 887 17640 902
rect 17578 853 17590 887
rect 17624 853 17640 887
rect 15878 717 15894 751
rect 15928 717 15940 751
rect 15878 702 15940 717
rect 17578 819 17640 853
rect 17578 785 17590 819
rect 17624 785 17640 819
rect 17578 751 17640 785
rect 17578 717 17590 751
rect 17624 717 17640 751
rect 17578 702 17640 717
rect 17670 887 17736 902
rect 17670 853 17686 887
rect 17720 853 17736 887
rect 17670 819 17736 853
rect 17670 785 17686 819
rect 17720 785 17736 819
rect 17670 751 17736 785
rect 17670 717 17686 751
rect 17720 717 17736 751
rect 17670 702 17736 717
rect 17766 887 17828 902
rect 17766 853 17782 887
rect 17816 853 17828 887
rect 18008 877 18020 911
rect 18054 877 18066 911
rect 18008 862 18066 877
rect 18096 1047 18154 1062
rect 18096 1013 18108 1047
rect 18142 1013 18154 1047
rect 18096 979 18154 1013
rect 18096 945 18108 979
rect 18142 945 18154 979
rect 18096 911 18154 945
rect 18096 877 18108 911
rect 18142 877 18154 911
rect 18290 1031 18298 1065
rect 18332 1031 18342 1065
rect 18290 997 18342 1031
rect 18290 963 18298 997
rect 18332 963 18342 997
rect 18290 929 18342 963
rect 18290 895 18298 929
rect 18332 895 18342 929
rect 18290 877 18342 895
rect 18372 1065 18424 1077
rect 18372 1031 18382 1065
rect 18416 1031 18424 1065
rect 18372 997 18424 1031
rect 18372 963 18382 997
rect 18416 963 18424 997
rect 18372 929 18424 963
rect 18372 895 18382 929
rect 18416 895 18424 929
rect 18595 1055 18647 1075
rect 18595 1021 18603 1055
rect 18637 1021 18647 1055
rect 18595 987 18647 1021
rect 18595 953 18603 987
rect 18637 953 18647 987
rect 18595 917 18647 953
rect 18677 1055 18735 1075
rect 18677 1021 18689 1055
rect 18723 1021 18735 1055
rect 18677 987 18735 1021
rect 18677 953 18689 987
rect 18723 953 18735 987
rect 18677 917 18735 953
rect 18765 1055 18817 1075
rect 18765 1021 18775 1055
rect 18809 1021 18817 1055
rect 18765 974 18817 1021
rect 18765 940 18775 974
rect 18809 940 18817 974
rect 18765 917 18817 940
rect 18982 1057 19034 1069
rect 18982 1023 18990 1057
rect 19024 1023 19034 1057
rect 18982 989 19034 1023
rect 18982 955 18990 989
rect 19024 955 19034 989
rect 18982 921 19034 955
rect 18372 877 18424 895
rect 18096 862 18154 877
rect 17766 819 17828 853
rect 17766 785 17782 819
rect 17816 785 17828 819
rect 17766 751 17828 785
rect 18982 887 18990 921
rect 19024 887 19034 921
rect 18982 869 19034 887
rect 19064 1057 19116 1069
rect 19064 1023 19074 1057
rect 19108 1023 19116 1057
rect 19064 989 19116 1023
rect 19064 955 19074 989
rect 19108 955 19116 989
rect 19064 921 19116 955
rect 19064 887 19074 921
rect 19108 887 19116 921
rect 19064 869 19116 887
rect 19250 1047 19308 1062
rect 19250 1013 19262 1047
rect 19296 1013 19308 1047
rect 19250 979 19308 1013
rect 19250 945 19262 979
rect 19296 945 19308 979
rect 19250 911 19308 945
rect 19250 877 19262 911
rect 19296 877 19308 911
rect 19250 862 19308 877
rect 19338 1047 19396 1062
rect 19338 1013 19350 1047
rect 19384 1013 19396 1047
rect 19338 979 19396 1013
rect 20178 1065 20230 1077
rect 19896 1047 19954 1062
rect 19896 1013 19908 1047
rect 19942 1013 19954 1047
rect 19338 945 19350 979
rect 19384 945 19396 979
rect 19338 911 19396 945
rect 19338 877 19350 911
rect 19384 877 19396 911
rect 19896 979 19954 1013
rect 19896 945 19908 979
rect 19942 945 19954 979
rect 19896 911 19954 945
rect 19338 862 19396 877
rect 19466 887 19528 902
rect 19466 853 19478 887
rect 19512 853 19528 887
rect 17766 717 17782 751
rect 17816 717 17828 751
rect 17766 702 17828 717
rect 19466 819 19528 853
rect 19466 785 19478 819
rect 19512 785 19528 819
rect 19466 751 19528 785
rect 19466 717 19478 751
rect 19512 717 19528 751
rect 19466 702 19528 717
rect 19558 887 19624 902
rect 19558 853 19574 887
rect 19608 853 19624 887
rect 19558 819 19624 853
rect 19558 785 19574 819
rect 19608 785 19624 819
rect 19558 751 19624 785
rect 19558 717 19574 751
rect 19608 717 19624 751
rect 19558 702 19624 717
rect 19654 887 19716 902
rect 19654 853 19670 887
rect 19704 853 19716 887
rect 19896 877 19908 911
rect 19942 877 19954 911
rect 19896 862 19954 877
rect 19984 1047 20042 1062
rect 19984 1013 19996 1047
rect 20030 1013 20042 1047
rect 19984 979 20042 1013
rect 19984 945 19996 979
rect 20030 945 20042 979
rect 19984 911 20042 945
rect 19984 877 19996 911
rect 20030 877 20042 911
rect 20178 1031 20186 1065
rect 20220 1031 20230 1065
rect 20178 997 20230 1031
rect 20178 963 20186 997
rect 20220 963 20230 997
rect 20178 929 20230 963
rect 20178 895 20186 929
rect 20220 895 20230 929
rect 20178 877 20230 895
rect 20260 1065 20312 1077
rect 20260 1031 20270 1065
rect 20304 1031 20312 1065
rect 20260 997 20312 1031
rect 20260 963 20270 997
rect 20304 963 20312 997
rect 20260 929 20312 963
rect 20260 895 20270 929
rect 20304 895 20312 929
rect 20483 1055 20535 1075
rect 20483 1021 20491 1055
rect 20525 1021 20535 1055
rect 20483 987 20535 1021
rect 20483 953 20491 987
rect 20525 953 20535 987
rect 20483 917 20535 953
rect 20565 1055 20623 1075
rect 20565 1021 20577 1055
rect 20611 1021 20623 1055
rect 20565 987 20623 1021
rect 20565 953 20577 987
rect 20611 953 20623 987
rect 20565 917 20623 953
rect 20653 1055 20705 1075
rect 20653 1021 20663 1055
rect 20697 1021 20705 1055
rect 20653 974 20705 1021
rect 20653 940 20663 974
rect 20697 940 20705 974
rect 20653 917 20705 940
rect 20870 1057 20922 1069
rect 20870 1023 20878 1057
rect 20912 1023 20922 1057
rect 20870 989 20922 1023
rect 20870 955 20878 989
rect 20912 955 20922 989
rect 20870 921 20922 955
rect 20260 877 20312 895
rect 19984 862 20042 877
rect 19654 819 19716 853
rect 19654 785 19670 819
rect 19704 785 19716 819
rect 19654 751 19716 785
rect 20870 887 20878 921
rect 20912 887 20922 921
rect 20870 869 20922 887
rect 20952 1057 21004 1069
rect 20952 1023 20962 1057
rect 20996 1023 21004 1057
rect 20952 989 21004 1023
rect 20952 955 20962 989
rect 20996 955 21004 989
rect 20952 921 21004 955
rect 20952 887 20962 921
rect 20996 887 21004 921
rect 20952 869 21004 887
rect 21138 1047 21196 1062
rect 21138 1013 21150 1047
rect 21184 1013 21196 1047
rect 21138 979 21196 1013
rect 21138 945 21150 979
rect 21184 945 21196 979
rect 21138 911 21196 945
rect 21138 877 21150 911
rect 21184 877 21196 911
rect 21138 862 21196 877
rect 21226 1047 21284 1062
rect 21226 1013 21238 1047
rect 21272 1013 21284 1047
rect 21226 979 21284 1013
rect 22066 1065 22118 1077
rect 21784 1047 21842 1062
rect 21784 1013 21796 1047
rect 21830 1013 21842 1047
rect 21226 945 21238 979
rect 21272 945 21284 979
rect 21226 911 21284 945
rect 21226 877 21238 911
rect 21272 877 21284 911
rect 21784 979 21842 1013
rect 21784 945 21796 979
rect 21830 945 21842 979
rect 21784 911 21842 945
rect 21226 862 21284 877
rect 21354 887 21416 902
rect 21354 853 21366 887
rect 21400 853 21416 887
rect 19654 717 19670 751
rect 19704 717 19716 751
rect 19654 702 19716 717
rect 21354 819 21416 853
rect 21354 785 21366 819
rect 21400 785 21416 819
rect 21354 751 21416 785
rect 21354 717 21366 751
rect 21400 717 21416 751
rect 21354 702 21416 717
rect 21446 887 21512 902
rect 21446 853 21462 887
rect 21496 853 21512 887
rect 21446 819 21512 853
rect 21446 785 21462 819
rect 21496 785 21512 819
rect 21446 751 21512 785
rect 21446 717 21462 751
rect 21496 717 21512 751
rect 21446 702 21512 717
rect 21542 887 21604 902
rect 21542 853 21558 887
rect 21592 853 21604 887
rect 21784 877 21796 911
rect 21830 877 21842 911
rect 21784 862 21842 877
rect 21872 1047 21930 1062
rect 21872 1013 21884 1047
rect 21918 1013 21930 1047
rect 21872 979 21930 1013
rect 21872 945 21884 979
rect 21918 945 21930 979
rect 21872 911 21930 945
rect 21872 877 21884 911
rect 21918 877 21930 911
rect 22066 1031 22074 1065
rect 22108 1031 22118 1065
rect 22066 997 22118 1031
rect 22066 963 22074 997
rect 22108 963 22118 997
rect 22066 929 22118 963
rect 22066 895 22074 929
rect 22108 895 22118 929
rect 22066 877 22118 895
rect 22148 1065 22200 1077
rect 22148 1031 22158 1065
rect 22192 1031 22200 1065
rect 22148 997 22200 1031
rect 22148 963 22158 997
rect 22192 963 22200 997
rect 22148 929 22200 963
rect 22148 895 22158 929
rect 22192 895 22200 929
rect 22371 1055 22423 1075
rect 22371 1021 22379 1055
rect 22413 1021 22423 1055
rect 22371 987 22423 1021
rect 22371 953 22379 987
rect 22413 953 22423 987
rect 22371 917 22423 953
rect 22453 1055 22511 1075
rect 22453 1021 22465 1055
rect 22499 1021 22511 1055
rect 22453 987 22511 1021
rect 22453 953 22465 987
rect 22499 953 22511 987
rect 22453 917 22511 953
rect 22541 1055 22593 1075
rect 22541 1021 22551 1055
rect 22585 1021 22593 1055
rect 22541 974 22593 1021
rect 22541 940 22551 974
rect 22585 940 22593 974
rect 22541 917 22593 940
rect 22758 1057 22810 1069
rect 22758 1023 22766 1057
rect 22800 1023 22810 1057
rect 22758 989 22810 1023
rect 22758 955 22766 989
rect 22800 955 22810 989
rect 22758 921 22810 955
rect 22148 877 22200 895
rect 21872 862 21930 877
rect 21542 819 21604 853
rect 21542 785 21558 819
rect 21592 785 21604 819
rect 21542 751 21604 785
rect 22758 887 22766 921
rect 22800 887 22810 921
rect 22758 869 22810 887
rect 22840 1057 22892 1069
rect 22840 1023 22850 1057
rect 22884 1023 22892 1057
rect 22840 989 22892 1023
rect 22840 955 22850 989
rect 22884 955 22892 989
rect 22840 921 22892 955
rect 22840 887 22850 921
rect 22884 887 22892 921
rect 22840 869 22892 887
rect 23026 1047 23084 1062
rect 23026 1013 23038 1047
rect 23072 1013 23084 1047
rect 23026 979 23084 1013
rect 23026 945 23038 979
rect 23072 945 23084 979
rect 23026 911 23084 945
rect 23026 877 23038 911
rect 23072 877 23084 911
rect 23026 862 23084 877
rect 23114 1047 23172 1062
rect 23114 1013 23126 1047
rect 23160 1013 23172 1047
rect 23114 979 23172 1013
rect 23954 1065 24006 1077
rect 23672 1047 23730 1062
rect 23672 1013 23684 1047
rect 23718 1013 23730 1047
rect 23114 945 23126 979
rect 23160 945 23172 979
rect 23114 911 23172 945
rect 23114 877 23126 911
rect 23160 877 23172 911
rect 23672 979 23730 1013
rect 23672 945 23684 979
rect 23718 945 23730 979
rect 23672 911 23730 945
rect 23114 862 23172 877
rect 23242 887 23304 902
rect 23242 853 23254 887
rect 23288 853 23304 887
rect 21542 717 21558 751
rect 21592 717 21604 751
rect 21542 702 21604 717
rect 23242 819 23304 853
rect 23242 785 23254 819
rect 23288 785 23304 819
rect 23242 751 23304 785
rect 23242 717 23254 751
rect 23288 717 23304 751
rect 23242 702 23304 717
rect 23334 887 23400 902
rect 23334 853 23350 887
rect 23384 853 23400 887
rect 23334 819 23400 853
rect 23334 785 23350 819
rect 23384 785 23400 819
rect 23334 751 23400 785
rect 23334 717 23350 751
rect 23384 717 23400 751
rect 23334 702 23400 717
rect 23430 887 23492 902
rect 23430 853 23446 887
rect 23480 853 23492 887
rect 23672 877 23684 911
rect 23718 877 23730 911
rect 23672 862 23730 877
rect 23760 1047 23818 1062
rect 23760 1013 23772 1047
rect 23806 1013 23818 1047
rect 23760 979 23818 1013
rect 23760 945 23772 979
rect 23806 945 23818 979
rect 23760 911 23818 945
rect 23760 877 23772 911
rect 23806 877 23818 911
rect 23954 1031 23962 1065
rect 23996 1031 24006 1065
rect 23954 997 24006 1031
rect 23954 963 23962 997
rect 23996 963 24006 997
rect 23954 929 24006 963
rect 23954 895 23962 929
rect 23996 895 24006 929
rect 23954 877 24006 895
rect 24036 1065 24088 1077
rect 24036 1031 24046 1065
rect 24080 1031 24088 1065
rect 24036 997 24088 1031
rect 24036 963 24046 997
rect 24080 963 24088 997
rect 24036 929 24088 963
rect 24036 895 24046 929
rect 24080 895 24088 929
rect 24259 1055 24311 1075
rect 24259 1021 24267 1055
rect 24301 1021 24311 1055
rect 24259 987 24311 1021
rect 24259 953 24267 987
rect 24301 953 24311 987
rect 24259 917 24311 953
rect 24341 1055 24399 1075
rect 24341 1021 24353 1055
rect 24387 1021 24399 1055
rect 24341 987 24399 1021
rect 24341 953 24353 987
rect 24387 953 24399 987
rect 24341 917 24399 953
rect 24429 1055 24481 1075
rect 24429 1021 24439 1055
rect 24473 1021 24481 1055
rect 24429 974 24481 1021
rect 24429 940 24439 974
rect 24473 940 24481 974
rect 24429 917 24481 940
rect 24646 1057 24698 1069
rect 24646 1023 24654 1057
rect 24688 1023 24698 1057
rect 24646 989 24698 1023
rect 24646 955 24654 989
rect 24688 955 24698 989
rect 24646 921 24698 955
rect 24036 877 24088 895
rect 23760 862 23818 877
rect 23430 819 23492 853
rect 23430 785 23446 819
rect 23480 785 23492 819
rect 23430 751 23492 785
rect 24646 887 24654 921
rect 24688 887 24698 921
rect 24646 869 24698 887
rect 24728 1057 24780 1069
rect 24728 1023 24738 1057
rect 24772 1023 24780 1057
rect 24728 989 24780 1023
rect 24728 955 24738 989
rect 24772 955 24780 989
rect 24728 921 24780 955
rect 24728 887 24738 921
rect 24772 887 24780 921
rect 24728 869 24780 887
rect 24914 1047 24972 1062
rect 24914 1013 24926 1047
rect 24960 1013 24972 1047
rect 24914 979 24972 1013
rect 24914 945 24926 979
rect 24960 945 24972 979
rect 24914 911 24972 945
rect 24914 877 24926 911
rect 24960 877 24972 911
rect 24914 862 24972 877
rect 25002 1047 25060 1062
rect 25002 1013 25014 1047
rect 25048 1013 25060 1047
rect 25002 979 25060 1013
rect 25842 1065 25894 1077
rect 25560 1047 25618 1062
rect 25560 1013 25572 1047
rect 25606 1013 25618 1047
rect 25002 945 25014 979
rect 25048 945 25060 979
rect 25002 911 25060 945
rect 25002 877 25014 911
rect 25048 877 25060 911
rect 25560 979 25618 1013
rect 25560 945 25572 979
rect 25606 945 25618 979
rect 25560 911 25618 945
rect 25002 862 25060 877
rect 25130 887 25192 902
rect 25130 853 25142 887
rect 25176 853 25192 887
rect 23430 717 23446 751
rect 23480 717 23492 751
rect 23430 702 23492 717
rect 25130 819 25192 853
rect 25130 785 25142 819
rect 25176 785 25192 819
rect 25130 751 25192 785
rect 25130 717 25142 751
rect 25176 717 25192 751
rect 25130 702 25192 717
rect 25222 887 25288 902
rect 25222 853 25238 887
rect 25272 853 25288 887
rect 25222 819 25288 853
rect 25222 785 25238 819
rect 25272 785 25288 819
rect 25222 751 25288 785
rect 25222 717 25238 751
rect 25272 717 25288 751
rect 25222 702 25288 717
rect 25318 887 25380 902
rect 25318 853 25334 887
rect 25368 853 25380 887
rect 25560 877 25572 911
rect 25606 877 25618 911
rect 25560 862 25618 877
rect 25648 1047 25706 1062
rect 25648 1013 25660 1047
rect 25694 1013 25706 1047
rect 25648 979 25706 1013
rect 25648 945 25660 979
rect 25694 945 25706 979
rect 25648 911 25706 945
rect 25648 877 25660 911
rect 25694 877 25706 911
rect 25842 1031 25850 1065
rect 25884 1031 25894 1065
rect 25842 997 25894 1031
rect 25842 963 25850 997
rect 25884 963 25894 997
rect 25842 929 25894 963
rect 25842 895 25850 929
rect 25884 895 25894 929
rect 25842 877 25894 895
rect 25924 1065 25976 1077
rect 25924 1031 25934 1065
rect 25968 1031 25976 1065
rect 25924 997 25976 1031
rect 25924 963 25934 997
rect 25968 963 25976 997
rect 25924 929 25976 963
rect 25924 895 25934 929
rect 25968 895 25976 929
rect 26147 1055 26199 1075
rect 26147 1021 26155 1055
rect 26189 1021 26199 1055
rect 26147 987 26199 1021
rect 26147 953 26155 987
rect 26189 953 26199 987
rect 26147 917 26199 953
rect 26229 1055 26287 1075
rect 26229 1021 26241 1055
rect 26275 1021 26287 1055
rect 26229 987 26287 1021
rect 26229 953 26241 987
rect 26275 953 26287 987
rect 26229 917 26287 953
rect 26317 1055 26369 1075
rect 26317 1021 26327 1055
rect 26361 1021 26369 1055
rect 26317 974 26369 1021
rect 26317 940 26327 974
rect 26361 940 26369 974
rect 26317 917 26369 940
rect 26534 1057 26586 1069
rect 26534 1023 26542 1057
rect 26576 1023 26586 1057
rect 26534 989 26586 1023
rect 26534 955 26542 989
rect 26576 955 26586 989
rect 26534 921 26586 955
rect 25924 877 25976 895
rect 25648 862 25706 877
rect 25318 819 25380 853
rect 25318 785 25334 819
rect 25368 785 25380 819
rect 25318 751 25380 785
rect 26534 887 26542 921
rect 26576 887 26586 921
rect 26534 869 26586 887
rect 26616 1057 26668 1069
rect 26616 1023 26626 1057
rect 26660 1023 26668 1057
rect 26616 989 26668 1023
rect 26616 955 26626 989
rect 26660 955 26668 989
rect 26616 921 26668 955
rect 26616 887 26626 921
rect 26660 887 26668 921
rect 26616 869 26668 887
rect 26802 1047 26860 1062
rect 26802 1013 26814 1047
rect 26848 1013 26860 1047
rect 26802 979 26860 1013
rect 26802 945 26814 979
rect 26848 945 26860 979
rect 26802 911 26860 945
rect 26802 877 26814 911
rect 26848 877 26860 911
rect 26802 862 26860 877
rect 26890 1047 26948 1062
rect 26890 1013 26902 1047
rect 26936 1013 26948 1047
rect 26890 979 26948 1013
rect 27730 1065 27782 1077
rect 27448 1047 27506 1062
rect 27448 1013 27460 1047
rect 27494 1013 27506 1047
rect 26890 945 26902 979
rect 26936 945 26948 979
rect 26890 911 26948 945
rect 26890 877 26902 911
rect 26936 877 26948 911
rect 27448 979 27506 1013
rect 27448 945 27460 979
rect 27494 945 27506 979
rect 27448 911 27506 945
rect 26890 862 26948 877
rect 27018 887 27080 902
rect 27018 853 27030 887
rect 27064 853 27080 887
rect 25318 717 25334 751
rect 25368 717 25380 751
rect 25318 702 25380 717
rect 27018 819 27080 853
rect 27018 785 27030 819
rect 27064 785 27080 819
rect 27018 751 27080 785
rect 27018 717 27030 751
rect 27064 717 27080 751
rect 27018 702 27080 717
rect 27110 887 27176 902
rect 27110 853 27126 887
rect 27160 853 27176 887
rect 27110 819 27176 853
rect 27110 785 27126 819
rect 27160 785 27176 819
rect 27110 751 27176 785
rect 27110 717 27126 751
rect 27160 717 27176 751
rect 27110 702 27176 717
rect 27206 887 27268 902
rect 27206 853 27222 887
rect 27256 853 27268 887
rect 27448 877 27460 911
rect 27494 877 27506 911
rect 27448 862 27506 877
rect 27536 1047 27594 1062
rect 27536 1013 27548 1047
rect 27582 1013 27594 1047
rect 27536 979 27594 1013
rect 27536 945 27548 979
rect 27582 945 27594 979
rect 27536 911 27594 945
rect 27536 877 27548 911
rect 27582 877 27594 911
rect 27730 1031 27738 1065
rect 27772 1031 27782 1065
rect 27730 997 27782 1031
rect 27730 963 27738 997
rect 27772 963 27782 997
rect 27730 929 27782 963
rect 27730 895 27738 929
rect 27772 895 27782 929
rect 27730 877 27782 895
rect 27812 1065 27864 1077
rect 27812 1031 27822 1065
rect 27856 1031 27864 1065
rect 27812 997 27864 1031
rect 27812 963 27822 997
rect 27856 963 27864 997
rect 27812 929 27864 963
rect 27812 895 27822 929
rect 27856 895 27864 929
rect 28035 1055 28087 1075
rect 28035 1021 28043 1055
rect 28077 1021 28087 1055
rect 28035 987 28087 1021
rect 28035 953 28043 987
rect 28077 953 28087 987
rect 28035 917 28087 953
rect 28117 1055 28175 1075
rect 28117 1021 28129 1055
rect 28163 1021 28175 1055
rect 28117 987 28175 1021
rect 28117 953 28129 987
rect 28163 953 28175 987
rect 28117 917 28175 953
rect 28205 1055 28257 1075
rect 28205 1021 28215 1055
rect 28249 1021 28257 1055
rect 28205 974 28257 1021
rect 28205 940 28215 974
rect 28249 940 28257 974
rect 28205 917 28257 940
rect 28422 1057 28474 1069
rect 28422 1023 28430 1057
rect 28464 1023 28474 1057
rect 28422 989 28474 1023
rect 28422 955 28430 989
rect 28464 955 28474 989
rect 28422 921 28474 955
rect 27812 877 27864 895
rect 27536 862 27594 877
rect 27206 819 27268 853
rect 27206 785 27222 819
rect 27256 785 27268 819
rect 27206 751 27268 785
rect 28422 887 28430 921
rect 28464 887 28474 921
rect 28422 869 28474 887
rect 28504 1057 28556 1069
rect 28504 1023 28514 1057
rect 28548 1023 28556 1057
rect 28504 989 28556 1023
rect 28504 955 28514 989
rect 28548 955 28556 989
rect 28504 921 28556 955
rect 28504 887 28514 921
rect 28548 887 28556 921
rect 28504 869 28556 887
rect 28690 1047 28748 1062
rect 28690 1013 28702 1047
rect 28736 1013 28748 1047
rect 28690 979 28748 1013
rect 28690 945 28702 979
rect 28736 945 28748 979
rect 28690 911 28748 945
rect 28690 877 28702 911
rect 28736 877 28748 911
rect 28690 862 28748 877
rect 28778 1047 28836 1062
rect 28778 1013 28790 1047
rect 28824 1013 28836 1047
rect 28778 979 28836 1013
rect 29618 1065 29670 1077
rect 29336 1047 29394 1062
rect 29336 1013 29348 1047
rect 29382 1013 29394 1047
rect 28778 945 28790 979
rect 28824 945 28836 979
rect 28778 911 28836 945
rect 28778 877 28790 911
rect 28824 877 28836 911
rect 29336 979 29394 1013
rect 29336 945 29348 979
rect 29382 945 29394 979
rect 29336 911 29394 945
rect 28778 862 28836 877
rect 28906 887 28968 902
rect 28906 853 28918 887
rect 28952 853 28968 887
rect 27206 717 27222 751
rect 27256 717 27268 751
rect 27206 702 27268 717
rect 28906 819 28968 853
rect 28906 785 28918 819
rect 28952 785 28968 819
rect 28906 751 28968 785
rect 28906 717 28918 751
rect 28952 717 28968 751
rect 28906 702 28968 717
rect 28998 887 29064 902
rect 28998 853 29014 887
rect 29048 853 29064 887
rect 28998 819 29064 853
rect 28998 785 29014 819
rect 29048 785 29064 819
rect 28998 751 29064 785
rect 28998 717 29014 751
rect 29048 717 29064 751
rect 28998 702 29064 717
rect 29094 887 29156 902
rect 29094 853 29110 887
rect 29144 853 29156 887
rect 29336 877 29348 911
rect 29382 877 29394 911
rect 29336 862 29394 877
rect 29424 1047 29482 1062
rect 29424 1013 29436 1047
rect 29470 1013 29482 1047
rect 29424 979 29482 1013
rect 29424 945 29436 979
rect 29470 945 29482 979
rect 29424 911 29482 945
rect 29424 877 29436 911
rect 29470 877 29482 911
rect 29618 1031 29626 1065
rect 29660 1031 29670 1065
rect 29618 997 29670 1031
rect 29618 963 29626 997
rect 29660 963 29670 997
rect 29618 929 29670 963
rect 29618 895 29626 929
rect 29660 895 29670 929
rect 29618 877 29670 895
rect 29700 1065 29752 1077
rect 29700 1031 29710 1065
rect 29744 1031 29752 1065
rect 29700 997 29752 1031
rect 29700 963 29710 997
rect 29744 963 29752 997
rect 29700 929 29752 963
rect 29700 895 29710 929
rect 29744 895 29752 929
rect 29923 1055 29975 1075
rect 29923 1021 29931 1055
rect 29965 1021 29975 1055
rect 29923 987 29975 1021
rect 29923 953 29931 987
rect 29965 953 29975 987
rect 29923 917 29975 953
rect 30005 1055 30063 1075
rect 30005 1021 30017 1055
rect 30051 1021 30063 1055
rect 30005 987 30063 1021
rect 30005 953 30017 987
rect 30051 953 30063 987
rect 30005 917 30063 953
rect 30093 1055 30145 1075
rect 30093 1021 30103 1055
rect 30137 1021 30145 1055
rect 30093 974 30145 1021
rect 30093 940 30103 974
rect 30137 940 30145 974
rect 30093 917 30145 940
rect 30310 1057 30362 1069
rect 30310 1023 30318 1057
rect 30352 1023 30362 1057
rect 30310 989 30362 1023
rect 30310 955 30318 989
rect 30352 955 30362 989
rect 30310 921 30362 955
rect 29700 877 29752 895
rect 29424 862 29482 877
rect 29094 819 29156 853
rect 29094 785 29110 819
rect 29144 785 29156 819
rect 29094 751 29156 785
rect 30310 887 30318 921
rect 30352 887 30362 921
rect 30310 869 30362 887
rect 30392 1057 30444 1069
rect 30392 1023 30402 1057
rect 30436 1023 30444 1057
rect 30392 989 30444 1023
rect 30392 955 30402 989
rect 30436 955 30444 989
rect 30392 921 30444 955
rect 30392 887 30402 921
rect 30436 887 30444 921
rect 30392 869 30444 887
rect 30578 1047 30636 1062
rect 30578 1013 30590 1047
rect 30624 1013 30636 1047
rect 30578 979 30636 1013
rect 30578 945 30590 979
rect 30624 945 30636 979
rect 30578 911 30636 945
rect 30578 877 30590 911
rect 30624 877 30636 911
rect 30578 862 30636 877
rect 30666 1047 30724 1062
rect 30666 1013 30678 1047
rect 30712 1013 30724 1047
rect 30666 979 30724 1013
rect 31506 1065 31558 1077
rect 31224 1047 31282 1062
rect 31224 1013 31236 1047
rect 31270 1013 31282 1047
rect 30666 945 30678 979
rect 30712 945 30724 979
rect 30666 911 30724 945
rect 30666 877 30678 911
rect 30712 877 30724 911
rect 31224 979 31282 1013
rect 31224 945 31236 979
rect 31270 945 31282 979
rect 31224 911 31282 945
rect 30666 862 30724 877
rect 30794 887 30856 902
rect 30794 853 30806 887
rect 30840 853 30856 887
rect 29094 717 29110 751
rect 29144 717 29156 751
rect 29094 702 29156 717
rect 30794 819 30856 853
rect 30794 785 30806 819
rect 30840 785 30856 819
rect 30794 751 30856 785
rect 30794 717 30806 751
rect 30840 717 30856 751
rect 30794 702 30856 717
rect 30886 887 30952 902
rect 30886 853 30902 887
rect 30936 853 30952 887
rect 30886 819 30952 853
rect 30886 785 30902 819
rect 30936 785 30952 819
rect 30886 751 30952 785
rect 30886 717 30902 751
rect 30936 717 30952 751
rect 30886 702 30952 717
rect 30982 887 31044 902
rect 30982 853 30998 887
rect 31032 853 31044 887
rect 31224 877 31236 911
rect 31270 877 31282 911
rect 31224 862 31282 877
rect 31312 1047 31370 1062
rect 31312 1013 31324 1047
rect 31358 1013 31370 1047
rect 31312 979 31370 1013
rect 31312 945 31324 979
rect 31358 945 31370 979
rect 31312 911 31370 945
rect 31312 877 31324 911
rect 31358 877 31370 911
rect 31506 1031 31514 1065
rect 31548 1031 31558 1065
rect 31506 997 31558 1031
rect 31506 963 31514 997
rect 31548 963 31558 997
rect 31506 929 31558 963
rect 31506 895 31514 929
rect 31548 895 31558 929
rect 31506 877 31558 895
rect 31588 1065 31640 1077
rect 31588 1031 31598 1065
rect 31632 1031 31640 1065
rect 31588 997 31640 1031
rect 31588 963 31598 997
rect 31632 963 31640 997
rect 31588 929 31640 963
rect 31588 895 31598 929
rect 31632 895 31640 929
rect 31811 1055 31863 1075
rect 31811 1021 31819 1055
rect 31853 1021 31863 1055
rect 31811 987 31863 1021
rect 31811 953 31819 987
rect 31853 953 31863 987
rect 31811 917 31863 953
rect 31893 1055 31951 1075
rect 31893 1021 31905 1055
rect 31939 1021 31951 1055
rect 31893 987 31951 1021
rect 31893 953 31905 987
rect 31939 953 31951 987
rect 31893 917 31951 953
rect 31981 1055 32033 1075
rect 31981 1021 31991 1055
rect 32025 1021 32033 1055
rect 31981 974 32033 1021
rect 31981 940 31991 974
rect 32025 940 32033 974
rect 31981 917 32033 940
rect 32198 1057 32250 1069
rect 32198 1023 32206 1057
rect 32240 1023 32250 1057
rect 32198 989 32250 1023
rect 32198 955 32206 989
rect 32240 955 32250 989
rect 32198 921 32250 955
rect 31588 877 31640 895
rect 31312 862 31370 877
rect 30982 819 31044 853
rect 30982 785 30998 819
rect 31032 785 31044 819
rect 30982 751 31044 785
rect 32198 887 32206 921
rect 32240 887 32250 921
rect 32198 869 32250 887
rect 32280 1057 32332 1069
rect 32280 1023 32290 1057
rect 32324 1023 32332 1057
rect 32280 989 32332 1023
rect 32280 955 32290 989
rect 32324 955 32332 989
rect 32280 921 32332 955
rect 32280 887 32290 921
rect 32324 887 32332 921
rect 32280 869 32332 887
rect 32466 1047 32524 1062
rect 32466 1013 32478 1047
rect 32512 1013 32524 1047
rect 32466 979 32524 1013
rect 32466 945 32478 979
rect 32512 945 32524 979
rect 32466 911 32524 945
rect 32466 877 32478 911
rect 32512 877 32524 911
rect 32466 862 32524 877
rect 32554 1047 32612 1062
rect 32554 1013 32566 1047
rect 32600 1013 32612 1047
rect 32554 979 32612 1013
rect 33394 1065 33446 1077
rect 33112 1047 33170 1062
rect 33112 1013 33124 1047
rect 33158 1013 33170 1047
rect 32554 945 32566 979
rect 32600 945 32612 979
rect 32554 911 32612 945
rect 32554 877 32566 911
rect 32600 877 32612 911
rect 33112 979 33170 1013
rect 33112 945 33124 979
rect 33158 945 33170 979
rect 33112 911 33170 945
rect 32554 862 32612 877
rect 32682 887 32744 902
rect 32682 853 32694 887
rect 32728 853 32744 887
rect 30982 717 30998 751
rect 31032 717 31044 751
rect 30982 702 31044 717
rect 32682 819 32744 853
rect 32682 785 32694 819
rect 32728 785 32744 819
rect 32682 751 32744 785
rect 32682 717 32694 751
rect 32728 717 32744 751
rect 32682 702 32744 717
rect 32774 887 32840 902
rect 32774 853 32790 887
rect 32824 853 32840 887
rect 32774 819 32840 853
rect 32774 785 32790 819
rect 32824 785 32840 819
rect 32774 751 32840 785
rect 32774 717 32790 751
rect 32824 717 32840 751
rect 32774 702 32840 717
rect 32870 887 32932 902
rect 32870 853 32886 887
rect 32920 853 32932 887
rect 33112 877 33124 911
rect 33158 877 33170 911
rect 33112 862 33170 877
rect 33200 1047 33258 1062
rect 33200 1013 33212 1047
rect 33246 1013 33258 1047
rect 33200 979 33258 1013
rect 33200 945 33212 979
rect 33246 945 33258 979
rect 33200 911 33258 945
rect 33200 877 33212 911
rect 33246 877 33258 911
rect 33394 1031 33402 1065
rect 33436 1031 33446 1065
rect 33394 997 33446 1031
rect 33394 963 33402 997
rect 33436 963 33446 997
rect 33394 929 33446 963
rect 33394 895 33402 929
rect 33436 895 33446 929
rect 33394 877 33446 895
rect 33476 1065 33528 1077
rect 33476 1031 33486 1065
rect 33520 1031 33528 1065
rect 33476 997 33528 1031
rect 33476 963 33486 997
rect 33520 963 33528 997
rect 33476 929 33528 963
rect 33476 895 33486 929
rect 33520 895 33528 929
rect 33699 1055 33751 1075
rect 33699 1021 33707 1055
rect 33741 1021 33751 1055
rect 33699 987 33751 1021
rect 33699 953 33707 987
rect 33741 953 33751 987
rect 33699 917 33751 953
rect 33781 1055 33839 1075
rect 33781 1021 33793 1055
rect 33827 1021 33839 1055
rect 33781 987 33839 1021
rect 33781 953 33793 987
rect 33827 953 33839 987
rect 33781 917 33839 953
rect 33869 1055 33921 1075
rect 33869 1021 33879 1055
rect 33913 1021 33921 1055
rect 33869 974 33921 1021
rect 33869 940 33879 974
rect 33913 940 33921 974
rect 33869 917 33921 940
rect 34086 1057 34138 1069
rect 34086 1023 34094 1057
rect 34128 1023 34138 1057
rect 34086 989 34138 1023
rect 34086 955 34094 989
rect 34128 955 34138 989
rect 34086 921 34138 955
rect 33476 877 33528 895
rect 33200 862 33258 877
rect 32870 819 32932 853
rect 32870 785 32886 819
rect 32920 785 32932 819
rect 32870 751 32932 785
rect 34086 887 34094 921
rect 34128 887 34138 921
rect 34086 869 34138 887
rect 34168 1057 34220 1069
rect 34168 1023 34178 1057
rect 34212 1023 34220 1057
rect 34168 989 34220 1023
rect 34168 955 34178 989
rect 34212 955 34220 989
rect 34168 921 34220 955
rect 34168 887 34178 921
rect 34212 887 34220 921
rect 34168 869 34220 887
rect 34354 1047 34412 1062
rect 34354 1013 34366 1047
rect 34400 1013 34412 1047
rect 34354 979 34412 1013
rect 34354 945 34366 979
rect 34400 945 34412 979
rect 34354 911 34412 945
rect 34354 877 34366 911
rect 34400 877 34412 911
rect 34354 862 34412 877
rect 34442 1047 34500 1062
rect 34442 1013 34454 1047
rect 34488 1013 34500 1047
rect 34442 979 34500 1013
rect 35282 1065 35334 1077
rect 35000 1047 35058 1062
rect 35000 1013 35012 1047
rect 35046 1013 35058 1047
rect 34442 945 34454 979
rect 34488 945 34500 979
rect 34442 911 34500 945
rect 34442 877 34454 911
rect 34488 877 34500 911
rect 35000 979 35058 1013
rect 35000 945 35012 979
rect 35046 945 35058 979
rect 35000 911 35058 945
rect 34442 862 34500 877
rect 34570 887 34632 902
rect 34570 853 34582 887
rect 34616 853 34632 887
rect 32870 717 32886 751
rect 32920 717 32932 751
rect 32870 702 32932 717
rect 34570 819 34632 853
rect 34570 785 34582 819
rect 34616 785 34632 819
rect 34570 751 34632 785
rect 34570 717 34582 751
rect 34616 717 34632 751
rect 34570 702 34632 717
rect 34662 887 34728 902
rect 34662 853 34678 887
rect 34712 853 34728 887
rect 34662 819 34728 853
rect 34662 785 34678 819
rect 34712 785 34728 819
rect 34662 751 34728 785
rect 34662 717 34678 751
rect 34712 717 34728 751
rect 34662 702 34728 717
rect 34758 887 34820 902
rect 34758 853 34774 887
rect 34808 853 34820 887
rect 35000 877 35012 911
rect 35046 877 35058 911
rect 35000 862 35058 877
rect 35088 1047 35146 1062
rect 35088 1013 35100 1047
rect 35134 1013 35146 1047
rect 35088 979 35146 1013
rect 35088 945 35100 979
rect 35134 945 35146 979
rect 35088 911 35146 945
rect 35088 877 35100 911
rect 35134 877 35146 911
rect 35282 1031 35290 1065
rect 35324 1031 35334 1065
rect 35282 997 35334 1031
rect 35282 963 35290 997
rect 35324 963 35334 997
rect 35282 929 35334 963
rect 35282 895 35290 929
rect 35324 895 35334 929
rect 35282 877 35334 895
rect 35364 1065 35416 1077
rect 35364 1031 35374 1065
rect 35408 1031 35416 1065
rect 35364 997 35416 1031
rect 35364 963 35374 997
rect 35408 963 35416 997
rect 35364 929 35416 963
rect 35364 895 35374 929
rect 35408 895 35416 929
rect 35587 1055 35639 1075
rect 35587 1021 35595 1055
rect 35629 1021 35639 1055
rect 35587 987 35639 1021
rect 35587 953 35595 987
rect 35629 953 35639 987
rect 35587 917 35639 953
rect 35669 1055 35727 1075
rect 35669 1021 35681 1055
rect 35715 1021 35727 1055
rect 35669 987 35727 1021
rect 35669 953 35681 987
rect 35715 953 35727 987
rect 35669 917 35727 953
rect 35757 1055 35809 1075
rect 35757 1021 35767 1055
rect 35801 1021 35809 1055
rect 35757 974 35809 1021
rect 35757 940 35767 974
rect 35801 940 35809 974
rect 35757 917 35809 940
rect 35974 1057 36026 1069
rect 35974 1023 35982 1057
rect 36016 1023 36026 1057
rect 35974 989 36026 1023
rect 35974 955 35982 989
rect 36016 955 36026 989
rect 35974 921 36026 955
rect 35364 877 35416 895
rect 35088 862 35146 877
rect 34758 819 34820 853
rect 34758 785 34774 819
rect 34808 785 34820 819
rect 34758 751 34820 785
rect 35974 887 35982 921
rect 36016 887 36026 921
rect 35974 869 36026 887
rect 36056 1057 36108 1069
rect 36056 1023 36066 1057
rect 36100 1023 36108 1057
rect 36056 989 36108 1023
rect 36056 955 36066 989
rect 36100 955 36108 989
rect 36056 921 36108 955
rect 36056 887 36066 921
rect 36100 887 36108 921
rect 36056 869 36108 887
rect 36242 1047 36300 1062
rect 36242 1013 36254 1047
rect 36288 1013 36300 1047
rect 36242 979 36300 1013
rect 36242 945 36254 979
rect 36288 945 36300 979
rect 36242 911 36300 945
rect 36242 877 36254 911
rect 36288 877 36300 911
rect 36242 862 36300 877
rect 36330 1047 36388 1062
rect 36330 1013 36342 1047
rect 36376 1013 36388 1047
rect 36330 979 36388 1013
rect 37170 1065 37222 1077
rect 36888 1047 36946 1062
rect 36888 1013 36900 1047
rect 36934 1013 36946 1047
rect 36330 945 36342 979
rect 36376 945 36388 979
rect 36330 911 36388 945
rect 36330 877 36342 911
rect 36376 877 36388 911
rect 36888 979 36946 1013
rect 36888 945 36900 979
rect 36934 945 36946 979
rect 36888 911 36946 945
rect 36330 862 36388 877
rect 36458 887 36520 902
rect 36458 853 36470 887
rect 36504 853 36520 887
rect 34758 717 34774 751
rect 34808 717 34820 751
rect 34758 702 34820 717
rect 36458 819 36520 853
rect 36458 785 36470 819
rect 36504 785 36520 819
rect 36458 751 36520 785
rect 36458 717 36470 751
rect 36504 717 36520 751
rect 36458 702 36520 717
rect 36550 887 36616 902
rect 36550 853 36566 887
rect 36600 853 36616 887
rect 36550 819 36616 853
rect 36550 785 36566 819
rect 36600 785 36616 819
rect 36550 751 36616 785
rect 36550 717 36566 751
rect 36600 717 36616 751
rect 36550 702 36616 717
rect 36646 887 36708 902
rect 36646 853 36662 887
rect 36696 853 36708 887
rect 36888 877 36900 911
rect 36934 877 36946 911
rect 36888 862 36946 877
rect 36976 1047 37034 1062
rect 36976 1013 36988 1047
rect 37022 1013 37034 1047
rect 36976 979 37034 1013
rect 36976 945 36988 979
rect 37022 945 37034 979
rect 36976 911 37034 945
rect 36976 877 36988 911
rect 37022 877 37034 911
rect 37170 1031 37178 1065
rect 37212 1031 37222 1065
rect 37170 997 37222 1031
rect 37170 963 37178 997
rect 37212 963 37222 997
rect 37170 929 37222 963
rect 37170 895 37178 929
rect 37212 895 37222 929
rect 37170 877 37222 895
rect 37252 1065 37304 1077
rect 37252 1031 37262 1065
rect 37296 1031 37304 1065
rect 37252 997 37304 1031
rect 37252 963 37262 997
rect 37296 963 37304 997
rect 37252 929 37304 963
rect 37252 895 37262 929
rect 37296 895 37304 929
rect 37475 1055 37527 1075
rect 37475 1021 37483 1055
rect 37517 1021 37527 1055
rect 37475 987 37527 1021
rect 37475 953 37483 987
rect 37517 953 37527 987
rect 37475 917 37527 953
rect 37557 1055 37615 1075
rect 37557 1021 37569 1055
rect 37603 1021 37615 1055
rect 37557 987 37615 1021
rect 37557 953 37569 987
rect 37603 953 37615 987
rect 37557 917 37615 953
rect 37645 1055 37697 1075
rect 37645 1021 37655 1055
rect 37689 1021 37697 1055
rect 37645 974 37697 1021
rect 37645 940 37655 974
rect 37689 940 37697 974
rect 37645 917 37697 940
rect 37862 1057 37914 1069
rect 37862 1023 37870 1057
rect 37904 1023 37914 1057
rect 37862 989 37914 1023
rect 37862 955 37870 989
rect 37904 955 37914 989
rect 37862 921 37914 955
rect 37252 877 37304 895
rect 36976 862 37034 877
rect 36646 819 36708 853
rect 36646 785 36662 819
rect 36696 785 36708 819
rect 36646 751 36708 785
rect 37862 887 37870 921
rect 37904 887 37914 921
rect 37862 869 37914 887
rect 37944 1057 37996 1069
rect 37944 1023 37954 1057
rect 37988 1023 37996 1057
rect 37944 989 37996 1023
rect 37944 955 37954 989
rect 37988 955 37996 989
rect 37944 921 37996 955
rect 37944 887 37954 921
rect 37988 887 37996 921
rect 37944 869 37996 887
rect 38130 1047 38188 1062
rect 38130 1013 38142 1047
rect 38176 1013 38188 1047
rect 38130 979 38188 1013
rect 38130 945 38142 979
rect 38176 945 38188 979
rect 38130 911 38188 945
rect 38130 877 38142 911
rect 38176 877 38188 911
rect 38130 862 38188 877
rect 38218 1047 38276 1062
rect 38218 1013 38230 1047
rect 38264 1013 38276 1047
rect 38218 979 38276 1013
rect 39058 1065 39110 1077
rect 38776 1047 38834 1062
rect 38776 1013 38788 1047
rect 38822 1013 38834 1047
rect 38218 945 38230 979
rect 38264 945 38276 979
rect 38218 911 38276 945
rect 38218 877 38230 911
rect 38264 877 38276 911
rect 38776 979 38834 1013
rect 38776 945 38788 979
rect 38822 945 38834 979
rect 38776 911 38834 945
rect 38218 862 38276 877
rect 38346 887 38408 902
rect 38346 853 38358 887
rect 38392 853 38408 887
rect 36646 717 36662 751
rect 36696 717 36708 751
rect 36646 702 36708 717
rect 38346 819 38408 853
rect 38346 785 38358 819
rect 38392 785 38408 819
rect 38346 751 38408 785
rect 38346 717 38358 751
rect 38392 717 38408 751
rect 38346 702 38408 717
rect 38438 887 38504 902
rect 38438 853 38454 887
rect 38488 853 38504 887
rect 38438 819 38504 853
rect 38438 785 38454 819
rect 38488 785 38504 819
rect 38438 751 38504 785
rect 38438 717 38454 751
rect 38488 717 38504 751
rect 38438 702 38504 717
rect 38534 887 38596 902
rect 38534 853 38550 887
rect 38584 853 38596 887
rect 38776 877 38788 911
rect 38822 877 38834 911
rect 38776 862 38834 877
rect 38864 1047 38922 1062
rect 38864 1013 38876 1047
rect 38910 1013 38922 1047
rect 38864 979 38922 1013
rect 38864 945 38876 979
rect 38910 945 38922 979
rect 38864 911 38922 945
rect 38864 877 38876 911
rect 38910 877 38922 911
rect 39058 1031 39066 1065
rect 39100 1031 39110 1065
rect 39058 997 39110 1031
rect 39058 963 39066 997
rect 39100 963 39110 997
rect 39058 929 39110 963
rect 39058 895 39066 929
rect 39100 895 39110 929
rect 39058 877 39110 895
rect 39140 1065 39192 1077
rect 39140 1031 39150 1065
rect 39184 1031 39192 1065
rect 39140 997 39192 1031
rect 39140 963 39150 997
rect 39184 963 39192 997
rect 39140 929 39192 963
rect 39140 895 39150 929
rect 39184 895 39192 929
rect 39363 1055 39415 1075
rect 39363 1021 39371 1055
rect 39405 1021 39415 1055
rect 39363 987 39415 1021
rect 39363 953 39371 987
rect 39405 953 39415 987
rect 39363 917 39415 953
rect 39445 1055 39503 1075
rect 39445 1021 39457 1055
rect 39491 1021 39503 1055
rect 39445 987 39503 1021
rect 39445 953 39457 987
rect 39491 953 39503 987
rect 39445 917 39503 953
rect 39533 1055 39585 1075
rect 39533 1021 39543 1055
rect 39577 1021 39585 1055
rect 39533 974 39585 1021
rect 39533 940 39543 974
rect 39577 940 39585 974
rect 39533 917 39585 940
rect 39750 1057 39802 1069
rect 39750 1023 39758 1057
rect 39792 1023 39802 1057
rect 39750 989 39802 1023
rect 39750 955 39758 989
rect 39792 955 39802 989
rect 39750 921 39802 955
rect 39140 877 39192 895
rect 38864 862 38922 877
rect 38534 819 38596 853
rect 38534 785 38550 819
rect 38584 785 38596 819
rect 38534 751 38596 785
rect 39750 887 39758 921
rect 39792 887 39802 921
rect 39750 869 39802 887
rect 39832 1057 39884 1069
rect 39832 1023 39842 1057
rect 39876 1023 39884 1057
rect 39832 989 39884 1023
rect 39832 955 39842 989
rect 39876 955 39884 989
rect 39832 921 39884 955
rect 39832 887 39842 921
rect 39876 887 39884 921
rect 39832 869 39884 887
rect 40018 1047 40076 1062
rect 40018 1013 40030 1047
rect 40064 1013 40076 1047
rect 40018 979 40076 1013
rect 40018 945 40030 979
rect 40064 945 40076 979
rect 40018 911 40076 945
rect 40018 877 40030 911
rect 40064 877 40076 911
rect 40018 862 40076 877
rect 40106 1047 40164 1062
rect 40106 1013 40118 1047
rect 40152 1013 40164 1047
rect 40106 979 40164 1013
rect 40946 1065 40998 1077
rect 40664 1047 40722 1062
rect 40664 1013 40676 1047
rect 40710 1013 40722 1047
rect 40106 945 40118 979
rect 40152 945 40164 979
rect 40106 911 40164 945
rect 40106 877 40118 911
rect 40152 877 40164 911
rect 40664 979 40722 1013
rect 40664 945 40676 979
rect 40710 945 40722 979
rect 40664 911 40722 945
rect 40106 862 40164 877
rect 40234 887 40296 902
rect 40234 853 40246 887
rect 40280 853 40296 887
rect 38534 717 38550 751
rect 38584 717 38596 751
rect 38534 702 38596 717
rect 40234 819 40296 853
rect 40234 785 40246 819
rect 40280 785 40296 819
rect 40234 751 40296 785
rect 40234 717 40246 751
rect 40280 717 40296 751
rect 40234 702 40296 717
rect 40326 887 40392 902
rect 40326 853 40342 887
rect 40376 853 40392 887
rect 40326 819 40392 853
rect 40326 785 40342 819
rect 40376 785 40392 819
rect 40326 751 40392 785
rect 40326 717 40342 751
rect 40376 717 40392 751
rect 40326 702 40392 717
rect 40422 887 40484 902
rect 40422 853 40438 887
rect 40472 853 40484 887
rect 40664 877 40676 911
rect 40710 877 40722 911
rect 40664 862 40722 877
rect 40752 1047 40810 1062
rect 40752 1013 40764 1047
rect 40798 1013 40810 1047
rect 40752 979 40810 1013
rect 40752 945 40764 979
rect 40798 945 40810 979
rect 40752 911 40810 945
rect 40752 877 40764 911
rect 40798 877 40810 911
rect 40946 1031 40954 1065
rect 40988 1031 40998 1065
rect 40946 997 40998 1031
rect 40946 963 40954 997
rect 40988 963 40998 997
rect 40946 929 40998 963
rect 40946 895 40954 929
rect 40988 895 40998 929
rect 40946 877 40998 895
rect 41028 1065 41080 1077
rect 41028 1031 41038 1065
rect 41072 1031 41080 1065
rect 41028 997 41080 1031
rect 41028 963 41038 997
rect 41072 963 41080 997
rect 41028 929 41080 963
rect 41028 895 41038 929
rect 41072 895 41080 929
rect 41251 1055 41303 1075
rect 41251 1021 41259 1055
rect 41293 1021 41303 1055
rect 41251 987 41303 1021
rect 41251 953 41259 987
rect 41293 953 41303 987
rect 41251 917 41303 953
rect 41333 1055 41391 1075
rect 41333 1021 41345 1055
rect 41379 1021 41391 1055
rect 41333 987 41391 1021
rect 41333 953 41345 987
rect 41379 953 41391 987
rect 41333 917 41391 953
rect 41421 1055 41473 1075
rect 41421 1021 41431 1055
rect 41465 1021 41473 1055
rect 41421 974 41473 1021
rect 41421 940 41431 974
rect 41465 940 41473 974
rect 41421 917 41473 940
rect 41638 1057 41690 1069
rect 41638 1023 41646 1057
rect 41680 1023 41690 1057
rect 41638 989 41690 1023
rect 41638 955 41646 989
rect 41680 955 41690 989
rect 41638 921 41690 955
rect 41028 877 41080 895
rect 40752 862 40810 877
rect 40422 819 40484 853
rect 40422 785 40438 819
rect 40472 785 40484 819
rect 40422 751 40484 785
rect 41638 887 41646 921
rect 41680 887 41690 921
rect 41638 869 41690 887
rect 41720 1057 41772 1069
rect 41720 1023 41730 1057
rect 41764 1023 41772 1057
rect 41720 989 41772 1023
rect 41720 955 41730 989
rect 41764 955 41772 989
rect 41720 921 41772 955
rect 41720 887 41730 921
rect 41764 887 41772 921
rect 41720 869 41772 887
rect 41906 1047 41964 1062
rect 41906 1013 41918 1047
rect 41952 1013 41964 1047
rect 41906 979 41964 1013
rect 41906 945 41918 979
rect 41952 945 41964 979
rect 41906 911 41964 945
rect 41906 877 41918 911
rect 41952 877 41964 911
rect 41906 862 41964 877
rect 41994 1047 42052 1062
rect 41994 1013 42006 1047
rect 42040 1013 42052 1047
rect 41994 979 42052 1013
rect 42834 1065 42886 1077
rect 42552 1047 42610 1062
rect 42552 1013 42564 1047
rect 42598 1013 42610 1047
rect 41994 945 42006 979
rect 42040 945 42052 979
rect 41994 911 42052 945
rect 41994 877 42006 911
rect 42040 877 42052 911
rect 42552 979 42610 1013
rect 42552 945 42564 979
rect 42598 945 42610 979
rect 42552 911 42610 945
rect 41994 862 42052 877
rect 42122 887 42184 902
rect 42122 853 42134 887
rect 42168 853 42184 887
rect 40422 717 40438 751
rect 40472 717 40484 751
rect 40422 702 40484 717
rect 42122 819 42184 853
rect 42122 785 42134 819
rect 42168 785 42184 819
rect 42122 751 42184 785
rect 42122 717 42134 751
rect 42168 717 42184 751
rect 42122 702 42184 717
rect 42214 887 42280 902
rect 42214 853 42230 887
rect 42264 853 42280 887
rect 42214 819 42280 853
rect 42214 785 42230 819
rect 42264 785 42280 819
rect 42214 751 42280 785
rect 42214 717 42230 751
rect 42264 717 42280 751
rect 42214 702 42280 717
rect 42310 887 42372 902
rect 42310 853 42326 887
rect 42360 853 42372 887
rect 42552 877 42564 911
rect 42598 877 42610 911
rect 42552 862 42610 877
rect 42640 1047 42698 1062
rect 42640 1013 42652 1047
rect 42686 1013 42698 1047
rect 42640 979 42698 1013
rect 42640 945 42652 979
rect 42686 945 42698 979
rect 42640 911 42698 945
rect 42640 877 42652 911
rect 42686 877 42698 911
rect 42834 1031 42842 1065
rect 42876 1031 42886 1065
rect 42834 997 42886 1031
rect 42834 963 42842 997
rect 42876 963 42886 997
rect 42834 929 42886 963
rect 42834 895 42842 929
rect 42876 895 42886 929
rect 42834 877 42886 895
rect 42916 1065 42968 1077
rect 42916 1031 42926 1065
rect 42960 1031 42968 1065
rect 42916 997 42968 1031
rect 42916 963 42926 997
rect 42960 963 42968 997
rect 42916 929 42968 963
rect 42916 895 42926 929
rect 42960 895 42968 929
rect 43139 1055 43191 1075
rect 43139 1021 43147 1055
rect 43181 1021 43191 1055
rect 43139 987 43191 1021
rect 43139 953 43147 987
rect 43181 953 43191 987
rect 43139 917 43191 953
rect 43221 1055 43279 1075
rect 43221 1021 43233 1055
rect 43267 1021 43279 1055
rect 43221 987 43279 1021
rect 43221 953 43233 987
rect 43267 953 43279 987
rect 43221 917 43279 953
rect 43309 1055 43361 1075
rect 43309 1021 43319 1055
rect 43353 1021 43361 1055
rect 43309 974 43361 1021
rect 43309 940 43319 974
rect 43353 940 43361 974
rect 43309 917 43361 940
rect 43526 1057 43578 1069
rect 43526 1023 43534 1057
rect 43568 1023 43578 1057
rect 43526 989 43578 1023
rect 43526 955 43534 989
rect 43568 955 43578 989
rect 43526 921 43578 955
rect 42916 877 42968 895
rect 42640 862 42698 877
rect 42310 819 42372 853
rect 42310 785 42326 819
rect 42360 785 42372 819
rect 42310 751 42372 785
rect 43526 887 43534 921
rect 43568 887 43578 921
rect 43526 869 43578 887
rect 43608 1057 43660 1069
rect 43608 1023 43618 1057
rect 43652 1023 43660 1057
rect 43608 989 43660 1023
rect 43608 955 43618 989
rect 43652 955 43660 989
rect 43608 921 43660 955
rect 43608 887 43618 921
rect 43652 887 43660 921
rect 43608 869 43660 887
rect 43794 1047 43852 1062
rect 43794 1013 43806 1047
rect 43840 1013 43852 1047
rect 43794 979 43852 1013
rect 43794 945 43806 979
rect 43840 945 43852 979
rect 43794 911 43852 945
rect 43794 877 43806 911
rect 43840 877 43852 911
rect 43794 862 43852 877
rect 43882 1047 43940 1062
rect 43882 1013 43894 1047
rect 43928 1013 43940 1047
rect 43882 979 43940 1013
rect 44722 1065 44774 1077
rect 44440 1047 44498 1062
rect 44440 1013 44452 1047
rect 44486 1013 44498 1047
rect 43882 945 43894 979
rect 43928 945 43940 979
rect 43882 911 43940 945
rect 43882 877 43894 911
rect 43928 877 43940 911
rect 44440 979 44498 1013
rect 44440 945 44452 979
rect 44486 945 44498 979
rect 44440 911 44498 945
rect 43882 862 43940 877
rect 44010 887 44072 902
rect 44010 853 44022 887
rect 44056 853 44072 887
rect 42310 717 42326 751
rect 42360 717 42372 751
rect 42310 702 42372 717
rect 44010 819 44072 853
rect 44010 785 44022 819
rect 44056 785 44072 819
rect 44010 751 44072 785
rect 44010 717 44022 751
rect 44056 717 44072 751
rect 44010 702 44072 717
rect 44102 887 44168 902
rect 44102 853 44118 887
rect 44152 853 44168 887
rect 44102 819 44168 853
rect 44102 785 44118 819
rect 44152 785 44168 819
rect 44102 751 44168 785
rect 44102 717 44118 751
rect 44152 717 44168 751
rect 44102 702 44168 717
rect 44198 887 44260 902
rect 44198 853 44214 887
rect 44248 853 44260 887
rect 44440 877 44452 911
rect 44486 877 44498 911
rect 44440 862 44498 877
rect 44528 1047 44586 1062
rect 44528 1013 44540 1047
rect 44574 1013 44586 1047
rect 44528 979 44586 1013
rect 44528 945 44540 979
rect 44574 945 44586 979
rect 44528 911 44586 945
rect 44528 877 44540 911
rect 44574 877 44586 911
rect 44722 1031 44730 1065
rect 44764 1031 44774 1065
rect 44722 997 44774 1031
rect 44722 963 44730 997
rect 44764 963 44774 997
rect 44722 929 44774 963
rect 44722 895 44730 929
rect 44764 895 44774 929
rect 44722 877 44774 895
rect 44804 1065 44856 1077
rect 44804 1031 44814 1065
rect 44848 1031 44856 1065
rect 44804 997 44856 1031
rect 44804 963 44814 997
rect 44848 963 44856 997
rect 44804 929 44856 963
rect 44804 895 44814 929
rect 44848 895 44856 929
rect 45027 1055 45079 1075
rect 45027 1021 45035 1055
rect 45069 1021 45079 1055
rect 45027 987 45079 1021
rect 45027 953 45035 987
rect 45069 953 45079 987
rect 45027 917 45079 953
rect 45109 1055 45167 1075
rect 45109 1021 45121 1055
rect 45155 1021 45167 1055
rect 45109 987 45167 1021
rect 45109 953 45121 987
rect 45155 953 45167 987
rect 45109 917 45167 953
rect 45197 1055 45249 1075
rect 45197 1021 45207 1055
rect 45241 1021 45249 1055
rect 45197 974 45249 1021
rect 45197 940 45207 974
rect 45241 940 45249 974
rect 45197 917 45249 940
rect 45408 1057 45460 1069
rect 45408 1023 45416 1057
rect 45450 1023 45460 1057
rect 45408 989 45460 1023
rect 45408 955 45416 989
rect 45450 955 45460 989
rect 45408 921 45460 955
rect 44804 877 44856 895
rect 44528 862 44586 877
rect 44198 819 44260 853
rect 44198 785 44214 819
rect 44248 785 44260 819
rect 44198 751 44260 785
rect 45408 887 45416 921
rect 45450 887 45460 921
rect 45408 869 45460 887
rect 45490 1057 45542 1069
rect 45490 1023 45500 1057
rect 45534 1023 45542 1057
rect 45490 989 45542 1023
rect 45490 955 45500 989
rect 45534 955 45542 989
rect 45490 921 45542 955
rect 45490 887 45500 921
rect 45534 887 45542 921
rect 45490 869 45542 887
rect 45676 1047 45734 1062
rect 45676 1013 45688 1047
rect 45722 1013 45734 1047
rect 45676 979 45734 1013
rect 45676 945 45688 979
rect 45722 945 45734 979
rect 45676 911 45734 945
rect 45676 877 45688 911
rect 45722 877 45734 911
rect 45676 862 45734 877
rect 45764 1047 45822 1062
rect 45764 1013 45776 1047
rect 45810 1013 45822 1047
rect 45764 979 45822 1013
rect 46604 1065 46656 1077
rect 46322 1047 46380 1062
rect 46322 1013 46334 1047
rect 46368 1013 46380 1047
rect 45764 945 45776 979
rect 45810 945 45822 979
rect 45764 911 45822 945
rect 45764 877 45776 911
rect 45810 877 45822 911
rect 46322 979 46380 1013
rect 46322 945 46334 979
rect 46368 945 46380 979
rect 46322 911 46380 945
rect 45764 862 45822 877
rect 45892 887 45954 902
rect 45892 853 45904 887
rect 45938 853 45954 887
rect 44198 717 44214 751
rect 44248 717 44260 751
rect 44198 702 44260 717
rect 45892 819 45954 853
rect 45892 785 45904 819
rect 45938 785 45954 819
rect 45892 751 45954 785
rect 45892 717 45904 751
rect 45938 717 45954 751
rect 45892 702 45954 717
rect 45984 887 46050 902
rect 45984 853 46000 887
rect 46034 853 46050 887
rect 45984 819 46050 853
rect 45984 785 46000 819
rect 46034 785 46050 819
rect 45984 751 46050 785
rect 45984 717 46000 751
rect 46034 717 46050 751
rect 45984 702 46050 717
rect 46080 887 46142 902
rect 46080 853 46096 887
rect 46130 853 46142 887
rect 46322 877 46334 911
rect 46368 877 46380 911
rect 46322 862 46380 877
rect 46410 1047 46468 1062
rect 46410 1013 46422 1047
rect 46456 1013 46468 1047
rect 46410 979 46468 1013
rect 46410 945 46422 979
rect 46456 945 46468 979
rect 46410 911 46468 945
rect 46410 877 46422 911
rect 46456 877 46468 911
rect 46604 1031 46612 1065
rect 46646 1031 46656 1065
rect 46604 997 46656 1031
rect 46604 963 46612 997
rect 46646 963 46656 997
rect 46604 929 46656 963
rect 46604 895 46612 929
rect 46646 895 46656 929
rect 46604 877 46656 895
rect 46686 1065 46738 1077
rect 46686 1031 46696 1065
rect 46730 1031 46738 1065
rect 46686 997 46738 1031
rect 46686 963 46696 997
rect 46730 963 46738 997
rect 46686 929 46738 963
rect 46686 895 46696 929
rect 46730 895 46738 929
rect 46909 1055 46961 1075
rect 46909 1021 46917 1055
rect 46951 1021 46961 1055
rect 46909 987 46961 1021
rect 46909 953 46917 987
rect 46951 953 46961 987
rect 46909 917 46961 953
rect 46991 1055 47049 1075
rect 46991 1021 47003 1055
rect 47037 1021 47049 1055
rect 46991 987 47049 1021
rect 46991 953 47003 987
rect 47037 953 47049 987
rect 46991 917 47049 953
rect 47079 1055 47131 1075
rect 47079 1021 47089 1055
rect 47123 1021 47131 1055
rect 47079 974 47131 1021
rect 47079 940 47089 974
rect 47123 940 47131 974
rect 47079 917 47131 940
rect 47296 1057 47348 1069
rect 47296 1023 47304 1057
rect 47338 1023 47348 1057
rect 47296 989 47348 1023
rect 47296 955 47304 989
rect 47338 955 47348 989
rect 47296 921 47348 955
rect 46686 877 46738 895
rect 46410 862 46468 877
rect 46080 819 46142 853
rect 46080 785 46096 819
rect 46130 785 46142 819
rect 46080 751 46142 785
rect 47296 887 47304 921
rect 47338 887 47348 921
rect 47296 869 47348 887
rect 47378 1057 47430 1069
rect 47378 1023 47388 1057
rect 47422 1023 47430 1057
rect 47378 989 47430 1023
rect 47378 955 47388 989
rect 47422 955 47430 989
rect 47378 921 47430 955
rect 47378 887 47388 921
rect 47422 887 47430 921
rect 47378 869 47430 887
rect 47564 1047 47622 1062
rect 47564 1013 47576 1047
rect 47610 1013 47622 1047
rect 47564 979 47622 1013
rect 47564 945 47576 979
rect 47610 945 47622 979
rect 47564 911 47622 945
rect 47564 877 47576 911
rect 47610 877 47622 911
rect 47564 862 47622 877
rect 47652 1047 47710 1062
rect 47652 1013 47664 1047
rect 47698 1013 47710 1047
rect 47652 979 47710 1013
rect 48492 1065 48544 1077
rect 48210 1047 48268 1062
rect 48210 1013 48222 1047
rect 48256 1013 48268 1047
rect 47652 945 47664 979
rect 47698 945 47710 979
rect 47652 911 47710 945
rect 47652 877 47664 911
rect 47698 877 47710 911
rect 48210 979 48268 1013
rect 48210 945 48222 979
rect 48256 945 48268 979
rect 48210 911 48268 945
rect 47652 862 47710 877
rect 47780 887 47842 902
rect 47780 853 47792 887
rect 47826 853 47842 887
rect 46080 717 46096 751
rect 46130 717 46142 751
rect 46080 702 46142 717
rect 47780 819 47842 853
rect 47780 785 47792 819
rect 47826 785 47842 819
rect 47780 751 47842 785
rect 47780 717 47792 751
rect 47826 717 47842 751
rect 47780 702 47842 717
rect 47872 887 47938 902
rect 47872 853 47888 887
rect 47922 853 47938 887
rect 47872 819 47938 853
rect 47872 785 47888 819
rect 47922 785 47938 819
rect 47872 751 47938 785
rect 47872 717 47888 751
rect 47922 717 47938 751
rect 47872 702 47938 717
rect 47968 887 48030 902
rect 47968 853 47984 887
rect 48018 853 48030 887
rect 48210 877 48222 911
rect 48256 877 48268 911
rect 48210 862 48268 877
rect 48298 1047 48356 1062
rect 48298 1013 48310 1047
rect 48344 1013 48356 1047
rect 48298 979 48356 1013
rect 48298 945 48310 979
rect 48344 945 48356 979
rect 48298 911 48356 945
rect 48298 877 48310 911
rect 48344 877 48356 911
rect 48492 1031 48500 1065
rect 48534 1031 48544 1065
rect 48492 997 48544 1031
rect 48492 963 48500 997
rect 48534 963 48544 997
rect 48492 929 48544 963
rect 48492 895 48500 929
rect 48534 895 48544 929
rect 48492 877 48544 895
rect 48574 1065 48626 1077
rect 48574 1031 48584 1065
rect 48618 1031 48626 1065
rect 48574 997 48626 1031
rect 48574 963 48584 997
rect 48618 963 48626 997
rect 48574 929 48626 963
rect 48574 895 48584 929
rect 48618 895 48626 929
rect 48797 1055 48849 1075
rect 48797 1021 48805 1055
rect 48839 1021 48849 1055
rect 48797 987 48849 1021
rect 48797 953 48805 987
rect 48839 953 48849 987
rect 48797 917 48849 953
rect 48879 1055 48937 1075
rect 48879 1021 48891 1055
rect 48925 1021 48937 1055
rect 48879 987 48937 1021
rect 48879 953 48891 987
rect 48925 953 48937 987
rect 48879 917 48937 953
rect 48967 1055 49019 1075
rect 48967 1021 48977 1055
rect 49011 1021 49019 1055
rect 48967 974 49019 1021
rect 48967 940 48977 974
rect 49011 940 49019 974
rect 48967 917 49019 940
rect 49184 1057 49236 1069
rect 49184 1023 49192 1057
rect 49226 1023 49236 1057
rect 49184 989 49236 1023
rect 49184 955 49192 989
rect 49226 955 49236 989
rect 49184 921 49236 955
rect 48574 877 48626 895
rect 48298 862 48356 877
rect 47968 819 48030 853
rect 47968 785 47984 819
rect 48018 785 48030 819
rect 47968 751 48030 785
rect 49184 887 49192 921
rect 49226 887 49236 921
rect 49184 869 49236 887
rect 49266 1057 49318 1069
rect 49266 1023 49276 1057
rect 49310 1023 49318 1057
rect 49266 989 49318 1023
rect 49266 955 49276 989
rect 49310 955 49318 989
rect 49266 921 49318 955
rect 49266 887 49276 921
rect 49310 887 49318 921
rect 49266 869 49318 887
rect 49452 1047 49510 1062
rect 49452 1013 49464 1047
rect 49498 1013 49510 1047
rect 49452 979 49510 1013
rect 49452 945 49464 979
rect 49498 945 49510 979
rect 49452 911 49510 945
rect 49452 877 49464 911
rect 49498 877 49510 911
rect 49452 862 49510 877
rect 49540 1047 49598 1062
rect 49540 1013 49552 1047
rect 49586 1013 49598 1047
rect 49540 979 49598 1013
rect 50380 1065 50432 1077
rect 50098 1047 50156 1062
rect 50098 1013 50110 1047
rect 50144 1013 50156 1047
rect 49540 945 49552 979
rect 49586 945 49598 979
rect 49540 911 49598 945
rect 49540 877 49552 911
rect 49586 877 49598 911
rect 50098 979 50156 1013
rect 50098 945 50110 979
rect 50144 945 50156 979
rect 50098 911 50156 945
rect 49540 862 49598 877
rect 49668 887 49730 902
rect 49668 853 49680 887
rect 49714 853 49730 887
rect 47968 717 47984 751
rect 48018 717 48030 751
rect 47968 702 48030 717
rect 49668 819 49730 853
rect 49668 785 49680 819
rect 49714 785 49730 819
rect 49668 751 49730 785
rect 49668 717 49680 751
rect 49714 717 49730 751
rect 49668 702 49730 717
rect 49760 887 49826 902
rect 49760 853 49776 887
rect 49810 853 49826 887
rect 49760 819 49826 853
rect 49760 785 49776 819
rect 49810 785 49826 819
rect 49760 751 49826 785
rect 49760 717 49776 751
rect 49810 717 49826 751
rect 49760 702 49826 717
rect 49856 887 49918 902
rect 49856 853 49872 887
rect 49906 853 49918 887
rect 50098 877 50110 911
rect 50144 877 50156 911
rect 50098 862 50156 877
rect 50186 1047 50244 1062
rect 50186 1013 50198 1047
rect 50232 1013 50244 1047
rect 50186 979 50244 1013
rect 50186 945 50198 979
rect 50232 945 50244 979
rect 50186 911 50244 945
rect 50186 877 50198 911
rect 50232 877 50244 911
rect 50380 1031 50388 1065
rect 50422 1031 50432 1065
rect 50380 997 50432 1031
rect 50380 963 50388 997
rect 50422 963 50432 997
rect 50380 929 50432 963
rect 50380 895 50388 929
rect 50422 895 50432 929
rect 50380 877 50432 895
rect 50462 1065 50514 1077
rect 50462 1031 50472 1065
rect 50506 1031 50514 1065
rect 50462 997 50514 1031
rect 50462 963 50472 997
rect 50506 963 50514 997
rect 50462 929 50514 963
rect 50462 895 50472 929
rect 50506 895 50514 929
rect 50685 1055 50737 1075
rect 50685 1021 50693 1055
rect 50727 1021 50737 1055
rect 50685 987 50737 1021
rect 50685 953 50693 987
rect 50727 953 50737 987
rect 50685 917 50737 953
rect 50767 1055 50825 1075
rect 50767 1021 50779 1055
rect 50813 1021 50825 1055
rect 50767 987 50825 1021
rect 50767 953 50779 987
rect 50813 953 50825 987
rect 50767 917 50825 953
rect 50855 1055 50907 1075
rect 50855 1021 50865 1055
rect 50899 1021 50907 1055
rect 50855 974 50907 1021
rect 50855 940 50865 974
rect 50899 940 50907 974
rect 50855 917 50907 940
rect 51072 1057 51124 1069
rect 51072 1023 51080 1057
rect 51114 1023 51124 1057
rect 51072 989 51124 1023
rect 51072 955 51080 989
rect 51114 955 51124 989
rect 51072 921 51124 955
rect 50462 877 50514 895
rect 50186 862 50244 877
rect 49856 819 49918 853
rect 49856 785 49872 819
rect 49906 785 49918 819
rect 49856 751 49918 785
rect 51072 887 51080 921
rect 51114 887 51124 921
rect 51072 869 51124 887
rect 51154 1057 51206 1069
rect 51154 1023 51164 1057
rect 51198 1023 51206 1057
rect 51154 989 51206 1023
rect 51154 955 51164 989
rect 51198 955 51206 989
rect 51154 921 51206 955
rect 51154 887 51164 921
rect 51198 887 51206 921
rect 51154 869 51206 887
rect 51340 1047 51398 1062
rect 51340 1013 51352 1047
rect 51386 1013 51398 1047
rect 51340 979 51398 1013
rect 51340 945 51352 979
rect 51386 945 51398 979
rect 51340 911 51398 945
rect 51340 877 51352 911
rect 51386 877 51398 911
rect 51340 862 51398 877
rect 51428 1047 51486 1062
rect 51428 1013 51440 1047
rect 51474 1013 51486 1047
rect 51428 979 51486 1013
rect 52268 1065 52320 1077
rect 51986 1047 52044 1062
rect 51986 1013 51998 1047
rect 52032 1013 52044 1047
rect 51428 945 51440 979
rect 51474 945 51486 979
rect 51428 911 51486 945
rect 51428 877 51440 911
rect 51474 877 51486 911
rect 51986 979 52044 1013
rect 51986 945 51998 979
rect 52032 945 52044 979
rect 51986 911 52044 945
rect 51428 862 51486 877
rect 51556 887 51618 902
rect 51556 853 51568 887
rect 51602 853 51618 887
rect 49856 717 49872 751
rect 49906 717 49918 751
rect 49856 702 49918 717
rect 51556 819 51618 853
rect 51556 785 51568 819
rect 51602 785 51618 819
rect 51556 751 51618 785
rect 51556 717 51568 751
rect 51602 717 51618 751
rect 51556 702 51618 717
rect 51648 887 51714 902
rect 51648 853 51664 887
rect 51698 853 51714 887
rect 51648 819 51714 853
rect 51648 785 51664 819
rect 51698 785 51714 819
rect 51648 751 51714 785
rect 51648 717 51664 751
rect 51698 717 51714 751
rect 51648 702 51714 717
rect 51744 887 51806 902
rect 51744 853 51760 887
rect 51794 853 51806 887
rect 51986 877 51998 911
rect 52032 877 52044 911
rect 51986 862 52044 877
rect 52074 1047 52132 1062
rect 52074 1013 52086 1047
rect 52120 1013 52132 1047
rect 52074 979 52132 1013
rect 52074 945 52086 979
rect 52120 945 52132 979
rect 52074 911 52132 945
rect 52074 877 52086 911
rect 52120 877 52132 911
rect 52268 1031 52276 1065
rect 52310 1031 52320 1065
rect 52268 997 52320 1031
rect 52268 963 52276 997
rect 52310 963 52320 997
rect 52268 929 52320 963
rect 52268 895 52276 929
rect 52310 895 52320 929
rect 52268 877 52320 895
rect 52350 1065 52402 1077
rect 52350 1031 52360 1065
rect 52394 1031 52402 1065
rect 52350 997 52402 1031
rect 52350 963 52360 997
rect 52394 963 52402 997
rect 52350 929 52402 963
rect 52350 895 52360 929
rect 52394 895 52402 929
rect 52573 1055 52625 1075
rect 52573 1021 52581 1055
rect 52615 1021 52625 1055
rect 52573 987 52625 1021
rect 52573 953 52581 987
rect 52615 953 52625 987
rect 52573 917 52625 953
rect 52655 1055 52713 1075
rect 52655 1021 52667 1055
rect 52701 1021 52713 1055
rect 52655 987 52713 1021
rect 52655 953 52667 987
rect 52701 953 52713 987
rect 52655 917 52713 953
rect 52743 1055 52795 1075
rect 52743 1021 52753 1055
rect 52787 1021 52795 1055
rect 52743 974 52795 1021
rect 52743 940 52753 974
rect 52787 940 52795 974
rect 52743 917 52795 940
rect 52960 1057 53012 1069
rect 52960 1023 52968 1057
rect 53002 1023 53012 1057
rect 52960 989 53012 1023
rect 52960 955 52968 989
rect 53002 955 53012 989
rect 52960 921 53012 955
rect 52350 877 52402 895
rect 52074 862 52132 877
rect 51744 819 51806 853
rect 51744 785 51760 819
rect 51794 785 51806 819
rect 51744 751 51806 785
rect 52960 887 52968 921
rect 53002 887 53012 921
rect 52960 869 53012 887
rect 53042 1057 53094 1069
rect 53042 1023 53052 1057
rect 53086 1023 53094 1057
rect 53042 989 53094 1023
rect 53042 955 53052 989
rect 53086 955 53094 989
rect 53042 921 53094 955
rect 53042 887 53052 921
rect 53086 887 53094 921
rect 53042 869 53094 887
rect 53228 1047 53286 1062
rect 53228 1013 53240 1047
rect 53274 1013 53286 1047
rect 53228 979 53286 1013
rect 53228 945 53240 979
rect 53274 945 53286 979
rect 53228 911 53286 945
rect 53228 877 53240 911
rect 53274 877 53286 911
rect 53228 862 53286 877
rect 53316 1047 53374 1062
rect 53316 1013 53328 1047
rect 53362 1013 53374 1047
rect 53316 979 53374 1013
rect 54156 1065 54208 1077
rect 53874 1047 53932 1062
rect 53874 1013 53886 1047
rect 53920 1013 53932 1047
rect 53316 945 53328 979
rect 53362 945 53374 979
rect 53316 911 53374 945
rect 53316 877 53328 911
rect 53362 877 53374 911
rect 53874 979 53932 1013
rect 53874 945 53886 979
rect 53920 945 53932 979
rect 53874 911 53932 945
rect 53316 862 53374 877
rect 53444 887 53506 902
rect 53444 853 53456 887
rect 53490 853 53506 887
rect 51744 717 51760 751
rect 51794 717 51806 751
rect 51744 702 51806 717
rect 53444 819 53506 853
rect 53444 785 53456 819
rect 53490 785 53506 819
rect 53444 751 53506 785
rect 53444 717 53456 751
rect 53490 717 53506 751
rect 53444 702 53506 717
rect 53536 887 53602 902
rect 53536 853 53552 887
rect 53586 853 53602 887
rect 53536 819 53602 853
rect 53536 785 53552 819
rect 53586 785 53602 819
rect 53536 751 53602 785
rect 53536 717 53552 751
rect 53586 717 53602 751
rect 53536 702 53602 717
rect 53632 887 53694 902
rect 53632 853 53648 887
rect 53682 853 53694 887
rect 53874 877 53886 911
rect 53920 877 53932 911
rect 53874 862 53932 877
rect 53962 1047 54020 1062
rect 53962 1013 53974 1047
rect 54008 1013 54020 1047
rect 53962 979 54020 1013
rect 53962 945 53974 979
rect 54008 945 54020 979
rect 53962 911 54020 945
rect 53962 877 53974 911
rect 54008 877 54020 911
rect 54156 1031 54164 1065
rect 54198 1031 54208 1065
rect 54156 997 54208 1031
rect 54156 963 54164 997
rect 54198 963 54208 997
rect 54156 929 54208 963
rect 54156 895 54164 929
rect 54198 895 54208 929
rect 54156 877 54208 895
rect 54238 1065 54290 1077
rect 54238 1031 54248 1065
rect 54282 1031 54290 1065
rect 54238 997 54290 1031
rect 54238 963 54248 997
rect 54282 963 54290 997
rect 54238 929 54290 963
rect 54238 895 54248 929
rect 54282 895 54290 929
rect 54461 1055 54513 1075
rect 54461 1021 54469 1055
rect 54503 1021 54513 1055
rect 54461 987 54513 1021
rect 54461 953 54469 987
rect 54503 953 54513 987
rect 54461 917 54513 953
rect 54543 1055 54601 1075
rect 54543 1021 54555 1055
rect 54589 1021 54601 1055
rect 54543 987 54601 1021
rect 54543 953 54555 987
rect 54589 953 54601 987
rect 54543 917 54601 953
rect 54631 1055 54683 1075
rect 54631 1021 54641 1055
rect 54675 1021 54683 1055
rect 54631 974 54683 1021
rect 54631 940 54641 974
rect 54675 940 54683 974
rect 54631 917 54683 940
rect 54848 1057 54900 1069
rect 54848 1023 54856 1057
rect 54890 1023 54900 1057
rect 54848 989 54900 1023
rect 54848 955 54856 989
rect 54890 955 54900 989
rect 54848 921 54900 955
rect 54238 877 54290 895
rect 53962 862 54020 877
rect 53632 819 53694 853
rect 53632 785 53648 819
rect 53682 785 53694 819
rect 53632 751 53694 785
rect 54848 887 54856 921
rect 54890 887 54900 921
rect 54848 869 54900 887
rect 54930 1057 54982 1069
rect 54930 1023 54940 1057
rect 54974 1023 54982 1057
rect 54930 989 54982 1023
rect 54930 955 54940 989
rect 54974 955 54982 989
rect 54930 921 54982 955
rect 54930 887 54940 921
rect 54974 887 54982 921
rect 54930 869 54982 887
rect 55116 1047 55174 1062
rect 55116 1013 55128 1047
rect 55162 1013 55174 1047
rect 55116 979 55174 1013
rect 55116 945 55128 979
rect 55162 945 55174 979
rect 55116 911 55174 945
rect 55116 877 55128 911
rect 55162 877 55174 911
rect 55116 862 55174 877
rect 55204 1047 55262 1062
rect 55204 1013 55216 1047
rect 55250 1013 55262 1047
rect 55204 979 55262 1013
rect 56044 1065 56096 1077
rect 55762 1047 55820 1062
rect 55762 1013 55774 1047
rect 55808 1013 55820 1047
rect 55204 945 55216 979
rect 55250 945 55262 979
rect 55204 911 55262 945
rect 55204 877 55216 911
rect 55250 877 55262 911
rect 55762 979 55820 1013
rect 55762 945 55774 979
rect 55808 945 55820 979
rect 55762 911 55820 945
rect 55204 862 55262 877
rect 55332 887 55394 902
rect 55332 853 55344 887
rect 55378 853 55394 887
rect 53632 717 53648 751
rect 53682 717 53694 751
rect 53632 702 53694 717
rect 55332 819 55394 853
rect 55332 785 55344 819
rect 55378 785 55394 819
rect 55332 751 55394 785
rect 55332 717 55344 751
rect 55378 717 55394 751
rect 55332 702 55394 717
rect 55424 887 55490 902
rect 55424 853 55440 887
rect 55474 853 55490 887
rect 55424 819 55490 853
rect 55424 785 55440 819
rect 55474 785 55490 819
rect 55424 751 55490 785
rect 55424 717 55440 751
rect 55474 717 55490 751
rect 55424 702 55490 717
rect 55520 887 55582 902
rect 55520 853 55536 887
rect 55570 853 55582 887
rect 55762 877 55774 911
rect 55808 877 55820 911
rect 55762 862 55820 877
rect 55850 1047 55908 1062
rect 55850 1013 55862 1047
rect 55896 1013 55908 1047
rect 55850 979 55908 1013
rect 55850 945 55862 979
rect 55896 945 55908 979
rect 55850 911 55908 945
rect 55850 877 55862 911
rect 55896 877 55908 911
rect 56044 1031 56052 1065
rect 56086 1031 56096 1065
rect 56044 997 56096 1031
rect 56044 963 56052 997
rect 56086 963 56096 997
rect 56044 929 56096 963
rect 56044 895 56052 929
rect 56086 895 56096 929
rect 56044 877 56096 895
rect 56126 1065 56178 1077
rect 56126 1031 56136 1065
rect 56170 1031 56178 1065
rect 56126 997 56178 1031
rect 56126 963 56136 997
rect 56170 963 56178 997
rect 56126 929 56178 963
rect 56126 895 56136 929
rect 56170 895 56178 929
rect 56349 1055 56401 1075
rect 56349 1021 56357 1055
rect 56391 1021 56401 1055
rect 56349 987 56401 1021
rect 56349 953 56357 987
rect 56391 953 56401 987
rect 56349 917 56401 953
rect 56431 1055 56489 1075
rect 56431 1021 56443 1055
rect 56477 1021 56489 1055
rect 56431 987 56489 1021
rect 56431 953 56443 987
rect 56477 953 56489 987
rect 56431 917 56489 953
rect 56519 1055 56571 1075
rect 56519 1021 56529 1055
rect 56563 1021 56571 1055
rect 56519 974 56571 1021
rect 56519 940 56529 974
rect 56563 940 56571 974
rect 56519 917 56571 940
rect 56736 1057 56788 1069
rect 56736 1023 56744 1057
rect 56778 1023 56788 1057
rect 56736 989 56788 1023
rect 56736 955 56744 989
rect 56778 955 56788 989
rect 56736 921 56788 955
rect 56126 877 56178 895
rect 55850 862 55908 877
rect 55520 819 55582 853
rect 55520 785 55536 819
rect 55570 785 55582 819
rect 55520 751 55582 785
rect 56736 887 56744 921
rect 56778 887 56788 921
rect 56736 869 56788 887
rect 56818 1057 56870 1069
rect 56818 1023 56828 1057
rect 56862 1023 56870 1057
rect 56818 989 56870 1023
rect 56818 955 56828 989
rect 56862 955 56870 989
rect 56818 921 56870 955
rect 56818 887 56828 921
rect 56862 887 56870 921
rect 56818 869 56870 887
rect 57004 1047 57062 1062
rect 57004 1013 57016 1047
rect 57050 1013 57062 1047
rect 57004 979 57062 1013
rect 57004 945 57016 979
rect 57050 945 57062 979
rect 57004 911 57062 945
rect 57004 877 57016 911
rect 57050 877 57062 911
rect 57004 862 57062 877
rect 57092 1047 57150 1062
rect 57092 1013 57104 1047
rect 57138 1013 57150 1047
rect 57092 979 57150 1013
rect 57932 1065 57984 1077
rect 57650 1047 57708 1062
rect 57650 1013 57662 1047
rect 57696 1013 57708 1047
rect 57092 945 57104 979
rect 57138 945 57150 979
rect 57092 911 57150 945
rect 57092 877 57104 911
rect 57138 877 57150 911
rect 57650 979 57708 1013
rect 57650 945 57662 979
rect 57696 945 57708 979
rect 57650 911 57708 945
rect 57092 862 57150 877
rect 57220 887 57282 902
rect 57220 853 57232 887
rect 57266 853 57282 887
rect 55520 717 55536 751
rect 55570 717 55582 751
rect 55520 702 55582 717
rect 57220 819 57282 853
rect 57220 785 57232 819
rect 57266 785 57282 819
rect 57220 751 57282 785
rect 57220 717 57232 751
rect 57266 717 57282 751
rect 57220 702 57282 717
rect 57312 887 57378 902
rect 57312 853 57328 887
rect 57362 853 57378 887
rect 57312 819 57378 853
rect 57312 785 57328 819
rect 57362 785 57378 819
rect 57312 751 57378 785
rect 57312 717 57328 751
rect 57362 717 57378 751
rect 57312 702 57378 717
rect 57408 887 57470 902
rect 57408 853 57424 887
rect 57458 853 57470 887
rect 57650 877 57662 911
rect 57696 877 57708 911
rect 57650 862 57708 877
rect 57738 1047 57796 1062
rect 57738 1013 57750 1047
rect 57784 1013 57796 1047
rect 57738 979 57796 1013
rect 57738 945 57750 979
rect 57784 945 57796 979
rect 57738 911 57796 945
rect 57738 877 57750 911
rect 57784 877 57796 911
rect 57932 1031 57940 1065
rect 57974 1031 57984 1065
rect 57932 997 57984 1031
rect 57932 963 57940 997
rect 57974 963 57984 997
rect 57932 929 57984 963
rect 57932 895 57940 929
rect 57974 895 57984 929
rect 57932 877 57984 895
rect 58014 1065 58066 1077
rect 58014 1031 58024 1065
rect 58058 1031 58066 1065
rect 58014 997 58066 1031
rect 58014 963 58024 997
rect 58058 963 58066 997
rect 58014 929 58066 963
rect 58014 895 58024 929
rect 58058 895 58066 929
rect 58237 1055 58289 1075
rect 58237 1021 58245 1055
rect 58279 1021 58289 1055
rect 58237 987 58289 1021
rect 58237 953 58245 987
rect 58279 953 58289 987
rect 58237 917 58289 953
rect 58319 1055 58377 1075
rect 58319 1021 58331 1055
rect 58365 1021 58377 1055
rect 58319 987 58377 1021
rect 58319 953 58331 987
rect 58365 953 58377 987
rect 58319 917 58377 953
rect 58407 1055 58459 1075
rect 58407 1021 58417 1055
rect 58451 1021 58459 1055
rect 58407 974 58459 1021
rect 58407 940 58417 974
rect 58451 940 58459 974
rect 58407 917 58459 940
rect 58624 1057 58676 1069
rect 58624 1023 58632 1057
rect 58666 1023 58676 1057
rect 58624 989 58676 1023
rect 58624 955 58632 989
rect 58666 955 58676 989
rect 58624 921 58676 955
rect 58014 877 58066 895
rect 57738 862 57796 877
rect 57408 819 57470 853
rect 57408 785 57424 819
rect 57458 785 57470 819
rect 57408 751 57470 785
rect 58624 887 58632 921
rect 58666 887 58676 921
rect 58624 869 58676 887
rect 58706 1057 58758 1069
rect 58706 1023 58716 1057
rect 58750 1023 58758 1057
rect 58706 989 58758 1023
rect 58706 955 58716 989
rect 58750 955 58758 989
rect 58706 921 58758 955
rect 58706 887 58716 921
rect 58750 887 58758 921
rect 58706 869 58758 887
rect 58892 1047 58950 1062
rect 58892 1013 58904 1047
rect 58938 1013 58950 1047
rect 58892 979 58950 1013
rect 58892 945 58904 979
rect 58938 945 58950 979
rect 58892 911 58950 945
rect 58892 877 58904 911
rect 58938 877 58950 911
rect 58892 862 58950 877
rect 58980 1047 59038 1062
rect 58980 1013 58992 1047
rect 59026 1013 59038 1047
rect 58980 979 59038 1013
rect 59820 1065 59872 1077
rect 59538 1047 59596 1062
rect 59538 1013 59550 1047
rect 59584 1013 59596 1047
rect 58980 945 58992 979
rect 59026 945 59038 979
rect 58980 911 59038 945
rect 58980 877 58992 911
rect 59026 877 59038 911
rect 59538 979 59596 1013
rect 59538 945 59550 979
rect 59584 945 59596 979
rect 59538 911 59596 945
rect 58980 862 59038 877
rect 59108 887 59170 902
rect 59108 853 59120 887
rect 59154 853 59170 887
rect 57408 717 57424 751
rect 57458 717 57470 751
rect 57408 702 57470 717
rect 59108 819 59170 853
rect 59108 785 59120 819
rect 59154 785 59170 819
rect 59108 751 59170 785
rect 59108 717 59120 751
rect 59154 717 59170 751
rect 59108 702 59170 717
rect 59200 887 59266 902
rect 59200 853 59216 887
rect 59250 853 59266 887
rect 59200 819 59266 853
rect 59200 785 59216 819
rect 59250 785 59266 819
rect 59200 751 59266 785
rect 59200 717 59216 751
rect 59250 717 59266 751
rect 59200 702 59266 717
rect 59296 887 59358 902
rect 59296 853 59312 887
rect 59346 853 59358 887
rect 59538 877 59550 911
rect 59584 877 59596 911
rect 59538 862 59596 877
rect 59626 1047 59684 1062
rect 59626 1013 59638 1047
rect 59672 1013 59684 1047
rect 59626 979 59684 1013
rect 59626 945 59638 979
rect 59672 945 59684 979
rect 59626 911 59684 945
rect 59626 877 59638 911
rect 59672 877 59684 911
rect 59820 1031 59828 1065
rect 59862 1031 59872 1065
rect 59820 997 59872 1031
rect 59820 963 59828 997
rect 59862 963 59872 997
rect 59820 929 59872 963
rect 59820 895 59828 929
rect 59862 895 59872 929
rect 59820 877 59872 895
rect 59902 1065 59954 1077
rect 59902 1031 59912 1065
rect 59946 1031 59954 1065
rect 59902 997 59954 1031
rect 59902 963 59912 997
rect 59946 963 59954 997
rect 59902 929 59954 963
rect 59902 895 59912 929
rect 59946 895 59954 929
rect 60125 1055 60177 1075
rect 60125 1021 60133 1055
rect 60167 1021 60177 1055
rect 60125 987 60177 1021
rect 60125 953 60133 987
rect 60167 953 60177 987
rect 60125 917 60177 953
rect 60207 1055 60265 1075
rect 60207 1021 60219 1055
rect 60253 1021 60265 1055
rect 60207 987 60265 1021
rect 60207 953 60219 987
rect 60253 953 60265 987
rect 60207 917 60265 953
rect 60295 1055 60347 1075
rect 60295 1021 60305 1055
rect 60339 1021 60347 1055
rect 60295 974 60347 1021
rect 60295 940 60305 974
rect 60339 940 60347 974
rect 60295 917 60347 940
rect 59902 877 59954 895
rect 59626 862 59684 877
rect 59296 819 59358 853
rect 59296 785 59312 819
rect 59346 785 59358 819
rect 59296 751 59358 785
rect 59296 717 59312 751
rect 59346 717 59358 751
rect 59296 702 59358 717
<< ndiffc >>
rect 620 7020 654 7054
rect 620 6952 654 6986
rect 716 7020 750 7054
rect 716 6952 750 6986
rect 812 7020 846 7054
rect 812 6952 846 6986
rect 2508 7020 2542 7054
rect 2508 6952 2542 6986
rect 2604 7020 2638 7054
rect 2604 6952 2638 6986
rect 2700 7020 2734 7054
rect 2700 6952 2734 6986
rect 4396 7020 4430 7054
rect 4396 6952 4430 6986
rect 4492 7020 4526 7054
rect 4492 6952 4526 6986
rect 4588 7020 4622 7054
rect 4588 6952 4622 6986
rect 6284 7020 6318 7054
rect 6284 6952 6318 6986
rect 6380 7020 6414 7054
rect 6380 6952 6414 6986
rect 6476 7020 6510 7054
rect 6476 6952 6510 6986
rect 8172 7020 8206 7054
rect 8172 6952 8206 6986
rect 8268 7020 8302 7054
rect 8268 6952 8302 6986
rect 8364 7020 8398 7054
rect 8364 6952 8398 6986
rect 10060 7020 10094 7054
rect 10060 6952 10094 6986
rect 10156 7020 10190 7054
rect 10156 6952 10190 6986
rect 10252 7020 10286 7054
rect 10252 6952 10286 6986
rect 11948 7020 11982 7054
rect 11948 6952 11982 6986
rect 12044 7020 12078 7054
rect 12044 6952 12078 6986
rect 12140 7020 12174 7054
rect 12140 6952 12174 6986
rect 13836 7020 13870 7054
rect 13836 6952 13870 6986
rect 13932 7020 13966 7054
rect 13932 6952 13966 6986
rect 14028 7020 14062 7054
rect 14028 6952 14062 6986
rect 15718 7020 15752 7054
rect 15718 6952 15752 6986
rect 15814 7020 15848 7054
rect 15814 6952 15848 6986
rect 15910 7020 15944 7054
rect 15910 6952 15944 6986
rect 17606 7020 17640 7054
rect 17606 6952 17640 6986
rect 17702 7020 17736 7054
rect 17702 6952 17736 6986
rect 17798 7020 17832 7054
rect 17798 6952 17832 6986
rect 19494 7020 19528 7054
rect 19494 6952 19528 6986
rect 19590 7020 19624 7054
rect 19590 6952 19624 6986
rect 19686 7020 19720 7054
rect 19686 6952 19720 6986
rect 21382 7020 21416 7054
rect 21382 6952 21416 6986
rect 21478 7020 21512 7054
rect 21478 6952 21512 6986
rect 21574 7020 21608 7054
rect 21574 6952 21608 6986
rect 23270 7020 23304 7054
rect 23270 6952 23304 6986
rect 23366 7020 23400 7054
rect 23366 6952 23400 6986
rect 23462 7020 23496 7054
rect 23462 6952 23496 6986
rect 25158 7020 25192 7054
rect 25158 6952 25192 6986
rect 25254 7020 25288 7054
rect 25254 6952 25288 6986
rect 25350 7020 25384 7054
rect 25350 6952 25384 6986
rect 27046 7020 27080 7054
rect 27046 6952 27080 6986
rect 27142 7020 27176 7054
rect 27142 6952 27176 6986
rect 27238 7020 27272 7054
rect 27238 6952 27272 6986
rect 28934 7020 28968 7054
rect 28934 6952 28968 6986
rect 29030 7020 29064 7054
rect 29030 6952 29064 6986
rect 29126 7020 29160 7054
rect 29126 6952 29160 6986
rect 30822 7020 30856 7054
rect 30822 6952 30856 6986
rect 30918 7020 30952 7054
rect 30918 6952 30952 6986
rect 31014 7020 31048 7054
rect 31014 6952 31048 6986
rect 32710 7020 32744 7054
rect 32710 6952 32744 6986
rect 32806 7020 32840 7054
rect 32806 6952 32840 6986
rect 32902 7020 32936 7054
rect 32902 6952 32936 6986
rect 34598 7020 34632 7054
rect 34598 6952 34632 6986
rect 34694 7020 34728 7054
rect 34694 6952 34728 6986
rect 34790 7020 34824 7054
rect 34790 6952 34824 6986
rect 36486 7020 36520 7054
rect 36486 6952 36520 6986
rect 36582 7020 36616 7054
rect 36582 6952 36616 6986
rect 36678 7020 36712 7054
rect 36678 6952 36712 6986
rect 38374 7020 38408 7054
rect 38374 6952 38408 6986
rect 38470 7020 38504 7054
rect 38470 6952 38504 6986
rect 38566 7020 38600 7054
rect 38566 6952 38600 6986
rect 40262 7020 40296 7054
rect 40262 6952 40296 6986
rect 40358 7020 40392 7054
rect 40358 6952 40392 6986
rect 40454 7020 40488 7054
rect 40454 6952 40488 6986
rect 42150 7020 42184 7054
rect 42150 6952 42184 6986
rect 42246 7020 42280 7054
rect 42246 6952 42280 6986
rect 42342 7020 42376 7054
rect 42342 6952 42376 6986
rect 44038 7020 44072 7054
rect 44038 6952 44072 6986
rect 44134 7020 44168 7054
rect 44134 6952 44168 6986
rect 44230 7020 44264 7054
rect 44230 6952 44264 6986
rect 45920 7020 45954 7054
rect 45920 6952 45954 6986
rect 46016 7020 46050 7054
rect 46016 6952 46050 6986
rect 46112 7020 46146 7054
rect 46112 6952 46146 6986
rect 47808 7020 47842 7054
rect 47808 6952 47842 6986
rect 47904 7020 47938 7054
rect 47904 6952 47938 6986
rect 48000 7020 48034 7054
rect 48000 6952 48034 6986
rect 49696 7020 49730 7054
rect 49696 6952 49730 6986
rect 49792 7020 49826 7054
rect 49792 6952 49826 6986
rect 49888 7020 49922 7054
rect 49888 6952 49922 6986
rect 51584 7020 51618 7054
rect 51584 6952 51618 6986
rect 51680 7020 51714 7054
rect 51680 6952 51714 6986
rect 51776 7020 51810 7054
rect 51776 6952 51810 6986
rect 53472 7020 53506 7054
rect 53472 6952 53506 6986
rect 53568 7020 53602 7054
rect 53568 6952 53602 6986
rect 53664 7020 53698 7054
rect 53664 6952 53698 6986
rect 55360 7020 55394 7054
rect 55360 6952 55394 6986
rect 55456 7020 55490 7054
rect 55456 6952 55490 6986
rect 55552 7020 55586 7054
rect 55552 6952 55586 6986
rect 57248 7020 57282 7054
rect 57248 6952 57282 6986
rect 57344 7020 57378 7054
rect 57344 6952 57378 6986
rect 57440 7020 57474 7054
rect 57440 6952 57474 6986
rect 59136 7020 59170 7054
rect 59136 6952 59170 6986
rect 59232 7020 59266 7054
rect 59232 6952 59266 6986
rect 59328 7020 59362 7054
rect 59328 6952 59362 6986
rect -357 6739 -323 6773
rect -271 6769 -237 6803
rect -185 6756 -151 6790
rect 36 6763 70 6797
rect 36 6695 70 6729
rect 120 6763 154 6797
rect 1232 6771 1266 6805
rect 120 6695 154 6729
rect 1232 6703 1266 6737
rect 1316 6771 1350 6805
rect 1316 6703 1350 6737
rect 1531 6739 1565 6773
rect 1617 6769 1651 6803
rect 1703 6756 1737 6790
rect 1924 6763 1958 6797
rect 1924 6695 1958 6729
rect 2008 6763 2042 6797
rect 3120 6771 3154 6805
rect 2008 6695 2042 6729
rect 3120 6703 3154 6737
rect 3204 6771 3238 6805
rect 3204 6703 3238 6737
rect 3419 6739 3453 6773
rect 3505 6769 3539 6803
rect 3591 6756 3625 6790
rect 3812 6763 3846 6797
rect 3812 6695 3846 6729
rect 3896 6763 3930 6797
rect 5008 6771 5042 6805
rect 3896 6695 3930 6729
rect 5008 6703 5042 6737
rect 5092 6771 5126 6805
rect 5092 6703 5126 6737
rect 5307 6739 5341 6773
rect 5393 6769 5427 6803
rect 5479 6756 5513 6790
rect 5700 6763 5734 6797
rect 5700 6695 5734 6729
rect 5784 6763 5818 6797
rect 6896 6771 6930 6805
rect 5784 6695 5818 6729
rect 6896 6703 6930 6737
rect 6980 6771 7014 6805
rect 6980 6703 7014 6737
rect 7195 6739 7229 6773
rect 7281 6769 7315 6803
rect 7367 6756 7401 6790
rect 7588 6763 7622 6797
rect 7588 6695 7622 6729
rect 7672 6763 7706 6797
rect 8784 6771 8818 6805
rect 7672 6695 7706 6729
rect 8784 6703 8818 6737
rect 8868 6771 8902 6805
rect 8868 6703 8902 6737
rect 9083 6739 9117 6773
rect 9169 6769 9203 6803
rect 9255 6756 9289 6790
rect 9476 6763 9510 6797
rect 9476 6695 9510 6729
rect 9560 6763 9594 6797
rect 10672 6771 10706 6805
rect 9560 6695 9594 6729
rect 10672 6703 10706 6737
rect 10756 6771 10790 6805
rect 10756 6703 10790 6737
rect 10971 6739 11005 6773
rect 11057 6769 11091 6803
rect 11143 6756 11177 6790
rect 11364 6763 11398 6797
rect 11364 6695 11398 6729
rect 11448 6763 11482 6797
rect 12560 6771 12594 6805
rect 11448 6695 11482 6729
rect 12560 6703 12594 6737
rect 12644 6771 12678 6805
rect 12644 6703 12678 6737
rect 12859 6739 12893 6773
rect 12945 6769 12979 6803
rect 13031 6756 13065 6790
rect 13252 6763 13286 6797
rect 13252 6695 13286 6729
rect 13336 6763 13370 6797
rect 14448 6771 14482 6805
rect 13336 6695 13370 6729
rect 14448 6703 14482 6737
rect 14532 6771 14566 6805
rect 14532 6703 14566 6737
rect 14741 6739 14775 6773
rect 14827 6769 14861 6803
rect 14913 6756 14947 6790
rect 15134 6763 15168 6797
rect 15134 6695 15168 6729
rect 15218 6763 15252 6797
rect 16330 6771 16364 6805
rect 15218 6695 15252 6729
rect 16330 6703 16364 6737
rect 16414 6771 16448 6805
rect 16414 6703 16448 6737
rect 16629 6739 16663 6773
rect 16715 6769 16749 6803
rect 16801 6756 16835 6790
rect 17022 6763 17056 6797
rect 17022 6695 17056 6729
rect 17106 6763 17140 6797
rect 18218 6771 18252 6805
rect 17106 6695 17140 6729
rect 18218 6703 18252 6737
rect 18302 6771 18336 6805
rect 18302 6703 18336 6737
rect 18517 6739 18551 6773
rect 18603 6769 18637 6803
rect 18689 6756 18723 6790
rect 18910 6763 18944 6797
rect 18910 6695 18944 6729
rect 18994 6763 19028 6797
rect 20106 6771 20140 6805
rect 18994 6695 19028 6729
rect 20106 6703 20140 6737
rect 20190 6771 20224 6805
rect 20190 6703 20224 6737
rect 20405 6739 20439 6773
rect 20491 6769 20525 6803
rect 20577 6756 20611 6790
rect 20798 6763 20832 6797
rect 20798 6695 20832 6729
rect 20882 6763 20916 6797
rect 21994 6771 22028 6805
rect 20882 6695 20916 6729
rect 21994 6703 22028 6737
rect 22078 6771 22112 6805
rect 22078 6703 22112 6737
rect 22293 6739 22327 6773
rect 22379 6769 22413 6803
rect 22465 6756 22499 6790
rect 22686 6763 22720 6797
rect 22686 6695 22720 6729
rect 22770 6763 22804 6797
rect 23882 6771 23916 6805
rect 22770 6695 22804 6729
rect 23882 6703 23916 6737
rect 23966 6771 24000 6805
rect 23966 6703 24000 6737
rect 24181 6739 24215 6773
rect 24267 6769 24301 6803
rect 24353 6756 24387 6790
rect 24574 6763 24608 6797
rect 24574 6695 24608 6729
rect 24658 6763 24692 6797
rect 25770 6771 25804 6805
rect 24658 6695 24692 6729
rect 25770 6703 25804 6737
rect 25854 6771 25888 6805
rect 25854 6703 25888 6737
rect 26069 6739 26103 6773
rect 26155 6769 26189 6803
rect 26241 6756 26275 6790
rect 26462 6763 26496 6797
rect 26462 6695 26496 6729
rect 26546 6763 26580 6797
rect 27658 6771 27692 6805
rect 26546 6695 26580 6729
rect 27658 6703 27692 6737
rect 27742 6771 27776 6805
rect 27742 6703 27776 6737
rect 27957 6739 27991 6773
rect 28043 6769 28077 6803
rect 28129 6756 28163 6790
rect 28350 6763 28384 6797
rect 28350 6695 28384 6729
rect 28434 6763 28468 6797
rect 29546 6771 29580 6805
rect 28434 6695 28468 6729
rect 29546 6703 29580 6737
rect 29630 6771 29664 6805
rect 29630 6703 29664 6737
rect 29845 6739 29879 6773
rect 29931 6769 29965 6803
rect 30017 6756 30051 6790
rect 30238 6763 30272 6797
rect 30238 6695 30272 6729
rect 30322 6763 30356 6797
rect 31434 6771 31468 6805
rect 30322 6695 30356 6729
rect 31434 6703 31468 6737
rect 31518 6771 31552 6805
rect 31518 6703 31552 6737
rect 31733 6739 31767 6773
rect 31819 6769 31853 6803
rect 31905 6756 31939 6790
rect 32126 6763 32160 6797
rect 32126 6695 32160 6729
rect 32210 6763 32244 6797
rect 33322 6771 33356 6805
rect 32210 6695 32244 6729
rect 33322 6703 33356 6737
rect 33406 6771 33440 6805
rect 33406 6703 33440 6737
rect 33621 6739 33655 6773
rect 33707 6769 33741 6803
rect 33793 6756 33827 6790
rect 34014 6763 34048 6797
rect 34014 6695 34048 6729
rect 34098 6763 34132 6797
rect 35210 6771 35244 6805
rect 34098 6695 34132 6729
rect 35210 6703 35244 6737
rect 35294 6771 35328 6805
rect 35294 6703 35328 6737
rect 35509 6739 35543 6773
rect 35595 6769 35629 6803
rect 35681 6756 35715 6790
rect 35902 6763 35936 6797
rect 35902 6695 35936 6729
rect 35986 6763 36020 6797
rect 37098 6771 37132 6805
rect 35986 6695 36020 6729
rect 37098 6703 37132 6737
rect 37182 6771 37216 6805
rect 37182 6703 37216 6737
rect 37397 6739 37431 6773
rect 37483 6769 37517 6803
rect 37569 6756 37603 6790
rect 37790 6763 37824 6797
rect 37790 6695 37824 6729
rect 37874 6763 37908 6797
rect 38986 6771 39020 6805
rect 37874 6695 37908 6729
rect 38986 6703 39020 6737
rect 39070 6771 39104 6805
rect 39070 6703 39104 6737
rect 39285 6739 39319 6773
rect 39371 6769 39405 6803
rect 39457 6756 39491 6790
rect 39678 6763 39712 6797
rect 39678 6695 39712 6729
rect 39762 6763 39796 6797
rect 40874 6771 40908 6805
rect 39762 6695 39796 6729
rect 40874 6703 40908 6737
rect 40958 6771 40992 6805
rect 40958 6703 40992 6737
rect 41173 6739 41207 6773
rect 41259 6769 41293 6803
rect 41345 6756 41379 6790
rect 41566 6763 41600 6797
rect 41566 6695 41600 6729
rect 41650 6763 41684 6797
rect 42762 6771 42796 6805
rect 41650 6695 41684 6729
rect 42762 6703 42796 6737
rect 42846 6771 42880 6805
rect 42846 6703 42880 6737
rect 43061 6739 43095 6773
rect 43147 6769 43181 6803
rect 43233 6756 43267 6790
rect 43454 6763 43488 6797
rect 43454 6695 43488 6729
rect 43538 6763 43572 6797
rect 44650 6771 44684 6805
rect 43538 6695 43572 6729
rect 44650 6703 44684 6737
rect 44734 6771 44768 6805
rect 44734 6703 44768 6737
rect 44943 6739 44977 6773
rect 45029 6769 45063 6803
rect 45115 6756 45149 6790
rect 45336 6763 45370 6797
rect 45336 6695 45370 6729
rect 45420 6763 45454 6797
rect 46532 6771 46566 6805
rect 45420 6695 45454 6729
rect 46532 6703 46566 6737
rect 46616 6771 46650 6805
rect 46616 6703 46650 6737
rect 46831 6739 46865 6773
rect 46917 6769 46951 6803
rect 47003 6756 47037 6790
rect 47224 6763 47258 6797
rect 47224 6695 47258 6729
rect 47308 6763 47342 6797
rect 48420 6771 48454 6805
rect 47308 6695 47342 6729
rect 48420 6703 48454 6737
rect 48504 6771 48538 6805
rect 48504 6703 48538 6737
rect 48719 6739 48753 6773
rect 48805 6769 48839 6803
rect 48891 6756 48925 6790
rect 49112 6763 49146 6797
rect 49112 6695 49146 6729
rect 49196 6763 49230 6797
rect 50308 6771 50342 6805
rect 49196 6695 49230 6729
rect 50308 6703 50342 6737
rect 50392 6771 50426 6805
rect 50392 6703 50426 6737
rect 50607 6739 50641 6773
rect 50693 6769 50727 6803
rect 50779 6756 50813 6790
rect 51000 6763 51034 6797
rect 51000 6695 51034 6729
rect 51084 6763 51118 6797
rect 52196 6771 52230 6805
rect 51084 6695 51118 6729
rect 52196 6703 52230 6737
rect 52280 6771 52314 6805
rect 52280 6703 52314 6737
rect 52495 6739 52529 6773
rect 52581 6769 52615 6803
rect 52667 6756 52701 6790
rect 52888 6763 52922 6797
rect 52888 6695 52922 6729
rect 52972 6763 53006 6797
rect 54084 6771 54118 6805
rect 52972 6695 53006 6729
rect 54084 6703 54118 6737
rect 54168 6771 54202 6805
rect 54168 6703 54202 6737
rect 54383 6739 54417 6773
rect 54469 6769 54503 6803
rect 54555 6756 54589 6790
rect 54776 6763 54810 6797
rect 54776 6695 54810 6729
rect 54860 6763 54894 6797
rect 55972 6771 56006 6805
rect 54860 6695 54894 6729
rect 55972 6703 56006 6737
rect 56056 6771 56090 6805
rect 56056 6703 56090 6737
rect 56271 6739 56305 6773
rect 56357 6769 56391 6803
rect 56443 6756 56477 6790
rect 56664 6763 56698 6797
rect 56664 6695 56698 6729
rect 56748 6763 56782 6797
rect 57860 6771 57894 6805
rect 56748 6695 56782 6729
rect 57860 6703 57894 6737
rect 57944 6771 57978 6805
rect 57944 6703 57978 6737
rect 58159 6739 58193 6773
rect 58245 6769 58279 6803
rect 58331 6756 58365 6790
rect 58552 6763 58586 6797
rect 58552 6695 58586 6729
rect 58636 6763 58670 6797
rect 59748 6771 59782 6805
rect 58636 6695 58670 6729
rect 59748 6703 59782 6737
rect 59832 6771 59866 6805
rect 59832 6703 59866 6737
rect 618 5964 652 5998
rect 618 5896 652 5930
rect 714 5964 748 5998
rect 714 5896 748 5930
rect 810 5964 844 5998
rect 810 5896 844 5930
rect 2506 5964 2540 5998
rect 2506 5896 2540 5930
rect 2602 5964 2636 5998
rect 2602 5896 2636 5930
rect 2698 5964 2732 5998
rect 2698 5896 2732 5930
rect 4394 5964 4428 5998
rect 4394 5896 4428 5930
rect 4490 5964 4524 5998
rect 4490 5896 4524 5930
rect 4586 5964 4620 5998
rect 4586 5896 4620 5930
rect 6282 5964 6316 5998
rect 6282 5896 6316 5930
rect 6378 5964 6412 5998
rect 6378 5896 6412 5930
rect 6474 5964 6508 5998
rect 6474 5896 6508 5930
rect 8170 5964 8204 5998
rect 8170 5896 8204 5930
rect 8266 5964 8300 5998
rect 8266 5896 8300 5930
rect 8362 5964 8396 5998
rect 8362 5896 8396 5930
rect 10058 5964 10092 5998
rect 10058 5896 10092 5930
rect 10154 5964 10188 5998
rect 10154 5896 10188 5930
rect 10250 5964 10284 5998
rect 10250 5896 10284 5930
rect 11946 5964 11980 5998
rect 11946 5896 11980 5930
rect 12042 5964 12076 5998
rect 12042 5896 12076 5930
rect 12138 5964 12172 5998
rect 12138 5896 12172 5930
rect 13834 5964 13868 5998
rect 13834 5896 13868 5930
rect 13930 5964 13964 5998
rect 13930 5896 13964 5930
rect 14026 5964 14060 5998
rect 14026 5896 14060 5930
rect 15716 5964 15750 5998
rect 15716 5896 15750 5930
rect 15812 5964 15846 5998
rect 15812 5896 15846 5930
rect 15908 5964 15942 5998
rect 15908 5896 15942 5930
rect 17604 5964 17638 5998
rect 17604 5896 17638 5930
rect 17700 5964 17734 5998
rect 17700 5896 17734 5930
rect 17796 5964 17830 5998
rect 17796 5896 17830 5930
rect 19492 5964 19526 5998
rect 19492 5896 19526 5930
rect 19588 5964 19622 5998
rect 19588 5896 19622 5930
rect 19684 5964 19718 5998
rect 19684 5896 19718 5930
rect 21380 5964 21414 5998
rect 21380 5896 21414 5930
rect 21476 5964 21510 5998
rect 21476 5896 21510 5930
rect 21572 5964 21606 5998
rect 21572 5896 21606 5930
rect 23268 5964 23302 5998
rect 23268 5896 23302 5930
rect 23364 5964 23398 5998
rect 23364 5896 23398 5930
rect 23460 5964 23494 5998
rect 23460 5896 23494 5930
rect 25156 5964 25190 5998
rect 25156 5896 25190 5930
rect 25252 5964 25286 5998
rect 25252 5896 25286 5930
rect 25348 5964 25382 5998
rect 25348 5896 25382 5930
rect 27044 5964 27078 5998
rect 27044 5896 27078 5930
rect 27140 5964 27174 5998
rect 27140 5896 27174 5930
rect 27236 5964 27270 5998
rect 27236 5896 27270 5930
rect 28932 5964 28966 5998
rect 28932 5896 28966 5930
rect 29028 5964 29062 5998
rect 29028 5896 29062 5930
rect 29124 5964 29158 5998
rect 29124 5896 29158 5930
rect 30820 5964 30854 5998
rect 30820 5896 30854 5930
rect 30916 5964 30950 5998
rect 30916 5896 30950 5930
rect 31012 5964 31046 5998
rect 31012 5896 31046 5930
rect 32708 5964 32742 5998
rect 32708 5896 32742 5930
rect 32804 5964 32838 5998
rect 32804 5896 32838 5930
rect 32900 5964 32934 5998
rect 32900 5896 32934 5930
rect 34596 5964 34630 5998
rect 34596 5896 34630 5930
rect 34692 5964 34726 5998
rect 34692 5896 34726 5930
rect 34788 5964 34822 5998
rect 34788 5896 34822 5930
rect 36484 5964 36518 5998
rect 36484 5896 36518 5930
rect 36580 5964 36614 5998
rect 36580 5896 36614 5930
rect 36676 5964 36710 5998
rect 36676 5896 36710 5930
rect 38372 5964 38406 5998
rect 38372 5896 38406 5930
rect 38468 5964 38502 5998
rect 38468 5896 38502 5930
rect 38564 5964 38598 5998
rect 38564 5896 38598 5930
rect 40260 5964 40294 5998
rect 40260 5896 40294 5930
rect 40356 5964 40390 5998
rect 40356 5896 40390 5930
rect 40452 5964 40486 5998
rect 40452 5896 40486 5930
rect 42148 5964 42182 5998
rect 42148 5896 42182 5930
rect 42244 5964 42278 5998
rect 42244 5896 42278 5930
rect 42340 5964 42374 5998
rect 42340 5896 42374 5930
rect 44036 5964 44070 5998
rect 44036 5896 44070 5930
rect 44132 5964 44166 5998
rect 44132 5896 44166 5930
rect 44228 5964 44262 5998
rect 44228 5896 44262 5930
rect 45918 5964 45952 5998
rect 45918 5896 45952 5930
rect 46014 5964 46048 5998
rect 46014 5896 46048 5930
rect 46110 5964 46144 5998
rect 46110 5896 46144 5930
rect 47806 5964 47840 5998
rect 47806 5896 47840 5930
rect 47902 5964 47936 5998
rect 47902 5896 47936 5930
rect 47998 5964 48032 5998
rect 47998 5896 48032 5930
rect 49694 5964 49728 5998
rect 49694 5896 49728 5930
rect 49790 5964 49824 5998
rect 49790 5896 49824 5930
rect 49886 5964 49920 5998
rect 49886 5896 49920 5930
rect 51582 5964 51616 5998
rect 51582 5896 51616 5930
rect 51678 5964 51712 5998
rect 51678 5896 51712 5930
rect 51774 5964 51808 5998
rect 51774 5896 51808 5930
rect 53470 5964 53504 5998
rect 53470 5896 53504 5930
rect 53566 5964 53600 5998
rect 53566 5896 53600 5930
rect 53662 5964 53696 5998
rect 53662 5896 53696 5930
rect 55358 5964 55392 5998
rect 55358 5896 55392 5930
rect 55454 5964 55488 5998
rect 55454 5896 55488 5930
rect 55550 5964 55584 5998
rect 55550 5896 55584 5930
rect 57246 5964 57280 5998
rect 57246 5896 57280 5930
rect 57342 5964 57376 5998
rect 57342 5896 57376 5930
rect 57438 5964 57472 5998
rect 57438 5896 57472 5930
rect 59134 5964 59168 5998
rect 59134 5896 59168 5930
rect 59230 5964 59264 5998
rect 59230 5896 59264 5930
rect 59326 5964 59360 5998
rect 59326 5896 59360 5930
rect 197 5719 231 5753
rect 197 5651 231 5685
rect 281 5719 315 5753
rect 281 5651 315 5685
rect 365 5719 399 5753
rect 1011 5719 1045 5753
rect 365 5651 399 5685
rect 1011 5651 1045 5685
rect 1095 5719 1129 5753
rect 1095 5651 1129 5685
rect 1179 5719 1213 5753
rect 1179 5651 1213 5685
rect 2085 5719 2119 5753
rect 2085 5651 2119 5685
rect 2169 5719 2203 5753
rect 2169 5651 2203 5685
rect 2253 5719 2287 5753
rect 2899 5719 2933 5753
rect 2253 5651 2287 5685
rect 2899 5651 2933 5685
rect 2983 5719 3017 5753
rect 2983 5651 3017 5685
rect 3067 5719 3101 5753
rect 3067 5651 3101 5685
rect 3973 5719 4007 5753
rect 3973 5651 4007 5685
rect 4057 5719 4091 5753
rect 4057 5651 4091 5685
rect 4141 5719 4175 5753
rect 4787 5719 4821 5753
rect 4141 5651 4175 5685
rect 4787 5651 4821 5685
rect 4871 5719 4905 5753
rect 4871 5651 4905 5685
rect 4955 5719 4989 5753
rect 4955 5651 4989 5685
rect 5861 5719 5895 5753
rect 5861 5651 5895 5685
rect 5945 5719 5979 5753
rect 5945 5651 5979 5685
rect 6029 5719 6063 5753
rect 6675 5719 6709 5753
rect 6029 5651 6063 5685
rect 6675 5651 6709 5685
rect 6759 5719 6793 5753
rect 6759 5651 6793 5685
rect 6843 5719 6877 5753
rect 6843 5651 6877 5685
rect 7749 5719 7783 5753
rect 7749 5651 7783 5685
rect 7833 5719 7867 5753
rect 7833 5651 7867 5685
rect 7917 5719 7951 5753
rect 8563 5719 8597 5753
rect 7917 5651 7951 5685
rect 8563 5651 8597 5685
rect 8647 5719 8681 5753
rect 8647 5651 8681 5685
rect 8731 5719 8765 5753
rect 8731 5651 8765 5685
rect 9637 5719 9671 5753
rect 9637 5651 9671 5685
rect 9721 5719 9755 5753
rect 9721 5651 9755 5685
rect 9805 5719 9839 5753
rect 10451 5719 10485 5753
rect 9805 5651 9839 5685
rect 10451 5651 10485 5685
rect 10535 5719 10569 5753
rect 10535 5651 10569 5685
rect 10619 5719 10653 5753
rect 10619 5651 10653 5685
rect 11525 5719 11559 5753
rect 11525 5651 11559 5685
rect 11609 5719 11643 5753
rect 11609 5651 11643 5685
rect 11693 5719 11727 5753
rect 12339 5719 12373 5753
rect 11693 5651 11727 5685
rect 12339 5651 12373 5685
rect 12423 5719 12457 5753
rect 12423 5651 12457 5685
rect 12507 5719 12541 5753
rect 12507 5651 12541 5685
rect 13413 5719 13447 5753
rect 13413 5651 13447 5685
rect 13497 5719 13531 5753
rect 13497 5651 13531 5685
rect 13581 5719 13615 5753
rect 14227 5719 14261 5753
rect 13581 5651 13615 5685
rect 14227 5651 14261 5685
rect 14311 5719 14345 5753
rect 14311 5651 14345 5685
rect 14395 5719 14429 5753
rect 14395 5651 14429 5685
rect 15295 5719 15329 5753
rect 15295 5651 15329 5685
rect 15379 5719 15413 5753
rect 15379 5651 15413 5685
rect 15463 5719 15497 5753
rect 16109 5719 16143 5753
rect 15463 5651 15497 5685
rect 16109 5651 16143 5685
rect 16193 5719 16227 5753
rect 16193 5651 16227 5685
rect 16277 5719 16311 5753
rect 16277 5651 16311 5685
rect 17183 5719 17217 5753
rect 17183 5651 17217 5685
rect 17267 5719 17301 5753
rect 17267 5651 17301 5685
rect 17351 5719 17385 5753
rect 17997 5719 18031 5753
rect 17351 5651 17385 5685
rect 17997 5651 18031 5685
rect 18081 5719 18115 5753
rect 18081 5651 18115 5685
rect 18165 5719 18199 5753
rect 18165 5651 18199 5685
rect 19071 5719 19105 5753
rect 19071 5651 19105 5685
rect 19155 5719 19189 5753
rect 19155 5651 19189 5685
rect 19239 5719 19273 5753
rect 19885 5719 19919 5753
rect 19239 5651 19273 5685
rect 19885 5651 19919 5685
rect 19969 5719 20003 5753
rect 19969 5651 20003 5685
rect 20053 5719 20087 5753
rect 20053 5651 20087 5685
rect 20959 5719 20993 5753
rect 20959 5651 20993 5685
rect 21043 5719 21077 5753
rect 21043 5651 21077 5685
rect 21127 5719 21161 5753
rect 21773 5719 21807 5753
rect 21127 5651 21161 5685
rect 21773 5651 21807 5685
rect 21857 5719 21891 5753
rect 21857 5651 21891 5685
rect 21941 5719 21975 5753
rect 21941 5651 21975 5685
rect 22847 5719 22881 5753
rect 22847 5651 22881 5685
rect 22931 5719 22965 5753
rect 22931 5651 22965 5685
rect 23015 5719 23049 5753
rect 23661 5719 23695 5753
rect 23015 5651 23049 5685
rect 23661 5651 23695 5685
rect 23745 5719 23779 5753
rect 23745 5651 23779 5685
rect 23829 5719 23863 5753
rect 23829 5651 23863 5685
rect 24735 5719 24769 5753
rect 24735 5651 24769 5685
rect 24819 5719 24853 5753
rect 24819 5651 24853 5685
rect 24903 5719 24937 5753
rect 25549 5719 25583 5753
rect 24903 5651 24937 5685
rect 25549 5651 25583 5685
rect 25633 5719 25667 5753
rect 25633 5651 25667 5685
rect 25717 5719 25751 5753
rect 25717 5651 25751 5685
rect 26623 5719 26657 5753
rect 26623 5651 26657 5685
rect 26707 5719 26741 5753
rect 26707 5651 26741 5685
rect 26791 5719 26825 5753
rect 27437 5719 27471 5753
rect 26791 5651 26825 5685
rect 27437 5651 27471 5685
rect 27521 5719 27555 5753
rect 27521 5651 27555 5685
rect 27605 5719 27639 5753
rect 27605 5651 27639 5685
rect 28511 5719 28545 5753
rect 28511 5651 28545 5685
rect 28595 5719 28629 5753
rect 28595 5651 28629 5685
rect 28679 5719 28713 5753
rect 29325 5719 29359 5753
rect 28679 5651 28713 5685
rect 29325 5651 29359 5685
rect 29409 5719 29443 5753
rect 29409 5651 29443 5685
rect 29493 5719 29527 5753
rect 29493 5651 29527 5685
rect 30399 5719 30433 5753
rect 30399 5651 30433 5685
rect 30483 5719 30517 5753
rect 30483 5651 30517 5685
rect 30567 5719 30601 5753
rect 31213 5719 31247 5753
rect 30567 5651 30601 5685
rect 31213 5651 31247 5685
rect 31297 5719 31331 5753
rect 31297 5651 31331 5685
rect 31381 5719 31415 5753
rect 31381 5651 31415 5685
rect 32287 5719 32321 5753
rect 32287 5651 32321 5685
rect 32371 5719 32405 5753
rect 32371 5651 32405 5685
rect 32455 5719 32489 5753
rect 33101 5719 33135 5753
rect 32455 5651 32489 5685
rect 33101 5651 33135 5685
rect 33185 5719 33219 5753
rect 33185 5651 33219 5685
rect 33269 5719 33303 5753
rect 33269 5651 33303 5685
rect 34175 5719 34209 5753
rect 34175 5651 34209 5685
rect 34259 5719 34293 5753
rect 34259 5651 34293 5685
rect 34343 5719 34377 5753
rect 34989 5719 35023 5753
rect 34343 5651 34377 5685
rect 34989 5651 35023 5685
rect 35073 5719 35107 5753
rect 35073 5651 35107 5685
rect 35157 5719 35191 5753
rect 35157 5651 35191 5685
rect 36063 5719 36097 5753
rect 36063 5651 36097 5685
rect 36147 5719 36181 5753
rect 36147 5651 36181 5685
rect 36231 5719 36265 5753
rect 36877 5719 36911 5753
rect 36231 5651 36265 5685
rect 36877 5651 36911 5685
rect 36961 5719 36995 5753
rect 36961 5651 36995 5685
rect 37045 5719 37079 5753
rect 37045 5651 37079 5685
rect 37951 5719 37985 5753
rect 37951 5651 37985 5685
rect 38035 5719 38069 5753
rect 38035 5651 38069 5685
rect 38119 5719 38153 5753
rect 38765 5719 38799 5753
rect 38119 5651 38153 5685
rect 38765 5651 38799 5685
rect 38849 5719 38883 5753
rect 38849 5651 38883 5685
rect 38933 5719 38967 5753
rect 38933 5651 38967 5685
rect 39839 5719 39873 5753
rect 39839 5651 39873 5685
rect 39923 5719 39957 5753
rect 39923 5651 39957 5685
rect 40007 5719 40041 5753
rect 40653 5719 40687 5753
rect 40007 5651 40041 5685
rect 40653 5651 40687 5685
rect 40737 5719 40771 5753
rect 40737 5651 40771 5685
rect 40821 5719 40855 5753
rect 40821 5651 40855 5685
rect 41727 5719 41761 5753
rect 41727 5651 41761 5685
rect 41811 5719 41845 5753
rect 41811 5651 41845 5685
rect 41895 5719 41929 5753
rect 42541 5719 42575 5753
rect 41895 5651 41929 5685
rect 42541 5651 42575 5685
rect 42625 5719 42659 5753
rect 42625 5651 42659 5685
rect 42709 5719 42743 5753
rect 42709 5651 42743 5685
rect 43615 5719 43649 5753
rect 43615 5651 43649 5685
rect 43699 5719 43733 5753
rect 43699 5651 43733 5685
rect 43783 5719 43817 5753
rect 44429 5719 44463 5753
rect 43783 5651 43817 5685
rect 44429 5651 44463 5685
rect 44513 5719 44547 5753
rect 44513 5651 44547 5685
rect 44597 5719 44631 5753
rect 44597 5651 44631 5685
rect 45497 5719 45531 5753
rect 45497 5651 45531 5685
rect 45581 5719 45615 5753
rect 45581 5651 45615 5685
rect 45665 5719 45699 5753
rect 46311 5719 46345 5753
rect 45665 5651 45699 5685
rect 46311 5651 46345 5685
rect 46395 5719 46429 5753
rect 46395 5651 46429 5685
rect 46479 5719 46513 5753
rect 46479 5651 46513 5685
rect 47385 5719 47419 5753
rect 47385 5651 47419 5685
rect 47469 5719 47503 5753
rect 47469 5651 47503 5685
rect 47553 5719 47587 5753
rect 48199 5719 48233 5753
rect 47553 5651 47587 5685
rect 48199 5651 48233 5685
rect 48283 5719 48317 5753
rect 48283 5651 48317 5685
rect 48367 5719 48401 5753
rect 48367 5651 48401 5685
rect 49273 5719 49307 5753
rect 49273 5651 49307 5685
rect 49357 5719 49391 5753
rect 49357 5651 49391 5685
rect 49441 5719 49475 5753
rect 50087 5719 50121 5753
rect 49441 5651 49475 5685
rect 50087 5651 50121 5685
rect 50171 5719 50205 5753
rect 50171 5651 50205 5685
rect 50255 5719 50289 5753
rect 50255 5651 50289 5685
rect 51161 5719 51195 5753
rect 51161 5651 51195 5685
rect 51245 5719 51279 5753
rect 51245 5651 51279 5685
rect 51329 5719 51363 5753
rect 51975 5719 52009 5753
rect 51329 5651 51363 5685
rect 51975 5651 52009 5685
rect 52059 5719 52093 5753
rect 52059 5651 52093 5685
rect 52143 5719 52177 5753
rect 52143 5651 52177 5685
rect 53049 5719 53083 5753
rect 53049 5651 53083 5685
rect 53133 5719 53167 5753
rect 53133 5651 53167 5685
rect 53217 5719 53251 5753
rect 53863 5719 53897 5753
rect 53217 5651 53251 5685
rect 53863 5651 53897 5685
rect 53947 5719 53981 5753
rect 53947 5651 53981 5685
rect 54031 5719 54065 5753
rect 54031 5651 54065 5685
rect 54937 5719 54971 5753
rect 54937 5651 54971 5685
rect 55021 5719 55055 5753
rect 55021 5651 55055 5685
rect 55105 5719 55139 5753
rect 55751 5719 55785 5753
rect 55105 5651 55139 5685
rect 55751 5651 55785 5685
rect 55835 5719 55869 5753
rect 55835 5651 55869 5685
rect 55919 5719 55953 5753
rect 55919 5651 55953 5685
rect 56825 5719 56859 5753
rect 56825 5651 56859 5685
rect 56909 5719 56943 5753
rect 56909 5651 56943 5685
rect 56993 5719 57027 5753
rect 57639 5719 57673 5753
rect 56993 5651 57027 5685
rect 57639 5651 57673 5685
rect 57723 5719 57757 5753
rect 57723 5651 57757 5685
rect 57807 5719 57841 5753
rect 57807 5651 57841 5685
rect 58713 5719 58747 5753
rect 58713 5651 58747 5685
rect 58797 5719 58831 5753
rect 58797 5651 58831 5685
rect 58881 5719 58915 5753
rect 59527 5719 59561 5753
rect 58881 5651 58915 5685
rect 59527 5651 59561 5685
rect 59611 5719 59645 5753
rect 59611 5651 59645 5685
rect 59695 5719 59729 5753
rect 59695 5651 59729 5685
rect 5710 4775 5744 4809
rect 5710 4707 5744 4741
rect 5794 4775 5828 4809
rect 5794 4707 5828 4741
rect 5878 4707 5912 4741
rect 5962 4775 5996 4809
rect 5962 4707 5996 4741
rect 6046 4707 6080 4741
rect 6130 4775 6164 4809
rect 6130 4707 6164 4741
rect 6214 4707 6248 4741
rect 6298 4775 6332 4809
rect 6298 4707 6332 4741
rect 6382 4707 6416 4741
rect 6466 4775 6500 4809
rect 6466 4707 6500 4741
rect 6550 4707 6584 4741
rect 6634 4775 6668 4809
rect 6634 4707 6668 4741
rect 6718 4707 6752 4741
rect 6802 4775 6836 4809
rect 6802 4707 6836 4741
rect 6886 4707 6920 4741
rect 6970 4775 7004 4809
rect 6970 4707 7004 4741
rect 7054 4775 7088 4809
rect 7054 4707 7088 4741
rect 7592 4773 7626 4807
rect 7592 4705 7626 4739
rect 7676 4773 7710 4807
rect 7676 4705 7710 4739
rect 7760 4705 7794 4739
rect 7844 4773 7878 4807
rect 7844 4705 7878 4739
rect 7928 4705 7962 4739
rect 8012 4773 8046 4807
rect 8012 4705 8046 4739
rect 8096 4705 8130 4739
rect 8180 4773 8214 4807
rect 8180 4705 8214 4739
rect 8264 4705 8298 4739
rect 8348 4773 8382 4807
rect 8348 4705 8382 4739
rect 8432 4705 8466 4739
rect 8516 4773 8550 4807
rect 8516 4705 8550 4739
rect 8600 4705 8634 4739
rect 8684 4773 8718 4807
rect 8684 4705 8718 4739
rect 8768 4705 8802 4739
rect 8852 4773 8886 4807
rect 8852 4705 8886 4739
rect 8936 4773 8970 4807
rect 8936 4705 8970 4739
rect 20808 4775 20842 4809
rect 20808 4707 20842 4741
rect 20892 4775 20926 4809
rect 20892 4707 20926 4741
rect 20976 4707 21010 4741
rect 21060 4775 21094 4809
rect 21060 4707 21094 4741
rect 21144 4707 21178 4741
rect 21228 4775 21262 4809
rect 21228 4707 21262 4741
rect 21312 4707 21346 4741
rect 21396 4775 21430 4809
rect 21396 4707 21430 4741
rect 21480 4707 21514 4741
rect 21564 4775 21598 4809
rect 21564 4707 21598 4741
rect 21648 4707 21682 4741
rect 21732 4775 21766 4809
rect 21732 4707 21766 4741
rect 21816 4707 21850 4741
rect 21900 4775 21934 4809
rect 21900 4707 21934 4741
rect 21984 4707 22018 4741
rect 22068 4775 22102 4809
rect 22068 4707 22102 4741
rect 22152 4775 22186 4809
rect 22152 4707 22186 4741
rect 22690 4773 22724 4807
rect 22690 4705 22724 4739
rect 22774 4773 22808 4807
rect 22774 4705 22808 4739
rect 22858 4705 22892 4739
rect 22942 4773 22976 4807
rect 22942 4705 22976 4739
rect 23026 4705 23060 4739
rect 23110 4773 23144 4807
rect 23110 4705 23144 4739
rect 23194 4705 23228 4739
rect 23278 4773 23312 4807
rect 23278 4705 23312 4739
rect 23362 4705 23396 4739
rect 23446 4773 23480 4807
rect 23446 4705 23480 4739
rect 23530 4705 23564 4739
rect 23614 4773 23648 4807
rect 23614 4705 23648 4739
rect 23698 4705 23732 4739
rect 23782 4773 23816 4807
rect 23782 4705 23816 4739
rect 23866 4705 23900 4739
rect 23950 4773 23984 4807
rect 23950 4705 23984 4739
rect 24034 4773 24068 4807
rect 24034 4705 24068 4739
rect 35912 4775 35946 4809
rect 35912 4707 35946 4741
rect 35996 4775 36030 4809
rect 35996 4707 36030 4741
rect 36080 4707 36114 4741
rect 36164 4775 36198 4809
rect 36164 4707 36198 4741
rect 36248 4707 36282 4741
rect 36332 4775 36366 4809
rect 36332 4707 36366 4741
rect 36416 4707 36450 4741
rect 36500 4775 36534 4809
rect 36500 4707 36534 4741
rect 36584 4707 36618 4741
rect 36668 4775 36702 4809
rect 36668 4707 36702 4741
rect 36752 4707 36786 4741
rect 36836 4775 36870 4809
rect 36836 4707 36870 4741
rect 36920 4707 36954 4741
rect 37004 4775 37038 4809
rect 37004 4707 37038 4741
rect 37088 4707 37122 4741
rect 37172 4775 37206 4809
rect 37172 4707 37206 4741
rect 37256 4775 37290 4809
rect 37256 4707 37290 4741
rect 37794 4773 37828 4807
rect 37794 4705 37828 4739
rect 37878 4773 37912 4807
rect 37878 4705 37912 4739
rect 37962 4705 37996 4739
rect 38046 4773 38080 4807
rect 38046 4705 38080 4739
rect 38130 4705 38164 4739
rect 38214 4773 38248 4807
rect 38214 4705 38248 4739
rect 38298 4705 38332 4739
rect 38382 4773 38416 4807
rect 38382 4705 38416 4739
rect 38466 4705 38500 4739
rect 38550 4773 38584 4807
rect 38550 4705 38584 4739
rect 38634 4705 38668 4739
rect 38718 4773 38752 4807
rect 38718 4705 38752 4739
rect 38802 4705 38836 4739
rect 38886 4773 38920 4807
rect 38886 4705 38920 4739
rect 38970 4705 39004 4739
rect 39054 4773 39088 4807
rect 39054 4705 39088 4739
rect 39138 4773 39172 4807
rect 39138 4705 39172 4739
rect 51010 4775 51044 4809
rect 51010 4707 51044 4741
rect 51094 4775 51128 4809
rect 51094 4707 51128 4741
rect 51178 4707 51212 4741
rect 51262 4775 51296 4809
rect 51262 4707 51296 4741
rect 51346 4707 51380 4741
rect 51430 4775 51464 4809
rect 51430 4707 51464 4741
rect 51514 4707 51548 4741
rect 51598 4775 51632 4809
rect 51598 4707 51632 4741
rect 51682 4707 51716 4741
rect 51766 4775 51800 4809
rect 51766 4707 51800 4741
rect 51850 4707 51884 4741
rect 51934 4775 51968 4809
rect 51934 4707 51968 4741
rect 52018 4707 52052 4741
rect 52102 4775 52136 4809
rect 52102 4707 52136 4741
rect 52186 4707 52220 4741
rect 52270 4775 52304 4809
rect 52270 4707 52304 4741
rect 52354 4775 52388 4809
rect 52354 4707 52388 4741
rect 52892 4773 52926 4807
rect 52892 4705 52926 4739
rect 52976 4773 53010 4807
rect 52976 4705 53010 4739
rect 53060 4705 53094 4739
rect 53144 4773 53178 4807
rect 53144 4705 53178 4739
rect 53228 4705 53262 4739
rect 53312 4773 53346 4807
rect 53312 4705 53346 4739
rect 53396 4705 53430 4739
rect 53480 4773 53514 4807
rect 53480 4705 53514 4739
rect 53564 4705 53598 4739
rect 53648 4773 53682 4807
rect 53648 4705 53682 4739
rect 53732 4705 53766 4739
rect 53816 4773 53850 4807
rect 53816 4705 53850 4739
rect 53900 4705 53934 4739
rect 53984 4773 54018 4807
rect 53984 4705 54018 4739
rect 54068 4705 54102 4739
rect 54152 4773 54186 4807
rect 54152 4705 54186 4739
rect 54236 4773 54270 4807
rect 54236 4705 54270 4739
rect 30072 3630 30106 3664
rect 30156 3638 30190 3672
rect 30240 3630 30274 3664
rect 30324 3638 30358 3672
rect 30408 3631 30442 3665
rect 30603 3698 30637 3732
rect 30603 3630 30637 3664
rect 30687 3698 30721 3732
rect 30687 3630 30721 3664
rect 30771 3630 30805 3664
rect 30855 3698 30889 3732
rect 30855 3630 30889 3664
rect 30939 3630 30973 3664
rect 31023 3698 31057 3732
rect 31023 3630 31057 3664
rect 31107 3630 31141 3664
rect 31191 3698 31225 3732
rect 31191 3630 31225 3664
rect 31275 3630 31309 3664
rect 31359 3698 31393 3732
rect 31359 3630 31393 3664
rect 31443 3630 31477 3664
rect 31527 3698 31561 3732
rect 31527 3630 31561 3664
rect 31611 3630 31645 3664
rect 31695 3698 31729 3732
rect 31695 3630 31729 3664
rect 31779 3630 31813 3664
rect 31863 3698 31897 3732
rect 31863 3630 31897 3664
rect 31947 3698 31981 3732
rect 31947 3630 31981 3664
rect 43429 3482 43463 3516
rect 43429 3414 43463 3448
rect 43513 3482 43547 3516
rect 43513 3414 43547 3448
rect 43597 3414 43631 3448
rect 43681 3482 43715 3516
rect 43681 3414 43715 3448
rect 43765 3414 43799 3448
rect 43849 3482 43883 3516
rect 43849 3414 43883 3448
rect 43933 3414 43967 3448
rect 44017 3482 44051 3516
rect 44017 3414 44051 3448
rect 44101 3414 44135 3448
rect 44185 3482 44219 3516
rect 44185 3414 44219 3448
rect 44269 3414 44303 3448
rect 44353 3482 44387 3516
rect 44353 3414 44387 3448
rect 44437 3414 44471 3448
rect 44521 3482 44555 3516
rect 44521 3414 44555 3448
rect 44605 3414 44639 3448
rect 44689 3482 44723 3516
rect 44689 3414 44723 3448
rect 44773 3482 44807 3516
rect 44773 3414 44807 3448
rect 45359 3482 45393 3516
rect 45359 3414 45393 3448
rect 45443 3482 45477 3516
rect 45443 3414 45477 3448
rect 45527 3414 45561 3448
rect 45611 3482 45645 3516
rect 45611 3414 45645 3448
rect 45695 3414 45729 3448
rect 45779 3482 45813 3516
rect 45779 3414 45813 3448
rect 45863 3414 45897 3448
rect 45947 3482 45981 3516
rect 45947 3414 45981 3448
rect 46031 3414 46065 3448
rect 46115 3482 46149 3516
rect 46115 3414 46149 3448
rect 46199 3414 46233 3448
rect 46283 3482 46317 3516
rect 46283 3414 46317 3448
rect 46367 3414 46401 3448
rect 46451 3482 46485 3516
rect 46451 3414 46485 3448
rect 46535 3414 46569 3448
rect 46619 3482 46653 3516
rect 46619 3414 46653 3448
rect 46703 3482 46737 3516
rect 46703 3414 46737 3448
rect 13287 3322 13321 3356
rect 13287 3254 13321 3288
rect 13371 3322 13405 3356
rect 13371 3254 13405 3288
rect 13455 3254 13489 3288
rect 13539 3322 13573 3356
rect 13539 3254 13573 3288
rect 13623 3254 13657 3288
rect 13707 3322 13741 3356
rect 13707 3254 13741 3288
rect 13791 3254 13825 3288
rect 13875 3322 13909 3356
rect 13875 3254 13909 3288
rect 13959 3254 13993 3288
rect 14043 3322 14077 3356
rect 14043 3254 14077 3288
rect 14127 3254 14161 3288
rect 14211 3322 14245 3356
rect 14211 3254 14245 3288
rect 14295 3254 14329 3288
rect 14379 3322 14413 3356
rect 14379 3254 14413 3288
rect 14463 3254 14497 3288
rect 14547 3322 14581 3356
rect 14547 3254 14581 3288
rect 14631 3322 14665 3356
rect 14631 3254 14665 3288
rect 15217 3322 15251 3356
rect 15217 3254 15251 3288
rect 15301 3322 15335 3356
rect 15301 3254 15335 3288
rect 15385 3254 15419 3288
rect 15469 3322 15503 3356
rect 15469 3254 15503 3288
rect 15553 3254 15587 3288
rect 15637 3322 15671 3356
rect 15637 3254 15671 3288
rect 15721 3254 15755 3288
rect 15805 3322 15839 3356
rect 15805 3254 15839 3288
rect 15889 3254 15923 3288
rect 15973 3322 16007 3356
rect 15973 3254 16007 3288
rect 16057 3254 16091 3288
rect 16141 3322 16175 3356
rect 16141 3254 16175 3288
rect 16225 3254 16259 3288
rect 16309 3322 16343 3356
rect 16309 3254 16343 3288
rect 16393 3254 16427 3288
rect 16477 3322 16511 3356
rect 16477 3254 16511 3288
rect 16561 3322 16595 3356
rect 16561 3254 16595 3288
rect 5712 2701 5746 2735
rect 5712 2633 5746 2667
rect 5796 2701 5830 2735
rect 5796 2633 5830 2667
rect 5880 2701 5914 2735
rect 5964 2701 5998 2735
rect 5964 2633 5998 2667
rect 6048 2701 6082 2735
rect 6132 2701 6166 2735
rect 6132 2633 6166 2667
rect 6216 2701 6250 2735
rect 6300 2701 6334 2735
rect 6300 2633 6334 2667
rect 6384 2701 6418 2735
rect 6468 2701 6502 2735
rect 6468 2633 6502 2667
rect 6552 2701 6586 2735
rect 6636 2701 6670 2735
rect 6636 2633 6670 2667
rect 6720 2701 6754 2735
rect 6804 2701 6838 2735
rect 6804 2633 6838 2667
rect 6888 2701 6922 2735
rect 6972 2701 7006 2735
rect 6972 2633 7006 2667
rect 7056 2701 7090 2735
rect 7056 2633 7090 2667
rect 7594 2699 7628 2733
rect 7594 2631 7628 2665
rect 7678 2699 7712 2733
rect 7678 2631 7712 2665
rect 7762 2699 7796 2733
rect 7846 2699 7880 2733
rect 7846 2631 7880 2665
rect 7930 2699 7964 2733
rect 8014 2699 8048 2733
rect 8014 2631 8048 2665
rect 8098 2699 8132 2733
rect 8182 2699 8216 2733
rect 8182 2631 8216 2665
rect 8266 2699 8300 2733
rect 8350 2699 8384 2733
rect 8350 2631 8384 2665
rect 8434 2699 8468 2733
rect 8518 2699 8552 2733
rect 8518 2631 8552 2665
rect 8602 2699 8636 2733
rect 8686 2699 8720 2733
rect 8686 2631 8720 2665
rect 8770 2699 8804 2733
rect 8854 2699 8888 2733
rect 8854 2631 8888 2665
rect 8938 2699 8972 2733
rect 8938 2631 8972 2665
rect 20810 2701 20844 2735
rect 20810 2633 20844 2667
rect 20894 2701 20928 2735
rect 20894 2633 20928 2667
rect 20978 2701 21012 2735
rect 21062 2701 21096 2735
rect 21062 2633 21096 2667
rect 21146 2701 21180 2735
rect 21230 2701 21264 2735
rect 21230 2633 21264 2667
rect 21314 2701 21348 2735
rect 21398 2701 21432 2735
rect 21398 2633 21432 2667
rect 21482 2701 21516 2735
rect 21566 2701 21600 2735
rect 21566 2633 21600 2667
rect 21650 2701 21684 2735
rect 21734 2701 21768 2735
rect 21734 2633 21768 2667
rect 21818 2701 21852 2735
rect 21902 2701 21936 2735
rect 21902 2633 21936 2667
rect 21986 2701 22020 2735
rect 22070 2701 22104 2735
rect 22070 2633 22104 2667
rect 22154 2701 22188 2735
rect 22154 2633 22188 2667
rect 22692 2699 22726 2733
rect 22692 2631 22726 2665
rect 22776 2699 22810 2733
rect 22776 2631 22810 2665
rect 22860 2699 22894 2733
rect 22944 2699 22978 2733
rect 22944 2631 22978 2665
rect 23028 2699 23062 2733
rect 23112 2699 23146 2733
rect 23112 2631 23146 2665
rect 23196 2699 23230 2733
rect 23280 2699 23314 2733
rect 23280 2631 23314 2665
rect 23364 2699 23398 2733
rect 23448 2699 23482 2733
rect 23448 2631 23482 2665
rect 23532 2699 23566 2733
rect 23616 2699 23650 2733
rect 23616 2631 23650 2665
rect 23700 2699 23734 2733
rect 23784 2699 23818 2733
rect 23784 2631 23818 2665
rect 23868 2699 23902 2733
rect 23952 2699 23986 2733
rect 23952 2631 23986 2665
rect 24036 2699 24070 2733
rect 24036 2631 24070 2665
rect 35914 2701 35948 2735
rect 35914 2633 35948 2667
rect 35998 2701 36032 2735
rect 35998 2633 36032 2667
rect 36082 2701 36116 2735
rect 36166 2701 36200 2735
rect 36166 2633 36200 2667
rect 36250 2701 36284 2735
rect 36334 2701 36368 2735
rect 36334 2633 36368 2667
rect 36418 2701 36452 2735
rect 36502 2701 36536 2735
rect 36502 2633 36536 2667
rect 36586 2701 36620 2735
rect 36670 2701 36704 2735
rect 36670 2633 36704 2667
rect 36754 2701 36788 2735
rect 36838 2701 36872 2735
rect 36838 2633 36872 2667
rect 36922 2701 36956 2735
rect 37006 2701 37040 2735
rect 37006 2633 37040 2667
rect 37090 2701 37124 2735
rect 37174 2701 37208 2735
rect 37174 2633 37208 2667
rect 37258 2701 37292 2735
rect 37258 2633 37292 2667
rect 37796 2699 37830 2733
rect 37796 2631 37830 2665
rect 37880 2699 37914 2733
rect 37880 2631 37914 2665
rect 37964 2699 37998 2733
rect 38048 2699 38082 2733
rect 38048 2631 38082 2665
rect 38132 2699 38166 2733
rect 38216 2699 38250 2733
rect 38216 2631 38250 2665
rect 38300 2699 38334 2733
rect 38384 2699 38418 2733
rect 38384 2631 38418 2665
rect 38468 2699 38502 2733
rect 38552 2699 38586 2733
rect 38552 2631 38586 2665
rect 38636 2699 38670 2733
rect 38720 2699 38754 2733
rect 38720 2631 38754 2665
rect 38804 2699 38838 2733
rect 38888 2699 38922 2733
rect 38888 2631 38922 2665
rect 38972 2699 39006 2733
rect 39056 2699 39090 2733
rect 39056 2631 39090 2665
rect 39140 2699 39174 2733
rect 39140 2631 39174 2665
rect 51012 2701 51046 2735
rect 51012 2633 51046 2667
rect 51096 2701 51130 2735
rect 51096 2633 51130 2667
rect 51180 2701 51214 2735
rect 51264 2701 51298 2735
rect 51264 2633 51298 2667
rect 51348 2701 51382 2735
rect 51432 2701 51466 2735
rect 51432 2633 51466 2667
rect 51516 2701 51550 2735
rect 51600 2701 51634 2735
rect 51600 2633 51634 2667
rect 51684 2701 51718 2735
rect 51768 2701 51802 2735
rect 51768 2633 51802 2667
rect 51852 2701 51886 2735
rect 51936 2701 51970 2735
rect 51936 2633 51970 2667
rect 52020 2701 52054 2735
rect 52104 2701 52138 2735
rect 52104 2633 52138 2667
rect 52188 2701 52222 2735
rect 52272 2701 52306 2735
rect 52272 2633 52306 2667
rect 52356 2701 52390 2735
rect 52356 2633 52390 2667
rect 52894 2699 52928 2733
rect 52894 2631 52928 2665
rect 52978 2699 53012 2733
rect 52978 2631 53012 2665
rect 53062 2699 53096 2733
rect 53146 2699 53180 2733
rect 53146 2631 53180 2665
rect 53230 2699 53264 2733
rect 53314 2699 53348 2733
rect 53314 2631 53348 2665
rect 53398 2699 53432 2733
rect 53482 2699 53516 2733
rect 53482 2631 53516 2665
rect 53566 2699 53600 2733
rect 53650 2699 53684 2733
rect 53650 2631 53684 2665
rect 53734 2699 53768 2733
rect 53818 2699 53852 2733
rect 53818 2631 53852 2665
rect 53902 2699 53936 2733
rect 53986 2699 54020 2733
rect 53986 2631 54020 2665
rect 54070 2699 54104 2733
rect 54154 2699 54188 2733
rect 54154 2631 54188 2665
rect 54238 2699 54272 2733
rect 54238 2631 54272 2665
rect 253 1755 287 1789
rect 253 1687 287 1721
rect 337 1755 371 1789
rect 337 1687 371 1721
rect 421 1755 455 1789
rect 1067 1755 1101 1789
rect 421 1687 455 1721
rect 1067 1687 1101 1721
rect 1151 1755 1185 1789
rect 1151 1687 1185 1721
rect 1235 1755 1269 1789
rect 1235 1687 1269 1721
rect 2141 1755 2175 1789
rect 2141 1687 2175 1721
rect 2225 1755 2259 1789
rect 2225 1687 2259 1721
rect 2309 1755 2343 1789
rect 2955 1755 2989 1789
rect 2309 1687 2343 1721
rect 2955 1687 2989 1721
rect 3039 1755 3073 1789
rect 3039 1687 3073 1721
rect 3123 1755 3157 1789
rect 3123 1687 3157 1721
rect 4029 1755 4063 1789
rect 4029 1687 4063 1721
rect 4113 1755 4147 1789
rect 4113 1687 4147 1721
rect 4197 1755 4231 1789
rect 4843 1755 4877 1789
rect 4197 1687 4231 1721
rect 4843 1687 4877 1721
rect 4927 1755 4961 1789
rect 4927 1687 4961 1721
rect 5011 1755 5045 1789
rect 5011 1687 5045 1721
rect 5917 1755 5951 1789
rect 5917 1687 5951 1721
rect 6001 1755 6035 1789
rect 6001 1687 6035 1721
rect 6085 1755 6119 1789
rect 6731 1755 6765 1789
rect 6085 1687 6119 1721
rect 6731 1687 6765 1721
rect 6815 1755 6849 1789
rect 6815 1687 6849 1721
rect 6899 1755 6933 1789
rect 6899 1687 6933 1721
rect 7805 1755 7839 1789
rect 7805 1687 7839 1721
rect 7889 1755 7923 1789
rect 7889 1687 7923 1721
rect 7973 1755 8007 1789
rect 8619 1755 8653 1789
rect 7973 1687 8007 1721
rect 8619 1687 8653 1721
rect 8703 1755 8737 1789
rect 8703 1687 8737 1721
rect 8787 1755 8821 1789
rect 8787 1687 8821 1721
rect 9693 1755 9727 1789
rect 9693 1687 9727 1721
rect 9777 1755 9811 1789
rect 9777 1687 9811 1721
rect 9861 1755 9895 1789
rect 10507 1755 10541 1789
rect 9861 1687 9895 1721
rect 10507 1687 10541 1721
rect 10591 1755 10625 1789
rect 10591 1687 10625 1721
rect 10675 1755 10709 1789
rect 10675 1687 10709 1721
rect 11581 1755 11615 1789
rect 11581 1687 11615 1721
rect 11665 1755 11699 1789
rect 11665 1687 11699 1721
rect 11749 1755 11783 1789
rect 12395 1755 12429 1789
rect 11749 1687 11783 1721
rect 12395 1687 12429 1721
rect 12479 1755 12513 1789
rect 12479 1687 12513 1721
rect 12563 1755 12597 1789
rect 12563 1687 12597 1721
rect 13469 1755 13503 1789
rect 13469 1687 13503 1721
rect 13553 1755 13587 1789
rect 13553 1687 13587 1721
rect 13637 1755 13671 1789
rect 14283 1755 14317 1789
rect 13637 1687 13671 1721
rect 14283 1687 14317 1721
rect 14367 1755 14401 1789
rect 14367 1687 14401 1721
rect 14451 1755 14485 1789
rect 14451 1687 14485 1721
rect 15351 1755 15385 1789
rect 15351 1687 15385 1721
rect 15435 1755 15469 1789
rect 15435 1687 15469 1721
rect 15519 1755 15553 1789
rect 16165 1755 16199 1789
rect 15519 1687 15553 1721
rect 16165 1687 16199 1721
rect 16249 1755 16283 1789
rect 16249 1687 16283 1721
rect 16333 1755 16367 1789
rect 16333 1687 16367 1721
rect 17239 1755 17273 1789
rect 17239 1687 17273 1721
rect 17323 1755 17357 1789
rect 17323 1687 17357 1721
rect 17407 1755 17441 1789
rect 18053 1755 18087 1789
rect 17407 1687 17441 1721
rect 18053 1687 18087 1721
rect 18137 1755 18171 1789
rect 18137 1687 18171 1721
rect 18221 1755 18255 1789
rect 18221 1687 18255 1721
rect 19127 1755 19161 1789
rect 19127 1687 19161 1721
rect 19211 1755 19245 1789
rect 19211 1687 19245 1721
rect 19295 1755 19329 1789
rect 19941 1755 19975 1789
rect 19295 1687 19329 1721
rect 19941 1687 19975 1721
rect 20025 1755 20059 1789
rect 20025 1687 20059 1721
rect 20109 1755 20143 1789
rect 20109 1687 20143 1721
rect 21015 1755 21049 1789
rect 21015 1687 21049 1721
rect 21099 1755 21133 1789
rect 21099 1687 21133 1721
rect 21183 1755 21217 1789
rect 21829 1755 21863 1789
rect 21183 1687 21217 1721
rect 21829 1687 21863 1721
rect 21913 1755 21947 1789
rect 21913 1687 21947 1721
rect 21997 1755 22031 1789
rect 21997 1687 22031 1721
rect 22903 1755 22937 1789
rect 22903 1687 22937 1721
rect 22987 1755 23021 1789
rect 22987 1687 23021 1721
rect 23071 1755 23105 1789
rect 23717 1755 23751 1789
rect 23071 1687 23105 1721
rect 23717 1687 23751 1721
rect 23801 1755 23835 1789
rect 23801 1687 23835 1721
rect 23885 1755 23919 1789
rect 23885 1687 23919 1721
rect 24791 1755 24825 1789
rect 24791 1687 24825 1721
rect 24875 1755 24909 1789
rect 24875 1687 24909 1721
rect 24959 1755 24993 1789
rect 25605 1755 25639 1789
rect 24959 1687 24993 1721
rect 25605 1687 25639 1721
rect 25689 1755 25723 1789
rect 25689 1687 25723 1721
rect 25773 1755 25807 1789
rect 25773 1687 25807 1721
rect 26679 1755 26713 1789
rect 26679 1687 26713 1721
rect 26763 1755 26797 1789
rect 26763 1687 26797 1721
rect 26847 1755 26881 1789
rect 27493 1755 27527 1789
rect 26847 1687 26881 1721
rect 27493 1687 27527 1721
rect 27577 1755 27611 1789
rect 27577 1687 27611 1721
rect 27661 1755 27695 1789
rect 27661 1687 27695 1721
rect 28567 1755 28601 1789
rect 28567 1687 28601 1721
rect 28651 1755 28685 1789
rect 28651 1687 28685 1721
rect 28735 1755 28769 1789
rect 29381 1755 29415 1789
rect 28735 1687 28769 1721
rect 29381 1687 29415 1721
rect 29465 1755 29499 1789
rect 29465 1687 29499 1721
rect 29549 1755 29583 1789
rect 29549 1687 29583 1721
rect 30455 1755 30489 1789
rect 30455 1687 30489 1721
rect 30539 1755 30573 1789
rect 30539 1687 30573 1721
rect 30623 1755 30657 1789
rect 31269 1755 31303 1789
rect 30623 1687 30657 1721
rect 31269 1687 31303 1721
rect 31353 1755 31387 1789
rect 31353 1687 31387 1721
rect 31437 1755 31471 1789
rect 31437 1687 31471 1721
rect 32343 1755 32377 1789
rect 32343 1687 32377 1721
rect 32427 1755 32461 1789
rect 32427 1687 32461 1721
rect 32511 1755 32545 1789
rect 33157 1755 33191 1789
rect 32511 1687 32545 1721
rect 33157 1687 33191 1721
rect 33241 1755 33275 1789
rect 33241 1687 33275 1721
rect 33325 1755 33359 1789
rect 33325 1687 33359 1721
rect 34231 1755 34265 1789
rect 34231 1687 34265 1721
rect 34315 1755 34349 1789
rect 34315 1687 34349 1721
rect 34399 1755 34433 1789
rect 35045 1755 35079 1789
rect 34399 1687 34433 1721
rect 35045 1687 35079 1721
rect 35129 1755 35163 1789
rect 35129 1687 35163 1721
rect 35213 1755 35247 1789
rect 35213 1687 35247 1721
rect 36119 1755 36153 1789
rect 36119 1687 36153 1721
rect 36203 1755 36237 1789
rect 36203 1687 36237 1721
rect 36287 1755 36321 1789
rect 36933 1755 36967 1789
rect 36287 1687 36321 1721
rect 36933 1687 36967 1721
rect 37017 1755 37051 1789
rect 37017 1687 37051 1721
rect 37101 1755 37135 1789
rect 37101 1687 37135 1721
rect 38007 1755 38041 1789
rect 38007 1687 38041 1721
rect 38091 1755 38125 1789
rect 38091 1687 38125 1721
rect 38175 1755 38209 1789
rect 38821 1755 38855 1789
rect 38175 1687 38209 1721
rect 38821 1687 38855 1721
rect 38905 1755 38939 1789
rect 38905 1687 38939 1721
rect 38989 1755 39023 1789
rect 38989 1687 39023 1721
rect 39895 1755 39929 1789
rect 39895 1687 39929 1721
rect 39979 1755 40013 1789
rect 39979 1687 40013 1721
rect 40063 1755 40097 1789
rect 40709 1755 40743 1789
rect 40063 1687 40097 1721
rect 40709 1687 40743 1721
rect 40793 1755 40827 1789
rect 40793 1687 40827 1721
rect 40877 1755 40911 1789
rect 40877 1687 40911 1721
rect 41783 1755 41817 1789
rect 41783 1687 41817 1721
rect 41867 1755 41901 1789
rect 41867 1687 41901 1721
rect 41951 1755 41985 1789
rect 42597 1755 42631 1789
rect 41951 1687 41985 1721
rect 42597 1687 42631 1721
rect 42681 1755 42715 1789
rect 42681 1687 42715 1721
rect 42765 1755 42799 1789
rect 42765 1687 42799 1721
rect 43671 1755 43705 1789
rect 43671 1687 43705 1721
rect 43755 1755 43789 1789
rect 43755 1687 43789 1721
rect 43839 1755 43873 1789
rect 44485 1755 44519 1789
rect 43839 1687 43873 1721
rect 44485 1687 44519 1721
rect 44569 1755 44603 1789
rect 44569 1687 44603 1721
rect 44653 1755 44687 1789
rect 44653 1687 44687 1721
rect 45553 1755 45587 1789
rect 45553 1687 45587 1721
rect 45637 1755 45671 1789
rect 45637 1687 45671 1721
rect 45721 1755 45755 1789
rect 46367 1755 46401 1789
rect 45721 1687 45755 1721
rect 46367 1687 46401 1721
rect 46451 1755 46485 1789
rect 46451 1687 46485 1721
rect 46535 1755 46569 1789
rect 46535 1687 46569 1721
rect 47441 1755 47475 1789
rect 47441 1687 47475 1721
rect 47525 1755 47559 1789
rect 47525 1687 47559 1721
rect 47609 1755 47643 1789
rect 48255 1755 48289 1789
rect 47609 1687 47643 1721
rect 48255 1687 48289 1721
rect 48339 1755 48373 1789
rect 48339 1687 48373 1721
rect 48423 1755 48457 1789
rect 48423 1687 48457 1721
rect 49329 1755 49363 1789
rect 49329 1687 49363 1721
rect 49413 1755 49447 1789
rect 49413 1687 49447 1721
rect 49497 1755 49531 1789
rect 50143 1755 50177 1789
rect 49497 1687 49531 1721
rect 50143 1687 50177 1721
rect 50227 1755 50261 1789
rect 50227 1687 50261 1721
rect 50311 1755 50345 1789
rect 50311 1687 50345 1721
rect 51217 1755 51251 1789
rect 51217 1687 51251 1721
rect 51301 1755 51335 1789
rect 51301 1687 51335 1721
rect 51385 1755 51419 1789
rect 52031 1755 52065 1789
rect 51385 1687 51419 1721
rect 52031 1687 52065 1721
rect 52115 1755 52149 1789
rect 52115 1687 52149 1721
rect 52199 1755 52233 1789
rect 52199 1687 52233 1721
rect 53105 1755 53139 1789
rect 53105 1687 53139 1721
rect 53189 1755 53223 1789
rect 53189 1687 53223 1721
rect 53273 1755 53307 1789
rect 53919 1755 53953 1789
rect 53273 1687 53307 1721
rect 53919 1687 53953 1721
rect 54003 1755 54037 1789
rect 54003 1687 54037 1721
rect 54087 1755 54121 1789
rect 54087 1687 54121 1721
rect 54993 1755 55027 1789
rect 54993 1687 55027 1721
rect 55077 1755 55111 1789
rect 55077 1687 55111 1721
rect 55161 1755 55195 1789
rect 55807 1755 55841 1789
rect 55161 1687 55195 1721
rect 55807 1687 55841 1721
rect 55891 1755 55925 1789
rect 55891 1687 55925 1721
rect 55975 1755 56009 1789
rect 55975 1687 56009 1721
rect 56881 1755 56915 1789
rect 56881 1687 56915 1721
rect 56965 1755 56999 1789
rect 56965 1687 56999 1721
rect 57049 1755 57083 1789
rect 57695 1755 57729 1789
rect 57049 1687 57083 1721
rect 57695 1687 57729 1721
rect 57779 1755 57813 1789
rect 57779 1687 57813 1721
rect 57863 1755 57897 1789
rect 57863 1687 57897 1721
rect 58769 1755 58803 1789
rect 58769 1687 58803 1721
rect 58853 1755 58887 1789
rect 58853 1687 58887 1721
rect 58937 1755 58971 1789
rect 59583 1755 59617 1789
rect 58937 1687 58971 1721
rect 59583 1687 59617 1721
rect 59667 1755 59701 1789
rect 59667 1687 59701 1721
rect 59751 1755 59785 1789
rect 59751 1687 59785 1721
rect 622 1510 656 1544
rect 622 1442 656 1476
rect 718 1510 752 1544
rect 718 1442 752 1476
rect 814 1510 848 1544
rect 814 1442 848 1476
rect 2510 1510 2544 1544
rect 2510 1442 2544 1476
rect 2606 1510 2640 1544
rect 2606 1442 2640 1476
rect 2702 1510 2736 1544
rect 2702 1442 2736 1476
rect 4398 1510 4432 1544
rect 4398 1442 4432 1476
rect 4494 1510 4528 1544
rect 4494 1442 4528 1476
rect 4590 1510 4624 1544
rect 4590 1442 4624 1476
rect 6286 1510 6320 1544
rect 6286 1442 6320 1476
rect 6382 1510 6416 1544
rect 6382 1442 6416 1476
rect 6478 1510 6512 1544
rect 6478 1442 6512 1476
rect 8174 1510 8208 1544
rect 8174 1442 8208 1476
rect 8270 1510 8304 1544
rect 8270 1442 8304 1476
rect 8366 1510 8400 1544
rect 8366 1442 8400 1476
rect 10062 1510 10096 1544
rect 10062 1442 10096 1476
rect 10158 1510 10192 1544
rect 10158 1442 10192 1476
rect 10254 1510 10288 1544
rect 10254 1442 10288 1476
rect 11950 1510 11984 1544
rect 11950 1442 11984 1476
rect 12046 1510 12080 1544
rect 12046 1442 12080 1476
rect 12142 1510 12176 1544
rect 12142 1442 12176 1476
rect 13838 1510 13872 1544
rect 13838 1442 13872 1476
rect 13934 1510 13968 1544
rect 13934 1442 13968 1476
rect 14030 1510 14064 1544
rect 14030 1442 14064 1476
rect 15720 1510 15754 1544
rect 15720 1442 15754 1476
rect 15816 1510 15850 1544
rect 15816 1442 15850 1476
rect 15912 1510 15946 1544
rect 15912 1442 15946 1476
rect 17608 1510 17642 1544
rect 17608 1442 17642 1476
rect 17704 1510 17738 1544
rect 17704 1442 17738 1476
rect 17800 1510 17834 1544
rect 17800 1442 17834 1476
rect 19496 1510 19530 1544
rect 19496 1442 19530 1476
rect 19592 1510 19626 1544
rect 19592 1442 19626 1476
rect 19688 1510 19722 1544
rect 19688 1442 19722 1476
rect 21384 1510 21418 1544
rect 21384 1442 21418 1476
rect 21480 1510 21514 1544
rect 21480 1442 21514 1476
rect 21576 1510 21610 1544
rect 21576 1442 21610 1476
rect 23272 1510 23306 1544
rect 23272 1442 23306 1476
rect 23368 1510 23402 1544
rect 23368 1442 23402 1476
rect 23464 1510 23498 1544
rect 23464 1442 23498 1476
rect 25160 1510 25194 1544
rect 25160 1442 25194 1476
rect 25256 1510 25290 1544
rect 25256 1442 25290 1476
rect 25352 1510 25386 1544
rect 25352 1442 25386 1476
rect 27048 1510 27082 1544
rect 27048 1442 27082 1476
rect 27144 1510 27178 1544
rect 27144 1442 27178 1476
rect 27240 1510 27274 1544
rect 27240 1442 27274 1476
rect 28936 1510 28970 1544
rect 28936 1442 28970 1476
rect 29032 1510 29066 1544
rect 29032 1442 29066 1476
rect 29128 1510 29162 1544
rect 29128 1442 29162 1476
rect 30824 1510 30858 1544
rect 30824 1442 30858 1476
rect 30920 1510 30954 1544
rect 30920 1442 30954 1476
rect 31016 1510 31050 1544
rect 31016 1442 31050 1476
rect 32712 1510 32746 1544
rect 32712 1442 32746 1476
rect 32808 1510 32842 1544
rect 32808 1442 32842 1476
rect 32904 1510 32938 1544
rect 32904 1442 32938 1476
rect 34600 1510 34634 1544
rect 34600 1442 34634 1476
rect 34696 1510 34730 1544
rect 34696 1442 34730 1476
rect 34792 1510 34826 1544
rect 34792 1442 34826 1476
rect 36488 1510 36522 1544
rect 36488 1442 36522 1476
rect 36584 1510 36618 1544
rect 36584 1442 36618 1476
rect 36680 1510 36714 1544
rect 36680 1442 36714 1476
rect 38376 1510 38410 1544
rect 38376 1442 38410 1476
rect 38472 1510 38506 1544
rect 38472 1442 38506 1476
rect 38568 1510 38602 1544
rect 38568 1442 38602 1476
rect 40264 1510 40298 1544
rect 40264 1442 40298 1476
rect 40360 1510 40394 1544
rect 40360 1442 40394 1476
rect 40456 1510 40490 1544
rect 40456 1442 40490 1476
rect 42152 1510 42186 1544
rect 42152 1442 42186 1476
rect 42248 1510 42282 1544
rect 42248 1442 42282 1476
rect 42344 1510 42378 1544
rect 42344 1442 42378 1476
rect 44040 1510 44074 1544
rect 44040 1442 44074 1476
rect 44136 1510 44170 1544
rect 44136 1442 44170 1476
rect 44232 1510 44266 1544
rect 44232 1442 44266 1476
rect 45922 1510 45956 1544
rect 45922 1442 45956 1476
rect 46018 1510 46052 1544
rect 46018 1442 46052 1476
rect 46114 1510 46148 1544
rect 46114 1442 46148 1476
rect 47810 1510 47844 1544
rect 47810 1442 47844 1476
rect 47906 1510 47940 1544
rect 47906 1442 47940 1476
rect 48002 1510 48036 1544
rect 48002 1442 48036 1476
rect 49698 1510 49732 1544
rect 49698 1442 49732 1476
rect 49794 1510 49828 1544
rect 49794 1442 49828 1476
rect 49890 1510 49924 1544
rect 49890 1442 49924 1476
rect 51586 1510 51620 1544
rect 51586 1442 51620 1476
rect 51682 1510 51716 1544
rect 51682 1442 51716 1476
rect 51778 1510 51812 1544
rect 51778 1442 51812 1476
rect 53474 1510 53508 1544
rect 53474 1442 53508 1476
rect 53570 1510 53604 1544
rect 53570 1442 53604 1476
rect 53666 1510 53700 1544
rect 53666 1442 53700 1476
rect 55362 1510 55396 1544
rect 55362 1442 55396 1476
rect 55458 1510 55492 1544
rect 55458 1442 55492 1476
rect 55554 1510 55588 1544
rect 55554 1442 55588 1476
rect 57250 1510 57284 1544
rect 57250 1442 57284 1476
rect 57346 1510 57380 1544
rect 57346 1442 57380 1476
rect 57442 1510 57476 1544
rect 57442 1442 57476 1476
rect 59138 1510 59172 1544
rect 59138 1442 59172 1476
rect 59234 1510 59268 1544
rect 59234 1442 59268 1476
rect 59330 1510 59364 1544
rect 59330 1442 59364 1476
rect 116 703 150 737
rect 116 635 150 669
rect 200 703 234 737
rect 1312 711 1346 745
rect 200 635 234 669
rect 1312 643 1346 677
rect 1396 711 1430 745
rect 1396 643 1430 677
rect 1617 650 1651 684
rect 1703 637 1737 671
rect 1789 667 1823 701
rect 2004 703 2038 737
rect 2004 635 2038 669
rect 2088 703 2122 737
rect 3200 711 3234 745
rect 2088 635 2122 669
rect 3200 643 3234 677
rect 3284 711 3318 745
rect 3284 643 3318 677
rect 3505 650 3539 684
rect 3591 637 3625 671
rect 3677 667 3711 701
rect 3892 703 3926 737
rect 3892 635 3926 669
rect 3976 703 4010 737
rect 5088 711 5122 745
rect 3976 635 4010 669
rect 5088 643 5122 677
rect 5172 711 5206 745
rect 5172 643 5206 677
rect 5393 650 5427 684
rect 5479 637 5513 671
rect 5565 667 5599 701
rect 5780 703 5814 737
rect 5780 635 5814 669
rect 5864 703 5898 737
rect 6976 711 7010 745
rect 5864 635 5898 669
rect 6976 643 7010 677
rect 7060 711 7094 745
rect 7060 643 7094 677
rect 7281 650 7315 684
rect 7367 637 7401 671
rect 7453 667 7487 701
rect 7668 703 7702 737
rect 7668 635 7702 669
rect 7752 703 7786 737
rect 8864 711 8898 745
rect 7752 635 7786 669
rect 8864 643 8898 677
rect 8948 711 8982 745
rect 8948 643 8982 677
rect 9169 650 9203 684
rect 9255 637 9289 671
rect 9341 667 9375 701
rect 9556 703 9590 737
rect 9556 635 9590 669
rect 9640 703 9674 737
rect 10752 711 10786 745
rect 9640 635 9674 669
rect 10752 643 10786 677
rect 10836 711 10870 745
rect 10836 643 10870 677
rect 11057 650 11091 684
rect 11143 637 11177 671
rect 11229 667 11263 701
rect 11444 703 11478 737
rect 11444 635 11478 669
rect 11528 703 11562 737
rect 12640 711 12674 745
rect 11528 635 11562 669
rect 12640 643 12674 677
rect 12724 711 12758 745
rect 12724 643 12758 677
rect 12945 650 12979 684
rect 13031 637 13065 671
rect 13117 667 13151 701
rect 13332 703 13366 737
rect 13332 635 13366 669
rect 13416 703 13450 737
rect 14528 711 14562 745
rect 13416 635 13450 669
rect 14528 643 14562 677
rect 14612 711 14646 745
rect 14612 643 14646 677
rect 14833 650 14867 684
rect 14919 637 14953 671
rect 15005 667 15039 701
rect 15214 703 15248 737
rect 15214 635 15248 669
rect 15298 703 15332 737
rect 16410 711 16444 745
rect 15298 635 15332 669
rect 16410 643 16444 677
rect 16494 711 16528 745
rect 16494 643 16528 677
rect 16715 650 16749 684
rect 16801 637 16835 671
rect 16887 667 16921 701
rect 17102 703 17136 737
rect 17102 635 17136 669
rect 17186 703 17220 737
rect 18298 711 18332 745
rect 17186 635 17220 669
rect 18298 643 18332 677
rect 18382 711 18416 745
rect 18382 643 18416 677
rect 18603 650 18637 684
rect 18689 637 18723 671
rect 18775 667 18809 701
rect 18990 703 19024 737
rect 18990 635 19024 669
rect 19074 703 19108 737
rect 20186 711 20220 745
rect 19074 635 19108 669
rect 20186 643 20220 677
rect 20270 711 20304 745
rect 20270 643 20304 677
rect 20491 650 20525 684
rect 20577 637 20611 671
rect 20663 667 20697 701
rect 20878 703 20912 737
rect 20878 635 20912 669
rect 20962 703 20996 737
rect 22074 711 22108 745
rect 20962 635 20996 669
rect 22074 643 22108 677
rect 22158 711 22192 745
rect 22158 643 22192 677
rect 22379 650 22413 684
rect 22465 637 22499 671
rect 22551 667 22585 701
rect 22766 703 22800 737
rect 22766 635 22800 669
rect 22850 703 22884 737
rect 23962 711 23996 745
rect 22850 635 22884 669
rect 23962 643 23996 677
rect 24046 711 24080 745
rect 24046 643 24080 677
rect 24267 650 24301 684
rect 24353 637 24387 671
rect 24439 667 24473 701
rect 24654 703 24688 737
rect 24654 635 24688 669
rect 24738 703 24772 737
rect 25850 711 25884 745
rect 24738 635 24772 669
rect 25850 643 25884 677
rect 25934 711 25968 745
rect 25934 643 25968 677
rect 26155 650 26189 684
rect 26241 637 26275 671
rect 26327 667 26361 701
rect 26542 703 26576 737
rect 26542 635 26576 669
rect 26626 703 26660 737
rect 27738 711 27772 745
rect 26626 635 26660 669
rect 27738 643 27772 677
rect 27822 711 27856 745
rect 27822 643 27856 677
rect 28043 650 28077 684
rect 28129 637 28163 671
rect 28215 667 28249 701
rect 28430 703 28464 737
rect 28430 635 28464 669
rect 28514 703 28548 737
rect 29626 711 29660 745
rect 28514 635 28548 669
rect 29626 643 29660 677
rect 29710 711 29744 745
rect 29710 643 29744 677
rect 29931 650 29965 684
rect 30017 637 30051 671
rect 30103 667 30137 701
rect 30318 703 30352 737
rect 30318 635 30352 669
rect 30402 703 30436 737
rect 31514 711 31548 745
rect 30402 635 30436 669
rect 31514 643 31548 677
rect 31598 711 31632 745
rect 31598 643 31632 677
rect 31819 650 31853 684
rect 31905 637 31939 671
rect 31991 667 32025 701
rect 32206 703 32240 737
rect 32206 635 32240 669
rect 32290 703 32324 737
rect 33402 711 33436 745
rect 32290 635 32324 669
rect 33402 643 33436 677
rect 33486 711 33520 745
rect 33486 643 33520 677
rect 33707 650 33741 684
rect 33793 637 33827 671
rect 33879 667 33913 701
rect 34094 703 34128 737
rect 34094 635 34128 669
rect 34178 703 34212 737
rect 35290 711 35324 745
rect 34178 635 34212 669
rect 35290 643 35324 677
rect 35374 711 35408 745
rect 35374 643 35408 677
rect 35595 650 35629 684
rect 35681 637 35715 671
rect 35767 667 35801 701
rect 35982 703 36016 737
rect 35982 635 36016 669
rect 36066 703 36100 737
rect 37178 711 37212 745
rect 36066 635 36100 669
rect 37178 643 37212 677
rect 37262 711 37296 745
rect 37262 643 37296 677
rect 37483 650 37517 684
rect 37569 637 37603 671
rect 37655 667 37689 701
rect 37870 703 37904 737
rect 37870 635 37904 669
rect 37954 703 37988 737
rect 39066 711 39100 745
rect 37954 635 37988 669
rect 39066 643 39100 677
rect 39150 711 39184 745
rect 39150 643 39184 677
rect 39371 650 39405 684
rect 39457 637 39491 671
rect 39543 667 39577 701
rect 39758 703 39792 737
rect 39758 635 39792 669
rect 39842 703 39876 737
rect 40954 711 40988 745
rect 39842 635 39876 669
rect 40954 643 40988 677
rect 41038 711 41072 745
rect 41038 643 41072 677
rect 41259 650 41293 684
rect 41345 637 41379 671
rect 41431 667 41465 701
rect 41646 703 41680 737
rect 41646 635 41680 669
rect 41730 703 41764 737
rect 42842 711 42876 745
rect 41730 635 41764 669
rect 42842 643 42876 677
rect 42926 711 42960 745
rect 42926 643 42960 677
rect 43147 650 43181 684
rect 43233 637 43267 671
rect 43319 667 43353 701
rect 43534 703 43568 737
rect 43534 635 43568 669
rect 43618 703 43652 737
rect 44730 711 44764 745
rect 43618 635 43652 669
rect 44730 643 44764 677
rect 44814 711 44848 745
rect 44814 643 44848 677
rect 45035 650 45069 684
rect 45121 637 45155 671
rect 45207 667 45241 701
rect 45416 703 45450 737
rect 45416 635 45450 669
rect 45500 703 45534 737
rect 46612 711 46646 745
rect 45500 635 45534 669
rect 46612 643 46646 677
rect 46696 711 46730 745
rect 46696 643 46730 677
rect 46917 650 46951 684
rect 47003 637 47037 671
rect 47089 667 47123 701
rect 47304 703 47338 737
rect 47304 635 47338 669
rect 47388 703 47422 737
rect 48500 711 48534 745
rect 47388 635 47422 669
rect 48500 643 48534 677
rect 48584 711 48618 745
rect 48584 643 48618 677
rect 48805 650 48839 684
rect 48891 637 48925 671
rect 48977 667 49011 701
rect 49192 703 49226 737
rect 49192 635 49226 669
rect 49276 703 49310 737
rect 50388 711 50422 745
rect 49276 635 49310 669
rect 50388 643 50422 677
rect 50472 711 50506 745
rect 50472 643 50506 677
rect 50693 650 50727 684
rect 50779 637 50813 671
rect 50865 667 50899 701
rect 51080 703 51114 737
rect 51080 635 51114 669
rect 51164 703 51198 737
rect 52276 711 52310 745
rect 51164 635 51198 669
rect 52276 643 52310 677
rect 52360 711 52394 745
rect 52360 643 52394 677
rect 52581 650 52615 684
rect 52667 637 52701 671
rect 52753 667 52787 701
rect 52968 703 53002 737
rect 52968 635 53002 669
rect 53052 703 53086 737
rect 54164 711 54198 745
rect 53052 635 53086 669
rect 54164 643 54198 677
rect 54248 711 54282 745
rect 54248 643 54282 677
rect 54469 650 54503 684
rect 54555 637 54589 671
rect 54641 667 54675 701
rect 54856 703 54890 737
rect 54856 635 54890 669
rect 54940 703 54974 737
rect 56052 711 56086 745
rect 54940 635 54974 669
rect 56052 643 56086 677
rect 56136 711 56170 745
rect 56136 643 56170 677
rect 56357 650 56391 684
rect 56443 637 56477 671
rect 56529 667 56563 701
rect 56744 703 56778 737
rect 56744 635 56778 669
rect 56828 703 56862 737
rect 57940 711 57974 745
rect 56828 635 56862 669
rect 57940 643 57974 677
rect 58024 711 58058 745
rect 58024 643 58058 677
rect 58245 650 58279 684
rect 58331 637 58365 671
rect 58417 667 58451 701
rect 58632 703 58666 737
rect 58632 635 58666 669
rect 58716 703 58750 737
rect 59828 711 59862 745
rect 58716 635 58750 669
rect 59828 643 59862 677
rect 59912 711 59946 745
rect 59912 643 59946 677
rect 60133 650 60167 684
rect 60219 637 60253 671
rect 60305 667 60339 701
rect 620 454 654 488
rect 620 386 654 420
rect 716 454 750 488
rect 716 386 750 420
rect 812 454 846 488
rect 812 386 846 420
rect 2508 454 2542 488
rect 2508 386 2542 420
rect 2604 454 2638 488
rect 2604 386 2638 420
rect 2700 454 2734 488
rect 2700 386 2734 420
rect 4396 454 4430 488
rect 4396 386 4430 420
rect 4492 454 4526 488
rect 4492 386 4526 420
rect 4588 454 4622 488
rect 4588 386 4622 420
rect 6284 454 6318 488
rect 6284 386 6318 420
rect 6380 454 6414 488
rect 6380 386 6414 420
rect 6476 454 6510 488
rect 6476 386 6510 420
rect 8172 454 8206 488
rect 8172 386 8206 420
rect 8268 454 8302 488
rect 8268 386 8302 420
rect 8364 454 8398 488
rect 8364 386 8398 420
rect 10060 454 10094 488
rect 10060 386 10094 420
rect 10156 454 10190 488
rect 10156 386 10190 420
rect 10252 454 10286 488
rect 10252 386 10286 420
rect 11948 454 11982 488
rect 11948 386 11982 420
rect 12044 454 12078 488
rect 12044 386 12078 420
rect 12140 454 12174 488
rect 12140 386 12174 420
rect 13836 454 13870 488
rect 13836 386 13870 420
rect 13932 454 13966 488
rect 13932 386 13966 420
rect 14028 454 14062 488
rect 14028 386 14062 420
rect 15718 454 15752 488
rect 15718 386 15752 420
rect 15814 454 15848 488
rect 15814 386 15848 420
rect 15910 454 15944 488
rect 15910 386 15944 420
rect 17606 454 17640 488
rect 17606 386 17640 420
rect 17702 454 17736 488
rect 17702 386 17736 420
rect 17798 454 17832 488
rect 17798 386 17832 420
rect 19494 454 19528 488
rect 19494 386 19528 420
rect 19590 454 19624 488
rect 19590 386 19624 420
rect 19686 454 19720 488
rect 19686 386 19720 420
rect 21382 454 21416 488
rect 21382 386 21416 420
rect 21478 454 21512 488
rect 21478 386 21512 420
rect 21574 454 21608 488
rect 21574 386 21608 420
rect 23270 454 23304 488
rect 23270 386 23304 420
rect 23366 454 23400 488
rect 23366 386 23400 420
rect 23462 454 23496 488
rect 23462 386 23496 420
rect 25158 454 25192 488
rect 25158 386 25192 420
rect 25254 454 25288 488
rect 25254 386 25288 420
rect 25350 454 25384 488
rect 25350 386 25384 420
rect 27046 454 27080 488
rect 27046 386 27080 420
rect 27142 454 27176 488
rect 27142 386 27176 420
rect 27238 454 27272 488
rect 27238 386 27272 420
rect 28934 454 28968 488
rect 28934 386 28968 420
rect 29030 454 29064 488
rect 29030 386 29064 420
rect 29126 454 29160 488
rect 29126 386 29160 420
rect 30822 454 30856 488
rect 30822 386 30856 420
rect 30918 454 30952 488
rect 30918 386 30952 420
rect 31014 454 31048 488
rect 31014 386 31048 420
rect 32710 454 32744 488
rect 32710 386 32744 420
rect 32806 454 32840 488
rect 32806 386 32840 420
rect 32902 454 32936 488
rect 32902 386 32936 420
rect 34598 454 34632 488
rect 34598 386 34632 420
rect 34694 454 34728 488
rect 34694 386 34728 420
rect 34790 454 34824 488
rect 34790 386 34824 420
rect 36486 454 36520 488
rect 36486 386 36520 420
rect 36582 454 36616 488
rect 36582 386 36616 420
rect 36678 454 36712 488
rect 36678 386 36712 420
rect 38374 454 38408 488
rect 38374 386 38408 420
rect 38470 454 38504 488
rect 38470 386 38504 420
rect 38566 454 38600 488
rect 38566 386 38600 420
rect 40262 454 40296 488
rect 40262 386 40296 420
rect 40358 454 40392 488
rect 40358 386 40392 420
rect 40454 454 40488 488
rect 40454 386 40488 420
rect 42150 454 42184 488
rect 42150 386 42184 420
rect 42246 454 42280 488
rect 42246 386 42280 420
rect 42342 454 42376 488
rect 42342 386 42376 420
rect 44038 454 44072 488
rect 44038 386 44072 420
rect 44134 454 44168 488
rect 44134 386 44168 420
rect 44230 454 44264 488
rect 44230 386 44264 420
rect 45920 454 45954 488
rect 45920 386 45954 420
rect 46016 454 46050 488
rect 46016 386 46050 420
rect 46112 454 46146 488
rect 46112 386 46146 420
rect 47808 454 47842 488
rect 47808 386 47842 420
rect 47904 454 47938 488
rect 47904 386 47938 420
rect 48000 454 48034 488
rect 48000 386 48034 420
rect 49696 454 49730 488
rect 49696 386 49730 420
rect 49792 454 49826 488
rect 49792 386 49826 420
rect 49888 454 49922 488
rect 49888 386 49922 420
rect 51584 454 51618 488
rect 51584 386 51618 420
rect 51680 454 51714 488
rect 51680 386 51714 420
rect 51776 454 51810 488
rect 51776 386 51810 420
rect 53472 454 53506 488
rect 53472 386 53506 420
rect 53568 454 53602 488
rect 53568 386 53602 420
rect 53664 454 53698 488
rect 53664 386 53698 420
rect 55360 454 55394 488
rect 55360 386 55394 420
rect 55456 454 55490 488
rect 55456 386 55490 420
rect 55552 454 55586 488
rect 55552 386 55586 420
rect 57248 454 57282 488
rect 57248 386 57282 420
rect 57344 454 57378 488
rect 57344 386 57378 420
rect 57440 454 57474 488
rect 57440 386 57474 420
rect 59136 454 59170 488
rect 59136 386 59170 420
rect 59232 454 59266 488
rect 59232 386 59266 420
rect 59328 454 59362 488
rect 59328 386 59362 420
<< pdiffc >>
rect 636 6689 670 6723
rect 636 6621 670 6655
rect -357 6466 -323 6500
rect -357 6385 -323 6419
rect -271 6453 -237 6487
rect -271 6385 -237 6419
rect -185 6453 -151 6487
rect -185 6385 -151 6419
rect 36 6511 70 6545
rect 36 6443 70 6477
rect 36 6375 70 6409
rect 120 6511 154 6545
rect 120 6443 154 6477
rect 120 6375 154 6409
rect 310 6529 344 6563
rect 310 6461 344 6495
rect 310 6393 344 6427
rect 398 6529 432 6563
rect 636 6553 670 6587
rect 732 6689 766 6723
rect 732 6621 766 6655
rect 732 6553 766 6587
rect 828 6689 862 6723
rect 828 6621 862 6655
rect 2524 6689 2558 6723
rect 828 6553 862 6587
rect 398 6461 432 6495
rect 956 6529 990 6563
rect 956 6461 990 6495
rect 398 6393 432 6427
rect 956 6393 990 6427
rect 1044 6529 1078 6563
rect 1044 6461 1078 6495
rect 1044 6393 1078 6427
rect 1232 6519 1266 6553
rect 1232 6451 1266 6485
rect 1232 6383 1266 6417
rect 1316 6519 1350 6553
rect 2524 6621 2558 6655
rect 1316 6451 1350 6485
rect 1316 6383 1350 6417
rect 1531 6466 1565 6500
rect 1531 6385 1565 6419
rect 1617 6453 1651 6487
rect 1617 6385 1651 6419
rect 1703 6453 1737 6487
rect 1703 6385 1737 6419
rect 1924 6511 1958 6545
rect 1924 6443 1958 6477
rect 1924 6375 1958 6409
rect 2008 6511 2042 6545
rect 2008 6443 2042 6477
rect 2008 6375 2042 6409
rect 2198 6529 2232 6563
rect 2198 6461 2232 6495
rect 2198 6393 2232 6427
rect 2286 6529 2320 6563
rect 2524 6553 2558 6587
rect 2620 6689 2654 6723
rect 2620 6621 2654 6655
rect 2620 6553 2654 6587
rect 2716 6689 2750 6723
rect 2716 6621 2750 6655
rect 4412 6689 4446 6723
rect 2716 6553 2750 6587
rect 2286 6461 2320 6495
rect 2844 6529 2878 6563
rect 2844 6461 2878 6495
rect 2286 6393 2320 6427
rect 2844 6393 2878 6427
rect 2932 6529 2966 6563
rect 2932 6461 2966 6495
rect 2932 6393 2966 6427
rect 3120 6519 3154 6553
rect 3120 6451 3154 6485
rect 3120 6383 3154 6417
rect 3204 6519 3238 6553
rect 4412 6621 4446 6655
rect 3204 6451 3238 6485
rect 3204 6383 3238 6417
rect 3419 6466 3453 6500
rect 3419 6385 3453 6419
rect 3505 6453 3539 6487
rect 3505 6385 3539 6419
rect 3591 6453 3625 6487
rect 3591 6385 3625 6419
rect 3812 6511 3846 6545
rect 3812 6443 3846 6477
rect 3812 6375 3846 6409
rect 3896 6511 3930 6545
rect 3896 6443 3930 6477
rect 3896 6375 3930 6409
rect 4086 6529 4120 6563
rect 4086 6461 4120 6495
rect 4086 6393 4120 6427
rect 4174 6529 4208 6563
rect 4412 6553 4446 6587
rect 4508 6689 4542 6723
rect 4508 6621 4542 6655
rect 4508 6553 4542 6587
rect 4604 6689 4638 6723
rect 4604 6621 4638 6655
rect 6300 6689 6334 6723
rect 4604 6553 4638 6587
rect 4174 6461 4208 6495
rect 4732 6529 4766 6563
rect 4732 6461 4766 6495
rect 4174 6393 4208 6427
rect 4732 6393 4766 6427
rect 4820 6529 4854 6563
rect 4820 6461 4854 6495
rect 4820 6393 4854 6427
rect 5008 6519 5042 6553
rect 5008 6451 5042 6485
rect 5008 6383 5042 6417
rect 5092 6519 5126 6553
rect 6300 6621 6334 6655
rect 5092 6451 5126 6485
rect 5092 6383 5126 6417
rect 5307 6466 5341 6500
rect 5307 6385 5341 6419
rect 5393 6453 5427 6487
rect 5393 6385 5427 6419
rect 5479 6453 5513 6487
rect 5479 6385 5513 6419
rect 5700 6511 5734 6545
rect 5700 6443 5734 6477
rect 5700 6375 5734 6409
rect 5784 6511 5818 6545
rect 5784 6443 5818 6477
rect 5784 6375 5818 6409
rect 5974 6529 6008 6563
rect 5974 6461 6008 6495
rect 5974 6393 6008 6427
rect 6062 6529 6096 6563
rect 6300 6553 6334 6587
rect 6396 6689 6430 6723
rect 6396 6621 6430 6655
rect 6396 6553 6430 6587
rect 6492 6689 6526 6723
rect 6492 6621 6526 6655
rect 8188 6689 8222 6723
rect 6492 6553 6526 6587
rect 6062 6461 6096 6495
rect 6620 6529 6654 6563
rect 6620 6461 6654 6495
rect 6062 6393 6096 6427
rect 6620 6393 6654 6427
rect 6708 6529 6742 6563
rect 6708 6461 6742 6495
rect 6708 6393 6742 6427
rect 6896 6519 6930 6553
rect 6896 6451 6930 6485
rect 6896 6383 6930 6417
rect 6980 6519 7014 6553
rect 8188 6621 8222 6655
rect 6980 6451 7014 6485
rect 6980 6383 7014 6417
rect 7195 6466 7229 6500
rect 7195 6385 7229 6419
rect 7281 6453 7315 6487
rect 7281 6385 7315 6419
rect 7367 6453 7401 6487
rect 7367 6385 7401 6419
rect 7588 6511 7622 6545
rect 7588 6443 7622 6477
rect 7588 6375 7622 6409
rect 7672 6511 7706 6545
rect 7672 6443 7706 6477
rect 7672 6375 7706 6409
rect 7862 6529 7896 6563
rect 7862 6461 7896 6495
rect 7862 6393 7896 6427
rect 7950 6529 7984 6563
rect 8188 6553 8222 6587
rect 8284 6689 8318 6723
rect 8284 6621 8318 6655
rect 8284 6553 8318 6587
rect 8380 6689 8414 6723
rect 8380 6621 8414 6655
rect 10076 6689 10110 6723
rect 8380 6553 8414 6587
rect 7950 6461 7984 6495
rect 8508 6529 8542 6563
rect 8508 6461 8542 6495
rect 7950 6393 7984 6427
rect 8508 6393 8542 6427
rect 8596 6529 8630 6563
rect 8596 6461 8630 6495
rect 8596 6393 8630 6427
rect 8784 6519 8818 6553
rect 8784 6451 8818 6485
rect 8784 6383 8818 6417
rect 8868 6519 8902 6553
rect 10076 6621 10110 6655
rect 8868 6451 8902 6485
rect 8868 6383 8902 6417
rect 9083 6466 9117 6500
rect 9083 6385 9117 6419
rect 9169 6453 9203 6487
rect 9169 6385 9203 6419
rect 9255 6453 9289 6487
rect 9255 6385 9289 6419
rect 9476 6511 9510 6545
rect 9476 6443 9510 6477
rect 9476 6375 9510 6409
rect 9560 6511 9594 6545
rect 9560 6443 9594 6477
rect 9560 6375 9594 6409
rect 9750 6529 9784 6563
rect 9750 6461 9784 6495
rect 9750 6393 9784 6427
rect 9838 6529 9872 6563
rect 10076 6553 10110 6587
rect 10172 6689 10206 6723
rect 10172 6621 10206 6655
rect 10172 6553 10206 6587
rect 10268 6689 10302 6723
rect 10268 6621 10302 6655
rect 11964 6689 11998 6723
rect 10268 6553 10302 6587
rect 9838 6461 9872 6495
rect 10396 6529 10430 6563
rect 10396 6461 10430 6495
rect 9838 6393 9872 6427
rect 10396 6393 10430 6427
rect 10484 6529 10518 6563
rect 10484 6461 10518 6495
rect 10484 6393 10518 6427
rect 10672 6519 10706 6553
rect 10672 6451 10706 6485
rect 10672 6383 10706 6417
rect 10756 6519 10790 6553
rect 11964 6621 11998 6655
rect 10756 6451 10790 6485
rect 10756 6383 10790 6417
rect 10971 6466 11005 6500
rect 10971 6385 11005 6419
rect 11057 6453 11091 6487
rect 11057 6385 11091 6419
rect 11143 6453 11177 6487
rect 11143 6385 11177 6419
rect 11364 6511 11398 6545
rect 11364 6443 11398 6477
rect 11364 6375 11398 6409
rect 11448 6511 11482 6545
rect 11448 6443 11482 6477
rect 11448 6375 11482 6409
rect 11638 6529 11672 6563
rect 11638 6461 11672 6495
rect 11638 6393 11672 6427
rect 11726 6529 11760 6563
rect 11964 6553 11998 6587
rect 12060 6689 12094 6723
rect 12060 6621 12094 6655
rect 12060 6553 12094 6587
rect 12156 6689 12190 6723
rect 12156 6621 12190 6655
rect 13852 6689 13886 6723
rect 12156 6553 12190 6587
rect 11726 6461 11760 6495
rect 12284 6529 12318 6563
rect 12284 6461 12318 6495
rect 11726 6393 11760 6427
rect 12284 6393 12318 6427
rect 12372 6529 12406 6563
rect 12372 6461 12406 6495
rect 12372 6393 12406 6427
rect 12560 6519 12594 6553
rect 12560 6451 12594 6485
rect 12560 6383 12594 6417
rect 12644 6519 12678 6553
rect 13852 6621 13886 6655
rect 12644 6451 12678 6485
rect 12644 6383 12678 6417
rect 12859 6466 12893 6500
rect 12859 6385 12893 6419
rect 12945 6453 12979 6487
rect 12945 6385 12979 6419
rect 13031 6453 13065 6487
rect 13031 6385 13065 6419
rect 13252 6511 13286 6545
rect 13252 6443 13286 6477
rect 13252 6375 13286 6409
rect 13336 6511 13370 6545
rect 13336 6443 13370 6477
rect 13336 6375 13370 6409
rect 13526 6529 13560 6563
rect 13526 6461 13560 6495
rect 13526 6393 13560 6427
rect 13614 6529 13648 6563
rect 13852 6553 13886 6587
rect 13948 6689 13982 6723
rect 13948 6621 13982 6655
rect 13948 6553 13982 6587
rect 14044 6689 14078 6723
rect 14044 6621 14078 6655
rect 15734 6689 15768 6723
rect 14044 6553 14078 6587
rect 13614 6461 13648 6495
rect 14172 6529 14206 6563
rect 14172 6461 14206 6495
rect 13614 6393 13648 6427
rect 14172 6393 14206 6427
rect 14260 6529 14294 6563
rect 14260 6461 14294 6495
rect 14260 6393 14294 6427
rect 14448 6519 14482 6553
rect 14448 6451 14482 6485
rect 14448 6383 14482 6417
rect 14532 6519 14566 6553
rect 15734 6621 15768 6655
rect 14532 6451 14566 6485
rect 14532 6383 14566 6417
rect 14741 6466 14775 6500
rect 14741 6385 14775 6419
rect 14827 6453 14861 6487
rect 14827 6385 14861 6419
rect 14913 6453 14947 6487
rect 14913 6385 14947 6419
rect 15134 6511 15168 6545
rect 15134 6443 15168 6477
rect 15134 6375 15168 6409
rect 15218 6511 15252 6545
rect 15218 6443 15252 6477
rect 15218 6375 15252 6409
rect 15408 6529 15442 6563
rect 15408 6461 15442 6495
rect 15408 6393 15442 6427
rect 15496 6529 15530 6563
rect 15734 6553 15768 6587
rect 15830 6689 15864 6723
rect 15830 6621 15864 6655
rect 15830 6553 15864 6587
rect 15926 6689 15960 6723
rect 15926 6621 15960 6655
rect 17622 6689 17656 6723
rect 15926 6553 15960 6587
rect 15496 6461 15530 6495
rect 16054 6529 16088 6563
rect 16054 6461 16088 6495
rect 15496 6393 15530 6427
rect 16054 6393 16088 6427
rect 16142 6529 16176 6563
rect 16142 6461 16176 6495
rect 16142 6393 16176 6427
rect 16330 6519 16364 6553
rect 16330 6451 16364 6485
rect 16330 6383 16364 6417
rect 16414 6519 16448 6553
rect 17622 6621 17656 6655
rect 16414 6451 16448 6485
rect 16414 6383 16448 6417
rect 16629 6466 16663 6500
rect 16629 6385 16663 6419
rect 16715 6453 16749 6487
rect 16715 6385 16749 6419
rect 16801 6453 16835 6487
rect 16801 6385 16835 6419
rect 17022 6511 17056 6545
rect 17022 6443 17056 6477
rect 17022 6375 17056 6409
rect 17106 6511 17140 6545
rect 17106 6443 17140 6477
rect 17106 6375 17140 6409
rect 17296 6529 17330 6563
rect 17296 6461 17330 6495
rect 17296 6393 17330 6427
rect 17384 6529 17418 6563
rect 17622 6553 17656 6587
rect 17718 6689 17752 6723
rect 17718 6621 17752 6655
rect 17718 6553 17752 6587
rect 17814 6689 17848 6723
rect 17814 6621 17848 6655
rect 19510 6689 19544 6723
rect 17814 6553 17848 6587
rect 17384 6461 17418 6495
rect 17942 6529 17976 6563
rect 17942 6461 17976 6495
rect 17384 6393 17418 6427
rect 17942 6393 17976 6427
rect 18030 6529 18064 6563
rect 18030 6461 18064 6495
rect 18030 6393 18064 6427
rect 18218 6519 18252 6553
rect 18218 6451 18252 6485
rect 18218 6383 18252 6417
rect 18302 6519 18336 6553
rect 19510 6621 19544 6655
rect 18302 6451 18336 6485
rect 18302 6383 18336 6417
rect 18517 6466 18551 6500
rect 18517 6385 18551 6419
rect 18603 6453 18637 6487
rect 18603 6385 18637 6419
rect 18689 6453 18723 6487
rect 18689 6385 18723 6419
rect 18910 6511 18944 6545
rect 18910 6443 18944 6477
rect 18910 6375 18944 6409
rect 18994 6511 19028 6545
rect 18994 6443 19028 6477
rect 18994 6375 19028 6409
rect 19184 6529 19218 6563
rect 19184 6461 19218 6495
rect 19184 6393 19218 6427
rect 19272 6529 19306 6563
rect 19510 6553 19544 6587
rect 19606 6689 19640 6723
rect 19606 6621 19640 6655
rect 19606 6553 19640 6587
rect 19702 6689 19736 6723
rect 19702 6621 19736 6655
rect 21398 6689 21432 6723
rect 19702 6553 19736 6587
rect 19272 6461 19306 6495
rect 19830 6529 19864 6563
rect 19830 6461 19864 6495
rect 19272 6393 19306 6427
rect 19830 6393 19864 6427
rect 19918 6529 19952 6563
rect 19918 6461 19952 6495
rect 19918 6393 19952 6427
rect 20106 6519 20140 6553
rect 20106 6451 20140 6485
rect 20106 6383 20140 6417
rect 20190 6519 20224 6553
rect 21398 6621 21432 6655
rect 20190 6451 20224 6485
rect 20190 6383 20224 6417
rect 20405 6466 20439 6500
rect 20405 6385 20439 6419
rect 20491 6453 20525 6487
rect 20491 6385 20525 6419
rect 20577 6453 20611 6487
rect 20577 6385 20611 6419
rect 20798 6511 20832 6545
rect 20798 6443 20832 6477
rect 20798 6375 20832 6409
rect 20882 6511 20916 6545
rect 20882 6443 20916 6477
rect 20882 6375 20916 6409
rect 21072 6529 21106 6563
rect 21072 6461 21106 6495
rect 21072 6393 21106 6427
rect 21160 6529 21194 6563
rect 21398 6553 21432 6587
rect 21494 6689 21528 6723
rect 21494 6621 21528 6655
rect 21494 6553 21528 6587
rect 21590 6689 21624 6723
rect 21590 6621 21624 6655
rect 23286 6689 23320 6723
rect 21590 6553 21624 6587
rect 21160 6461 21194 6495
rect 21718 6529 21752 6563
rect 21718 6461 21752 6495
rect 21160 6393 21194 6427
rect 21718 6393 21752 6427
rect 21806 6529 21840 6563
rect 21806 6461 21840 6495
rect 21806 6393 21840 6427
rect 21994 6519 22028 6553
rect 21994 6451 22028 6485
rect 21994 6383 22028 6417
rect 22078 6519 22112 6553
rect 23286 6621 23320 6655
rect 22078 6451 22112 6485
rect 22078 6383 22112 6417
rect 22293 6466 22327 6500
rect 22293 6385 22327 6419
rect 22379 6453 22413 6487
rect 22379 6385 22413 6419
rect 22465 6453 22499 6487
rect 22465 6385 22499 6419
rect 22686 6511 22720 6545
rect 22686 6443 22720 6477
rect 22686 6375 22720 6409
rect 22770 6511 22804 6545
rect 22770 6443 22804 6477
rect 22770 6375 22804 6409
rect 22960 6529 22994 6563
rect 22960 6461 22994 6495
rect 22960 6393 22994 6427
rect 23048 6529 23082 6563
rect 23286 6553 23320 6587
rect 23382 6689 23416 6723
rect 23382 6621 23416 6655
rect 23382 6553 23416 6587
rect 23478 6689 23512 6723
rect 23478 6621 23512 6655
rect 25174 6689 25208 6723
rect 23478 6553 23512 6587
rect 23048 6461 23082 6495
rect 23606 6529 23640 6563
rect 23606 6461 23640 6495
rect 23048 6393 23082 6427
rect 23606 6393 23640 6427
rect 23694 6529 23728 6563
rect 23694 6461 23728 6495
rect 23694 6393 23728 6427
rect 23882 6519 23916 6553
rect 23882 6451 23916 6485
rect 23882 6383 23916 6417
rect 23966 6519 24000 6553
rect 25174 6621 25208 6655
rect 23966 6451 24000 6485
rect 23966 6383 24000 6417
rect 24181 6466 24215 6500
rect 24181 6385 24215 6419
rect 24267 6453 24301 6487
rect 24267 6385 24301 6419
rect 24353 6453 24387 6487
rect 24353 6385 24387 6419
rect 24574 6511 24608 6545
rect 24574 6443 24608 6477
rect 24574 6375 24608 6409
rect 24658 6511 24692 6545
rect 24658 6443 24692 6477
rect 24658 6375 24692 6409
rect 24848 6529 24882 6563
rect 24848 6461 24882 6495
rect 24848 6393 24882 6427
rect 24936 6529 24970 6563
rect 25174 6553 25208 6587
rect 25270 6689 25304 6723
rect 25270 6621 25304 6655
rect 25270 6553 25304 6587
rect 25366 6689 25400 6723
rect 25366 6621 25400 6655
rect 27062 6689 27096 6723
rect 25366 6553 25400 6587
rect 24936 6461 24970 6495
rect 25494 6529 25528 6563
rect 25494 6461 25528 6495
rect 24936 6393 24970 6427
rect 25494 6393 25528 6427
rect 25582 6529 25616 6563
rect 25582 6461 25616 6495
rect 25582 6393 25616 6427
rect 25770 6519 25804 6553
rect 25770 6451 25804 6485
rect 25770 6383 25804 6417
rect 25854 6519 25888 6553
rect 27062 6621 27096 6655
rect 25854 6451 25888 6485
rect 25854 6383 25888 6417
rect 26069 6466 26103 6500
rect 26069 6385 26103 6419
rect 26155 6453 26189 6487
rect 26155 6385 26189 6419
rect 26241 6453 26275 6487
rect 26241 6385 26275 6419
rect 26462 6511 26496 6545
rect 26462 6443 26496 6477
rect 26462 6375 26496 6409
rect 26546 6511 26580 6545
rect 26546 6443 26580 6477
rect 26546 6375 26580 6409
rect 26736 6529 26770 6563
rect 26736 6461 26770 6495
rect 26736 6393 26770 6427
rect 26824 6529 26858 6563
rect 27062 6553 27096 6587
rect 27158 6689 27192 6723
rect 27158 6621 27192 6655
rect 27158 6553 27192 6587
rect 27254 6689 27288 6723
rect 27254 6621 27288 6655
rect 28950 6689 28984 6723
rect 27254 6553 27288 6587
rect 26824 6461 26858 6495
rect 27382 6529 27416 6563
rect 27382 6461 27416 6495
rect 26824 6393 26858 6427
rect 27382 6393 27416 6427
rect 27470 6529 27504 6563
rect 27470 6461 27504 6495
rect 27470 6393 27504 6427
rect 27658 6519 27692 6553
rect 27658 6451 27692 6485
rect 27658 6383 27692 6417
rect 27742 6519 27776 6553
rect 28950 6621 28984 6655
rect 27742 6451 27776 6485
rect 27742 6383 27776 6417
rect 27957 6466 27991 6500
rect 27957 6385 27991 6419
rect 28043 6453 28077 6487
rect 28043 6385 28077 6419
rect 28129 6453 28163 6487
rect 28129 6385 28163 6419
rect 28350 6511 28384 6545
rect 28350 6443 28384 6477
rect 28350 6375 28384 6409
rect 28434 6511 28468 6545
rect 28434 6443 28468 6477
rect 28434 6375 28468 6409
rect 28624 6529 28658 6563
rect 28624 6461 28658 6495
rect 28624 6393 28658 6427
rect 28712 6529 28746 6563
rect 28950 6553 28984 6587
rect 29046 6689 29080 6723
rect 29046 6621 29080 6655
rect 29046 6553 29080 6587
rect 29142 6689 29176 6723
rect 29142 6621 29176 6655
rect 30838 6689 30872 6723
rect 29142 6553 29176 6587
rect 28712 6461 28746 6495
rect 29270 6529 29304 6563
rect 29270 6461 29304 6495
rect 28712 6393 28746 6427
rect 29270 6393 29304 6427
rect 29358 6529 29392 6563
rect 29358 6461 29392 6495
rect 29358 6393 29392 6427
rect 29546 6519 29580 6553
rect 29546 6451 29580 6485
rect 29546 6383 29580 6417
rect 29630 6519 29664 6553
rect 30838 6621 30872 6655
rect 29630 6451 29664 6485
rect 29630 6383 29664 6417
rect 29845 6466 29879 6500
rect 29845 6385 29879 6419
rect 29931 6453 29965 6487
rect 29931 6385 29965 6419
rect 30017 6453 30051 6487
rect 30017 6385 30051 6419
rect 30238 6511 30272 6545
rect 30238 6443 30272 6477
rect 30238 6375 30272 6409
rect 30322 6511 30356 6545
rect 30322 6443 30356 6477
rect 30322 6375 30356 6409
rect 30512 6529 30546 6563
rect 30512 6461 30546 6495
rect 30512 6393 30546 6427
rect 30600 6529 30634 6563
rect 30838 6553 30872 6587
rect 30934 6689 30968 6723
rect 30934 6621 30968 6655
rect 30934 6553 30968 6587
rect 31030 6689 31064 6723
rect 31030 6621 31064 6655
rect 32726 6689 32760 6723
rect 31030 6553 31064 6587
rect 30600 6461 30634 6495
rect 31158 6529 31192 6563
rect 31158 6461 31192 6495
rect 30600 6393 30634 6427
rect 31158 6393 31192 6427
rect 31246 6529 31280 6563
rect 31246 6461 31280 6495
rect 31246 6393 31280 6427
rect 31434 6519 31468 6553
rect 31434 6451 31468 6485
rect 31434 6383 31468 6417
rect 31518 6519 31552 6553
rect 32726 6621 32760 6655
rect 31518 6451 31552 6485
rect 31518 6383 31552 6417
rect 31733 6466 31767 6500
rect 31733 6385 31767 6419
rect 31819 6453 31853 6487
rect 31819 6385 31853 6419
rect 31905 6453 31939 6487
rect 31905 6385 31939 6419
rect 32126 6511 32160 6545
rect 32126 6443 32160 6477
rect 32126 6375 32160 6409
rect 32210 6511 32244 6545
rect 32210 6443 32244 6477
rect 32210 6375 32244 6409
rect 32400 6529 32434 6563
rect 32400 6461 32434 6495
rect 32400 6393 32434 6427
rect 32488 6529 32522 6563
rect 32726 6553 32760 6587
rect 32822 6689 32856 6723
rect 32822 6621 32856 6655
rect 32822 6553 32856 6587
rect 32918 6689 32952 6723
rect 32918 6621 32952 6655
rect 34614 6689 34648 6723
rect 32918 6553 32952 6587
rect 32488 6461 32522 6495
rect 33046 6529 33080 6563
rect 33046 6461 33080 6495
rect 32488 6393 32522 6427
rect 33046 6393 33080 6427
rect 33134 6529 33168 6563
rect 33134 6461 33168 6495
rect 33134 6393 33168 6427
rect 33322 6519 33356 6553
rect 33322 6451 33356 6485
rect 33322 6383 33356 6417
rect 33406 6519 33440 6553
rect 34614 6621 34648 6655
rect 33406 6451 33440 6485
rect 33406 6383 33440 6417
rect 33621 6466 33655 6500
rect 33621 6385 33655 6419
rect 33707 6453 33741 6487
rect 33707 6385 33741 6419
rect 33793 6453 33827 6487
rect 33793 6385 33827 6419
rect 34014 6511 34048 6545
rect 34014 6443 34048 6477
rect 34014 6375 34048 6409
rect 34098 6511 34132 6545
rect 34098 6443 34132 6477
rect 34098 6375 34132 6409
rect 34288 6529 34322 6563
rect 34288 6461 34322 6495
rect 34288 6393 34322 6427
rect 34376 6529 34410 6563
rect 34614 6553 34648 6587
rect 34710 6689 34744 6723
rect 34710 6621 34744 6655
rect 34710 6553 34744 6587
rect 34806 6689 34840 6723
rect 34806 6621 34840 6655
rect 36502 6689 36536 6723
rect 34806 6553 34840 6587
rect 34376 6461 34410 6495
rect 34934 6529 34968 6563
rect 34934 6461 34968 6495
rect 34376 6393 34410 6427
rect 34934 6393 34968 6427
rect 35022 6529 35056 6563
rect 35022 6461 35056 6495
rect 35022 6393 35056 6427
rect 35210 6519 35244 6553
rect 35210 6451 35244 6485
rect 35210 6383 35244 6417
rect 35294 6519 35328 6553
rect 36502 6621 36536 6655
rect 35294 6451 35328 6485
rect 35294 6383 35328 6417
rect 35509 6466 35543 6500
rect 35509 6385 35543 6419
rect 35595 6453 35629 6487
rect 35595 6385 35629 6419
rect 35681 6453 35715 6487
rect 35681 6385 35715 6419
rect 35902 6511 35936 6545
rect 35902 6443 35936 6477
rect 35902 6375 35936 6409
rect 35986 6511 36020 6545
rect 35986 6443 36020 6477
rect 35986 6375 36020 6409
rect 36176 6529 36210 6563
rect 36176 6461 36210 6495
rect 36176 6393 36210 6427
rect 36264 6529 36298 6563
rect 36502 6553 36536 6587
rect 36598 6689 36632 6723
rect 36598 6621 36632 6655
rect 36598 6553 36632 6587
rect 36694 6689 36728 6723
rect 36694 6621 36728 6655
rect 38390 6689 38424 6723
rect 36694 6553 36728 6587
rect 36264 6461 36298 6495
rect 36822 6529 36856 6563
rect 36822 6461 36856 6495
rect 36264 6393 36298 6427
rect 36822 6393 36856 6427
rect 36910 6529 36944 6563
rect 36910 6461 36944 6495
rect 36910 6393 36944 6427
rect 37098 6519 37132 6553
rect 37098 6451 37132 6485
rect 37098 6383 37132 6417
rect 37182 6519 37216 6553
rect 38390 6621 38424 6655
rect 37182 6451 37216 6485
rect 37182 6383 37216 6417
rect 37397 6466 37431 6500
rect 37397 6385 37431 6419
rect 37483 6453 37517 6487
rect 37483 6385 37517 6419
rect 37569 6453 37603 6487
rect 37569 6385 37603 6419
rect 37790 6511 37824 6545
rect 37790 6443 37824 6477
rect 37790 6375 37824 6409
rect 37874 6511 37908 6545
rect 37874 6443 37908 6477
rect 37874 6375 37908 6409
rect 38064 6529 38098 6563
rect 38064 6461 38098 6495
rect 38064 6393 38098 6427
rect 38152 6529 38186 6563
rect 38390 6553 38424 6587
rect 38486 6689 38520 6723
rect 38486 6621 38520 6655
rect 38486 6553 38520 6587
rect 38582 6689 38616 6723
rect 38582 6621 38616 6655
rect 40278 6689 40312 6723
rect 38582 6553 38616 6587
rect 38152 6461 38186 6495
rect 38710 6529 38744 6563
rect 38710 6461 38744 6495
rect 38152 6393 38186 6427
rect 38710 6393 38744 6427
rect 38798 6529 38832 6563
rect 38798 6461 38832 6495
rect 38798 6393 38832 6427
rect 38986 6519 39020 6553
rect 38986 6451 39020 6485
rect 38986 6383 39020 6417
rect 39070 6519 39104 6553
rect 40278 6621 40312 6655
rect 39070 6451 39104 6485
rect 39070 6383 39104 6417
rect 39285 6466 39319 6500
rect 39285 6385 39319 6419
rect 39371 6453 39405 6487
rect 39371 6385 39405 6419
rect 39457 6453 39491 6487
rect 39457 6385 39491 6419
rect 39678 6511 39712 6545
rect 39678 6443 39712 6477
rect 39678 6375 39712 6409
rect 39762 6511 39796 6545
rect 39762 6443 39796 6477
rect 39762 6375 39796 6409
rect 39952 6529 39986 6563
rect 39952 6461 39986 6495
rect 39952 6393 39986 6427
rect 40040 6529 40074 6563
rect 40278 6553 40312 6587
rect 40374 6689 40408 6723
rect 40374 6621 40408 6655
rect 40374 6553 40408 6587
rect 40470 6689 40504 6723
rect 40470 6621 40504 6655
rect 42166 6689 42200 6723
rect 40470 6553 40504 6587
rect 40040 6461 40074 6495
rect 40598 6529 40632 6563
rect 40598 6461 40632 6495
rect 40040 6393 40074 6427
rect 40598 6393 40632 6427
rect 40686 6529 40720 6563
rect 40686 6461 40720 6495
rect 40686 6393 40720 6427
rect 40874 6519 40908 6553
rect 40874 6451 40908 6485
rect 40874 6383 40908 6417
rect 40958 6519 40992 6553
rect 42166 6621 42200 6655
rect 40958 6451 40992 6485
rect 40958 6383 40992 6417
rect 41173 6466 41207 6500
rect 41173 6385 41207 6419
rect 41259 6453 41293 6487
rect 41259 6385 41293 6419
rect 41345 6453 41379 6487
rect 41345 6385 41379 6419
rect 41566 6511 41600 6545
rect 41566 6443 41600 6477
rect 41566 6375 41600 6409
rect 41650 6511 41684 6545
rect 41650 6443 41684 6477
rect 41650 6375 41684 6409
rect 41840 6529 41874 6563
rect 41840 6461 41874 6495
rect 41840 6393 41874 6427
rect 41928 6529 41962 6563
rect 42166 6553 42200 6587
rect 42262 6689 42296 6723
rect 42262 6621 42296 6655
rect 42262 6553 42296 6587
rect 42358 6689 42392 6723
rect 42358 6621 42392 6655
rect 44054 6689 44088 6723
rect 42358 6553 42392 6587
rect 41928 6461 41962 6495
rect 42486 6529 42520 6563
rect 42486 6461 42520 6495
rect 41928 6393 41962 6427
rect 42486 6393 42520 6427
rect 42574 6529 42608 6563
rect 42574 6461 42608 6495
rect 42574 6393 42608 6427
rect 42762 6519 42796 6553
rect 42762 6451 42796 6485
rect 42762 6383 42796 6417
rect 42846 6519 42880 6553
rect 44054 6621 44088 6655
rect 42846 6451 42880 6485
rect 42846 6383 42880 6417
rect 43061 6466 43095 6500
rect 43061 6385 43095 6419
rect 43147 6453 43181 6487
rect 43147 6385 43181 6419
rect 43233 6453 43267 6487
rect 43233 6385 43267 6419
rect 43454 6511 43488 6545
rect 43454 6443 43488 6477
rect 43454 6375 43488 6409
rect 43538 6511 43572 6545
rect 43538 6443 43572 6477
rect 43538 6375 43572 6409
rect 43728 6529 43762 6563
rect 43728 6461 43762 6495
rect 43728 6393 43762 6427
rect 43816 6529 43850 6563
rect 44054 6553 44088 6587
rect 44150 6689 44184 6723
rect 44150 6621 44184 6655
rect 44150 6553 44184 6587
rect 44246 6689 44280 6723
rect 44246 6621 44280 6655
rect 45936 6689 45970 6723
rect 44246 6553 44280 6587
rect 43816 6461 43850 6495
rect 44374 6529 44408 6563
rect 44374 6461 44408 6495
rect 43816 6393 43850 6427
rect 44374 6393 44408 6427
rect 44462 6529 44496 6563
rect 44462 6461 44496 6495
rect 44462 6393 44496 6427
rect 44650 6519 44684 6553
rect 44650 6451 44684 6485
rect 44650 6383 44684 6417
rect 44734 6519 44768 6553
rect 45936 6621 45970 6655
rect 44734 6451 44768 6485
rect 44734 6383 44768 6417
rect 44943 6466 44977 6500
rect 44943 6385 44977 6419
rect 45029 6453 45063 6487
rect 45029 6385 45063 6419
rect 45115 6453 45149 6487
rect 45115 6385 45149 6419
rect 45336 6511 45370 6545
rect 45336 6443 45370 6477
rect 45336 6375 45370 6409
rect 45420 6511 45454 6545
rect 45420 6443 45454 6477
rect 45420 6375 45454 6409
rect 45610 6529 45644 6563
rect 45610 6461 45644 6495
rect 45610 6393 45644 6427
rect 45698 6529 45732 6563
rect 45936 6553 45970 6587
rect 46032 6689 46066 6723
rect 46032 6621 46066 6655
rect 46032 6553 46066 6587
rect 46128 6689 46162 6723
rect 46128 6621 46162 6655
rect 47824 6689 47858 6723
rect 46128 6553 46162 6587
rect 45698 6461 45732 6495
rect 46256 6529 46290 6563
rect 46256 6461 46290 6495
rect 45698 6393 45732 6427
rect 46256 6393 46290 6427
rect 46344 6529 46378 6563
rect 46344 6461 46378 6495
rect 46344 6393 46378 6427
rect 46532 6519 46566 6553
rect 46532 6451 46566 6485
rect 46532 6383 46566 6417
rect 46616 6519 46650 6553
rect 47824 6621 47858 6655
rect 46616 6451 46650 6485
rect 46616 6383 46650 6417
rect 46831 6466 46865 6500
rect 46831 6385 46865 6419
rect 46917 6453 46951 6487
rect 46917 6385 46951 6419
rect 47003 6453 47037 6487
rect 47003 6385 47037 6419
rect 47224 6511 47258 6545
rect 47224 6443 47258 6477
rect 47224 6375 47258 6409
rect 47308 6511 47342 6545
rect 47308 6443 47342 6477
rect 47308 6375 47342 6409
rect 47498 6529 47532 6563
rect 47498 6461 47532 6495
rect 47498 6393 47532 6427
rect 47586 6529 47620 6563
rect 47824 6553 47858 6587
rect 47920 6689 47954 6723
rect 47920 6621 47954 6655
rect 47920 6553 47954 6587
rect 48016 6689 48050 6723
rect 48016 6621 48050 6655
rect 49712 6689 49746 6723
rect 48016 6553 48050 6587
rect 47586 6461 47620 6495
rect 48144 6529 48178 6563
rect 48144 6461 48178 6495
rect 47586 6393 47620 6427
rect 48144 6393 48178 6427
rect 48232 6529 48266 6563
rect 48232 6461 48266 6495
rect 48232 6393 48266 6427
rect 48420 6519 48454 6553
rect 48420 6451 48454 6485
rect 48420 6383 48454 6417
rect 48504 6519 48538 6553
rect 49712 6621 49746 6655
rect 48504 6451 48538 6485
rect 48504 6383 48538 6417
rect 48719 6466 48753 6500
rect 48719 6385 48753 6419
rect 48805 6453 48839 6487
rect 48805 6385 48839 6419
rect 48891 6453 48925 6487
rect 48891 6385 48925 6419
rect 49112 6511 49146 6545
rect 49112 6443 49146 6477
rect 49112 6375 49146 6409
rect 49196 6511 49230 6545
rect 49196 6443 49230 6477
rect 49196 6375 49230 6409
rect 49386 6529 49420 6563
rect 49386 6461 49420 6495
rect 49386 6393 49420 6427
rect 49474 6529 49508 6563
rect 49712 6553 49746 6587
rect 49808 6689 49842 6723
rect 49808 6621 49842 6655
rect 49808 6553 49842 6587
rect 49904 6689 49938 6723
rect 49904 6621 49938 6655
rect 51600 6689 51634 6723
rect 49904 6553 49938 6587
rect 49474 6461 49508 6495
rect 50032 6529 50066 6563
rect 50032 6461 50066 6495
rect 49474 6393 49508 6427
rect 50032 6393 50066 6427
rect 50120 6529 50154 6563
rect 50120 6461 50154 6495
rect 50120 6393 50154 6427
rect 50308 6519 50342 6553
rect 50308 6451 50342 6485
rect 50308 6383 50342 6417
rect 50392 6519 50426 6553
rect 51600 6621 51634 6655
rect 50392 6451 50426 6485
rect 50392 6383 50426 6417
rect 50607 6466 50641 6500
rect 50607 6385 50641 6419
rect 50693 6453 50727 6487
rect 50693 6385 50727 6419
rect 50779 6453 50813 6487
rect 50779 6385 50813 6419
rect 51000 6511 51034 6545
rect 51000 6443 51034 6477
rect 51000 6375 51034 6409
rect 51084 6511 51118 6545
rect 51084 6443 51118 6477
rect 51084 6375 51118 6409
rect 51274 6529 51308 6563
rect 51274 6461 51308 6495
rect 51274 6393 51308 6427
rect 51362 6529 51396 6563
rect 51600 6553 51634 6587
rect 51696 6689 51730 6723
rect 51696 6621 51730 6655
rect 51696 6553 51730 6587
rect 51792 6689 51826 6723
rect 51792 6621 51826 6655
rect 53488 6689 53522 6723
rect 51792 6553 51826 6587
rect 51362 6461 51396 6495
rect 51920 6529 51954 6563
rect 51920 6461 51954 6495
rect 51362 6393 51396 6427
rect 51920 6393 51954 6427
rect 52008 6529 52042 6563
rect 52008 6461 52042 6495
rect 52008 6393 52042 6427
rect 52196 6519 52230 6553
rect 52196 6451 52230 6485
rect 52196 6383 52230 6417
rect 52280 6519 52314 6553
rect 53488 6621 53522 6655
rect 52280 6451 52314 6485
rect 52280 6383 52314 6417
rect 52495 6466 52529 6500
rect 52495 6385 52529 6419
rect 52581 6453 52615 6487
rect 52581 6385 52615 6419
rect 52667 6453 52701 6487
rect 52667 6385 52701 6419
rect 52888 6511 52922 6545
rect 52888 6443 52922 6477
rect 52888 6375 52922 6409
rect 52972 6511 53006 6545
rect 52972 6443 53006 6477
rect 52972 6375 53006 6409
rect 53162 6529 53196 6563
rect 53162 6461 53196 6495
rect 53162 6393 53196 6427
rect 53250 6529 53284 6563
rect 53488 6553 53522 6587
rect 53584 6689 53618 6723
rect 53584 6621 53618 6655
rect 53584 6553 53618 6587
rect 53680 6689 53714 6723
rect 53680 6621 53714 6655
rect 55376 6689 55410 6723
rect 53680 6553 53714 6587
rect 53250 6461 53284 6495
rect 53808 6529 53842 6563
rect 53808 6461 53842 6495
rect 53250 6393 53284 6427
rect 53808 6393 53842 6427
rect 53896 6529 53930 6563
rect 53896 6461 53930 6495
rect 53896 6393 53930 6427
rect 54084 6519 54118 6553
rect 54084 6451 54118 6485
rect 54084 6383 54118 6417
rect 54168 6519 54202 6553
rect 55376 6621 55410 6655
rect 54168 6451 54202 6485
rect 54168 6383 54202 6417
rect 54383 6466 54417 6500
rect 54383 6385 54417 6419
rect 54469 6453 54503 6487
rect 54469 6385 54503 6419
rect 54555 6453 54589 6487
rect 54555 6385 54589 6419
rect 54776 6511 54810 6545
rect 54776 6443 54810 6477
rect 54776 6375 54810 6409
rect 54860 6511 54894 6545
rect 54860 6443 54894 6477
rect 54860 6375 54894 6409
rect 55050 6529 55084 6563
rect 55050 6461 55084 6495
rect 55050 6393 55084 6427
rect 55138 6529 55172 6563
rect 55376 6553 55410 6587
rect 55472 6689 55506 6723
rect 55472 6621 55506 6655
rect 55472 6553 55506 6587
rect 55568 6689 55602 6723
rect 55568 6621 55602 6655
rect 57264 6689 57298 6723
rect 55568 6553 55602 6587
rect 55138 6461 55172 6495
rect 55696 6529 55730 6563
rect 55696 6461 55730 6495
rect 55138 6393 55172 6427
rect 55696 6393 55730 6427
rect 55784 6529 55818 6563
rect 55784 6461 55818 6495
rect 55784 6393 55818 6427
rect 55972 6519 56006 6553
rect 55972 6451 56006 6485
rect 55972 6383 56006 6417
rect 56056 6519 56090 6553
rect 57264 6621 57298 6655
rect 56056 6451 56090 6485
rect 56056 6383 56090 6417
rect 56271 6466 56305 6500
rect 56271 6385 56305 6419
rect 56357 6453 56391 6487
rect 56357 6385 56391 6419
rect 56443 6453 56477 6487
rect 56443 6385 56477 6419
rect 56664 6511 56698 6545
rect 56664 6443 56698 6477
rect 56664 6375 56698 6409
rect 56748 6511 56782 6545
rect 56748 6443 56782 6477
rect 56748 6375 56782 6409
rect 56938 6529 56972 6563
rect 56938 6461 56972 6495
rect 56938 6393 56972 6427
rect 57026 6529 57060 6563
rect 57264 6553 57298 6587
rect 57360 6689 57394 6723
rect 57360 6621 57394 6655
rect 57360 6553 57394 6587
rect 57456 6689 57490 6723
rect 57456 6621 57490 6655
rect 59152 6689 59186 6723
rect 57456 6553 57490 6587
rect 57026 6461 57060 6495
rect 57584 6529 57618 6563
rect 57584 6461 57618 6495
rect 57026 6393 57060 6427
rect 57584 6393 57618 6427
rect 57672 6529 57706 6563
rect 57672 6461 57706 6495
rect 57672 6393 57706 6427
rect 57860 6519 57894 6553
rect 57860 6451 57894 6485
rect 57860 6383 57894 6417
rect 57944 6519 57978 6553
rect 59152 6621 59186 6655
rect 57944 6451 57978 6485
rect 57944 6383 57978 6417
rect 58159 6466 58193 6500
rect 58159 6385 58193 6419
rect 58245 6453 58279 6487
rect 58245 6385 58279 6419
rect 58331 6453 58365 6487
rect 58331 6385 58365 6419
rect 58552 6511 58586 6545
rect 58552 6443 58586 6477
rect 58552 6375 58586 6409
rect 58636 6511 58670 6545
rect 58636 6443 58670 6477
rect 58636 6375 58670 6409
rect 58826 6529 58860 6563
rect 58826 6461 58860 6495
rect 58826 6393 58860 6427
rect 58914 6529 58948 6563
rect 59152 6553 59186 6587
rect 59248 6689 59282 6723
rect 59248 6621 59282 6655
rect 59248 6553 59282 6587
rect 59344 6689 59378 6723
rect 59344 6621 59378 6655
rect 59344 6553 59378 6587
rect 58914 6461 58948 6495
rect 59472 6529 59506 6563
rect 59472 6461 59506 6495
rect 58914 6393 58948 6427
rect 59472 6393 59506 6427
rect 59560 6529 59594 6563
rect 59560 6461 59594 6495
rect 59560 6393 59594 6427
rect 59748 6519 59782 6553
rect 59748 6451 59782 6485
rect 59748 6383 59782 6417
rect 59832 6519 59866 6553
rect 59832 6451 59866 6485
rect 59832 6383 59866 6417
rect 634 5633 668 5667
rect 634 5565 668 5599
rect 209 5465 243 5499
rect 209 5397 243 5431
rect 209 5329 243 5363
rect 365 5465 399 5499
rect 634 5497 668 5531
rect 730 5633 764 5667
rect 730 5565 764 5599
rect 730 5497 764 5531
rect 826 5633 860 5667
rect 826 5565 860 5599
rect 826 5497 860 5531
rect 2522 5633 2556 5667
rect 2522 5565 2556 5599
rect 1023 5465 1057 5499
rect 365 5397 399 5431
rect 1023 5397 1057 5431
rect 365 5329 399 5363
rect 1023 5329 1057 5363
rect 1179 5465 1213 5499
rect 1179 5397 1213 5431
rect 1179 5329 1213 5363
rect 2097 5465 2131 5499
rect 2097 5397 2131 5431
rect 2097 5329 2131 5363
rect 2253 5465 2287 5499
rect 2522 5497 2556 5531
rect 2618 5633 2652 5667
rect 2618 5565 2652 5599
rect 2618 5497 2652 5531
rect 2714 5633 2748 5667
rect 2714 5565 2748 5599
rect 2714 5497 2748 5531
rect 4410 5633 4444 5667
rect 4410 5565 4444 5599
rect 2911 5465 2945 5499
rect 2253 5397 2287 5431
rect 2911 5397 2945 5431
rect 2253 5329 2287 5363
rect 2911 5329 2945 5363
rect 3067 5465 3101 5499
rect 3067 5397 3101 5431
rect 3067 5329 3101 5363
rect 3985 5465 4019 5499
rect 3985 5397 4019 5431
rect 3985 5329 4019 5363
rect 4141 5465 4175 5499
rect 4410 5497 4444 5531
rect 4506 5633 4540 5667
rect 4506 5565 4540 5599
rect 4506 5497 4540 5531
rect 4602 5633 4636 5667
rect 4602 5565 4636 5599
rect 4602 5497 4636 5531
rect 6298 5633 6332 5667
rect 6298 5565 6332 5599
rect 4799 5465 4833 5499
rect 4141 5397 4175 5431
rect 4799 5397 4833 5431
rect 4141 5329 4175 5363
rect 4799 5329 4833 5363
rect 4955 5465 4989 5499
rect 4955 5397 4989 5431
rect 4955 5329 4989 5363
rect 5873 5465 5907 5499
rect 5873 5397 5907 5431
rect 5873 5329 5907 5363
rect 6029 5465 6063 5499
rect 6298 5497 6332 5531
rect 6394 5633 6428 5667
rect 6394 5565 6428 5599
rect 6394 5497 6428 5531
rect 6490 5633 6524 5667
rect 6490 5565 6524 5599
rect 6490 5497 6524 5531
rect 8186 5633 8220 5667
rect 8186 5565 8220 5599
rect 6687 5465 6721 5499
rect 6029 5397 6063 5431
rect 6687 5397 6721 5431
rect 6029 5329 6063 5363
rect 6687 5329 6721 5363
rect 6843 5465 6877 5499
rect 6843 5397 6877 5431
rect 6843 5329 6877 5363
rect 7761 5465 7795 5499
rect 7761 5397 7795 5431
rect 7761 5329 7795 5363
rect 7917 5465 7951 5499
rect 8186 5497 8220 5531
rect 8282 5633 8316 5667
rect 8282 5565 8316 5599
rect 8282 5497 8316 5531
rect 8378 5633 8412 5667
rect 8378 5565 8412 5599
rect 8378 5497 8412 5531
rect 10074 5633 10108 5667
rect 10074 5565 10108 5599
rect 8575 5465 8609 5499
rect 7917 5397 7951 5431
rect 8575 5397 8609 5431
rect 7917 5329 7951 5363
rect 8575 5329 8609 5363
rect 8731 5465 8765 5499
rect 8731 5397 8765 5431
rect 8731 5329 8765 5363
rect 9649 5465 9683 5499
rect 9649 5397 9683 5431
rect 9649 5329 9683 5363
rect 9805 5465 9839 5499
rect 10074 5497 10108 5531
rect 10170 5633 10204 5667
rect 10170 5565 10204 5599
rect 10170 5497 10204 5531
rect 10266 5633 10300 5667
rect 10266 5565 10300 5599
rect 10266 5497 10300 5531
rect 11962 5633 11996 5667
rect 11962 5565 11996 5599
rect 10463 5465 10497 5499
rect 9805 5397 9839 5431
rect 10463 5397 10497 5431
rect 9805 5329 9839 5363
rect 10463 5329 10497 5363
rect 10619 5465 10653 5499
rect 10619 5397 10653 5431
rect 10619 5329 10653 5363
rect 11537 5465 11571 5499
rect 11537 5397 11571 5431
rect 11537 5329 11571 5363
rect 11693 5465 11727 5499
rect 11962 5497 11996 5531
rect 12058 5633 12092 5667
rect 12058 5565 12092 5599
rect 12058 5497 12092 5531
rect 12154 5633 12188 5667
rect 12154 5565 12188 5599
rect 12154 5497 12188 5531
rect 13850 5633 13884 5667
rect 13850 5565 13884 5599
rect 12351 5465 12385 5499
rect 11693 5397 11727 5431
rect 12351 5397 12385 5431
rect 11693 5329 11727 5363
rect 12351 5329 12385 5363
rect 12507 5465 12541 5499
rect 12507 5397 12541 5431
rect 12507 5329 12541 5363
rect 13425 5465 13459 5499
rect 13425 5397 13459 5431
rect 13425 5329 13459 5363
rect 13581 5465 13615 5499
rect 13850 5497 13884 5531
rect 13946 5633 13980 5667
rect 13946 5565 13980 5599
rect 13946 5497 13980 5531
rect 14042 5633 14076 5667
rect 14042 5565 14076 5599
rect 14042 5497 14076 5531
rect 15732 5633 15766 5667
rect 15732 5565 15766 5599
rect 14239 5465 14273 5499
rect 13581 5397 13615 5431
rect 14239 5397 14273 5431
rect 13581 5329 13615 5363
rect 14239 5329 14273 5363
rect 14395 5465 14429 5499
rect 14395 5397 14429 5431
rect 14395 5329 14429 5363
rect 15307 5465 15341 5499
rect 15307 5397 15341 5431
rect 15307 5329 15341 5363
rect 15463 5465 15497 5499
rect 15732 5497 15766 5531
rect 15828 5633 15862 5667
rect 15828 5565 15862 5599
rect 15828 5497 15862 5531
rect 15924 5633 15958 5667
rect 15924 5565 15958 5599
rect 15924 5497 15958 5531
rect 17620 5633 17654 5667
rect 17620 5565 17654 5599
rect 16121 5465 16155 5499
rect 15463 5397 15497 5431
rect 16121 5397 16155 5431
rect 15463 5329 15497 5363
rect 16121 5329 16155 5363
rect 16277 5465 16311 5499
rect 16277 5397 16311 5431
rect 16277 5329 16311 5363
rect 17195 5465 17229 5499
rect 17195 5397 17229 5431
rect 17195 5329 17229 5363
rect 17351 5465 17385 5499
rect 17620 5497 17654 5531
rect 17716 5633 17750 5667
rect 17716 5565 17750 5599
rect 17716 5497 17750 5531
rect 17812 5633 17846 5667
rect 17812 5565 17846 5599
rect 17812 5497 17846 5531
rect 19508 5633 19542 5667
rect 19508 5565 19542 5599
rect 18009 5465 18043 5499
rect 17351 5397 17385 5431
rect 18009 5397 18043 5431
rect 17351 5329 17385 5363
rect 18009 5329 18043 5363
rect 18165 5465 18199 5499
rect 18165 5397 18199 5431
rect 18165 5329 18199 5363
rect 19083 5465 19117 5499
rect 19083 5397 19117 5431
rect 19083 5329 19117 5363
rect 19239 5465 19273 5499
rect 19508 5497 19542 5531
rect 19604 5633 19638 5667
rect 19604 5565 19638 5599
rect 19604 5497 19638 5531
rect 19700 5633 19734 5667
rect 19700 5565 19734 5599
rect 19700 5497 19734 5531
rect 21396 5633 21430 5667
rect 21396 5565 21430 5599
rect 19897 5465 19931 5499
rect 19239 5397 19273 5431
rect 19897 5397 19931 5431
rect 19239 5329 19273 5363
rect 19897 5329 19931 5363
rect 20053 5465 20087 5499
rect 20053 5397 20087 5431
rect 20053 5329 20087 5363
rect 20971 5465 21005 5499
rect 20971 5397 21005 5431
rect 20971 5329 21005 5363
rect 21127 5465 21161 5499
rect 21396 5497 21430 5531
rect 21492 5633 21526 5667
rect 21492 5565 21526 5599
rect 21492 5497 21526 5531
rect 21588 5633 21622 5667
rect 21588 5565 21622 5599
rect 21588 5497 21622 5531
rect 23284 5633 23318 5667
rect 23284 5565 23318 5599
rect 21785 5465 21819 5499
rect 21127 5397 21161 5431
rect 21785 5397 21819 5431
rect 21127 5329 21161 5363
rect 21785 5329 21819 5363
rect 21941 5465 21975 5499
rect 21941 5397 21975 5431
rect 21941 5329 21975 5363
rect 22859 5465 22893 5499
rect 22859 5397 22893 5431
rect 22859 5329 22893 5363
rect 23015 5465 23049 5499
rect 23284 5497 23318 5531
rect 23380 5633 23414 5667
rect 23380 5565 23414 5599
rect 23380 5497 23414 5531
rect 23476 5633 23510 5667
rect 23476 5565 23510 5599
rect 23476 5497 23510 5531
rect 25172 5633 25206 5667
rect 25172 5565 25206 5599
rect 23673 5465 23707 5499
rect 23015 5397 23049 5431
rect 23673 5397 23707 5431
rect 23015 5329 23049 5363
rect 23673 5329 23707 5363
rect 23829 5465 23863 5499
rect 23829 5397 23863 5431
rect 23829 5329 23863 5363
rect 24747 5465 24781 5499
rect 24747 5397 24781 5431
rect 24747 5329 24781 5363
rect 24903 5465 24937 5499
rect 25172 5497 25206 5531
rect 25268 5633 25302 5667
rect 25268 5565 25302 5599
rect 25268 5497 25302 5531
rect 25364 5633 25398 5667
rect 25364 5565 25398 5599
rect 25364 5497 25398 5531
rect 27060 5633 27094 5667
rect 27060 5565 27094 5599
rect 25561 5465 25595 5499
rect 24903 5397 24937 5431
rect 25561 5397 25595 5431
rect 24903 5329 24937 5363
rect 25561 5329 25595 5363
rect 25717 5465 25751 5499
rect 25717 5397 25751 5431
rect 25717 5329 25751 5363
rect 26635 5465 26669 5499
rect 26635 5397 26669 5431
rect 26635 5329 26669 5363
rect 26791 5465 26825 5499
rect 27060 5497 27094 5531
rect 27156 5633 27190 5667
rect 27156 5565 27190 5599
rect 27156 5497 27190 5531
rect 27252 5633 27286 5667
rect 27252 5565 27286 5599
rect 27252 5497 27286 5531
rect 28948 5633 28982 5667
rect 28948 5565 28982 5599
rect 27449 5465 27483 5499
rect 26791 5397 26825 5431
rect 27449 5397 27483 5431
rect 26791 5329 26825 5363
rect 27449 5329 27483 5363
rect 27605 5465 27639 5499
rect 27605 5397 27639 5431
rect 27605 5329 27639 5363
rect 28523 5465 28557 5499
rect 28523 5397 28557 5431
rect 28523 5329 28557 5363
rect 28679 5465 28713 5499
rect 28948 5497 28982 5531
rect 29044 5633 29078 5667
rect 29044 5565 29078 5599
rect 29044 5497 29078 5531
rect 29140 5633 29174 5667
rect 29140 5565 29174 5599
rect 29140 5497 29174 5531
rect 30836 5633 30870 5667
rect 30836 5565 30870 5599
rect 29337 5465 29371 5499
rect 28679 5397 28713 5431
rect 29337 5397 29371 5431
rect 28679 5329 28713 5363
rect 29337 5329 29371 5363
rect 29493 5465 29527 5499
rect 29493 5397 29527 5431
rect 29493 5329 29527 5363
rect 30411 5465 30445 5499
rect 30411 5397 30445 5431
rect 30411 5329 30445 5363
rect 30567 5465 30601 5499
rect 30836 5497 30870 5531
rect 30932 5633 30966 5667
rect 30932 5565 30966 5599
rect 30932 5497 30966 5531
rect 31028 5633 31062 5667
rect 31028 5565 31062 5599
rect 31028 5497 31062 5531
rect 32724 5633 32758 5667
rect 32724 5565 32758 5599
rect 31225 5465 31259 5499
rect 30567 5397 30601 5431
rect 31225 5397 31259 5431
rect 30567 5329 30601 5363
rect 31225 5329 31259 5363
rect 31381 5465 31415 5499
rect 31381 5397 31415 5431
rect 31381 5329 31415 5363
rect 32299 5465 32333 5499
rect 32299 5397 32333 5431
rect 32299 5329 32333 5363
rect 32455 5465 32489 5499
rect 32724 5497 32758 5531
rect 32820 5633 32854 5667
rect 32820 5565 32854 5599
rect 32820 5497 32854 5531
rect 32916 5633 32950 5667
rect 32916 5565 32950 5599
rect 32916 5497 32950 5531
rect 34612 5633 34646 5667
rect 34612 5565 34646 5599
rect 33113 5465 33147 5499
rect 32455 5397 32489 5431
rect 33113 5397 33147 5431
rect 32455 5329 32489 5363
rect 33113 5329 33147 5363
rect 33269 5465 33303 5499
rect 33269 5397 33303 5431
rect 33269 5329 33303 5363
rect 34187 5465 34221 5499
rect 34187 5397 34221 5431
rect 34187 5329 34221 5363
rect 34343 5465 34377 5499
rect 34612 5497 34646 5531
rect 34708 5633 34742 5667
rect 34708 5565 34742 5599
rect 34708 5497 34742 5531
rect 34804 5633 34838 5667
rect 34804 5565 34838 5599
rect 34804 5497 34838 5531
rect 36500 5633 36534 5667
rect 36500 5565 36534 5599
rect 35001 5465 35035 5499
rect 34343 5397 34377 5431
rect 35001 5397 35035 5431
rect 34343 5329 34377 5363
rect 35001 5329 35035 5363
rect 35157 5465 35191 5499
rect 35157 5397 35191 5431
rect 35157 5329 35191 5363
rect 36075 5465 36109 5499
rect 36075 5397 36109 5431
rect 36075 5329 36109 5363
rect 36231 5465 36265 5499
rect 36500 5497 36534 5531
rect 36596 5633 36630 5667
rect 36596 5565 36630 5599
rect 36596 5497 36630 5531
rect 36692 5633 36726 5667
rect 36692 5565 36726 5599
rect 36692 5497 36726 5531
rect 38388 5633 38422 5667
rect 38388 5565 38422 5599
rect 36889 5465 36923 5499
rect 36231 5397 36265 5431
rect 36889 5397 36923 5431
rect 36231 5329 36265 5363
rect 36889 5329 36923 5363
rect 37045 5465 37079 5499
rect 37045 5397 37079 5431
rect 37045 5329 37079 5363
rect 37963 5465 37997 5499
rect 37963 5397 37997 5431
rect 37963 5329 37997 5363
rect 38119 5465 38153 5499
rect 38388 5497 38422 5531
rect 38484 5633 38518 5667
rect 38484 5565 38518 5599
rect 38484 5497 38518 5531
rect 38580 5633 38614 5667
rect 38580 5565 38614 5599
rect 38580 5497 38614 5531
rect 40276 5633 40310 5667
rect 40276 5565 40310 5599
rect 38777 5465 38811 5499
rect 38119 5397 38153 5431
rect 38777 5397 38811 5431
rect 38119 5329 38153 5363
rect 38777 5329 38811 5363
rect 38933 5465 38967 5499
rect 38933 5397 38967 5431
rect 38933 5329 38967 5363
rect 39851 5465 39885 5499
rect 39851 5397 39885 5431
rect 39851 5329 39885 5363
rect 40007 5465 40041 5499
rect 40276 5497 40310 5531
rect 40372 5633 40406 5667
rect 40372 5565 40406 5599
rect 40372 5497 40406 5531
rect 40468 5633 40502 5667
rect 40468 5565 40502 5599
rect 40468 5497 40502 5531
rect 42164 5633 42198 5667
rect 42164 5565 42198 5599
rect 40665 5465 40699 5499
rect 40007 5397 40041 5431
rect 40665 5397 40699 5431
rect 40007 5329 40041 5363
rect 40665 5329 40699 5363
rect 40821 5465 40855 5499
rect 40821 5397 40855 5431
rect 40821 5329 40855 5363
rect 41739 5465 41773 5499
rect 41739 5397 41773 5431
rect 41739 5329 41773 5363
rect 41895 5465 41929 5499
rect 42164 5497 42198 5531
rect 42260 5633 42294 5667
rect 42260 5565 42294 5599
rect 42260 5497 42294 5531
rect 42356 5633 42390 5667
rect 42356 5565 42390 5599
rect 42356 5497 42390 5531
rect 44052 5633 44086 5667
rect 44052 5565 44086 5599
rect 42553 5465 42587 5499
rect 41895 5397 41929 5431
rect 42553 5397 42587 5431
rect 41895 5329 41929 5363
rect 42553 5329 42587 5363
rect 42709 5465 42743 5499
rect 42709 5397 42743 5431
rect 42709 5329 42743 5363
rect 43627 5465 43661 5499
rect 43627 5397 43661 5431
rect 43627 5329 43661 5363
rect 43783 5465 43817 5499
rect 44052 5497 44086 5531
rect 44148 5633 44182 5667
rect 44148 5565 44182 5599
rect 44148 5497 44182 5531
rect 44244 5633 44278 5667
rect 44244 5565 44278 5599
rect 44244 5497 44278 5531
rect 45934 5633 45968 5667
rect 45934 5565 45968 5599
rect 44441 5465 44475 5499
rect 43783 5397 43817 5431
rect 44441 5397 44475 5431
rect 43783 5329 43817 5363
rect 44441 5329 44475 5363
rect 44597 5465 44631 5499
rect 44597 5397 44631 5431
rect 44597 5329 44631 5363
rect 45509 5465 45543 5499
rect 45509 5397 45543 5431
rect 45509 5329 45543 5363
rect 45665 5465 45699 5499
rect 45934 5497 45968 5531
rect 46030 5633 46064 5667
rect 46030 5565 46064 5599
rect 46030 5497 46064 5531
rect 46126 5633 46160 5667
rect 46126 5565 46160 5599
rect 46126 5497 46160 5531
rect 47822 5633 47856 5667
rect 47822 5565 47856 5599
rect 46323 5465 46357 5499
rect 45665 5397 45699 5431
rect 46323 5397 46357 5431
rect 45665 5329 45699 5363
rect 46323 5329 46357 5363
rect 46479 5465 46513 5499
rect 46479 5397 46513 5431
rect 46479 5329 46513 5363
rect 47397 5465 47431 5499
rect 47397 5397 47431 5431
rect 47397 5329 47431 5363
rect 47553 5465 47587 5499
rect 47822 5497 47856 5531
rect 47918 5633 47952 5667
rect 47918 5565 47952 5599
rect 47918 5497 47952 5531
rect 48014 5633 48048 5667
rect 48014 5565 48048 5599
rect 48014 5497 48048 5531
rect 49710 5633 49744 5667
rect 49710 5565 49744 5599
rect 48211 5465 48245 5499
rect 47553 5397 47587 5431
rect 48211 5397 48245 5431
rect 47553 5329 47587 5363
rect 48211 5329 48245 5363
rect 48367 5465 48401 5499
rect 48367 5397 48401 5431
rect 48367 5329 48401 5363
rect 49285 5465 49319 5499
rect 49285 5397 49319 5431
rect 49285 5329 49319 5363
rect 49441 5465 49475 5499
rect 49710 5497 49744 5531
rect 49806 5633 49840 5667
rect 49806 5565 49840 5599
rect 49806 5497 49840 5531
rect 49902 5633 49936 5667
rect 49902 5565 49936 5599
rect 49902 5497 49936 5531
rect 51598 5633 51632 5667
rect 51598 5565 51632 5599
rect 50099 5465 50133 5499
rect 49441 5397 49475 5431
rect 50099 5397 50133 5431
rect 49441 5329 49475 5363
rect 50099 5329 50133 5363
rect 50255 5465 50289 5499
rect 50255 5397 50289 5431
rect 50255 5329 50289 5363
rect 51173 5465 51207 5499
rect 51173 5397 51207 5431
rect 51173 5329 51207 5363
rect 51329 5465 51363 5499
rect 51598 5497 51632 5531
rect 51694 5633 51728 5667
rect 51694 5565 51728 5599
rect 51694 5497 51728 5531
rect 51790 5633 51824 5667
rect 51790 5565 51824 5599
rect 51790 5497 51824 5531
rect 53486 5633 53520 5667
rect 53486 5565 53520 5599
rect 51987 5465 52021 5499
rect 51329 5397 51363 5431
rect 51987 5397 52021 5431
rect 51329 5329 51363 5363
rect 51987 5329 52021 5363
rect 52143 5465 52177 5499
rect 52143 5397 52177 5431
rect 52143 5329 52177 5363
rect 53061 5465 53095 5499
rect 53061 5397 53095 5431
rect 53061 5329 53095 5363
rect 53217 5465 53251 5499
rect 53486 5497 53520 5531
rect 53582 5633 53616 5667
rect 53582 5565 53616 5599
rect 53582 5497 53616 5531
rect 53678 5633 53712 5667
rect 53678 5565 53712 5599
rect 53678 5497 53712 5531
rect 55374 5633 55408 5667
rect 55374 5565 55408 5599
rect 53875 5465 53909 5499
rect 53217 5397 53251 5431
rect 53875 5397 53909 5431
rect 53217 5329 53251 5363
rect 53875 5329 53909 5363
rect 54031 5465 54065 5499
rect 54031 5397 54065 5431
rect 54031 5329 54065 5363
rect 54949 5465 54983 5499
rect 54949 5397 54983 5431
rect 54949 5329 54983 5363
rect 55105 5465 55139 5499
rect 55374 5497 55408 5531
rect 55470 5633 55504 5667
rect 55470 5565 55504 5599
rect 55470 5497 55504 5531
rect 55566 5633 55600 5667
rect 55566 5565 55600 5599
rect 55566 5497 55600 5531
rect 57262 5633 57296 5667
rect 57262 5565 57296 5599
rect 55763 5465 55797 5499
rect 55105 5397 55139 5431
rect 55763 5397 55797 5431
rect 55105 5329 55139 5363
rect 55763 5329 55797 5363
rect 55919 5465 55953 5499
rect 55919 5397 55953 5431
rect 55919 5329 55953 5363
rect 56837 5465 56871 5499
rect 56837 5397 56871 5431
rect 56837 5329 56871 5363
rect 56993 5465 57027 5499
rect 57262 5497 57296 5531
rect 57358 5633 57392 5667
rect 57358 5565 57392 5599
rect 57358 5497 57392 5531
rect 57454 5633 57488 5667
rect 57454 5565 57488 5599
rect 57454 5497 57488 5531
rect 59150 5633 59184 5667
rect 59150 5565 59184 5599
rect 57651 5465 57685 5499
rect 56993 5397 57027 5431
rect 57651 5397 57685 5431
rect 56993 5329 57027 5363
rect 57651 5329 57685 5363
rect 57807 5465 57841 5499
rect 57807 5397 57841 5431
rect 57807 5329 57841 5363
rect 58725 5465 58759 5499
rect 58725 5397 58759 5431
rect 58725 5329 58759 5363
rect 58881 5465 58915 5499
rect 59150 5497 59184 5531
rect 59246 5633 59280 5667
rect 59246 5565 59280 5599
rect 59246 5497 59280 5531
rect 59342 5633 59376 5667
rect 59342 5565 59376 5599
rect 59342 5497 59376 5531
rect 59539 5465 59573 5499
rect 58881 5397 58915 5431
rect 59539 5397 59573 5431
rect 58881 5329 58915 5363
rect 59539 5329 59573 5363
rect 59695 5465 59729 5499
rect 59695 5397 59729 5431
rect 59695 5329 59729 5363
rect 5710 5099 5744 5133
rect 5710 5031 5744 5065
rect 5794 5099 5828 5133
rect 5794 5031 5828 5065
rect 5794 4961 5828 4995
rect 5878 5099 5912 5133
rect 5878 5031 5912 5065
rect 5962 5099 5996 5133
rect 5962 5031 5996 5065
rect 5962 4961 5996 4995
rect 6046 5099 6080 5133
rect 6046 5031 6080 5065
rect 6130 5099 6164 5133
rect 6130 5031 6164 5065
rect 6130 4961 6164 4995
rect 6214 5099 6248 5133
rect 6214 5031 6248 5065
rect 6298 5099 6332 5133
rect 6298 5031 6332 5065
rect 6298 4961 6332 4995
rect 6382 5099 6416 5133
rect 6382 5031 6416 5065
rect 6466 5099 6500 5133
rect 6466 5031 6500 5065
rect 6466 4961 6500 4995
rect 6550 5099 6584 5133
rect 6550 5031 6584 5065
rect 6634 5099 6668 5133
rect 6634 5031 6668 5065
rect 6634 4961 6668 4995
rect 6718 5099 6752 5133
rect 6718 5031 6752 5065
rect 6802 5099 6836 5133
rect 6802 5031 6836 5065
rect 6802 4961 6836 4995
rect 6886 5099 6920 5133
rect 6886 5031 6920 5065
rect 6970 5099 7004 5133
rect 6970 5031 7004 5065
rect 6970 4961 7004 4995
rect 7054 5099 7088 5133
rect 7054 5031 7088 5065
rect 7054 4961 7088 4995
rect 7592 5097 7626 5131
rect 7592 5029 7626 5063
rect 7676 5097 7710 5131
rect 7676 5029 7710 5063
rect 7676 4959 7710 4993
rect 7760 5097 7794 5131
rect 7760 5029 7794 5063
rect 7844 5097 7878 5131
rect 7844 5029 7878 5063
rect 7844 4959 7878 4993
rect 7928 5097 7962 5131
rect 7928 5029 7962 5063
rect 8012 5097 8046 5131
rect 8012 5029 8046 5063
rect 8012 4959 8046 4993
rect 8096 5097 8130 5131
rect 8096 5029 8130 5063
rect 8180 5097 8214 5131
rect 8180 5029 8214 5063
rect 8180 4959 8214 4993
rect 8264 5097 8298 5131
rect 8264 5029 8298 5063
rect 8348 5097 8382 5131
rect 8348 5029 8382 5063
rect 8348 4959 8382 4993
rect 8432 5097 8466 5131
rect 8432 5029 8466 5063
rect 8516 5097 8550 5131
rect 8516 5029 8550 5063
rect 8516 4959 8550 4993
rect 8600 5097 8634 5131
rect 8600 5029 8634 5063
rect 8684 5097 8718 5131
rect 8684 5029 8718 5063
rect 8684 4959 8718 4993
rect 8768 5097 8802 5131
rect 8768 5029 8802 5063
rect 8852 5097 8886 5131
rect 8852 5029 8886 5063
rect 8852 4959 8886 4993
rect 8936 5097 8970 5131
rect 8936 5029 8970 5063
rect 8936 4959 8970 4993
rect 20808 5099 20842 5133
rect 20808 5031 20842 5065
rect 20892 5099 20926 5133
rect 20892 5031 20926 5065
rect 20892 4961 20926 4995
rect 20976 5099 21010 5133
rect 20976 5031 21010 5065
rect 21060 5099 21094 5133
rect 21060 5031 21094 5065
rect 21060 4961 21094 4995
rect 21144 5099 21178 5133
rect 21144 5031 21178 5065
rect 21228 5099 21262 5133
rect 21228 5031 21262 5065
rect 21228 4961 21262 4995
rect 21312 5099 21346 5133
rect 21312 5031 21346 5065
rect 21396 5099 21430 5133
rect 21396 5031 21430 5065
rect 21396 4961 21430 4995
rect 21480 5099 21514 5133
rect 21480 5031 21514 5065
rect 21564 5099 21598 5133
rect 21564 5031 21598 5065
rect 21564 4961 21598 4995
rect 21648 5099 21682 5133
rect 21648 5031 21682 5065
rect 21732 5099 21766 5133
rect 21732 5031 21766 5065
rect 21732 4961 21766 4995
rect 21816 5099 21850 5133
rect 21816 5031 21850 5065
rect 21900 5099 21934 5133
rect 21900 5031 21934 5065
rect 21900 4961 21934 4995
rect 21984 5099 22018 5133
rect 21984 5031 22018 5065
rect 22068 5099 22102 5133
rect 22068 5031 22102 5065
rect 22068 4961 22102 4995
rect 22152 5099 22186 5133
rect 22152 5031 22186 5065
rect 22152 4961 22186 4995
rect 22690 5097 22724 5131
rect 22690 5029 22724 5063
rect 22774 5097 22808 5131
rect 22774 5029 22808 5063
rect 22774 4959 22808 4993
rect 22858 5097 22892 5131
rect 22858 5029 22892 5063
rect 22942 5097 22976 5131
rect 22942 5029 22976 5063
rect 22942 4959 22976 4993
rect 23026 5097 23060 5131
rect 23026 5029 23060 5063
rect 23110 5097 23144 5131
rect 23110 5029 23144 5063
rect 23110 4959 23144 4993
rect 23194 5097 23228 5131
rect 23194 5029 23228 5063
rect 23278 5097 23312 5131
rect 23278 5029 23312 5063
rect 23278 4959 23312 4993
rect 23362 5097 23396 5131
rect 23362 5029 23396 5063
rect 23446 5097 23480 5131
rect 23446 5029 23480 5063
rect 23446 4959 23480 4993
rect 23530 5097 23564 5131
rect 23530 5029 23564 5063
rect 23614 5097 23648 5131
rect 23614 5029 23648 5063
rect 23614 4959 23648 4993
rect 23698 5097 23732 5131
rect 23698 5029 23732 5063
rect 23782 5097 23816 5131
rect 23782 5029 23816 5063
rect 23782 4959 23816 4993
rect 23866 5097 23900 5131
rect 23866 5029 23900 5063
rect 23950 5097 23984 5131
rect 23950 5029 23984 5063
rect 23950 4959 23984 4993
rect 24034 5097 24068 5131
rect 24034 5029 24068 5063
rect 24034 4959 24068 4993
rect 35912 5099 35946 5133
rect 35912 5031 35946 5065
rect 35996 5099 36030 5133
rect 35996 5031 36030 5065
rect 35996 4961 36030 4995
rect 36080 5099 36114 5133
rect 36080 5031 36114 5065
rect 36164 5099 36198 5133
rect 36164 5031 36198 5065
rect 36164 4961 36198 4995
rect 36248 5099 36282 5133
rect 36248 5031 36282 5065
rect 36332 5099 36366 5133
rect 36332 5031 36366 5065
rect 36332 4961 36366 4995
rect 36416 5099 36450 5133
rect 36416 5031 36450 5065
rect 36500 5099 36534 5133
rect 36500 5031 36534 5065
rect 36500 4961 36534 4995
rect 36584 5099 36618 5133
rect 36584 5031 36618 5065
rect 36668 5099 36702 5133
rect 36668 5031 36702 5065
rect 36668 4961 36702 4995
rect 36752 5099 36786 5133
rect 36752 5031 36786 5065
rect 36836 5099 36870 5133
rect 36836 5031 36870 5065
rect 36836 4961 36870 4995
rect 36920 5099 36954 5133
rect 36920 5031 36954 5065
rect 37004 5099 37038 5133
rect 37004 5031 37038 5065
rect 37004 4961 37038 4995
rect 37088 5099 37122 5133
rect 37088 5031 37122 5065
rect 37172 5099 37206 5133
rect 37172 5031 37206 5065
rect 37172 4961 37206 4995
rect 37256 5099 37290 5133
rect 37256 5031 37290 5065
rect 37256 4961 37290 4995
rect 37794 5097 37828 5131
rect 37794 5029 37828 5063
rect 37878 5097 37912 5131
rect 37878 5029 37912 5063
rect 37878 4959 37912 4993
rect 37962 5097 37996 5131
rect 37962 5029 37996 5063
rect 38046 5097 38080 5131
rect 38046 5029 38080 5063
rect 38046 4959 38080 4993
rect 38130 5097 38164 5131
rect 38130 5029 38164 5063
rect 38214 5097 38248 5131
rect 38214 5029 38248 5063
rect 38214 4959 38248 4993
rect 38298 5097 38332 5131
rect 38298 5029 38332 5063
rect 38382 5097 38416 5131
rect 38382 5029 38416 5063
rect 38382 4959 38416 4993
rect 38466 5097 38500 5131
rect 38466 5029 38500 5063
rect 38550 5097 38584 5131
rect 38550 5029 38584 5063
rect 38550 4959 38584 4993
rect 38634 5097 38668 5131
rect 38634 5029 38668 5063
rect 38718 5097 38752 5131
rect 38718 5029 38752 5063
rect 38718 4959 38752 4993
rect 38802 5097 38836 5131
rect 38802 5029 38836 5063
rect 38886 5097 38920 5131
rect 38886 5029 38920 5063
rect 38886 4959 38920 4993
rect 38970 5097 39004 5131
rect 38970 5029 39004 5063
rect 39054 5097 39088 5131
rect 39054 5029 39088 5063
rect 39054 4959 39088 4993
rect 39138 5097 39172 5131
rect 39138 5029 39172 5063
rect 39138 4959 39172 4993
rect 51010 5099 51044 5133
rect 51010 5031 51044 5065
rect 51094 5099 51128 5133
rect 51094 5031 51128 5065
rect 51094 4961 51128 4995
rect 51178 5099 51212 5133
rect 51178 5031 51212 5065
rect 51262 5099 51296 5133
rect 51262 5031 51296 5065
rect 51262 4961 51296 4995
rect 51346 5099 51380 5133
rect 51346 5031 51380 5065
rect 51430 5099 51464 5133
rect 51430 5031 51464 5065
rect 51430 4961 51464 4995
rect 51514 5099 51548 5133
rect 51514 5031 51548 5065
rect 51598 5099 51632 5133
rect 51598 5031 51632 5065
rect 51598 4961 51632 4995
rect 51682 5099 51716 5133
rect 51682 5031 51716 5065
rect 51766 5099 51800 5133
rect 51766 5031 51800 5065
rect 51766 4961 51800 4995
rect 51850 5099 51884 5133
rect 51850 5031 51884 5065
rect 51934 5099 51968 5133
rect 51934 5031 51968 5065
rect 51934 4961 51968 4995
rect 52018 5099 52052 5133
rect 52018 5031 52052 5065
rect 52102 5099 52136 5133
rect 52102 5031 52136 5065
rect 52102 4961 52136 4995
rect 52186 5099 52220 5133
rect 52186 5031 52220 5065
rect 52270 5099 52304 5133
rect 52270 5031 52304 5065
rect 52270 4961 52304 4995
rect 52354 5099 52388 5133
rect 52354 5031 52388 5065
rect 52354 4961 52388 4995
rect 52892 5097 52926 5131
rect 52892 5029 52926 5063
rect 52976 5097 53010 5131
rect 52976 5029 53010 5063
rect 52976 4959 53010 4993
rect 53060 5097 53094 5131
rect 53060 5029 53094 5063
rect 53144 5097 53178 5131
rect 53144 5029 53178 5063
rect 53144 4959 53178 4993
rect 53228 5097 53262 5131
rect 53228 5029 53262 5063
rect 53312 5097 53346 5131
rect 53312 5029 53346 5063
rect 53312 4959 53346 4993
rect 53396 5097 53430 5131
rect 53396 5029 53430 5063
rect 53480 5097 53514 5131
rect 53480 5029 53514 5063
rect 53480 4959 53514 4993
rect 53564 5097 53598 5131
rect 53564 5029 53598 5063
rect 53648 5097 53682 5131
rect 53648 5029 53682 5063
rect 53648 4959 53682 4993
rect 53732 5097 53766 5131
rect 53732 5029 53766 5063
rect 53816 5097 53850 5131
rect 53816 5029 53850 5063
rect 53816 4959 53850 4993
rect 53900 5097 53934 5131
rect 53900 5029 53934 5063
rect 53984 5097 54018 5131
rect 53984 5029 54018 5063
rect 53984 4959 54018 4993
rect 54068 5097 54102 5131
rect 54068 5029 54102 5063
rect 54152 5097 54186 5131
rect 54152 5029 54186 5063
rect 54152 4959 54186 4993
rect 54236 5097 54270 5131
rect 54236 5029 54270 5063
rect 54236 4959 54270 4993
rect 30072 4022 30106 4056
rect 30072 3954 30106 3988
rect 30072 3886 30106 3920
rect 30156 4022 30190 4056
rect 30156 3954 30190 3988
rect 30156 3886 30190 3920
rect 30240 4022 30274 4056
rect 30240 3954 30274 3988
rect 30324 4022 30358 4056
rect 30324 3954 30358 3988
rect 30324 3886 30358 3920
rect 30408 4022 30442 4056
rect 30603 4022 30637 4056
rect 30603 3954 30637 3988
rect 30603 3884 30637 3918
rect 30687 4022 30721 4056
rect 30687 3954 30721 3988
rect 30687 3884 30721 3918
rect 30771 4022 30805 4056
rect 30771 3954 30805 3988
rect 30855 4022 30889 4056
rect 30855 3954 30889 3988
rect 30855 3884 30889 3918
rect 30939 4022 30973 4056
rect 30939 3954 30973 3988
rect 31023 4022 31057 4056
rect 31023 3954 31057 3988
rect 31023 3884 31057 3918
rect 31107 4022 31141 4056
rect 31107 3954 31141 3988
rect 31191 4022 31225 4056
rect 31191 3954 31225 3988
rect 31191 3884 31225 3918
rect 31275 4022 31309 4056
rect 31275 3954 31309 3988
rect 31359 4022 31393 4056
rect 31359 3954 31393 3988
rect 31359 3884 31393 3918
rect 31443 4022 31477 4056
rect 31443 3954 31477 3988
rect 31527 4022 31561 4056
rect 31527 3954 31561 3988
rect 31527 3884 31561 3918
rect 31611 4022 31645 4056
rect 31611 3954 31645 3988
rect 31695 4022 31729 4056
rect 31695 3954 31729 3988
rect 31695 3884 31729 3918
rect 31779 4022 31813 4056
rect 31779 3954 31813 3988
rect 31863 4022 31897 4056
rect 31863 3954 31897 3988
rect 31863 3884 31897 3918
rect 31947 4022 31981 4056
rect 31947 3954 31981 3988
rect 43429 3806 43463 3840
rect 13287 3646 13321 3680
rect 13287 3578 13321 3612
rect 13287 3508 13321 3542
rect 13371 3646 13405 3680
rect 13371 3578 13405 3612
rect 13371 3508 13405 3542
rect 13455 3646 13489 3680
rect 13455 3578 13489 3612
rect 13539 3646 13573 3680
rect 13539 3578 13573 3612
rect 13539 3508 13573 3542
rect 13623 3646 13657 3680
rect 13623 3578 13657 3612
rect 13707 3646 13741 3680
rect 13707 3578 13741 3612
rect 13707 3508 13741 3542
rect 13791 3646 13825 3680
rect 13791 3578 13825 3612
rect 13875 3646 13909 3680
rect 13875 3578 13909 3612
rect 13875 3508 13909 3542
rect 13959 3646 13993 3680
rect 13959 3578 13993 3612
rect 14043 3646 14077 3680
rect 14043 3578 14077 3612
rect 14043 3508 14077 3542
rect 14127 3646 14161 3680
rect 14127 3578 14161 3612
rect 14211 3646 14245 3680
rect 14211 3578 14245 3612
rect 14211 3508 14245 3542
rect 14295 3646 14329 3680
rect 14295 3578 14329 3612
rect 14379 3646 14413 3680
rect 14379 3578 14413 3612
rect 14379 3508 14413 3542
rect 14463 3646 14497 3680
rect 14463 3578 14497 3612
rect 14547 3646 14581 3680
rect 14547 3578 14581 3612
rect 14547 3508 14581 3542
rect 14631 3646 14665 3680
rect 14631 3578 14665 3612
rect 15217 3646 15251 3680
rect 15217 3578 15251 3612
rect 15217 3508 15251 3542
rect 15301 3646 15335 3680
rect 15301 3578 15335 3612
rect 15301 3508 15335 3542
rect 15385 3646 15419 3680
rect 15385 3578 15419 3612
rect 15469 3646 15503 3680
rect 15469 3578 15503 3612
rect 15469 3508 15503 3542
rect 15553 3646 15587 3680
rect 15553 3578 15587 3612
rect 15637 3646 15671 3680
rect 15637 3578 15671 3612
rect 15637 3508 15671 3542
rect 15721 3646 15755 3680
rect 15721 3578 15755 3612
rect 15805 3646 15839 3680
rect 15805 3578 15839 3612
rect 15805 3508 15839 3542
rect 15889 3646 15923 3680
rect 15889 3578 15923 3612
rect 15973 3646 16007 3680
rect 15973 3578 16007 3612
rect 15973 3508 16007 3542
rect 16057 3646 16091 3680
rect 16057 3578 16091 3612
rect 16141 3646 16175 3680
rect 16141 3578 16175 3612
rect 16141 3508 16175 3542
rect 16225 3646 16259 3680
rect 16225 3578 16259 3612
rect 16309 3646 16343 3680
rect 16309 3578 16343 3612
rect 16309 3508 16343 3542
rect 16393 3646 16427 3680
rect 16393 3578 16427 3612
rect 16477 3646 16511 3680
rect 16477 3578 16511 3612
rect 16477 3508 16511 3542
rect 16561 3646 16595 3680
rect 43429 3738 43463 3772
rect 43429 3668 43463 3702
rect 43513 3806 43547 3840
rect 43513 3738 43547 3772
rect 43513 3668 43547 3702
rect 43597 3806 43631 3840
rect 43597 3738 43631 3772
rect 43681 3806 43715 3840
rect 43681 3738 43715 3772
rect 43681 3668 43715 3702
rect 43765 3806 43799 3840
rect 43765 3738 43799 3772
rect 43849 3806 43883 3840
rect 43849 3738 43883 3772
rect 43849 3668 43883 3702
rect 43933 3806 43967 3840
rect 43933 3738 43967 3772
rect 44017 3806 44051 3840
rect 44017 3738 44051 3772
rect 44017 3668 44051 3702
rect 44101 3806 44135 3840
rect 44101 3738 44135 3772
rect 44185 3806 44219 3840
rect 44185 3738 44219 3772
rect 44185 3668 44219 3702
rect 44269 3806 44303 3840
rect 44269 3738 44303 3772
rect 44353 3806 44387 3840
rect 44353 3738 44387 3772
rect 44353 3668 44387 3702
rect 44437 3806 44471 3840
rect 44437 3738 44471 3772
rect 44521 3806 44555 3840
rect 44521 3738 44555 3772
rect 44521 3668 44555 3702
rect 44605 3806 44639 3840
rect 44605 3738 44639 3772
rect 44689 3806 44723 3840
rect 44689 3738 44723 3772
rect 44689 3668 44723 3702
rect 44773 3806 44807 3840
rect 44773 3738 44807 3772
rect 45359 3806 45393 3840
rect 45359 3738 45393 3772
rect 45359 3668 45393 3702
rect 45443 3806 45477 3840
rect 45443 3738 45477 3772
rect 45443 3668 45477 3702
rect 45527 3806 45561 3840
rect 45527 3738 45561 3772
rect 45611 3806 45645 3840
rect 45611 3738 45645 3772
rect 45611 3668 45645 3702
rect 45695 3806 45729 3840
rect 45695 3738 45729 3772
rect 45779 3806 45813 3840
rect 45779 3738 45813 3772
rect 45779 3668 45813 3702
rect 45863 3806 45897 3840
rect 45863 3738 45897 3772
rect 45947 3806 45981 3840
rect 45947 3738 45981 3772
rect 45947 3668 45981 3702
rect 46031 3806 46065 3840
rect 46031 3738 46065 3772
rect 46115 3806 46149 3840
rect 46115 3738 46149 3772
rect 46115 3668 46149 3702
rect 46199 3806 46233 3840
rect 46199 3738 46233 3772
rect 46283 3806 46317 3840
rect 46283 3738 46317 3772
rect 46283 3668 46317 3702
rect 46367 3806 46401 3840
rect 46367 3738 46401 3772
rect 46451 3806 46485 3840
rect 46451 3738 46485 3772
rect 46451 3668 46485 3702
rect 46535 3806 46569 3840
rect 46535 3738 46569 3772
rect 46619 3806 46653 3840
rect 46619 3738 46653 3772
rect 46619 3668 46653 3702
rect 46703 3806 46737 3840
rect 46703 3738 46737 3772
rect 16561 3578 16595 3612
rect 5712 2447 5746 2481
rect 5712 2377 5746 2411
rect 5712 2309 5746 2343
rect 5796 2447 5830 2481
rect 5796 2377 5830 2411
rect 5796 2309 5830 2343
rect 5880 2377 5914 2411
rect 5880 2309 5914 2343
rect 5964 2447 5998 2481
rect 5964 2377 5998 2411
rect 5964 2309 5998 2343
rect 6048 2377 6082 2411
rect 6048 2309 6082 2343
rect 6132 2447 6166 2481
rect 6132 2377 6166 2411
rect 6132 2309 6166 2343
rect 6216 2377 6250 2411
rect 6216 2309 6250 2343
rect 6300 2447 6334 2481
rect 6300 2377 6334 2411
rect 6300 2309 6334 2343
rect 6384 2377 6418 2411
rect 6384 2309 6418 2343
rect 6468 2447 6502 2481
rect 6468 2377 6502 2411
rect 6468 2309 6502 2343
rect 6552 2377 6586 2411
rect 6552 2309 6586 2343
rect 6636 2447 6670 2481
rect 6636 2377 6670 2411
rect 6636 2309 6670 2343
rect 6720 2377 6754 2411
rect 6720 2309 6754 2343
rect 6804 2447 6838 2481
rect 6804 2377 6838 2411
rect 6804 2309 6838 2343
rect 6888 2377 6922 2411
rect 6888 2309 6922 2343
rect 6972 2447 7006 2481
rect 6972 2377 7006 2411
rect 6972 2309 7006 2343
rect 7056 2377 7090 2411
rect 7056 2309 7090 2343
rect 7594 2445 7628 2479
rect 7594 2375 7628 2409
rect 7594 2307 7628 2341
rect 7678 2445 7712 2479
rect 7678 2375 7712 2409
rect 7678 2307 7712 2341
rect 7762 2375 7796 2409
rect 7762 2307 7796 2341
rect 7846 2445 7880 2479
rect 7846 2375 7880 2409
rect 7846 2307 7880 2341
rect 7930 2375 7964 2409
rect 7930 2307 7964 2341
rect 8014 2445 8048 2479
rect 8014 2375 8048 2409
rect 8014 2307 8048 2341
rect 8098 2375 8132 2409
rect 8098 2307 8132 2341
rect 8182 2445 8216 2479
rect 8182 2375 8216 2409
rect 8182 2307 8216 2341
rect 8266 2375 8300 2409
rect 8266 2307 8300 2341
rect 8350 2445 8384 2479
rect 8350 2375 8384 2409
rect 8350 2307 8384 2341
rect 8434 2375 8468 2409
rect 8434 2307 8468 2341
rect 8518 2445 8552 2479
rect 8518 2375 8552 2409
rect 8518 2307 8552 2341
rect 8602 2375 8636 2409
rect 8602 2307 8636 2341
rect 8686 2445 8720 2479
rect 8686 2375 8720 2409
rect 8686 2307 8720 2341
rect 8770 2375 8804 2409
rect 8770 2307 8804 2341
rect 8854 2445 8888 2479
rect 8854 2375 8888 2409
rect 8854 2307 8888 2341
rect 8938 2375 8972 2409
rect 8938 2307 8972 2341
rect 20810 2447 20844 2481
rect 20810 2377 20844 2411
rect 20810 2309 20844 2343
rect 20894 2447 20928 2481
rect 20894 2377 20928 2411
rect 20894 2309 20928 2343
rect 20978 2377 21012 2411
rect 20978 2309 21012 2343
rect 21062 2447 21096 2481
rect 21062 2377 21096 2411
rect 21062 2309 21096 2343
rect 21146 2377 21180 2411
rect 21146 2309 21180 2343
rect 21230 2447 21264 2481
rect 21230 2377 21264 2411
rect 21230 2309 21264 2343
rect 21314 2377 21348 2411
rect 21314 2309 21348 2343
rect 21398 2447 21432 2481
rect 21398 2377 21432 2411
rect 21398 2309 21432 2343
rect 21482 2377 21516 2411
rect 21482 2309 21516 2343
rect 21566 2447 21600 2481
rect 21566 2377 21600 2411
rect 21566 2309 21600 2343
rect 21650 2377 21684 2411
rect 21650 2309 21684 2343
rect 21734 2447 21768 2481
rect 21734 2377 21768 2411
rect 21734 2309 21768 2343
rect 21818 2377 21852 2411
rect 21818 2309 21852 2343
rect 21902 2447 21936 2481
rect 21902 2377 21936 2411
rect 21902 2309 21936 2343
rect 21986 2377 22020 2411
rect 21986 2309 22020 2343
rect 22070 2447 22104 2481
rect 22070 2377 22104 2411
rect 22070 2309 22104 2343
rect 22154 2377 22188 2411
rect 22154 2309 22188 2343
rect 22692 2445 22726 2479
rect 22692 2375 22726 2409
rect 22692 2307 22726 2341
rect 22776 2445 22810 2479
rect 22776 2375 22810 2409
rect 22776 2307 22810 2341
rect 22860 2375 22894 2409
rect 22860 2307 22894 2341
rect 22944 2445 22978 2479
rect 22944 2375 22978 2409
rect 22944 2307 22978 2341
rect 23028 2375 23062 2409
rect 23028 2307 23062 2341
rect 23112 2445 23146 2479
rect 23112 2375 23146 2409
rect 23112 2307 23146 2341
rect 23196 2375 23230 2409
rect 23196 2307 23230 2341
rect 23280 2445 23314 2479
rect 23280 2375 23314 2409
rect 23280 2307 23314 2341
rect 23364 2375 23398 2409
rect 23364 2307 23398 2341
rect 23448 2445 23482 2479
rect 23448 2375 23482 2409
rect 23448 2307 23482 2341
rect 23532 2375 23566 2409
rect 23532 2307 23566 2341
rect 23616 2445 23650 2479
rect 23616 2375 23650 2409
rect 23616 2307 23650 2341
rect 23700 2375 23734 2409
rect 23700 2307 23734 2341
rect 23784 2445 23818 2479
rect 23784 2375 23818 2409
rect 23784 2307 23818 2341
rect 23868 2375 23902 2409
rect 23868 2307 23902 2341
rect 23952 2445 23986 2479
rect 23952 2375 23986 2409
rect 23952 2307 23986 2341
rect 24036 2375 24070 2409
rect 24036 2307 24070 2341
rect 35914 2447 35948 2481
rect 35914 2377 35948 2411
rect 35914 2309 35948 2343
rect 35998 2447 36032 2481
rect 35998 2377 36032 2411
rect 35998 2309 36032 2343
rect 36082 2377 36116 2411
rect 36082 2309 36116 2343
rect 36166 2447 36200 2481
rect 36166 2377 36200 2411
rect 36166 2309 36200 2343
rect 36250 2377 36284 2411
rect 36250 2309 36284 2343
rect 36334 2447 36368 2481
rect 36334 2377 36368 2411
rect 36334 2309 36368 2343
rect 36418 2377 36452 2411
rect 36418 2309 36452 2343
rect 36502 2447 36536 2481
rect 36502 2377 36536 2411
rect 36502 2309 36536 2343
rect 36586 2377 36620 2411
rect 36586 2309 36620 2343
rect 36670 2447 36704 2481
rect 36670 2377 36704 2411
rect 36670 2309 36704 2343
rect 36754 2377 36788 2411
rect 36754 2309 36788 2343
rect 36838 2447 36872 2481
rect 36838 2377 36872 2411
rect 36838 2309 36872 2343
rect 36922 2377 36956 2411
rect 36922 2309 36956 2343
rect 37006 2447 37040 2481
rect 37006 2377 37040 2411
rect 37006 2309 37040 2343
rect 37090 2377 37124 2411
rect 37090 2309 37124 2343
rect 37174 2447 37208 2481
rect 37174 2377 37208 2411
rect 37174 2309 37208 2343
rect 37258 2377 37292 2411
rect 37258 2309 37292 2343
rect 37796 2445 37830 2479
rect 37796 2375 37830 2409
rect 37796 2307 37830 2341
rect 37880 2445 37914 2479
rect 37880 2375 37914 2409
rect 37880 2307 37914 2341
rect 37964 2375 37998 2409
rect 37964 2307 37998 2341
rect 38048 2445 38082 2479
rect 38048 2375 38082 2409
rect 38048 2307 38082 2341
rect 38132 2375 38166 2409
rect 38132 2307 38166 2341
rect 38216 2445 38250 2479
rect 38216 2375 38250 2409
rect 38216 2307 38250 2341
rect 38300 2375 38334 2409
rect 38300 2307 38334 2341
rect 38384 2445 38418 2479
rect 38384 2375 38418 2409
rect 38384 2307 38418 2341
rect 38468 2375 38502 2409
rect 38468 2307 38502 2341
rect 38552 2445 38586 2479
rect 38552 2375 38586 2409
rect 38552 2307 38586 2341
rect 38636 2375 38670 2409
rect 38636 2307 38670 2341
rect 38720 2445 38754 2479
rect 38720 2375 38754 2409
rect 38720 2307 38754 2341
rect 38804 2375 38838 2409
rect 38804 2307 38838 2341
rect 38888 2445 38922 2479
rect 38888 2375 38922 2409
rect 38888 2307 38922 2341
rect 38972 2375 39006 2409
rect 38972 2307 39006 2341
rect 39056 2445 39090 2479
rect 39056 2375 39090 2409
rect 39056 2307 39090 2341
rect 39140 2375 39174 2409
rect 39140 2307 39174 2341
rect 51012 2447 51046 2481
rect 51012 2377 51046 2411
rect 51012 2309 51046 2343
rect 51096 2447 51130 2481
rect 51096 2377 51130 2411
rect 51096 2309 51130 2343
rect 51180 2377 51214 2411
rect 51180 2309 51214 2343
rect 51264 2447 51298 2481
rect 51264 2377 51298 2411
rect 51264 2309 51298 2343
rect 51348 2377 51382 2411
rect 51348 2309 51382 2343
rect 51432 2447 51466 2481
rect 51432 2377 51466 2411
rect 51432 2309 51466 2343
rect 51516 2377 51550 2411
rect 51516 2309 51550 2343
rect 51600 2447 51634 2481
rect 51600 2377 51634 2411
rect 51600 2309 51634 2343
rect 51684 2377 51718 2411
rect 51684 2309 51718 2343
rect 51768 2447 51802 2481
rect 51768 2377 51802 2411
rect 51768 2309 51802 2343
rect 51852 2377 51886 2411
rect 51852 2309 51886 2343
rect 51936 2447 51970 2481
rect 51936 2377 51970 2411
rect 51936 2309 51970 2343
rect 52020 2377 52054 2411
rect 52020 2309 52054 2343
rect 52104 2447 52138 2481
rect 52104 2377 52138 2411
rect 52104 2309 52138 2343
rect 52188 2377 52222 2411
rect 52188 2309 52222 2343
rect 52272 2447 52306 2481
rect 52272 2377 52306 2411
rect 52272 2309 52306 2343
rect 52356 2377 52390 2411
rect 52356 2309 52390 2343
rect 52894 2445 52928 2479
rect 52894 2375 52928 2409
rect 52894 2307 52928 2341
rect 52978 2445 53012 2479
rect 52978 2375 53012 2409
rect 52978 2307 53012 2341
rect 53062 2375 53096 2409
rect 53062 2307 53096 2341
rect 53146 2445 53180 2479
rect 53146 2375 53180 2409
rect 53146 2307 53180 2341
rect 53230 2375 53264 2409
rect 53230 2307 53264 2341
rect 53314 2445 53348 2479
rect 53314 2375 53348 2409
rect 53314 2307 53348 2341
rect 53398 2375 53432 2409
rect 53398 2307 53432 2341
rect 53482 2445 53516 2479
rect 53482 2375 53516 2409
rect 53482 2307 53516 2341
rect 53566 2375 53600 2409
rect 53566 2307 53600 2341
rect 53650 2445 53684 2479
rect 53650 2375 53684 2409
rect 53650 2307 53684 2341
rect 53734 2375 53768 2409
rect 53734 2307 53768 2341
rect 53818 2445 53852 2479
rect 53818 2375 53852 2409
rect 53818 2307 53852 2341
rect 53902 2375 53936 2409
rect 53902 2307 53936 2341
rect 53986 2445 54020 2479
rect 53986 2375 54020 2409
rect 53986 2307 54020 2341
rect 54070 2375 54104 2409
rect 54070 2307 54104 2341
rect 54154 2445 54188 2479
rect 54154 2375 54188 2409
rect 54154 2307 54188 2341
rect 54238 2375 54272 2409
rect 54238 2307 54272 2341
rect 253 2077 287 2111
rect 253 2009 287 2043
rect 253 1941 287 1975
rect 409 2077 443 2111
rect 1067 2077 1101 2111
rect 409 2009 443 2043
rect 1067 2009 1101 2043
rect 409 1941 443 1975
rect 606 1909 640 1943
rect 606 1841 640 1875
rect 606 1773 640 1807
rect 702 1909 736 1943
rect 702 1841 736 1875
rect 702 1773 736 1807
rect 798 1909 832 1943
rect 1067 1941 1101 1975
rect 1223 2077 1257 2111
rect 1223 2009 1257 2043
rect 1223 1941 1257 1975
rect 2141 2077 2175 2111
rect 2141 2009 2175 2043
rect 2141 1941 2175 1975
rect 2297 2077 2331 2111
rect 2955 2077 2989 2111
rect 2297 2009 2331 2043
rect 2955 2009 2989 2043
rect 2297 1941 2331 1975
rect 798 1841 832 1875
rect 798 1773 832 1807
rect 2494 1909 2528 1943
rect 2494 1841 2528 1875
rect 2494 1773 2528 1807
rect 2590 1909 2624 1943
rect 2590 1841 2624 1875
rect 2590 1773 2624 1807
rect 2686 1909 2720 1943
rect 2955 1941 2989 1975
rect 3111 2077 3145 2111
rect 3111 2009 3145 2043
rect 3111 1941 3145 1975
rect 4029 2077 4063 2111
rect 4029 2009 4063 2043
rect 4029 1941 4063 1975
rect 4185 2077 4219 2111
rect 4843 2077 4877 2111
rect 4185 2009 4219 2043
rect 4843 2009 4877 2043
rect 4185 1941 4219 1975
rect 2686 1841 2720 1875
rect 2686 1773 2720 1807
rect 4382 1909 4416 1943
rect 4382 1841 4416 1875
rect 4382 1773 4416 1807
rect 4478 1909 4512 1943
rect 4478 1841 4512 1875
rect 4478 1773 4512 1807
rect 4574 1909 4608 1943
rect 4843 1941 4877 1975
rect 4999 2077 5033 2111
rect 4999 2009 5033 2043
rect 4999 1941 5033 1975
rect 5917 2077 5951 2111
rect 5917 2009 5951 2043
rect 5917 1941 5951 1975
rect 6073 2077 6107 2111
rect 6731 2077 6765 2111
rect 6073 2009 6107 2043
rect 6731 2009 6765 2043
rect 6073 1941 6107 1975
rect 4574 1841 4608 1875
rect 4574 1773 4608 1807
rect 6270 1909 6304 1943
rect 6270 1841 6304 1875
rect 6270 1773 6304 1807
rect 6366 1909 6400 1943
rect 6366 1841 6400 1875
rect 6366 1773 6400 1807
rect 6462 1909 6496 1943
rect 6731 1941 6765 1975
rect 6887 2077 6921 2111
rect 6887 2009 6921 2043
rect 6887 1941 6921 1975
rect 7805 2077 7839 2111
rect 7805 2009 7839 2043
rect 7805 1941 7839 1975
rect 7961 2077 7995 2111
rect 8619 2077 8653 2111
rect 7961 2009 7995 2043
rect 8619 2009 8653 2043
rect 7961 1941 7995 1975
rect 6462 1841 6496 1875
rect 6462 1773 6496 1807
rect 8158 1909 8192 1943
rect 8158 1841 8192 1875
rect 8158 1773 8192 1807
rect 8254 1909 8288 1943
rect 8254 1841 8288 1875
rect 8254 1773 8288 1807
rect 8350 1909 8384 1943
rect 8619 1941 8653 1975
rect 8775 2077 8809 2111
rect 8775 2009 8809 2043
rect 8775 1941 8809 1975
rect 9693 2077 9727 2111
rect 9693 2009 9727 2043
rect 9693 1941 9727 1975
rect 9849 2077 9883 2111
rect 10507 2077 10541 2111
rect 9849 2009 9883 2043
rect 10507 2009 10541 2043
rect 9849 1941 9883 1975
rect 8350 1841 8384 1875
rect 8350 1773 8384 1807
rect 10046 1909 10080 1943
rect 10046 1841 10080 1875
rect 10046 1773 10080 1807
rect 10142 1909 10176 1943
rect 10142 1841 10176 1875
rect 10142 1773 10176 1807
rect 10238 1909 10272 1943
rect 10507 1941 10541 1975
rect 10663 2077 10697 2111
rect 10663 2009 10697 2043
rect 10663 1941 10697 1975
rect 11581 2077 11615 2111
rect 11581 2009 11615 2043
rect 11581 1941 11615 1975
rect 11737 2077 11771 2111
rect 12395 2077 12429 2111
rect 11737 2009 11771 2043
rect 12395 2009 12429 2043
rect 11737 1941 11771 1975
rect 10238 1841 10272 1875
rect 10238 1773 10272 1807
rect 11934 1909 11968 1943
rect 11934 1841 11968 1875
rect 11934 1773 11968 1807
rect 12030 1909 12064 1943
rect 12030 1841 12064 1875
rect 12030 1773 12064 1807
rect 12126 1909 12160 1943
rect 12395 1941 12429 1975
rect 12551 2077 12585 2111
rect 12551 2009 12585 2043
rect 12551 1941 12585 1975
rect 13469 2077 13503 2111
rect 13469 2009 13503 2043
rect 13469 1941 13503 1975
rect 13625 2077 13659 2111
rect 14283 2077 14317 2111
rect 13625 2009 13659 2043
rect 14283 2009 14317 2043
rect 13625 1941 13659 1975
rect 12126 1841 12160 1875
rect 12126 1773 12160 1807
rect 13822 1909 13856 1943
rect 13822 1841 13856 1875
rect 13822 1773 13856 1807
rect 13918 1909 13952 1943
rect 13918 1841 13952 1875
rect 13918 1773 13952 1807
rect 14014 1909 14048 1943
rect 14283 1941 14317 1975
rect 14439 2077 14473 2111
rect 14439 2009 14473 2043
rect 14439 1941 14473 1975
rect 15351 2077 15385 2111
rect 15351 2009 15385 2043
rect 15351 1941 15385 1975
rect 15507 2077 15541 2111
rect 16165 2077 16199 2111
rect 15507 2009 15541 2043
rect 16165 2009 16199 2043
rect 15507 1941 15541 1975
rect 14014 1841 14048 1875
rect 14014 1773 14048 1807
rect 15704 1909 15738 1943
rect 15704 1841 15738 1875
rect 15704 1773 15738 1807
rect 15800 1909 15834 1943
rect 15800 1841 15834 1875
rect 15800 1773 15834 1807
rect 15896 1909 15930 1943
rect 16165 1941 16199 1975
rect 16321 2077 16355 2111
rect 16321 2009 16355 2043
rect 16321 1941 16355 1975
rect 17239 2077 17273 2111
rect 17239 2009 17273 2043
rect 17239 1941 17273 1975
rect 17395 2077 17429 2111
rect 18053 2077 18087 2111
rect 17395 2009 17429 2043
rect 18053 2009 18087 2043
rect 17395 1941 17429 1975
rect 15896 1841 15930 1875
rect 15896 1773 15930 1807
rect 17592 1909 17626 1943
rect 17592 1841 17626 1875
rect 17592 1773 17626 1807
rect 17688 1909 17722 1943
rect 17688 1841 17722 1875
rect 17688 1773 17722 1807
rect 17784 1909 17818 1943
rect 18053 1941 18087 1975
rect 18209 2077 18243 2111
rect 18209 2009 18243 2043
rect 18209 1941 18243 1975
rect 19127 2077 19161 2111
rect 19127 2009 19161 2043
rect 19127 1941 19161 1975
rect 19283 2077 19317 2111
rect 19941 2077 19975 2111
rect 19283 2009 19317 2043
rect 19941 2009 19975 2043
rect 19283 1941 19317 1975
rect 17784 1841 17818 1875
rect 17784 1773 17818 1807
rect 19480 1909 19514 1943
rect 19480 1841 19514 1875
rect 19480 1773 19514 1807
rect 19576 1909 19610 1943
rect 19576 1841 19610 1875
rect 19576 1773 19610 1807
rect 19672 1909 19706 1943
rect 19941 1941 19975 1975
rect 20097 2077 20131 2111
rect 20097 2009 20131 2043
rect 20097 1941 20131 1975
rect 21015 2077 21049 2111
rect 21015 2009 21049 2043
rect 21015 1941 21049 1975
rect 21171 2077 21205 2111
rect 21829 2077 21863 2111
rect 21171 2009 21205 2043
rect 21829 2009 21863 2043
rect 21171 1941 21205 1975
rect 19672 1841 19706 1875
rect 19672 1773 19706 1807
rect 21368 1909 21402 1943
rect 21368 1841 21402 1875
rect 21368 1773 21402 1807
rect 21464 1909 21498 1943
rect 21464 1841 21498 1875
rect 21464 1773 21498 1807
rect 21560 1909 21594 1943
rect 21829 1941 21863 1975
rect 21985 2077 22019 2111
rect 21985 2009 22019 2043
rect 21985 1941 22019 1975
rect 22903 2077 22937 2111
rect 22903 2009 22937 2043
rect 22903 1941 22937 1975
rect 23059 2077 23093 2111
rect 23717 2077 23751 2111
rect 23059 2009 23093 2043
rect 23717 2009 23751 2043
rect 23059 1941 23093 1975
rect 21560 1841 21594 1875
rect 21560 1773 21594 1807
rect 23256 1909 23290 1943
rect 23256 1841 23290 1875
rect 23256 1773 23290 1807
rect 23352 1909 23386 1943
rect 23352 1841 23386 1875
rect 23352 1773 23386 1807
rect 23448 1909 23482 1943
rect 23717 1941 23751 1975
rect 23873 2077 23907 2111
rect 23873 2009 23907 2043
rect 23873 1941 23907 1975
rect 24791 2077 24825 2111
rect 24791 2009 24825 2043
rect 24791 1941 24825 1975
rect 24947 2077 24981 2111
rect 25605 2077 25639 2111
rect 24947 2009 24981 2043
rect 25605 2009 25639 2043
rect 24947 1941 24981 1975
rect 23448 1841 23482 1875
rect 23448 1773 23482 1807
rect 25144 1909 25178 1943
rect 25144 1841 25178 1875
rect 25144 1773 25178 1807
rect 25240 1909 25274 1943
rect 25240 1841 25274 1875
rect 25240 1773 25274 1807
rect 25336 1909 25370 1943
rect 25605 1941 25639 1975
rect 25761 2077 25795 2111
rect 25761 2009 25795 2043
rect 25761 1941 25795 1975
rect 26679 2077 26713 2111
rect 26679 2009 26713 2043
rect 26679 1941 26713 1975
rect 26835 2077 26869 2111
rect 27493 2077 27527 2111
rect 26835 2009 26869 2043
rect 27493 2009 27527 2043
rect 26835 1941 26869 1975
rect 25336 1841 25370 1875
rect 25336 1773 25370 1807
rect 27032 1909 27066 1943
rect 27032 1841 27066 1875
rect 27032 1773 27066 1807
rect 27128 1909 27162 1943
rect 27128 1841 27162 1875
rect 27128 1773 27162 1807
rect 27224 1909 27258 1943
rect 27493 1941 27527 1975
rect 27649 2077 27683 2111
rect 27649 2009 27683 2043
rect 27649 1941 27683 1975
rect 28567 2077 28601 2111
rect 28567 2009 28601 2043
rect 28567 1941 28601 1975
rect 28723 2077 28757 2111
rect 29381 2077 29415 2111
rect 28723 2009 28757 2043
rect 29381 2009 29415 2043
rect 28723 1941 28757 1975
rect 27224 1841 27258 1875
rect 27224 1773 27258 1807
rect 28920 1909 28954 1943
rect 28920 1841 28954 1875
rect 28920 1773 28954 1807
rect 29016 1909 29050 1943
rect 29016 1841 29050 1875
rect 29016 1773 29050 1807
rect 29112 1909 29146 1943
rect 29381 1941 29415 1975
rect 29537 2077 29571 2111
rect 29537 2009 29571 2043
rect 29537 1941 29571 1975
rect 30455 2077 30489 2111
rect 30455 2009 30489 2043
rect 30455 1941 30489 1975
rect 30611 2077 30645 2111
rect 31269 2077 31303 2111
rect 30611 2009 30645 2043
rect 31269 2009 31303 2043
rect 30611 1941 30645 1975
rect 29112 1841 29146 1875
rect 29112 1773 29146 1807
rect 30808 1909 30842 1943
rect 30808 1841 30842 1875
rect 30808 1773 30842 1807
rect 30904 1909 30938 1943
rect 30904 1841 30938 1875
rect 30904 1773 30938 1807
rect 31000 1909 31034 1943
rect 31269 1941 31303 1975
rect 31425 2077 31459 2111
rect 31425 2009 31459 2043
rect 31425 1941 31459 1975
rect 32343 2077 32377 2111
rect 32343 2009 32377 2043
rect 32343 1941 32377 1975
rect 32499 2077 32533 2111
rect 33157 2077 33191 2111
rect 32499 2009 32533 2043
rect 33157 2009 33191 2043
rect 32499 1941 32533 1975
rect 31000 1841 31034 1875
rect 31000 1773 31034 1807
rect 32696 1909 32730 1943
rect 32696 1841 32730 1875
rect 32696 1773 32730 1807
rect 32792 1909 32826 1943
rect 32792 1841 32826 1875
rect 32792 1773 32826 1807
rect 32888 1909 32922 1943
rect 33157 1941 33191 1975
rect 33313 2077 33347 2111
rect 33313 2009 33347 2043
rect 33313 1941 33347 1975
rect 34231 2077 34265 2111
rect 34231 2009 34265 2043
rect 34231 1941 34265 1975
rect 34387 2077 34421 2111
rect 35045 2077 35079 2111
rect 34387 2009 34421 2043
rect 35045 2009 35079 2043
rect 34387 1941 34421 1975
rect 32888 1841 32922 1875
rect 32888 1773 32922 1807
rect 34584 1909 34618 1943
rect 34584 1841 34618 1875
rect 34584 1773 34618 1807
rect 34680 1909 34714 1943
rect 34680 1841 34714 1875
rect 34680 1773 34714 1807
rect 34776 1909 34810 1943
rect 35045 1941 35079 1975
rect 35201 2077 35235 2111
rect 35201 2009 35235 2043
rect 35201 1941 35235 1975
rect 36119 2077 36153 2111
rect 36119 2009 36153 2043
rect 36119 1941 36153 1975
rect 36275 2077 36309 2111
rect 36933 2077 36967 2111
rect 36275 2009 36309 2043
rect 36933 2009 36967 2043
rect 36275 1941 36309 1975
rect 34776 1841 34810 1875
rect 34776 1773 34810 1807
rect 36472 1909 36506 1943
rect 36472 1841 36506 1875
rect 36472 1773 36506 1807
rect 36568 1909 36602 1943
rect 36568 1841 36602 1875
rect 36568 1773 36602 1807
rect 36664 1909 36698 1943
rect 36933 1941 36967 1975
rect 37089 2077 37123 2111
rect 37089 2009 37123 2043
rect 37089 1941 37123 1975
rect 38007 2077 38041 2111
rect 38007 2009 38041 2043
rect 38007 1941 38041 1975
rect 38163 2077 38197 2111
rect 38821 2077 38855 2111
rect 38163 2009 38197 2043
rect 38821 2009 38855 2043
rect 38163 1941 38197 1975
rect 36664 1841 36698 1875
rect 36664 1773 36698 1807
rect 38360 1909 38394 1943
rect 38360 1841 38394 1875
rect 38360 1773 38394 1807
rect 38456 1909 38490 1943
rect 38456 1841 38490 1875
rect 38456 1773 38490 1807
rect 38552 1909 38586 1943
rect 38821 1941 38855 1975
rect 38977 2077 39011 2111
rect 38977 2009 39011 2043
rect 38977 1941 39011 1975
rect 39895 2077 39929 2111
rect 39895 2009 39929 2043
rect 39895 1941 39929 1975
rect 40051 2077 40085 2111
rect 40709 2077 40743 2111
rect 40051 2009 40085 2043
rect 40709 2009 40743 2043
rect 40051 1941 40085 1975
rect 38552 1841 38586 1875
rect 38552 1773 38586 1807
rect 40248 1909 40282 1943
rect 40248 1841 40282 1875
rect 40248 1773 40282 1807
rect 40344 1909 40378 1943
rect 40344 1841 40378 1875
rect 40344 1773 40378 1807
rect 40440 1909 40474 1943
rect 40709 1941 40743 1975
rect 40865 2077 40899 2111
rect 40865 2009 40899 2043
rect 40865 1941 40899 1975
rect 41783 2077 41817 2111
rect 41783 2009 41817 2043
rect 41783 1941 41817 1975
rect 41939 2077 41973 2111
rect 42597 2077 42631 2111
rect 41939 2009 41973 2043
rect 42597 2009 42631 2043
rect 41939 1941 41973 1975
rect 40440 1841 40474 1875
rect 40440 1773 40474 1807
rect 42136 1909 42170 1943
rect 42136 1841 42170 1875
rect 42136 1773 42170 1807
rect 42232 1909 42266 1943
rect 42232 1841 42266 1875
rect 42232 1773 42266 1807
rect 42328 1909 42362 1943
rect 42597 1941 42631 1975
rect 42753 2077 42787 2111
rect 42753 2009 42787 2043
rect 42753 1941 42787 1975
rect 43671 2077 43705 2111
rect 43671 2009 43705 2043
rect 43671 1941 43705 1975
rect 43827 2077 43861 2111
rect 44485 2077 44519 2111
rect 43827 2009 43861 2043
rect 44485 2009 44519 2043
rect 43827 1941 43861 1975
rect 42328 1841 42362 1875
rect 42328 1773 42362 1807
rect 44024 1909 44058 1943
rect 44024 1841 44058 1875
rect 44024 1773 44058 1807
rect 44120 1909 44154 1943
rect 44120 1841 44154 1875
rect 44120 1773 44154 1807
rect 44216 1909 44250 1943
rect 44485 1941 44519 1975
rect 44641 2077 44675 2111
rect 44641 2009 44675 2043
rect 44641 1941 44675 1975
rect 45553 2077 45587 2111
rect 45553 2009 45587 2043
rect 45553 1941 45587 1975
rect 45709 2077 45743 2111
rect 46367 2077 46401 2111
rect 45709 2009 45743 2043
rect 46367 2009 46401 2043
rect 45709 1941 45743 1975
rect 44216 1841 44250 1875
rect 44216 1773 44250 1807
rect 45906 1909 45940 1943
rect 45906 1841 45940 1875
rect 45906 1773 45940 1807
rect 46002 1909 46036 1943
rect 46002 1841 46036 1875
rect 46002 1773 46036 1807
rect 46098 1909 46132 1943
rect 46367 1941 46401 1975
rect 46523 2077 46557 2111
rect 46523 2009 46557 2043
rect 46523 1941 46557 1975
rect 47441 2077 47475 2111
rect 47441 2009 47475 2043
rect 47441 1941 47475 1975
rect 47597 2077 47631 2111
rect 48255 2077 48289 2111
rect 47597 2009 47631 2043
rect 48255 2009 48289 2043
rect 47597 1941 47631 1975
rect 46098 1841 46132 1875
rect 46098 1773 46132 1807
rect 47794 1909 47828 1943
rect 47794 1841 47828 1875
rect 47794 1773 47828 1807
rect 47890 1909 47924 1943
rect 47890 1841 47924 1875
rect 47890 1773 47924 1807
rect 47986 1909 48020 1943
rect 48255 1941 48289 1975
rect 48411 2077 48445 2111
rect 48411 2009 48445 2043
rect 48411 1941 48445 1975
rect 49329 2077 49363 2111
rect 49329 2009 49363 2043
rect 49329 1941 49363 1975
rect 49485 2077 49519 2111
rect 50143 2077 50177 2111
rect 49485 2009 49519 2043
rect 50143 2009 50177 2043
rect 49485 1941 49519 1975
rect 47986 1841 48020 1875
rect 47986 1773 48020 1807
rect 49682 1909 49716 1943
rect 49682 1841 49716 1875
rect 49682 1773 49716 1807
rect 49778 1909 49812 1943
rect 49778 1841 49812 1875
rect 49778 1773 49812 1807
rect 49874 1909 49908 1943
rect 50143 1941 50177 1975
rect 50299 2077 50333 2111
rect 50299 2009 50333 2043
rect 50299 1941 50333 1975
rect 51217 2077 51251 2111
rect 51217 2009 51251 2043
rect 51217 1941 51251 1975
rect 51373 2077 51407 2111
rect 52031 2077 52065 2111
rect 51373 2009 51407 2043
rect 52031 2009 52065 2043
rect 51373 1941 51407 1975
rect 49874 1841 49908 1875
rect 49874 1773 49908 1807
rect 51570 1909 51604 1943
rect 51570 1841 51604 1875
rect 51570 1773 51604 1807
rect 51666 1909 51700 1943
rect 51666 1841 51700 1875
rect 51666 1773 51700 1807
rect 51762 1909 51796 1943
rect 52031 1941 52065 1975
rect 52187 2077 52221 2111
rect 52187 2009 52221 2043
rect 52187 1941 52221 1975
rect 53105 2077 53139 2111
rect 53105 2009 53139 2043
rect 53105 1941 53139 1975
rect 53261 2077 53295 2111
rect 53919 2077 53953 2111
rect 53261 2009 53295 2043
rect 53919 2009 53953 2043
rect 53261 1941 53295 1975
rect 51762 1841 51796 1875
rect 51762 1773 51796 1807
rect 53458 1909 53492 1943
rect 53458 1841 53492 1875
rect 53458 1773 53492 1807
rect 53554 1909 53588 1943
rect 53554 1841 53588 1875
rect 53554 1773 53588 1807
rect 53650 1909 53684 1943
rect 53919 1941 53953 1975
rect 54075 2077 54109 2111
rect 54075 2009 54109 2043
rect 54075 1941 54109 1975
rect 54993 2077 55027 2111
rect 54993 2009 55027 2043
rect 54993 1941 55027 1975
rect 55149 2077 55183 2111
rect 55807 2077 55841 2111
rect 55149 2009 55183 2043
rect 55807 2009 55841 2043
rect 55149 1941 55183 1975
rect 53650 1841 53684 1875
rect 53650 1773 53684 1807
rect 55346 1909 55380 1943
rect 55346 1841 55380 1875
rect 55346 1773 55380 1807
rect 55442 1909 55476 1943
rect 55442 1841 55476 1875
rect 55442 1773 55476 1807
rect 55538 1909 55572 1943
rect 55807 1941 55841 1975
rect 55963 2077 55997 2111
rect 55963 2009 55997 2043
rect 55963 1941 55997 1975
rect 56881 2077 56915 2111
rect 56881 2009 56915 2043
rect 56881 1941 56915 1975
rect 57037 2077 57071 2111
rect 57695 2077 57729 2111
rect 57037 2009 57071 2043
rect 57695 2009 57729 2043
rect 57037 1941 57071 1975
rect 55538 1841 55572 1875
rect 55538 1773 55572 1807
rect 57234 1909 57268 1943
rect 57234 1841 57268 1875
rect 57234 1773 57268 1807
rect 57330 1909 57364 1943
rect 57330 1841 57364 1875
rect 57330 1773 57364 1807
rect 57426 1909 57460 1943
rect 57695 1941 57729 1975
rect 57851 2077 57885 2111
rect 57851 2009 57885 2043
rect 57851 1941 57885 1975
rect 58769 2077 58803 2111
rect 58769 2009 58803 2043
rect 58769 1941 58803 1975
rect 58925 2077 58959 2111
rect 59583 2077 59617 2111
rect 58925 2009 58959 2043
rect 59583 2009 59617 2043
rect 58925 1941 58959 1975
rect 57426 1841 57460 1875
rect 57426 1773 57460 1807
rect 59122 1909 59156 1943
rect 59122 1841 59156 1875
rect 59122 1773 59156 1807
rect 59218 1909 59252 1943
rect 59218 1841 59252 1875
rect 59218 1773 59252 1807
rect 59314 1909 59348 1943
rect 59583 1941 59617 1975
rect 59739 2077 59773 2111
rect 59739 2009 59773 2043
rect 59739 1941 59773 1975
rect 59314 1841 59348 1875
rect 59314 1773 59348 1807
rect 116 1023 150 1057
rect 116 955 150 989
rect 116 887 150 921
rect 200 1023 234 1057
rect 200 955 234 989
rect 200 887 234 921
rect 388 1013 422 1047
rect 388 945 422 979
rect 388 877 422 911
rect 476 1013 510 1047
rect 1034 1013 1068 1047
rect 476 945 510 979
rect 476 877 510 911
rect 1034 945 1068 979
rect 604 853 638 887
rect 604 785 638 819
rect 604 717 638 751
rect 700 853 734 887
rect 700 785 734 819
rect 700 717 734 751
rect 796 853 830 887
rect 1034 877 1068 911
rect 1122 1013 1156 1047
rect 1122 945 1156 979
rect 1122 877 1156 911
rect 1312 1031 1346 1065
rect 1312 963 1346 997
rect 1312 895 1346 929
rect 1396 1031 1430 1065
rect 1396 963 1430 997
rect 1396 895 1430 929
rect 1617 1021 1651 1055
rect 1617 953 1651 987
rect 1703 1021 1737 1055
rect 1703 953 1737 987
rect 1789 1021 1823 1055
rect 1789 940 1823 974
rect 2004 1023 2038 1057
rect 2004 955 2038 989
rect 796 785 830 819
rect 2004 887 2038 921
rect 2088 1023 2122 1057
rect 2088 955 2122 989
rect 2088 887 2122 921
rect 2276 1013 2310 1047
rect 2276 945 2310 979
rect 2276 877 2310 911
rect 2364 1013 2398 1047
rect 2922 1013 2956 1047
rect 2364 945 2398 979
rect 2364 877 2398 911
rect 2922 945 2956 979
rect 2492 853 2526 887
rect 796 717 830 751
rect 2492 785 2526 819
rect 2492 717 2526 751
rect 2588 853 2622 887
rect 2588 785 2622 819
rect 2588 717 2622 751
rect 2684 853 2718 887
rect 2922 877 2956 911
rect 3010 1013 3044 1047
rect 3010 945 3044 979
rect 3010 877 3044 911
rect 3200 1031 3234 1065
rect 3200 963 3234 997
rect 3200 895 3234 929
rect 3284 1031 3318 1065
rect 3284 963 3318 997
rect 3284 895 3318 929
rect 3505 1021 3539 1055
rect 3505 953 3539 987
rect 3591 1021 3625 1055
rect 3591 953 3625 987
rect 3677 1021 3711 1055
rect 3677 940 3711 974
rect 3892 1023 3926 1057
rect 3892 955 3926 989
rect 2684 785 2718 819
rect 3892 887 3926 921
rect 3976 1023 4010 1057
rect 3976 955 4010 989
rect 3976 887 4010 921
rect 4164 1013 4198 1047
rect 4164 945 4198 979
rect 4164 877 4198 911
rect 4252 1013 4286 1047
rect 4810 1013 4844 1047
rect 4252 945 4286 979
rect 4252 877 4286 911
rect 4810 945 4844 979
rect 4380 853 4414 887
rect 2684 717 2718 751
rect 4380 785 4414 819
rect 4380 717 4414 751
rect 4476 853 4510 887
rect 4476 785 4510 819
rect 4476 717 4510 751
rect 4572 853 4606 887
rect 4810 877 4844 911
rect 4898 1013 4932 1047
rect 4898 945 4932 979
rect 4898 877 4932 911
rect 5088 1031 5122 1065
rect 5088 963 5122 997
rect 5088 895 5122 929
rect 5172 1031 5206 1065
rect 5172 963 5206 997
rect 5172 895 5206 929
rect 5393 1021 5427 1055
rect 5393 953 5427 987
rect 5479 1021 5513 1055
rect 5479 953 5513 987
rect 5565 1021 5599 1055
rect 5565 940 5599 974
rect 5780 1023 5814 1057
rect 5780 955 5814 989
rect 4572 785 4606 819
rect 5780 887 5814 921
rect 5864 1023 5898 1057
rect 5864 955 5898 989
rect 5864 887 5898 921
rect 6052 1013 6086 1047
rect 6052 945 6086 979
rect 6052 877 6086 911
rect 6140 1013 6174 1047
rect 6698 1013 6732 1047
rect 6140 945 6174 979
rect 6140 877 6174 911
rect 6698 945 6732 979
rect 6268 853 6302 887
rect 4572 717 4606 751
rect 6268 785 6302 819
rect 6268 717 6302 751
rect 6364 853 6398 887
rect 6364 785 6398 819
rect 6364 717 6398 751
rect 6460 853 6494 887
rect 6698 877 6732 911
rect 6786 1013 6820 1047
rect 6786 945 6820 979
rect 6786 877 6820 911
rect 6976 1031 7010 1065
rect 6976 963 7010 997
rect 6976 895 7010 929
rect 7060 1031 7094 1065
rect 7060 963 7094 997
rect 7060 895 7094 929
rect 7281 1021 7315 1055
rect 7281 953 7315 987
rect 7367 1021 7401 1055
rect 7367 953 7401 987
rect 7453 1021 7487 1055
rect 7453 940 7487 974
rect 7668 1023 7702 1057
rect 7668 955 7702 989
rect 6460 785 6494 819
rect 7668 887 7702 921
rect 7752 1023 7786 1057
rect 7752 955 7786 989
rect 7752 887 7786 921
rect 7940 1013 7974 1047
rect 7940 945 7974 979
rect 7940 877 7974 911
rect 8028 1013 8062 1047
rect 8586 1013 8620 1047
rect 8028 945 8062 979
rect 8028 877 8062 911
rect 8586 945 8620 979
rect 8156 853 8190 887
rect 6460 717 6494 751
rect 8156 785 8190 819
rect 8156 717 8190 751
rect 8252 853 8286 887
rect 8252 785 8286 819
rect 8252 717 8286 751
rect 8348 853 8382 887
rect 8586 877 8620 911
rect 8674 1013 8708 1047
rect 8674 945 8708 979
rect 8674 877 8708 911
rect 8864 1031 8898 1065
rect 8864 963 8898 997
rect 8864 895 8898 929
rect 8948 1031 8982 1065
rect 8948 963 8982 997
rect 8948 895 8982 929
rect 9169 1021 9203 1055
rect 9169 953 9203 987
rect 9255 1021 9289 1055
rect 9255 953 9289 987
rect 9341 1021 9375 1055
rect 9341 940 9375 974
rect 9556 1023 9590 1057
rect 9556 955 9590 989
rect 8348 785 8382 819
rect 9556 887 9590 921
rect 9640 1023 9674 1057
rect 9640 955 9674 989
rect 9640 887 9674 921
rect 9828 1013 9862 1047
rect 9828 945 9862 979
rect 9828 877 9862 911
rect 9916 1013 9950 1047
rect 10474 1013 10508 1047
rect 9916 945 9950 979
rect 9916 877 9950 911
rect 10474 945 10508 979
rect 10044 853 10078 887
rect 8348 717 8382 751
rect 10044 785 10078 819
rect 10044 717 10078 751
rect 10140 853 10174 887
rect 10140 785 10174 819
rect 10140 717 10174 751
rect 10236 853 10270 887
rect 10474 877 10508 911
rect 10562 1013 10596 1047
rect 10562 945 10596 979
rect 10562 877 10596 911
rect 10752 1031 10786 1065
rect 10752 963 10786 997
rect 10752 895 10786 929
rect 10836 1031 10870 1065
rect 10836 963 10870 997
rect 10836 895 10870 929
rect 11057 1021 11091 1055
rect 11057 953 11091 987
rect 11143 1021 11177 1055
rect 11143 953 11177 987
rect 11229 1021 11263 1055
rect 11229 940 11263 974
rect 11444 1023 11478 1057
rect 11444 955 11478 989
rect 10236 785 10270 819
rect 11444 887 11478 921
rect 11528 1023 11562 1057
rect 11528 955 11562 989
rect 11528 887 11562 921
rect 11716 1013 11750 1047
rect 11716 945 11750 979
rect 11716 877 11750 911
rect 11804 1013 11838 1047
rect 12362 1013 12396 1047
rect 11804 945 11838 979
rect 11804 877 11838 911
rect 12362 945 12396 979
rect 11932 853 11966 887
rect 10236 717 10270 751
rect 11932 785 11966 819
rect 11932 717 11966 751
rect 12028 853 12062 887
rect 12028 785 12062 819
rect 12028 717 12062 751
rect 12124 853 12158 887
rect 12362 877 12396 911
rect 12450 1013 12484 1047
rect 12450 945 12484 979
rect 12450 877 12484 911
rect 12640 1031 12674 1065
rect 12640 963 12674 997
rect 12640 895 12674 929
rect 12724 1031 12758 1065
rect 12724 963 12758 997
rect 12724 895 12758 929
rect 12945 1021 12979 1055
rect 12945 953 12979 987
rect 13031 1021 13065 1055
rect 13031 953 13065 987
rect 13117 1021 13151 1055
rect 13117 940 13151 974
rect 13332 1023 13366 1057
rect 13332 955 13366 989
rect 12124 785 12158 819
rect 13332 887 13366 921
rect 13416 1023 13450 1057
rect 13416 955 13450 989
rect 13416 887 13450 921
rect 13604 1013 13638 1047
rect 13604 945 13638 979
rect 13604 877 13638 911
rect 13692 1013 13726 1047
rect 14250 1013 14284 1047
rect 13692 945 13726 979
rect 13692 877 13726 911
rect 14250 945 14284 979
rect 13820 853 13854 887
rect 12124 717 12158 751
rect 13820 785 13854 819
rect 13820 717 13854 751
rect 13916 853 13950 887
rect 13916 785 13950 819
rect 13916 717 13950 751
rect 14012 853 14046 887
rect 14250 877 14284 911
rect 14338 1013 14372 1047
rect 14338 945 14372 979
rect 14338 877 14372 911
rect 14528 1031 14562 1065
rect 14528 963 14562 997
rect 14528 895 14562 929
rect 14612 1031 14646 1065
rect 14612 963 14646 997
rect 14612 895 14646 929
rect 14833 1021 14867 1055
rect 14833 953 14867 987
rect 14919 1021 14953 1055
rect 14919 953 14953 987
rect 15005 1021 15039 1055
rect 15005 940 15039 974
rect 15214 1023 15248 1057
rect 15214 955 15248 989
rect 14012 785 14046 819
rect 15214 887 15248 921
rect 15298 1023 15332 1057
rect 15298 955 15332 989
rect 15298 887 15332 921
rect 15486 1013 15520 1047
rect 15486 945 15520 979
rect 15486 877 15520 911
rect 15574 1013 15608 1047
rect 16132 1013 16166 1047
rect 15574 945 15608 979
rect 15574 877 15608 911
rect 16132 945 16166 979
rect 15702 853 15736 887
rect 14012 717 14046 751
rect 15702 785 15736 819
rect 15702 717 15736 751
rect 15798 853 15832 887
rect 15798 785 15832 819
rect 15798 717 15832 751
rect 15894 853 15928 887
rect 16132 877 16166 911
rect 16220 1013 16254 1047
rect 16220 945 16254 979
rect 16220 877 16254 911
rect 16410 1031 16444 1065
rect 16410 963 16444 997
rect 16410 895 16444 929
rect 16494 1031 16528 1065
rect 16494 963 16528 997
rect 16494 895 16528 929
rect 16715 1021 16749 1055
rect 16715 953 16749 987
rect 16801 1021 16835 1055
rect 16801 953 16835 987
rect 16887 1021 16921 1055
rect 16887 940 16921 974
rect 17102 1023 17136 1057
rect 17102 955 17136 989
rect 15894 785 15928 819
rect 17102 887 17136 921
rect 17186 1023 17220 1057
rect 17186 955 17220 989
rect 17186 887 17220 921
rect 17374 1013 17408 1047
rect 17374 945 17408 979
rect 17374 877 17408 911
rect 17462 1013 17496 1047
rect 18020 1013 18054 1047
rect 17462 945 17496 979
rect 17462 877 17496 911
rect 18020 945 18054 979
rect 17590 853 17624 887
rect 15894 717 15928 751
rect 17590 785 17624 819
rect 17590 717 17624 751
rect 17686 853 17720 887
rect 17686 785 17720 819
rect 17686 717 17720 751
rect 17782 853 17816 887
rect 18020 877 18054 911
rect 18108 1013 18142 1047
rect 18108 945 18142 979
rect 18108 877 18142 911
rect 18298 1031 18332 1065
rect 18298 963 18332 997
rect 18298 895 18332 929
rect 18382 1031 18416 1065
rect 18382 963 18416 997
rect 18382 895 18416 929
rect 18603 1021 18637 1055
rect 18603 953 18637 987
rect 18689 1021 18723 1055
rect 18689 953 18723 987
rect 18775 1021 18809 1055
rect 18775 940 18809 974
rect 18990 1023 19024 1057
rect 18990 955 19024 989
rect 17782 785 17816 819
rect 18990 887 19024 921
rect 19074 1023 19108 1057
rect 19074 955 19108 989
rect 19074 887 19108 921
rect 19262 1013 19296 1047
rect 19262 945 19296 979
rect 19262 877 19296 911
rect 19350 1013 19384 1047
rect 19908 1013 19942 1047
rect 19350 945 19384 979
rect 19350 877 19384 911
rect 19908 945 19942 979
rect 19478 853 19512 887
rect 17782 717 17816 751
rect 19478 785 19512 819
rect 19478 717 19512 751
rect 19574 853 19608 887
rect 19574 785 19608 819
rect 19574 717 19608 751
rect 19670 853 19704 887
rect 19908 877 19942 911
rect 19996 1013 20030 1047
rect 19996 945 20030 979
rect 19996 877 20030 911
rect 20186 1031 20220 1065
rect 20186 963 20220 997
rect 20186 895 20220 929
rect 20270 1031 20304 1065
rect 20270 963 20304 997
rect 20270 895 20304 929
rect 20491 1021 20525 1055
rect 20491 953 20525 987
rect 20577 1021 20611 1055
rect 20577 953 20611 987
rect 20663 1021 20697 1055
rect 20663 940 20697 974
rect 20878 1023 20912 1057
rect 20878 955 20912 989
rect 19670 785 19704 819
rect 20878 887 20912 921
rect 20962 1023 20996 1057
rect 20962 955 20996 989
rect 20962 887 20996 921
rect 21150 1013 21184 1047
rect 21150 945 21184 979
rect 21150 877 21184 911
rect 21238 1013 21272 1047
rect 21796 1013 21830 1047
rect 21238 945 21272 979
rect 21238 877 21272 911
rect 21796 945 21830 979
rect 21366 853 21400 887
rect 19670 717 19704 751
rect 21366 785 21400 819
rect 21366 717 21400 751
rect 21462 853 21496 887
rect 21462 785 21496 819
rect 21462 717 21496 751
rect 21558 853 21592 887
rect 21796 877 21830 911
rect 21884 1013 21918 1047
rect 21884 945 21918 979
rect 21884 877 21918 911
rect 22074 1031 22108 1065
rect 22074 963 22108 997
rect 22074 895 22108 929
rect 22158 1031 22192 1065
rect 22158 963 22192 997
rect 22158 895 22192 929
rect 22379 1021 22413 1055
rect 22379 953 22413 987
rect 22465 1021 22499 1055
rect 22465 953 22499 987
rect 22551 1021 22585 1055
rect 22551 940 22585 974
rect 22766 1023 22800 1057
rect 22766 955 22800 989
rect 21558 785 21592 819
rect 22766 887 22800 921
rect 22850 1023 22884 1057
rect 22850 955 22884 989
rect 22850 887 22884 921
rect 23038 1013 23072 1047
rect 23038 945 23072 979
rect 23038 877 23072 911
rect 23126 1013 23160 1047
rect 23684 1013 23718 1047
rect 23126 945 23160 979
rect 23126 877 23160 911
rect 23684 945 23718 979
rect 23254 853 23288 887
rect 21558 717 21592 751
rect 23254 785 23288 819
rect 23254 717 23288 751
rect 23350 853 23384 887
rect 23350 785 23384 819
rect 23350 717 23384 751
rect 23446 853 23480 887
rect 23684 877 23718 911
rect 23772 1013 23806 1047
rect 23772 945 23806 979
rect 23772 877 23806 911
rect 23962 1031 23996 1065
rect 23962 963 23996 997
rect 23962 895 23996 929
rect 24046 1031 24080 1065
rect 24046 963 24080 997
rect 24046 895 24080 929
rect 24267 1021 24301 1055
rect 24267 953 24301 987
rect 24353 1021 24387 1055
rect 24353 953 24387 987
rect 24439 1021 24473 1055
rect 24439 940 24473 974
rect 24654 1023 24688 1057
rect 24654 955 24688 989
rect 23446 785 23480 819
rect 24654 887 24688 921
rect 24738 1023 24772 1057
rect 24738 955 24772 989
rect 24738 887 24772 921
rect 24926 1013 24960 1047
rect 24926 945 24960 979
rect 24926 877 24960 911
rect 25014 1013 25048 1047
rect 25572 1013 25606 1047
rect 25014 945 25048 979
rect 25014 877 25048 911
rect 25572 945 25606 979
rect 25142 853 25176 887
rect 23446 717 23480 751
rect 25142 785 25176 819
rect 25142 717 25176 751
rect 25238 853 25272 887
rect 25238 785 25272 819
rect 25238 717 25272 751
rect 25334 853 25368 887
rect 25572 877 25606 911
rect 25660 1013 25694 1047
rect 25660 945 25694 979
rect 25660 877 25694 911
rect 25850 1031 25884 1065
rect 25850 963 25884 997
rect 25850 895 25884 929
rect 25934 1031 25968 1065
rect 25934 963 25968 997
rect 25934 895 25968 929
rect 26155 1021 26189 1055
rect 26155 953 26189 987
rect 26241 1021 26275 1055
rect 26241 953 26275 987
rect 26327 1021 26361 1055
rect 26327 940 26361 974
rect 26542 1023 26576 1057
rect 26542 955 26576 989
rect 25334 785 25368 819
rect 26542 887 26576 921
rect 26626 1023 26660 1057
rect 26626 955 26660 989
rect 26626 887 26660 921
rect 26814 1013 26848 1047
rect 26814 945 26848 979
rect 26814 877 26848 911
rect 26902 1013 26936 1047
rect 27460 1013 27494 1047
rect 26902 945 26936 979
rect 26902 877 26936 911
rect 27460 945 27494 979
rect 27030 853 27064 887
rect 25334 717 25368 751
rect 27030 785 27064 819
rect 27030 717 27064 751
rect 27126 853 27160 887
rect 27126 785 27160 819
rect 27126 717 27160 751
rect 27222 853 27256 887
rect 27460 877 27494 911
rect 27548 1013 27582 1047
rect 27548 945 27582 979
rect 27548 877 27582 911
rect 27738 1031 27772 1065
rect 27738 963 27772 997
rect 27738 895 27772 929
rect 27822 1031 27856 1065
rect 27822 963 27856 997
rect 27822 895 27856 929
rect 28043 1021 28077 1055
rect 28043 953 28077 987
rect 28129 1021 28163 1055
rect 28129 953 28163 987
rect 28215 1021 28249 1055
rect 28215 940 28249 974
rect 28430 1023 28464 1057
rect 28430 955 28464 989
rect 27222 785 27256 819
rect 28430 887 28464 921
rect 28514 1023 28548 1057
rect 28514 955 28548 989
rect 28514 887 28548 921
rect 28702 1013 28736 1047
rect 28702 945 28736 979
rect 28702 877 28736 911
rect 28790 1013 28824 1047
rect 29348 1013 29382 1047
rect 28790 945 28824 979
rect 28790 877 28824 911
rect 29348 945 29382 979
rect 28918 853 28952 887
rect 27222 717 27256 751
rect 28918 785 28952 819
rect 28918 717 28952 751
rect 29014 853 29048 887
rect 29014 785 29048 819
rect 29014 717 29048 751
rect 29110 853 29144 887
rect 29348 877 29382 911
rect 29436 1013 29470 1047
rect 29436 945 29470 979
rect 29436 877 29470 911
rect 29626 1031 29660 1065
rect 29626 963 29660 997
rect 29626 895 29660 929
rect 29710 1031 29744 1065
rect 29710 963 29744 997
rect 29710 895 29744 929
rect 29931 1021 29965 1055
rect 29931 953 29965 987
rect 30017 1021 30051 1055
rect 30017 953 30051 987
rect 30103 1021 30137 1055
rect 30103 940 30137 974
rect 30318 1023 30352 1057
rect 30318 955 30352 989
rect 29110 785 29144 819
rect 30318 887 30352 921
rect 30402 1023 30436 1057
rect 30402 955 30436 989
rect 30402 887 30436 921
rect 30590 1013 30624 1047
rect 30590 945 30624 979
rect 30590 877 30624 911
rect 30678 1013 30712 1047
rect 31236 1013 31270 1047
rect 30678 945 30712 979
rect 30678 877 30712 911
rect 31236 945 31270 979
rect 30806 853 30840 887
rect 29110 717 29144 751
rect 30806 785 30840 819
rect 30806 717 30840 751
rect 30902 853 30936 887
rect 30902 785 30936 819
rect 30902 717 30936 751
rect 30998 853 31032 887
rect 31236 877 31270 911
rect 31324 1013 31358 1047
rect 31324 945 31358 979
rect 31324 877 31358 911
rect 31514 1031 31548 1065
rect 31514 963 31548 997
rect 31514 895 31548 929
rect 31598 1031 31632 1065
rect 31598 963 31632 997
rect 31598 895 31632 929
rect 31819 1021 31853 1055
rect 31819 953 31853 987
rect 31905 1021 31939 1055
rect 31905 953 31939 987
rect 31991 1021 32025 1055
rect 31991 940 32025 974
rect 32206 1023 32240 1057
rect 32206 955 32240 989
rect 30998 785 31032 819
rect 32206 887 32240 921
rect 32290 1023 32324 1057
rect 32290 955 32324 989
rect 32290 887 32324 921
rect 32478 1013 32512 1047
rect 32478 945 32512 979
rect 32478 877 32512 911
rect 32566 1013 32600 1047
rect 33124 1013 33158 1047
rect 32566 945 32600 979
rect 32566 877 32600 911
rect 33124 945 33158 979
rect 32694 853 32728 887
rect 30998 717 31032 751
rect 32694 785 32728 819
rect 32694 717 32728 751
rect 32790 853 32824 887
rect 32790 785 32824 819
rect 32790 717 32824 751
rect 32886 853 32920 887
rect 33124 877 33158 911
rect 33212 1013 33246 1047
rect 33212 945 33246 979
rect 33212 877 33246 911
rect 33402 1031 33436 1065
rect 33402 963 33436 997
rect 33402 895 33436 929
rect 33486 1031 33520 1065
rect 33486 963 33520 997
rect 33486 895 33520 929
rect 33707 1021 33741 1055
rect 33707 953 33741 987
rect 33793 1021 33827 1055
rect 33793 953 33827 987
rect 33879 1021 33913 1055
rect 33879 940 33913 974
rect 34094 1023 34128 1057
rect 34094 955 34128 989
rect 32886 785 32920 819
rect 34094 887 34128 921
rect 34178 1023 34212 1057
rect 34178 955 34212 989
rect 34178 887 34212 921
rect 34366 1013 34400 1047
rect 34366 945 34400 979
rect 34366 877 34400 911
rect 34454 1013 34488 1047
rect 35012 1013 35046 1047
rect 34454 945 34488 979
rect 34454 877 34488 911
rect 35012 945 35046 979
rect 34582 853 34616 887
rect 32886 717 32920 751
rect 34582 785 34616 819
rect 34582 717 34616 751
rect 34678 853 34712 887
rect 34678 785 34712 819
rect 34678 717 34712 751
rect 34774 853 34808 887
rect 35012 877 35046 911
rect 35100 1013 35134 1047
rect 35100 945 35134 979
rect 35100 877 35134 911
rect 35290 1031 35324 1065
rect 35290 963 35324 997
rect 35290 895 35324 929
rect 35374 1031 35408 1065
rect 35374 963 35408 997
rect 35374 895 35408 929
rect 35595 1021 35629 1055
rect 35595 953 35629 987
rect 35681 1021 35715 1055
rect 35681 953 35715 987
rect 35767 1021 35801 1055
rect 35767 940 35801 974
rect 35982 1023 36016 1057
rect 35982 955 36016 989
rect 34774 785 34808 819
rect 35982 887 36016 921
rect 36066 1023 36100 1057
rect 36066 955 36100 989
rect 36066 887 36100 921
rect 36254 1013 36288 1047
rect 36254 945 36288 979
rect 36254 877 36288 911
rect 36342 1013 36376 1047
rect 36900 1013 36934 1047
rect 36342 945 36376 979
rect 36342 877 36376 911
rect 36900 945 36934 979
rect 36470 853 36504 887
rect 34774 717 34808 751
rect 36470 785 36504 819
rect 36470 717 36504 751
rect 36566 853 36600 887
rect 36566 785 36600 819
rect 36566 717 36600 751
rect 36662 853 36696 887
rect 36900 877 36934 911
rect 36988 1013 37022 1047
rect 36988 945 37022 979
rect 36988 877 37022 911
rect 37178 1031 37212 1065
rect 37178 963 37212 997
rect 37178 895 37212 929
rect 37262 1031 37296 1065
rect 37262 963 37296 997
rect 37262 895 37296 929
rect 37483 1021 37517 1055
rect 37483 953 37517 987
rect 37569 1021 37603 1055
rect 37569 953 37603 987
rect 37655 1021 37689 1055
rect 37655 940 37689 974
rect 37870 1023 37904 1057
rect 37870 955 37904 989
rect 36662 785 36696 819
rect 37870 887 37904 921
rect 37954 1023 37988 1057
rect 37954 955 37988 989
rect 37954 887 37988 921
rect 38142 1013 38176 1047
rect 38142 945 38176 979
rect 38142 877 38176 911
rect 38230 1013 38264 1047
rect 38788 1013 38822 1047
rect 38230 945 38264 979
rect 38230 877 38264 911
rect 38788 945 38822 979
rect 38358 853 38392 887
rect 36662 717 36696 751
rect 38358 785 38392 819
rect 38358 717 38392 751
rect 38454 853 38488 887
rect 38454 785 38488 819
rect 38454 717 38488 751
rect 38550 853 38584 887
rect 38788 877 38822 911
rect 38876 1013 38910 1047
rect 38876 945 38910 979
rect 38876 877 38910 911
rect 39066 1031 39100 1065
rect 39066 963 39100 997
rect 39066 895 39100 929
rect 39150 1031 39184 1065
rect 39150 963 39184 997
rect 39150 895 39184 929
rect 39371 1021 39405 1055
rect 39371 953 39405 987
rect 39457 1021 39491 1055
rect 39457 953 39491 987
rect 39543 1021 39577 1055
rect 39543 940 39577 974
rect 39758 1023 39792 1057
rect 39758 955 39792 989
rect 38550 785 38584 819
rect 39758 887 39792 921
rect 39842 1023 39876 1057
rect 39842 955 39876 989
rect 39842 887 39876 921
rect 40030 1013 40064 1047
rect 40030 945 40064 979
rect 40030 877 40064 911
rect 40118 1013 40152 1047
rect 40676 1013 40710 1047
rect 40118 945 40152 979
rect 40118 877 40152 911
rect 40676 945 40710 979
rect 40246 853 40280 887
rect 38550 717 38584 751
rect 40246 785 40280 819
rect 40246 717 40280 751
rect 40342 853 40376 887
rect 40342 785 40376 819
rect 40342 717 40376 751
rect 40438 853 40472 887
rect 40676 877 40710 911
rect 40764 1013 40798 1047
rect 40764 945 40798 979
rect 40764 877 40798 911
rect 40954 1031 40988 1065
rect 40954 963 40988 997
rect 40954 895 40988 929
rect 41038 1031 41072 1065
rect 41038 963 41072 997
rect 41038 895 41072 929
rect 41259 1021 41293 1055
rect 41259 953 41293 987
rect 41345 1021 41379 1055
rect 41345 953 41379 987
rect 41431 1021 41465 1055
rect 41431 940 41465 974
rect 41646 1023 41680 1057
rect 41646 955 41680 989
rect 40438 785 40472 819
rect 41646 887 41680 921
rect 41730 1023 41764 1057
rect 41730 955 41764 989
rect 41730 887 41764 921
rect 41918 1013 41952 1047
rect 41918 945 41952 979
rect 41918 877 41952 911
rect 42006 1013 42040 1047
rect 42564 1013 42598 1047
rect 42006 945 42040 979
rect 42006 877 42040 911
rect 42564 945 42598 979
rect 42134 853 42168 887
rect 40438 717 40472 751
rect 42134 785 42168 819
rect 42134 717 42168 751
rect 42230 853 42264 887
rect 42230 785 42264 819
rect 42230 717 42264 751
rect 42326 853 42360 887
rect 42564 877 42598 911
rect 42652 1013 42686 1047
rect 42652 945 42686 979
rect 42652 877 42686 911
rect 42842 1031 42876 1065
rect 42842 963 42876 997
rect 42842 895 42876 929
rect 42926 1031 42960 1065
rect 42926 963 42960 997
rect 42926 895 42960 929
rect 43147 1021 43181 1055
rect 43147 953 43181 987
rect 43233 1021 43267 1055
rect 43233 953 43267 987
rect 43319 1021 43353 1055
rect 43319 940 43353 974
rect 43534 1023 43568 1057
rect 43534 955 43568 989
rect 42326 785 42360 819
rect 43534 887 43568 921
rect 43618 1023 43652 1057
rect 43618 955 43652 989
rect 43618 887 43652 921
rect 43806 1013 43840 1047
rect 43806 945 43840 979
rect 43806 877 43840 911
rect 43894 1013 43928 1047
rect 44452 1013 44486 1047
rect 43894 945 43928 979
rect 43894 877 43928 911
rect 44452 945 44486 979
rect 44022 853 44056 887
rect 42326 717 42360 751
rect 44022 785 44056 819
rect 44022 717 44056 751
rect 44118 853 44152 887
rect 44118 785 44152 819
rect 44118 717 44152 751
rect 44214 853 44248 887
rect 44452 877 44486 911
rect 44540 1013 44574 1047
rect 44540 945 44574 979
rect 44540 877 44574 911
rect 44730 1031 44764 1065
rect 44730 963 44764 997
rect 44730 895 44764 929
rect 44814 1031 44848 1065
rect 44814 963 44848 997
rect 44814 895 44848 929
rect 45035 1021 45069 1055
rect 45035 953 45069 987
rect 45121 1021 45155 1055
rect 45121 953 45155 987
rect 45207 1021 45241 1055
rect 45207 940 45241 974
rect 45416 1023 45450 1057
rect 45416 955 45450 989
rect 44214 785 44248 819
rect 45416 887 45450 921
rect 45500 1023 45534 1057
rect 45500 955 45534 989
rect 45500 887 45534 921
rect 45688 1013 45722 1047
rect 45688 945 45722 979
rect 45688 877 45722 911
rect 45776 1013 45810 1047
rect 46334 1013 46368 1047
rect 45776 945 45810 979
rect 45776 877 45810 911
rect 46334 945 46368 979
rect 45904 853 45938 887
rect 44214 717 44248 751
rect 45904 785 45938 819
rect 45904 717 45938 751
rect 46000 853 46034 887
rect 46000 785 46034 819
rect 46000 717 46034 751
rect 46096 853 46130 887
rect 46334 877 46368 911
rect 46422 1013 46456 1047
rect 46422 945 46456 979
rect 46422 877 46456 911
rect 46612 1031 46646 1065
rect 46612 963 46646 997
rect 46612 895 46646 929
rect 46696 1031 46730 1065
rect 46696 963 46730 997
rect 46696 895 46730 929
rect 46917 1021 46951 1055
rect 46917 953 46951 987
rect 47003 1021 47037 1055
rect 47003 953 47037 987
rect 47089 1021 47123 1055
rect 47089 940 47123 974
rect 47304 1023 47338 1057
rect 47304 955 47338 989
rect 46096 785 46130 819
rect 47304 887 47338 921
rect 47388 1023 47422 1057
rect 47388 955 47422 989
rect 47388 887 47422 921
rect 47576 1013 47610 1047
rect 47576 945 47610 979
rect 47576 877 47610 911
rect 47664 1013 47698 1047
rect 48222 1013 48256 1047
rect 47664 945 47698 979
rect 47664 877 47698 911
rect 48222 945 48256 979
rect 47792 853 47826 887
rect 46096 717 46130 751
rect 47792 785 47826 819
rect 47792 717 47826 751
rect 47888 853 47922 887
rect 47888 785 47922 819
rect 47888 717 47922 751
rect 47984 853 48018 887
rect 48222 877 48256 911
rect 48310 1013 48344 1047
rect 48310 945 48344 979
rect 48310 877 48344 911
rect 48500 1031 48534 1065
rect 48500 963 48534 997
rect 48500 895 48534 929
rect 48584 1031 48618 1065
rect 48584 963 48618 997
rect 48584 895 48618 929
rect 48805 1021 48839 1055
rect 48805 953 48839 987
rect 48891 1021 48925 1055
rect 48891 953 48925 987
rect 48977 1021 49011 1055
rect 48977 940 49011 974
rect 49192 1023 49226 1057
rect 49192 955 49226 989
rect 47984 785 48018 819
rect 49192 887 49226 921
rect 49276 1023 49310 1057
rect 49276 955 49310 989
rect 49276 887 49310 921
rect 49464 1013 49498 1047
rect 49464 945 49498 979
rect 49464 877 49498 911
rect 49552 1013 49586 1047
rect 50110 1013 50144 1047
rect 49552 945 49586 979
rect 49552 877 49586 911
rect 50110 945 50144 979
rect 49680 853 49714 887
rect 47984 717 48018 751
rect 49680 785 49714 819
rect 49680 717 49714 751
rect 49776 853 49810 887
rect 49776 785 49810 819
rect 49776 717 49810 751
rect 49872 853 49906 887
rect 50110 877 50144 911
rect 50198 1013 50232 1047
rect 50198 945 50232 979
rect 50198 877 50232 911
rect 50388 1031 50422 1065
rect 50388 963 50422 997
rect 50388 895 50422 929
rect 50472 1031 50506 1065
rect 50472 963 50506 997
rect 50472 895 50506 929
rect 50693 1021 50727 1055
rect 50693 953 50727 987
rect 50779 1021 50813 1055
rect 50779 953 50813 987
rect 50865 1021 50899 1055
rect 50865 940 50899 974
rect 51080 1023 51114 1057
rect 51080 955 51114 989
rect 49872 785 49906 819
rect 51080 887 51114 921
rect 51164 1023 51198 1057
rect 51164 955 51198 989
rect 51164 887 51198 921
rect 51352 1013 51386 1047
rect 51352 945 51386 979
rect 51352 877 51386 911
rect 51440 1013 51474 1047
rect 51998 1013 52032 1047
rect 51440 945 51474 979
rect 51440 877 51474 911
rect 51998 945 52032 979
rect 51568 853 51602 887
rect 49872 717 49906 751
rect 51568 785 51602 819
rect 51568 717 51602 751
rect 51664 853 51698 887
rect 51664 785 51698 819
rect 51664 717 51698 751
rect 51760 853 51794 887
rect 51998 877 52032 911
rect 52086 1013 52120 1047
rect 52086 945 52120 979
rect 52086 877 52120 911
rect 52276 1031 52310 1065
rect 52276 963 52310 997
rect 52276 895 52310 929
rect 52360 1031 52394 1065
rect 52360 963 52394 997
rect 52360 895 52394 929
rect 52581 1021 52615 1055
rect 52581 953 52615 987
rect 52667 1021 52701 1055
rect 52667 953 52701 987
rect 52753 1021 52787 1055
rect 52753 940 52787 974
rect 52968 1023 53002 1057
rect 52968 955 53002 989
rect 51760 785 51794 819
rect 52968 887 53002 921
rect 53052 1023 53086 1057
rect 53052 955 53086 989
rect 53052 887 53086 921
rect 53240 1013 53274 1047
rect 53240 945 53274 979
rect 53240 877 53274 911
rect 53328 1013 53362 1047
rect 53886 1013 53920 1047
rect 53328 945 53362 979
rect 53328 877 53362 911
rect 53886 945 53920 979
rect 53456 853 53490 887
rect 51760 717 51794 751
rect 53456 785 53490 819
rect 53456 717 53490 751
rect 53552 853 53586 887
rect 53552 785 53586 819
rect 53552 717 53586 751
rect 53648 853 53682 887
rect 53886 877 53920 911
rect 53974 1013 54008 1047
rect 53974 945 54008 979
rect 53974 877 54008 911
rect 54164 1031 54198 1065
rect 54164 963 54198 997
rect 54164 895 54198 929
rect 54248 1031 54282 1065
rect 54248 963 54282 997
rect 54248 895 54282 929
rect 54469 1021 54503 1055
rect 54469 953 54503 987
rect 54555 1021 54589 1055
rect 54555 953 54589 987
rect 54641 1021 54675 1055
rect 54641 940 54675 974
rect 54856 1023 54890 1057
rect 54856 955 54890 989
rect 53648 785 53682 819
rect 54856 887 54890 921
rect 54940 1023 54974 1057
rect 54940 955 54974 989
rect 54940 887 54974 921
rect 55128 1013 55162 1047
rect 55128 945 55162 979
rect 55128 877 55162 911
rect 55216 1013 55250 1047
rect 55774 1013 55808 1047
rect 55216 945 55250 979
rect 55216 877 55250 911
rect 55774 945 55808 979
rect 55344 853 55378 887
rect 53648 717 53682 751
rect 55344 785 55378 819
rect 55344 717 55378 751
rect 55440 853 55474 887
rect 55440 785 55474 819
rect 55440 717 55474 751
rect 55536 853 55570 887
rect 55774 877 55808 911
rect 55862 1013 55896 1047
rect 55862 945 55896 979
rect 55862 877 55896 911
rect 56052 1031 56086 1065
rect 56052 963 56086 997
rect 56052 895 56086 929
rect 56136 1031 56170 1065
rect 56136 963 56170 997
rect 56136 895 56170 929
rect 56357 1021 56391 1055
rect 56357 953 56391 987
rect 56443 1021 56477 1055
rect 56443 953 56477 987
rect 56529 1021 56563 1055
rect 56529 940 56563 974
rect 56744 1023 56778 1057
rect 56744 955 56778 989
rect 55536 785 55570 819
rect 56744 887 56778 921
rect 56828 1023 56862 1057
rect 56828 955 56862 989
rect 56828 887 56862 921
rect 57016 1013 57050 1047
rect 57016 945 57050 979
rect 57016 877 57050 911
rect 57104 1013 57138 1047
rect 57662 1013 57696 1047
rect 57104 945 57138 979
rect 57104 877 57138 911
rect 57662 945 57696 979
rect 57232 853 57266 887
rect 55536 717 55570 751
rect 57232 785 57266 819
rect 57232 717 57266 751
rect 57328 853 57362 887
rect 57328 785 57362 819
rect 57328 717 57362 751
rect 57424 853 57458 887
rect 57662 877 57696 911
rect 57750 1013 57784 1047
rect 57750 945 57784 979
rect 57750 877 57784 911
rect 57940 1031 57974 1065
rect 57940 963 57974 997
rect 57940 895 57974 929
rect 58024 1031 58058 1065
rect 58024 963 58058 997
rect 58024 895 58058 929
rect 58245 1021 58279 1055
rect 58245 953 58279 987
rect 58331 1021 58365 1055
rect 58331 953 58365 987
rect 58417 1021 58451 1055
rect 58417 940 58451 974
rect 58632 1023 58666 1057
rect 58632 955 58666 989
rect 57424 785 57458 819
rect 58632 887 58666 921
rect 58716 1023 58750 1057
rect 58716 955 58750 989
rect 58716 887 58750 921
rect 58904 1013 58938 1047
rect 58904 945 58938 979
rect 58904 877 58938 911
rect 58992 1013 59026 1047
rect 59550 1013 59584 1047
rect 58992 945 59026 979
rect 58992 877 59026 911
rect 59550 945 59584 979
rect 59120 853 59154 887
rect 57424 717 57458 751
rect 59120 785 59154 819
rect 59120 717 59154 751
rect 59216 853 59250 887
rect 59216 785 59250 819
rect 59216 717 59250 751
rect 59312 853 59346 887
rect 59550 877 59584 911
rect 59638 1013 59672 1047
rect 59638 945 59672 979
rect 59638 877 59672 911
rect 59828 1031 59862 1065
rect 59828 963 59862 997
rect 59828 895 59862 929
rect 59912 1031 59946 1065
rect 59912 963 59946 997
rect 59912 895 59946 929
rect 60133 1021 60167 1055
rect 60133 953 60167 987
rect 60219 1021 60253 1055
rect 60219 953 60253 987
rect 60305 1021 60339 1055
rect 60305 940 60339 974
rect 59312 785 59346 819
rect 59312 717 59346 751
<< psubdiff >>
rect 654 7244 814 7252
rect 654 7210 723 7244
rect 757 7210 814 7244
rect 654 7204 814 7210
rect 2542 7244 2702 7252
rect 2542 7210 2611 7244
rect 2645 7210 2702 7244
rect 2542 7204 2702 7210
rect 4430 7244 4590 7252
rect 4430 7210 4499 7244
rect 4533 7210 4590 7244
rect 4430 7204 4590 7210
rect 6318 7244 6478 7252
rect 6318 7210 6387 7244
rect 6421 7210 6478 7244
rect 6318 7204 6478 7210
rect 8206 7244 8366 7252
rect 8206 7210 8275 7244
rect 8309 7210 8366 7244
rect 8206 7204 8366 7210
rect 10094 7244 10254 7252
rect 10094 7210 10163 7244
rect 10197 7210 10254 7244
rect 10094 7204 10254 7210
rect 11982 7244 12142 7252
rect 11982 7210 12051 7244
rect 12085 7210 12142 7244
rect 11982 7204 12142 7210
rect 13870 7244 14030 7252
rect 13870 7210 13939 7244
rect 13973 7210 14030 7244
rect 13870 7204 14030 7210
rect 15752 7244 15912 7252
rect 15752 7210 15821 7244
rect 15855 7210 15912 7244
rect 15752 7204 15912 7210
rect 17640 7244 17800 7252
rect 17640 7210 17709 7244
rect 17743 7210 17800 7244
rect 17640 7204 17800 7210
rect 19528 7244 19688 7252
rect 19528 7210 19597 7244
rect 19631 7210 19688 7244
rect 19528 7204 19688 7210
rect 21416 7244 21576 7252
rect 21416 7210 21485 7244
rect 21519 7210 21576 7244
rect 21416 7204 21576 7210
rect 23304 7244 23464 7252
rect 23304 7210 23373 7244
rect 23407 7210 23464 7244
rect 23304 7204 23464 7210
rect 25192 7244 25352 7252
rect 25192 7210 25261 7244
rect 25295 7210 25352 7244
rect 25192 7204 25352 7210
rect 27080 7244 27240 7252
rect 27080 7210 27149 7244
rect 27183 7210 27240 7244
rect 27080 7204 27240 7210
rect 28968 7244 29128 7252
rect 28968 7210 29037 7244
rect 29071 7210 29128 7244
rect 28968 7204 29128 7210
rect 30856 7244 31016 7252
rect 30856 7210 30925 7244
rect 30959 7210 31016 7244
rect 30856 7204 31016 7210
rect 32744 7244 32904 7252
rect 32744 7210 32813 7244
rect 32847 7210 32904 7244
rect 32744 7204 32904 7210
rect 34632 7244 34792 7252
rect 34632 7210 34701 7244
rect 34735 7210 34792 7244
rect 34632 7204 34792 7210
rect 36520 7244 36680 7252
rect 36520 7210 36589 7244
rect 36623 7210 36680 7244
rect 36520 7204 36680 7210
rect 38408 7244 38568 7252
rect 38408 7210 38477 7244
rect 38511 7210 38568 7244
rect 38408 7204 38568 7210
rect 40296 7244 40456 7252
rect 40296 7210 40365 7244
rect 40399 7210 40456 7244
rect 40296 7204 40456 7210
rect 42184 7244 42344 7252
rect 42184 7210 42253 7244
rect 42287 7210 42344 7244
rect 42184 7204 42344 7210
rect 44072 7244 44232 7252
rect 44072 7210 44141 7244
rect 44175 7210 44232 7244
rect 44072 7204 44232 7210
rect 45954 7244 46114 7252
rect 45954 7210 46023 7244
rect 46057 7210 46114 7244
rect 45954 7204 46114 7210
rect 47842 7244 48002 7252
rect 47842 7210 47911 7244
rect 47945 7210 48002 7244
rect 47842 7204 48002 7210
rect 49730 7244 49890 7252
rect 49730 7210 49799 7244
rect 49833 7210 49890 7244
rect 49730 7204 49890 7210
rect 51618 7244 51778 7252
rect 51618 7210 51687 7244
rect 51721 7210 51778 7244
rect 51618 7204 51778 7210
rect 53506 7244 53666 7252
rect 53506 7210 53575 7244
rect 53609 7210 53666 7244
rect 53506 7204 53666 7210
rect 55394 7244 55554 7252
rect 55394 7210 55463 7244
rect 55497 7210 55554 7244
rect 55394 7204 55554 7210
rect 57282 7244 57442 7252
rect 57282 7210 57351 7244
rect 57385 7210 57442 7244
rect 57282 7204 57442 7210
rect 59170 7244 59330 7252
rect 59170 7210 59239 7244
rect 59273 7210 59330 7244
rect 59170 7204 59330 7210
rect 652 6188 812 6196
rect 652 6154 721 6188
rect 755 6154 812 6188
rect 652 6148 812 6154
rect 2540 6188 2700 6196
rect 2540 6154 2609 6188
rect 2643 6154 2700 6188
rect 2540 6148 2700 6154
rect 4428 6188 4588 6196
rect 4428 6154 4497 6188
rect 4531 6154 4588 6188
rect 4428 6148 4588 6154
rect 6316 6188 6476 6196
rect 6316 6154 6385 6188
rect 6419 6154 6476 6188
rect 6316 6148 6476 6154
rect 8204 6188 8364 6196
rect 8204 6154 8273 6188
rect 8307 6154 8364 6188
rect 8204 6148 8364 6154
rect 10092 6188 10252 6196
rect 10092 6154 10161 6188
rect 10195 6154 10252 6188
rect 10092 6148 10252 6154
rect 11980 6188 12140 6196
rect 11980 6154 12049 6188
rect 12083 6154 12140 6188
rect 11980 6148 12140 6154
rect 13868 6188 14028 6196
rect 13868 6154 13937 6188
rect 13971 6154 14028 6188
rect 13868 6148 14028 6154
rect 15750 6188 15910 6196
rect 15750 6154 15819 6188
rect 15853 6154 15910 6188
rect 15750 6148 15910 6154
rect 17638 6188 17798 6196
rect 17638 6154 17707 6188
rect 17741 6154 17798 6188
rect 17638 6148 17798 6154
rect 19526 6188 19686 6196
rect 19526 6154 19595 6188
rect 19629 6154 19686 6188
rect 19526 6148 19686 6154
rect 21414 6188 21574 6196
rect 21414 6154 21483 6188
rect 21517 6154 21574 6188
rect 21414 6148 21574 6154
rect 23302 6188 23462 6196
rect 23302 6154 23371 6188
rect 23405 6154 23462 6188
rect 23302 6148 23462 6154
rect 25190 6188 25350 6196
rect 25190 6154 25259 6188
rect 25293 6154 25350 6188
rect 25190 6148 25350 6154
rect 27078 6188 27238 6196
rect 27078 6154 27147 6188
rect 27181 6154 27238 6188
rect 27078 6148 27238 6154
rect 28966 6188 29126 6196
rect 28966 6154 29035 6188
rect 29069 6154 29126 6188
rect 28966 6148 29126 6154
rect 30854 6188 31014 6196
rect 30854 6154 30923 6188
rect 30957 6154 31014 6188
rect 30854 6148 31014 6154
rect 32742 6188 32902 6196
rect 32742 6154 32811 6188
rect 32845 6154 32902 6188
rect 32742 6148 32902 6154
rect 34630 6188 34790 6196
rect 34630 6154 34699 6188
rect 34733 6154 34790 6188
rect 34630 6148 34790 6154
rect 36518 6188 36678 6196
rect 36518 6154 36587 6188
rect 36621 6154 36678 6188
rect 36518 6148 36678 6154
rect 38406 6188 38566 6196
rect 38406 6154 38475 6188
rect 38509 6154 38566 6188
rect 38406 6148 38566 6154
rect 40294 6188 40454 6196
rect 40294 6154 40363 6188
rect 40397 6154 40454 6188
rect 40294 6148 40454 6154
rect 42182 6188 42342 6196
rect 42182 6154 42251 6188
rect 42285 6154 42342 6188
rect 42182 6148 42342 6154
rect 44070 6188 44230 6196
rect 44070 6154 44139 6188
rect 44173 6154 44230 6188
rect 44070 6148 44230 6154
rect 45952 6188 46112 6196
rect 45952 6154 46021 6188
rect 46055 6154 46112 6188
rect 45952 6148 46112 6154
rect 47840 6188 48000 6196
rect 47840 6154 47909 6188
rect 47943 6154 48000 6188
rect 47840 6148 48000 6154
rect 49728 6188 49888 6196
rect 49728 6154 49797 6188
rect 49831 6154 49888 6188
rect 49728 6148 49888 6154
rect 51616 6188 51776 6196
rect 51616 6154 51685 6188
rect 51719 6154 51776 6188
rect 51616 6148 51776 6154
rect 53504 6188 53664 6196
rect 53504 6154 53573 6188
rect 53607 6154 53664 6188
rect 53504 6148 53664 6154
rect 55392 6188 55552 6196
rect 55392 6154 55461 6188
rect 55495 6154 55552 6188
rect 55392 6148 55552 6154
rect 57280 6188 57440 6196
rect 57280 6154 57349 6188
rect 57383 6154 57440 6188
rect 57280 6148 57440 6154
rect 59168 6188 59328 6196
rect 59168 6154 59237 6188
rect 59271 6154 59328 6188
rect 59168 6148 59328 6154
rect 654 1286 814 1292
rect 654 1252 711 1286
rect 745 1252 814 1286
rect 654 1244 814 1252
rect 2542 1286 2702 1292
rect 2542 1252 2599 1286
rect 2633 1252 2702 1286
rect 2542 1244 2702 1252
rect 4430 1286 4590 1292
rect 4430 1252 4487 1286
rect 4521 1252 4590 1286
rect 4430 1244 4590 1252
rect 6318 1286 6478 1292
rect 6318 1252 6375 1286
rect 6409 1252 6478 1286
rect 6318 1244 6478 1252
rect 8206 1286 8366 1292
rect 8206 1252 8263 1286
rect 8297 1252 8366 1286
rect 8206 1244 8366 1252
rect 10094 1286 10254 1292
rect 10094 1252 10151 1286
rect 10185 1252 10254 1286
rect 10094 1244 10254 1252
rect 11982 1286 12142 1292
rect 11982 1252 12039 1286
rect 12073 1252 12142 1286
rect 11982 1244 12142 1252
rect 13870 1286 14030 1292
rect 13870 1252 13927 1286
rect 13961 1252 14030 1286
rect 13870 1244 14030 1252
rect 15752 1286 15912 1292
rect 15752 1252 15809 1286
rect 15843 1252 15912 1286
rect 15752 1244 15912 1252
rect 17640 1286 17800 1292
rect 17640 1252 17697 1286
rect 17731 1252 17800 1286
rect 17640 1244 17800 1252
rect 19528 1286 19688 1292
rect 19528 1252 19585 1286
rect 19619 1252 19688 1286
rect 19528 1244 19688 1252
rect 21416 1286 21576 1292
rect 21416 1252 21473 1286
rect 21507 1252 21576 1286
rect 21416 1244 21576 1252
rect 23304 1286 23464 1292
rect 23304 1252 23361 1286
rect 23395 1252 23464 1286
rect 23304 1244 23464 1252
rect 25192 1286 25352 1292
rect 25192 1252 25249 1286
rect 25283 1252 25352 1286
rect 25192 1244 25352 1252
rect 27080 1286 27240 1292
rect 27080 1252 27137 1286
rect 27171 1252 27240 1286
rect 27080 1244 27240 1252
rect 28968 1286 29128 1292
rect 28968 1252 29025 1286
rect 29059 1252 29128 1286
rect 28968 1244 29128 1252
rect 30856 1286 31016 1292
rect 30856 1252 30913 1286
rect 30947 1252 31016 1286
rect 30856 1244 31016 1252
rect 32744 1286 32904 1292
rect 32744 1252 32801 1286
rect 32835 1252 32904 1286
rect 32744 1244 32904 1252
rect 34632 1286 34792 1292
rect 34632 1252 34689 1286
rect 34723 1252 34792 1286
rect 34632 1244 34792 1252
rect 36520 1286 36680 1292
rect 36520 1252 36577 1286
rect 36611 1252 36680 1286
rect 36520 1244 36680 1252
rect 38408 1286 38568 1292
rect 38408 1252 38465 1286
rect 38499 1252 38568 1286
rect 38408 1244 38568 1252
rect 40296 1286 40456 1292
rect 40296 1252 40353 1286
rect 40387 1252 40456 1286
rect 40296 1244 40456 1252
rect 42184 1286 42344 1292
rect 42184 1252 42241 1286
rect 42275 1252 42344 1286
rect 42184 1244 42344 1252
rect 44072 1286 44232 1292
rect 44072 1252 44129 1286
rect 44163 1252 44232 1286
rect 44072 1244 44232 1252
rect 45954 1286 46114 1292
rect 45954 1252 46011 1286
rect 46045 1252 46114 1286
rect 45954 1244 46114 1252
rect 47842 1286 48002 1292
rect 47842 1252 47899 1286
rect 47933 1252 48002 1286
rect 47842 1244 48002 1252
rect 49730 1286 49890 1292
rect 49730 1252 49787 1286
rect 49821 1252 49890 1286
rect 49730 1244 49890 1252
rect 51618 1286 51778 1292
rect 51618 1252 51675 1286
rect 51709 1252 51778 1286
rect 51618 1244 51778 1252
rect 53506 1286 53666 1292
rect 53506 1252 53563 1286
rect 53597 1252 53666 1286
rect 53506 1244 53666 1252
rect 55394 1286 55554 1292
rect 55394 1252 55451 1286
rect 55485 1252 55554 1286
rect 55394 1244 55554 1252
rect 57282 1286 57442 1292
rect 57282 1252 57339 1286
rect 57373 1252 57442 1286
rect 57282 1244 57442 1252
rect 59170 1286 59330 1292
rect 59170 1252 59227 1286
rect 59261 1252 59330 1286
rect 59170 1244 59330 1252
rect 652 230 812 236
rect 652 196 709 230
rect 743 196 812 230
rect 652 188 812 196
rect 2540 230 2700 236
rect 2540 196 2597 230
rect 2631 196 2700 230
rect 2540 188 2700 196
rect 4428 230 4588 236
rect 4428 196 4485 230
rect 4519 196 4588 230
rect 4428 188 4588 196
rect 6316 230 6476 236
rect 6316 196 6373 230
rect 6407 196 6476 230
rect 6316 188 6476 196
rect 8204 230 8364 236
rect 8204 196 8261 230
rect 8295 196 8364 230
rect 8204 188 8364 196
rect 10092 230 10252 236
rect 10092 196 10149 230
rect 10183 196 10252 230
rect 10092 188 10252 196
rect 11980 230 12140 236
rect 11980 196 12037 230
rect 12071 196 12140 230
rect 11980 188 12140 196
rect 13868 230 14028 236
rect 13868 196 13925 230
rect 13959 196 14028 230
rect 13868 188 14028 196
rect 15750 230 15910 236
rect 15750 196 15807 230
rect 15841 196 15910 230
rect 15750 188 15910 196
rect 17638 230 17798 236
rect 17638 196 17695 230
rect 17729 196 17798 230
rect 17638 188 17798 196
rect 19526 230 19686 236
rect 19526 196 19583 230
rect 19617 196 19686 230
rect 19526 188 19686 196
rect 21414 230 21574 236
rect 21414 196 21471 230
rect 21505 196 21574 230
rect 21414 188 21574 196
rect 23302 230 23462 236
rect 23302 196 23359 230
rect 23393 196 23462 230
rect 23302 188 23462 196
rect 25190 230 25350 236
rect 25190 196 25247 230
rect 25281 196 25350 230
rect 25190 188 25350 196
rect 27078 230 27238 236
rect 27078 196 27135 230
rect 27169 196 27238 230
rect 27078 188 27238 196
rect 28966 230 29126 236
rect 28966 196 29023 230
rect 29057 196 29126 230
rect 28966 188 29126 196
rect 30854 230 31014 236
rect 30854 196 30911 230
rect 30945 196 31014 230
rect 30854 188 31014 196
rect 32742 230 32902 236
rect 32742 196 32799 230
rect 32833 196 32902 230
rect 32742 188 32902 196
rect 34630 230 34790 236
rect 34630 196 34687 230
rect 34721 196 34790 230
rect 34630 188 34790 196
rect 36518 230 36678 236
rect 36518 196 36575 230
rect 36609 196 36678 230
rect 36518 188 36678 196
rect 38406 230 38566 236
rect 38406 196 38463 230
rect 38497 196 38566 230
rect 38406 188 38566 196
rect 40294 230 40454 236
rect 40294 196 40351 230
rect 40385 196 40454 230
rect 40294 188 40454 196
rect 42182 230 42342 236
rect 42182 196 42239 230
rect 42273 196 42342 230
rect 42182 188 42342 196
rect 44070 230 44230 236
rect 44070 196 44127 230
rect 44161 196 44230 230
rect 44070 188 44230 196
rect 45952 230 46112 236
rect 45952 196 46009 230
rect 46043 196 46112 230
rect 45952 188 46112 196
rect 47840 230 48000 236
rect 47840 196 47897 230
rect 47931 196 48000 230
rect 47840 188 48000 196
rect 49728 230 49888 236
rect 49728 196 49785 230
rect 49819 196 49888 230
rect 49728 188 49888 196
rect 51616 230 51776 236
rect 51616 196 51673 230
rect 51707 196 51776 230
rect 51616 188 51776 196
rect 53504 230 53664 236
rect 53504 196 53561 230
rect 53595 196 53664 230
rect 53504 188 53664 196
rect 55392 230 55552 236
rect 55392 196 55449 230
rect 55483 196 55552 230
rect 55392 188 55552 196
rect 57280 230 57440 236
rect 57280 196 57337 230
rect 57371 196 57440 230
rect 57280 188 57440 196
rect 59168 230 59328 236
rect 59168 196 59225 230
rect 59259 196 59328 230
rect 59168 188 59328 196
<< nsubdiff >>
rect 562 6385 696 6404
rect 562 6351 634 6385
rect 668 6351 696 6385
rect 562 6334 696 6351
rect 2450 6385 2584 6404
rect 2450 6351 2522 6385
rect 2556 6351 2584 6385
rect 2450 6334 2584 6351
rect 4338 6385 4472 6404
rect 4338 6351 4410 6385
rect 4444 6351 4472 6385
rect 4338 6334 4472 6351
rect 6226 6385 6360 6404
rect 6226 6351 6298 6385
rect 6332 6351 6360 6385
rect 6226 6334 6360 6351
rect 8114 6385 8248 6404
rect 8114 6351 8186 6385
rect 8220 6351 8248 6385
rect 8114 6334 8248 6351
rect 10002 6385 10136 6404
rect 10002 6351 10074 6385
rect 10108 6351 10136 6385
rect 10002 6334 10136 6351
rect 11890 6385 12024 6404
rect 11890 6351 11962 6385
rect 11996 6351 12024 6385
rect 11890 6334 12024 6351
rect 13778 6385 13912 6404
rect 13778 6351 13850 6385
rect 13884 6351 13912 6385
rect 13778 6334 13912 6351
rect 15660 6385 15794 6404
rect 15660 6351 15732 6385
rect 15766 6351 15794 6385
rect 15660 6334 15794 6351
rect 17548 6385 17682 6404
rect 17548 6351 17620 6385
rect 17654 6351 17682 6385
rect 17548 6334 17682 6351
rect 19436 6385 19570 6404
rect 19436 6351 19508 6385
rect 19542 6351 19570 6385
rect 19436 6334 19570 6351
rect 21324 6385 21458 6404
rect 21324 6351 21396 6385
rect 21430 6351 21458 6385
rect 21324 6334 21458 6351
rect 23212 6385 23346 6404
rect 23212 6351 23284 6385
rect 23318 6351 23346 6385
rect 23212 6334 23346 6351
rect 25100 6385 25234 6404
rect 25100 6351 25172 6385
rect 25206 6351 25234 6385
rect 25100 6334 25234 6351
rect 26988 6385 27122 6404
rect 26988 6351 27060 6385
rect 27094 6351 27122 6385
rect 26988 6334 27122 6351
rect 28876 6385 29010 6404
rect 28876 6351 28948 6385
rect 28982 6351 29010 6385
rect 28876 6334 29010 6351
rect 30764 6385 30898 6404
rect 30764 6351 30836 6385
rect 30870 6351 30898 6385
rect 30764 6334 30898 6351
rect 32652 6385 32786 6404
rect 32652 6351 32724 6385
rect 32758 6351 32786 6385
rect 32652 6334 32786 6351
rect 34540 6385 34674 6404
rect 34540 6351 34612 6385
rect 34646 6351 34674 6385
rect 34540 6334 34674 6351
rect 36428 6385 36562 6404
rect 36428 6351 36500 6385
rect 36534 6351 36562 6385
rect 36428 6334 36562 6351
rect 38316 6385 38450 6404
rect 38316 6351 38388 6385
rect 38422 6351 38450 6385
rect 38316 6334 38450 6351
rect 40204 6385 40338 6404
rect 40204 6351 40276 6385
rect 40310 6351 40338 6385
rect 40204 6334 40338 6351
rect 42092 6385 42226 6404
rect 42092 6351 42164 6385
rect 42198 6351 42226 6385
rect 42092 6334 42226 6351
rect 43980 6385 44114 6404
rect 43980 6351 44052 6385
rect 44086 6351 44114 6385
rect 43980 6334 44114 6351
rect 45862 6385 45996 6404
rect 45862 6351 45934 6385
rect 45968 6351 45996 6385
rect 45862 6334 45996 6351
rect 47750 6385 47884 6404
rect 47750 6351 47822 6385
rect 47856 6351 47884 6385
rect 47750 6334 47884 6351
rect 49638 6385 49772 6404
rect 49638 6351 49710 6385
rect 49744 6351 49772 6385
rect 49638 6334 49772 6351
rect 51526 6385 51660 6404
rect 51526 6351 51598 6385
rect 51632 6351 51660 6385
rect 51526 6334 51660 6351
rect 53414 6385 53548 6404
rect 53414 6351 53486 6385
rect 53520 6351 53548 6385
rect 53414 6334 53548 6351
rect 55302 6385 55436 6404
rect 55302 6351 55374 6385
rect 55408 6351 55436 6385
rect 55302 6334 55436 6351
rect 57190 6385 57324 6404
rect 57190 6351 57262 6385
rect 57296 6351 57324 6385
rect 57190 6334 57324 6351
rect 59078 6385 59212 6404
rect 59078 6351 59150 6385
rect 59184 6351 59212 6385
rect 59078 6334 59212 6351
rect 560 5329 694 5348
rect 560 5295 632 5329
rect 666 5295 694 5329
rect 2448 5329 2582 5348
rect 560 5278 694 5295
rect 2448 5295 2520 5329
rect 2554 5295 2582 5329
rect 4336 5329 4470 5348
rect 2448 5278 2582 5295
rect 4336 5295 4408 5329
rect 4442 5295 4470 5329
rect 6224 5329 6358 5348
rect 4336 5278 4470 5295
rect 6224 5295 6296 5329
rect 6330 5295 6358 5329
rect 8112 5329 8246 5348
rect 6224 5278 6358 5295
rect 8112 5295 8184 5329
rect 8218 5295 8246 5329
rect 10000 5329 10134 5348
rect 8112 5278 8246 5295
rect 10000 5295 10072 5329
rect 10106 5295 10134 5329
rect 11888 5329 12022 5348
rect 10000 5278 10134 5295
rect 11888 5295 11960 5329
rect 11994 5295 12022 5329
rect 13776 5329 13910 5348
rect 11888 5278 12022 5295
rect 13776 5295 13848 5329
rect 13882 5295 13910 5329
rect 15658 5329 15792 5348
rect 13776 5278 13910 5295
rect 15658 5295 15730 5329
rect 15764 5295 15792 5329
rect 17546 5329 17680 5348
rect 15658 5278 15792 5295
rect 17546 5295 17618 5329
rect 17652 5295 17680 5329
rect 19434 5329 19568 5348
rect 17546 5278 17680 5295
rect 19434 5295 19506 5329
rect 19540 5295 19568 5329
rect 21322 5329 21456 5348
rect 19434 5278 19568 5295
rect 21322 5295 21394 5329
rect 21428 5295 21456 5329
rect 23210 5329 23344 5348
rect 21322 5278 21456 5295
rect 23210 5295 23282 5329
rect 23316 5295 23344 5329
rect 25098 5329 25232 5348
rect 23210 5278 23344 5295
rect 25098 5295 25170 5329
rect 25204 5295 25232 5329
rect 26986 5329 27120 5348
rect 25098 5278 25232 5295
rect 26986 5295 27058 5329
rect 27092 5295 27120 5329
rect 28874 5329 29008 5348
rect 26986 5278 27120 5295
rect 28874 5295 28946 5329
rect 28980 5295 29008 5329
rect 30762 5329 30896 5348
rect 28874 5278 29008 5295
rect 30762 5295 30834 5329
rect 30868 5295 30896 5329
rect 32650 5329 32784 5348
rect 30762 5278 30896 5295
rect 32650 5295 32722 5329
rect 32756 5295 32784 5329
rect 34538 5329 34672 5348
rect 32650 5278 32784 5295
rect 34538 5295 34610 5329
rect 34644 5295 34672 5329
rect 36426 5329 36560 5348
rect 34538 5278 34672 5295
rect 36426 5295 36498 5329
rect 36532 5295 36560 5329
rect 38314 5329 38448 5348
rect 36426 5278 36560 5295
rect 38314 5295 38386 5329
rect 38420 5295 38448 5329
rect 40202 5329 40336 5348
rect 38314 5278 38448 5295
rect 40202 5295 40274 5329
rect 40308 5295 40336 5329
rect 42090 5329 42224 5348
rect 40202 5278 40336 5295
rect 42090 5295 42162 5329
rect 42196 5295 42224 5329
rect 43978 5329 44112 5348
rect 42090 5278 42224 5295
rect 43978 5295 44050 5329
rect 44084 5295 44112 5329
rect 45860 5329 45994 5348
rect 43978 5278 44112 5295
rect 45860 5295 45932 5329
rect 45966 5295 45994 5329
rect 47748 5329 47882 5348
rect 45860 5278 45994 5295
rect 47748 5295 47820 5329
rect 47854 5295 47882 5329
rect 49636 5329 49770 5348
rect 47748 5278 47882 5295
rect 49636 5295 49708 5329
rect 49742 5295 49770 5329
rect 51524 5329 51658 5348
rect 49636 5278 49770 5295
rect 51524 5295 51596 5329
rect 51630 5295 51658 5329
rect 53412 5329 53546 5348
rect 51524 5278 51658 5295
rect 53412 5295 53484 5329
rect 53518 5295 53546 5329
rect 55300 5329 55434 5348
rect 53412 5278 53546 5295
rect 55300 5295 55372 5329
rect 55406 5295 55434 5329
rect 57188 5329 57322 5348
rect 55300 5278 55434 5295
rect 57188 5295 57260 5329
rect 57294 5295 57322 5329
rect 59076 5329 59210 5348
rect 57188 5278 57322 5295
rect 59076 5295 59148 5329
rect 59182 5295 59210 5329
rect 59076 5278 59210 5295
rect 14874 3629 15008 3648
rect 14874 3595 14946 3629
rect 14980 3595 15008 3629
rect 14874 3578 15008 3595
rect 45016 3789 45150 3808
rect 45016 3755 45088 3789
rect 45122 3755 45150 3789
rect 45016 3738 45150 3755
rect 772 2145 906 2162
rect 772 2111 800 2145
rect 834 2111 906 2145
rect 2660 2145 2794 2162
rect 772 2092 906 2111
rect 2660 2111 2688 2145
rect 2722 2111 2794 2145
rect 4548 2145 4682 2162
rect 2660 2092 2794 2111
rect 4548 2111 4576 2145
rect 4610 2111 4682 2145
rect 6436 2145 6570 2162
rect 4548 2092 4682 2111
rect 6436 2111 6464 2145
rect 6498 2111 6570 2145
rect 8324 2145 8458 2162
rect 6436 2092 6570 2111
rect 8324 2111 8352 2145
rect 8386 2111 8458 2145
rect 10212 2145 10346 2162
rect 8324 2092 8458 2111
rect 10212 2111 10240 2145
rect 10274 2111 10346 2145
rect 12100 2145 12234 2162
rect 10212 2092 10346 2111
rect 12100 2111 12128 2145
rect 12162 2111 12234 2145
rect 13988 2145 14122 2162
rect 12100 2092 12234 2111
rect 13988 2111 14016 2145
rect 14050 2111 14122 2145
rect 15870 2145 16004 2162
rect 13988 2092 14122 2111
rect 15870 2111 15898 2145
rect 15932 2111 16004 2145
rect 17758 2145 17892 2162
rect 15870 2092 16004 2111
rect 17758 2111 17786 2145
rect 17820 2111 17892 2145
rect 19646 2145 19780 2162
rect 17758 2092 17892 2111
rect 19646 2111 19674 2145
rect 19708 2111 19780 2145
rect 21534 2145 21668 2162
rect 19646 2092 19780 2111
rect 21534 2111 21562 2145
rect 21596 2111 21668 2145
rect 23422 2145 23556 2162
rect 21534 2092 21668 2111
rect 23422 2111 23450 2145
rect 23484 2111 23556 2145
rect 25310 2145 25444 2162
rect 23422 2092 23556 2111
rect 25310 2111 25338 2145
rect 25372 2111 25444 2145
rect 27198 2145 27332 2162
rect 25310 2092 25444 2111
rect 27198 2111 27226 2145
rect 27260 2111 27332 2145
rect 29086 2145 29220 2162
rect 27198 2092 27332 2111
rect 29086 2111 29114 2145
rect 29148 2111 29220 2145
rect 30974 2145 31108 2162
rect 29086 2092 29220 2111
rect 30974 2111 31002 2145
rect 31036 2111 31108 2145
rect 32862 2145 32996 2162
rect 30974 2092 31108 2111
rect 32862 2111 32890 2145
rect 32924 2111 32996 2145
rect 34750 2145 34884 2162
rect 32862 2092 32996 2111
rect 34750 2111 34778 2145
rect 34812 2111 34884 2145
rect 36638 2145 36772 2162
rect 34750 2092 34884 2111
rect 36638 2111 36666 2145
rect 36700 2111 36772 2145
rect 38526 2145 38660 2162
rect 36638 2092 36772 2111
rect 38526 2111 38554 2145
rect 38588 2111 38660 2145
rect 40414 2145 40548 2162
rect 38526 2092 38660 2111
rect 40414 2111 40442 2145
rect 40476 2111 40548 2145
rect 42302 2145 42436 2162
rect 40414 2092 40548 2111
rect 42302 2111 42330 2145
rect 42364 2111 42436 2145
rect 44190 2145 44324 2162
rect 42302 2092 42436 2111
rect 44190 2111 44218 2145
rect 44252 2111 44324 2145
rect 46072 2145 46206 2162
rect 44190 2092 44324 2111
rect 46072 2111 46100 2145
rect 46134 2111 46206 2145
rect 47960 2145 48094 2162
rect 46072 2092 46206 2111
rect 47960 2111 47988 2145
rect 48022 2111 48094 2145
rect 49848 2145 49982 2162
rect 47960 2092 48094 2111
rect 49848 2111 49876 2145
rect 49910 2111 49982 2145
rect 51736 2145 51870 2162
rect 49848 2092 49982 2111
rect 51736 2111 51764 2145
rect 51798 2111 51870 2145
rect 53624 2145 53758 2162
rect 51736 2092 51870 2111
rect 53624 2111 53652 2145
rect 53686 2111 53758 2145
rect 55512 2145 55646 2162
rect 53624 2092 53758 2111
rect 55512 2111 55540 2145
rect 55574 2111 55646 2145
rect 57400 2145 57534 2162
rect 55512 2092 55646 2111
rect 57400 2111 57428 2145
rect 57462 2111 57534 2145
rect 59288 2145 59422 2162
rect 57400 2092 57534 2111
rect 59288 2111 59316 2145
rect 59350 2111 59422 2145
rect 59288 2092 59422 2111
rect 770 1089 904 1106
rect 770 1055 798 1089
rect 832 1055 904 1089
rect 770 1036 904 1055
rect 2658 1089 2792 1106
rect 2658 1055 2686 1089
rect 2720 1055 2792 1089
rect 2658 1036 2792 1055
rect 4546 1089 4680 1106
rect 4546 1055 4574 1089
rect 4608 1055 4680 1089
rect 4546 1036 4680 1055
rect 6434 1089 6568 1106
rect 6434 1055 6462 1089
rect 6496 1055 6568 1089
rect 6434 1036 6568 1055
rect 8322 1089 8456 1106
rect 8322 1055 8350 1089
rect 8384 1055 8456 1089
rect 8322 1036 8456 1055
rect 10210 1089 10344 1106
rect 10210 1055 10238 1089
rect 10272 1055 10344 1089
rect 10210 1036 10344 1055
rect 12098 1089 12232 1106
rect 12098 1055 12126 1089
rect 12160 1055 12232 1089
rect 12098 1036 12232 1055
rect 13986 1089 14120 1106
rect 13986 1055 14014 1089
rect 14048 1055 14120 1089
rect 13986 1036 14120 1055
rect 15868 1089 16002 1106
rect 15868 1055 15896 1089
rect 15930 1055 16002 1089
rect 15868 1036 16002 1055
rect 17756 1089 17890 1106
rect 17756 1055 17784 1089
rect 17818 1055 17890 1089
rect 17756 1036 17890 1055
rect 19644 1089 19778 1106
rect 19644 1055 19672 1089
rect 19706 1055 19778 1089
rect 19644 1036 19778 1055
rect 21532 1089 21666 1106
rect 21532 1055 21560 1089
rect 21594 1055 21666 1089
rect 21532 1036 21666 1055
rect 23420 1089 23554 1106
rect 23420 1055 23448 1089
rect 23482 1055 23554 1089
rect 23420 1036 23554 1055
rect 25308 1089 25442 1106
rect 25308 1055 25336 1089
rect 25370 1055 25442 1089
rect 25308 1036 25442 1055
rect 27196 1089 27330 1106
rect 27196 1055 27224 1089
rect 27258 1055 27330 1089
rect 27196 1036 27330 1055
rect 29084 1089 29218 1106
rect 29084 1055 29112 1089
rect 29146 1055 29218 1089
rect 29084 1036 29218 1055
rect 30972 1089 31106 1106
rect 30972 1055 31000 1089
rect 31034 1055 31106 1089
rect 30972 1036 31106 1055
rect 32860 1089 32994 1106
rect 32860 1055 32888 1089
rect 32922 1055 32994 1089
rect 32860 1036 32994 1055
rect 34748 1089 34882 1106
rect 34748 1055 34776 1089
rect 34810 1055 34882 1089
rect 34748 1036 34882 1055
rect 36636 1089 36770 1106
rect 36636 1055 36664 1089
rect 36698 1055 36770 1089
rect 36636 1036 36770 1055
rect 38524 1089 38658 1106
rect 38524 1055 38552 1089
rect 38586 1055 38658 1089
rect 38524 1036 38658 1055
rect 40412 1089 40546 1106
rect 40412 1055 40440 1089
rect 40474 1055 40546 1089
rect 40412 1036 40546 1055
rect 42300 1089 42434 1106
rect 42300 1055 42328 1089
rect 42362 1055 42434 1089
rect 42300 1036 42434 1055
rect 44188 1089 44322 1106
rect 44188 1055 44216 1089
rect 44250 1055 44322 1089
rect 44188 1036 44322 1055
rect 46070 1089 46204 1106
rect 46070 1055 46098 1089
rect 46132 1055 46204 1089
rect 46070 1036 46204 1055
rect 47958 1089 48092 1106
rect 47958 1055 47986 1089
rect 48020 1055 48092 1089
rect 47958 1036 48092 1055
rect 49846 1089 49980 1106
rect 49846 1055 49874 1089
rect 49908 1055 49980 1089
rect 49846 1036 49980 1055
rect 51734 1089 51868 1106
rect 51734 1055 51762 1089
rect 51796 1055 51868 1089
rect 51734 1036 51868 1055
rect 53622 1089 53756 1106
rect 53622 1055 53650 1089
rect 53684 1055 53756 1089
rect 53622 1036 53756 1055
rect 55510 1089 55644 1106
rect 55510 1055 55538 1089
rect 55572 1055 55644 1089
rect 55510 1036 55644 1055
rect 57398 1089 57532 1106
rect 57398 1055 57426 1089
rect 57460 1055 57532 1089
rect 57398 1036 57532 1055
rect 59286 1089 59420 1106
rect 59286 1055 59314 1089
rect 59348 1055 59420 1089
rect 59286 1036 59420 1055
<< psubdiffcont >>
rect 723 7210 757 7244
rect 2611 7210 2645 7244
rect 4499 7210 4533 7244
rect 6387 7210 6421 7244
rect 8275 7210 8309 7244
rect 10163 7210 10197 7244
rect 12051 7210 12085 7244
rect 13939 7210 13973 7244
rect 15821 7210 15855 7244
rect 17709 7210 17743 7244
rect 19597 7210 19631 7244
rect 21485 7210 21519 7244
rect 23373 7210 23407 7244
rect 25261 7210 25295 7244
rect 27149 7210 27183 7244
rect 29037 7210 29071 7244
rect 30925 7210 30959 7244
rect 32813 7210 32847 7244
rect 34701 7210 34735 7244
rect 36589 7210 36623 7244
rect 38477 7210 38511 7244
rect 40365 7210 40399 7244
rect 42253 7210 42287 7244
rect 44141 7210 44175 7244
rect 46023 7210 46057 7244
rect 47911 7210 47945 7244
rect 49799 7210 49833 7244
rect 51687 7210 51721 7244
rect 53575 7210 53609 7244
rect 55463 7210 55497 7244
rect 57351 7210 57385 7244
rect 59239 7210 59273 7244
rect 721 6154 755 6188
rect 2609 6154 2643 6188
rect 4497 6154 4531 6188
rect 6385 6154 6419 6188
rect 8273 6154 8307 6188
rect 10161 6154 10195 6188
rect 12049 6154 12083 6188
rect 13937 6154 13971 6188
rect 15819 6154 15853 6188
rect 17707 6154 17741 6188
rect 19595 6154 19629 6188
rect 21483 6154 21517 6188
rect 23371 6154 23405 6188
rect 25259 6154 25293 6188
rect 27147 6154 27181 6188
rect 29035 6154 29069 6188
rect 30923 6154 30957 6188
rect 32811 6154 32845 6188
rect 34699 6154 34733 6188
rect 36587 6154 36621 6188
rect 38475 6154 38509 6188
rect 40363 6154 40397 6188
rect 42251 6154 42285 6188
rect 44139 6154 44173 6188
rect 46021 6154 46055 6188
rect 47909 6154 47943 6188
rect 49797 6154 49831 6188
rect 51685 6154 51719 6188
rect 53573 6154 53607 6188
rect 55461 6154 55495 6188
rect 57349 6154 57383 6188
rect 59237 6154 59271 6188
rect 711 1252 745 1286
rect 2599 1252 2633 1286
rect 4487 1252 4521 1286
rect 6375 1252 6409 1286
rect 8263 1252 8297 1286
rect 10151 1252 10185 1286
rect 12039 1252 12073 1286
rect 13927 1252 13961 1286
rect 15809 1252 15843 1286
rect 17697 1252 17731 1286
rect 19585 1252 19619 1286
rect 21473 1252 21507 1286
rect 23361 1252 23395 1286
rect 25249 1252 25283 1286
rect 27137 1252 27171 1286
rect 29025 1252 29059 1286
rect 30913 1252 30947 1286
rect 32801 1252 32835 1286
rect 34689 1252 34723 1286
rect 36577 1252 36611 1286
rect 38465 1252 38499 1286
rect 40353 1252 40387 1286
rect 42241 1252 42275 1286
rect 44129 1252 44163 1286
rect 46011 1252 46045 1286
rect 47899 1252 47933 1286
rect 49787 1252 49821 1286
rect 51675 1252 51709 1286
rect 53563 1252 53597 1286
rect 55451 1252 55485 1286
rect 57339 1252 57373 1286
rect 59227 1252 59261 1286
rect 709 196 743 230
rect 2597 196 2631 230
rect 4485 196 4519 230
rect 6373 196 6407 230
rect 8261 196 8295 230
rect 10149 196 10183 230
rect 12037 196 12071 230
rect 13925 196 13959 230
rect 15807 196 15841 230
rect 17695 196 17729 230
rect 19583 196 19617 230
rect 21471 196 21505 230
rect 23359 196 23393 230
rect 25247 196 25281 230
rect 27135 196 27169 230
rect 29023 196 29057 230
rect 30911 196 30945 230
rect 32799 196 32833 230
rect 34687 196 34721 230
rect 36575 196 36609 230
rect 38463 196 38497 230
rect 40351 196 40385 230
rect 42239 196 42273 230
rect 44127 196 44161 230
rect 46009 196 46043 230
rect 47897 196 47931 230
rect 49785 196 49819 230
rect 51673 196 51707 230
rect 53561 196 53595 230
rect 55449 196 55483 230
rect 57337 196 57371 230
rect 59225 196 59259 230
<< nsubdiffcont >>
rect 634 6351 668 6385
rect 2522 6351 2556 6385
rect 4410 6351 4444 6385
rect 6298 6351 6332 6385
rect 8186 6351 8220 6385
rect 10074 6351 10108 6385
rect 11962 6351 11996 6385
rect 13850 6351 13884 6385
rect 15732 6351 15766 6385
rect 17620 6351 17654 6385
rect 19508 6351 19542 6385
rect 21396 6351 21430 6385
rect 23284 6351 23318 6385
rect 25172 6351 25206 6385
rect 27060 6351 27094 6385
rect 28948 6351 28982 6385
rect 30836 6351 30870 6385
rect 32724 6351 32758 6385
rect 34612 6351 34646 6385
rect 36500 6351 36534 6385
rect 38388 6351 38422 6385
rect 40276 6351 40310 6385
rect 42164 6351 42198 6385
rect 44052 6351 44086 6385
rect 45934 6351 45968 6385
rect 47822 6351 47856 6385
rect 49710 6351 49744 6385
rect 51598 6351 51632 6385
rect 53486 6351 53520 6385
rect 55374 6351 55408 6385
rect 57262 6351 57296 6385
rect 59150 6351 59184 6385
rect 632 5295 666 5329
rect 2520 5295 2554 5329
rect 4408 5295 4442 5329
rect 6296 5295 6330 5329
rect 8184 5295 8218 5329
rect 10072 5295 10106 5329
rect 11960 5295 11994 5329
rect 13848 5295 13882 5329
rect 15730 5295 15764 5329
rect 17618 5295 17652 5329
rect 19506 5295 19540 5329
rect 21394 5295 21428 5329
rect 23282 5295 23316 5329
rect 25170 5295 25204 5329
rect 27058 5295 27092 5329
rect 28946 5295 28980 5329
rect 30834 5295 30868 5329
rect 32722 5295 32756 5329
rect 34610 5295 34644 5329
rect 36498 5295 36532 5329
rect 38386 5295 38420 5329
rect 40274 5295 40308 5329
rect 42162 5295 42196 5329
rect 44050 5295 44084 5329
rect 45932 5295 45966 5329
rect 47820 5295 47854 5329
rect 49708 5295 49742 5329
rect 51596 5295 51630 5329
rect 53484 5295 53518 5329
rect 55372 5295 55406 5329
rect 57260 5295 57294 5329
rect 59148 5295 59182 5329
rect 14946 3595 14980 3629
rect 45088 3755 45122 3789
rect 800 2111 834 2145
rect 2688 2111 2722 2145
rect 4576 2111 4610 2145
rect 6464 2111 6498 2145
rect 8352 2111 8386 2145
rect 10240 2111 10274 2145
rect 12128 2111 12162 2145
rect 14016 2111 14050 2145
rect 15898 2111 15932 2145
rect 17786 2111 17820 2145
rect 19674 2111 19708 2145
rect 21562 2111 21596 2145
rect 23450 2111 23484 2145
rect 25338 2111 25372 2145
rect 27226 2111 27260 2145
rect 29114 2111 29148 2145
rect 31002 2111 31036 2145
rect 32890 2111 32924 2145
rect 34778 2111 34812 2145
rect 36666 2111 36700 2145
rect 38554 2111 38588 2145
rect 40442 2111 40476 2145
rect 42330 2111 42364 2145
rect 44218 2111 44252 2145
rect 46100 2111 46134 2145
rect 47988 2111 48022 2145
rect 49876 2111 49910 2145
rect 51764 2111 51798 2145
rect 53652 2111 53686 2145
rect 55540 2111 55574 2145
rect 57428 2111 57462 2145
rect 59316 2111 59350 2145
rect 798 1055 832 1089
rect 2686 1055 2720 1089
rect 4574 1055 4608 1089
rect 6462 1055 6496 1089
rect 8350 1055 8384 1089
rect 10238 1055 10272 1089
rect 12126 1055 12160 1089
rect 14014 1055 14048 1089
rect 15896 1055 15930 1089
rect 17784 1055 17818 1089
rect 19672 1055 19706 1089
rect 21560 1055 21594 1089
rect 23448 1055 23482 1089
rect 25336 1055 25370 1089
rect 27224 1055 27258 1089
rect 29112 1055 29146 1089
rect 31000 1055 31034 1089
rect 32888 1055 32922 1089
rect 34776 1055 34810 1089
rect 36664 1055 36698 1089
rect 38552 1055 38586 1089
rect 40440 1055 40474 1089
rect 42328 1055 42362 1089
rect 44216 1055 44250 1089
rect 46098 1055 46132 1089
rect 47986 1055 48020 1089
rect 49874 1055 49908 1089
rect 51762 1055 51796 1089
rect 53650 1055 53684 1089
rect 55538 1055 55572 1089
rect 57426 1055 57460 1089
rect 59314 1055 59348 1089
<< poly >>
rect 748 7140 814 7156
rect 748 7106 764 7140
rect 798 7106 814 7140
rect 670 7068 700 7094
rect 748 7090 814 7106
rect 2636 7140 2702 7156
rect 2636 7106 2652 7140
rect 2686 7106 2702 7140
rect 766 7068 796 7090
rect 2558 7068 2588 7094
rect 2636 7090 2702 7106
rect 4524 7140 4590 7156
rect 4524 7106 4540 7140
rect 4574 7106 4590 7140
rect 2654 7068 2684 7090
rect 4446 7068 4476 7094
rect 4524 7090 4590 7106
rect 6412 7140 6478 7156
rect 6412 7106 6428 7140
rect 6462 7106 6478 7140
rect 4542 7068 4572 7090
rect 6334 7068 6364 7094
rect 6412 7090 6478 7106
rect 8300 7140 8366 7156
rect 8300 7106 8316 7140
rect 8350 7106 8366 7140
rect 6430 7068 6460 7090
rect 8222 7068 8252 7094
rect 8300 7090 8366 7106
rect 10188 7140 10254 7156
rect 10188 7106 10204 7140
rect 10238 7106 10254 7140
rect 8318 7068 8348 7090
rect 10110 7068 10140 7094
rect 10188 7090 10254 7106
rect 12076 7140 12142 7156
rect 12076 7106 12092 7140
rect 12126 7106 12142 7140
rect 10206 7068 10236 7090
rect 11998 7068 12028 7094
rect 12076 7090 12142 7106
rect 13964 7140 14030 7156
rect 13964 7106 13980 7140
rect 14014 7106 14030 7140
rect 12094 7068 12124 7090
rect 13886 7068 13916 7094
rect 13964 7090 14030 7106
rect 15846 7140 15912 7156
rect 15846 7106 15862 7140
rect 15896 7106 15912 7140
rect 13982 7068 14012 7090
rect 15768 7068 15798 7094
rect 15846 7090 15912 7106
rect 17734 7140 17800 7156
rect 17734 7106 17750 7140
rect 17784 7106 17800 7140
rect 15864 7068 15894 7090
rect 17656 7068 17686 7094
rect 17734 7090 17800 7106
rect 19622 7140 19688 7156
rect 19622 7106 19638 7140
rect 19672 7106 19688 7140
rect 17752 7068 17782 7090
rect 19544 7068 19574 7094
rect 19622 7090 19688 7106
rect 21510 7140 21576 7156
rect 21510 7106 21526 7140
rect 21560 7106 21576 7140
rect 19640 7068 19670 7090
rect 21432 7068 21462 7094
rect 21510 7090 21576 7106
rect 23398 7140 23464 7156
rect 23398 7106 23414 7140
rect 23448 7106 23464 7140
rect 21528 7068 21558 7090
rect 23320 7068 23350 7094
rect 23398 7090 23464 7106
rect 25286 7140 25352 7156
rect 25286 7106 25302 7140
rect 25336 7106 25352 7140
rect 23416 7068 23446 7090
rect 25208 7068 25238 7094
rect 25286 7090 25352 7106
rect 27174 7140 27240 7156
rect 27174 7106 27190 7140
rect 27224 7106 27240 7140
rect 25304 7068 25334 7090
rect 27096 7068 27126 7094
rect 27174 7090 27240 7106
rect 29062 7140 29128 7156
rect 29062 7106 29078 7140
rect 29112 7106 29128 7140
rect 27192 7068 27222 7090
rect 28984 7068 29014 7094
rect 29062 7090 29128 7106
rect 30950 7140 31016 7156
rect 30950 7106 30966 7140
rect 31000 7106 31016 7140
rect 29080 7068 29110 7090
rect 30872 7068 30902 7094
rect 30950 7090 31016 7106
rect 32838 7140 32904 7156
rect 32838 7106 32854 7140
rect 32888 7106 32904 7140
rect 30968 7068 30998 7090
rect 32760 7068 32790 7094
rect 32838 7090 32904 7106
rect 34726 7140 34792 7156
rect 34726 7106 34742 7140
rect 34776 7106 34792 7140
rect 32856 7068 32886 7090
rect 34648 7068 34678 7094
rect 34726 7090 34792 7106
rect 36614 7140 36680 7156
rect 36614 7106 36630 7140
rect 36664 7106 36680 7140
rect 34744 7068 34774 7090
rect 36536 7068 36566 7094
rect 36614 7090 36680 7106
rect 38502 7140 38568 7156
rect 38502 7106 38518 7140
rect 38552 7106 38568 7140
rect 36632 7068 36662 7090
rect 38424 7068 38454 7094
rect 38502 7090 38568 7106
rect 40390 7140 40456 7156
rect 40390 7106 40406 7140
rect 40440 7106 40456 7140
rect 38520 7068 38550 7090
rect 40312 7068 40342 7094
rect 40390 7090 40456 7106
rect 42278 7140 42344 7156
rect 42278 7106 42294 7140
rect 42328 7106 42344 7140
rect 40408 7068 40438 7090
rect 42200 7068 42230 7094
rect 42278 7090 42344 7106
rect 44166 7140 44232 7156
rect 44166 7106 44182 7140
rect 44216 7106 44232 7140
rect 42296 7068 42326 7090
rect 44088 7068 44118 7094
rect 44166 7090 44232 7106
rect 46048 7140 46114 7156
rect 46048 7106 46064 7140
rect 46098 7106 46114 7140
rect 44184 7068 44214 7090
rect 45970 7068 46000 7094
rect 46048 7090 46114 7106
rect 47936 7140 48002 7156
rect 47936 7106 47952 7140
rect 47986 7106 48002 7140
rect 46066 7068 46096 7090
rect 47858 7068 47888 7094
rect 47936 7090 48002 7106
rect 49824 7140 49890 7156
rect 49824 7106 49840 7140
rect 49874 7106 49890 7140
rect 47954 7068 47984 7090
rect 49746 7068 49776 7094
rect 49824 7090 49890 7106
rect 51712 7140 51778 7156
rect 51712 7106 51728 7140
rect 51762 7106 51778 7140
rect 49842 7068 49872 7090
rect 51634 7068 51664 7094
rect 51712 7090 51778 7106
rect 53600 7140 53666 7156
rect 53600 7106 53616 7140
rect 53650 7106 53666 7140
rect 51730 7068 51760 7090
rect 53522 7068 53552 7094
rect 53600 7090 53666 7106
rect 55488 7140 55554 7156
rect 55488 7106 55504 7140
rect 55538 7106 55554 7140
rect 53618 7068 53648 7090
rect 55410 7068 55440 7094
rect 55488 7090 55554 7106
rect 57376 7140 57442 7156
rect 57376 7106 57392 7140
rect 57426 7106 57442 7140
rect 55506 7068 55536 7090
rect 57298 7068 57328 7094
rect 57376 7090 57442 7106
rect 59264 7140 59330 7156
rect 59264 7106 59280 7140
rect 59314 7106 59330 7140
rect 57394 7068 57424 7090
rect 59186 7068 59216 7094
rect 59264 7090 59330 7106
rect 59282 7068 59312 7090
rect 670 6916 700 6938
rect 652 6900 718 6916
rect 766 6912 796 6938
rect 2558 6916 2588 6938
rect 652 6866 668 6900
rect 702 6866 718 6900
rect -313 6815 -283 6841
rect -225 6815 -195 6841
rect 80 6813 110 6839
rect 652 6838 718 6866
rect 2540 6900 2606 6916
rect 2654 6912 2684 6938
rect 4446 6916 4476 6938
rect 2540 6866 2556 6900
rect 2590 6866 2606 6900
rect 652 6819 830 6838
rect 1276 6821 1306 6847
rect -313 6650 -283 6711
rect -225 6696 -195 6711
rect -225 6672 -189 6696
rect 652 6806 780 6819
rect 764 6785 780 6806
rect 814 6785 830 6819
rect 764 6769 830 6785
rect 686 6738 716 6764
rect 782 6738 812 6769
rect -219 6663 -189 6672
rect -315 6634 -261 6650
rect -315 6600 -305 6634
rect -271 6600 -261 6634
rect -315 6584 -261 6600
rect -219 6647 -143 6663
rect -219 6613 -187 6647
rect -153 6613 -143 6647
rect -219 6597 -143 6613
rect 80 6661 110 6683
rect 80 6645 166 6661
rect 80 6611 116 6645
rect 150 6611 166 6645
rect -313 6523 -283 6584
rect -219 6562 -189 6597
rect 80 6595 166 6611
rect 338 6659 404 6675
rect 338 6625 354 6659
rect 388 6625 404 6659
rect 338 6609 404 6625
rect 80 6563 110 6595
rect 356 6578 386 6609
rect -225 6538 -189 6562
rect -225 6523 -195 6538
rect -313 6339 -283 6365
rect -225 6339 -195 6365
rect 1575 6815 1605 6841
rect 1663 6815 1693 6841
rect 1968 6813 1998 6839
rect 2540 6838 2606 6866
rect 4428 6900 4494 6916
rect 4542 6912 4572 6938
rect 6334 6916 6364 6938
rect 4428 6866 4444 6900
rect 4478 6866 4494 6900
rect 2540 6819 2718 6838
rect 3164 6821 3194 6847
rect 984 6659 1050 6675
rect 984 6625 1000 6659
rect 1034 6625 1050 6659
rect 984 6609 1050 6625
rect 1276 6669 1306 6691
rect 1276 6653 1362 6669
rect 1276 6619 1312 6653
rect 1346 6619 1362 6653
rect 1575 6650 1605 6711
rect 1663 6696 1693 6711
rect 1663 6672 1699 6696
rect 2540 6806 2668 6819
rect 2652 6785 2668 6806
rect 2702 6785 2718 6819
rect 2652 6769 2718 6785
rect 2574 6738 2604 6764
rect 2670 6738 2700 6769
rect 1669 6663 1699 6672
rect 1002 6578 1032 6609
rect 1276 6603 1362 6619
rect 1573 6634 1627 6650
rect 686 6507 716 6538
rect 668 6491 734 6507
rect 668 6457 684 6491
rect 718 6457 734 6491
rect 668 6441 734 6457
rect 782 6454 812 6538
rect 782 6424 868 6454
rect 80 6337 110 6363
rect 356 6348 386 6378
rect 356 6347 418 6348
rect 338 6331 418 6347
rect 338 6297 354 6331
rect 388 6297 418 6331
rect 338 6281 418 6297
rect 386 6266 418 6281
rect 838 6266 868 6424
rect 1276 6571 1306 6603
rect 1573 6600 1583 6634
rect 1617 6600 1627 6634
rect 1573 6584 1627 6600
rect 1669 6647 1745 6663
rect 1669 6613 1701 6647
rect 1735 6613 1745 6647
rect 1669 6597 1745 6613
rect 1968 6661 1998 6683
rect 1968 6645 2054 6661
rect 1968 6611 2004 6645
rect 2038 6611 2054 6645
rect 1002 6347 1032 6378
rect 1575 6523 1605 6584
rect 1669 6562 1699 6597
rect 1968 6595 2054 6611
rect 2226 6659 2292 6675
rect 2226 6625 2242 6659
rect 2276 6625 2292 6659
rect 2226 6609 2292 6625
rect 1968 6563 1998 6595
rect 2244 6578 2274 6609
rect 1663 6538 1699 6562
rect 1663 6523 1693 6538
rect 984 6331 1050 6347
rect 1276 6345 1306 6371
rect 1575 6339 1605 6365
rect 1663 6339 1693 6365
rect 3463 6815 3493 6841
rect 3551 6815 3581 6841
rect 3856 6813 3886 6839
rect 4428 6838 4494 6866
rect 6316 6900 6382 6916
rect 6430 6912 6460 6938
rect 8222 6916 8252 6938
rect 6316 6866 6332 6900
rect 6366 6866 6382 6900
rect 4428 6819 4606 6838
rect 5052 6821 5082 6847
rect 2872 6659 2938 6675
rect 2872 6625 2888 6659
rect 2922 6625 2938 6659
rect 2872 6609 2938 6625
rect 3164 6669 3194 6691
rect 3164 6653 3250 6669
rect 3164 6619 3200 6653
rect 3234 6619 3250 6653
rect 3463 6650 3493 6711
rect 3551 6696 3581 6711
rect 3551 6672 3587 6696
rect 4428 6806 4556 6819
rect 4540 6785 4556 6806
rect 4590 6785 4606 6819
rect 4540 6769 4606 6785
rect 4462 6738 4492 6764
rect 4558 6738 4588 6769
rect 3557 6663 3587 6672
rect 2890 6578 2920 6609
rect 3164 6603 3250 6619
rect 3461 6634 3515 6650
rect 2574 6507 2604 6538
rect 2556 6491 2622 6507
rect 2556 6457 2572 6491
rect 2606 6457 2622 6491
rect 2556 6441 2622 6457
rect 2670 6454 2700 6538
rect 2670 6424 2756 6454
rect 1968 6337 1998 6363
rect 2244 6348 2274 6378
rect 2244 6347 2306 6348
rect 984 6297 1000 6331
rect 1034 6297 1050 6331
rect 984 6281 1050 6297
rect 2226 6331 2306 6347
rect 2226 6297 2242 6331
rect 2276 6297 2306 6331
rect 2226 6281 2306 6297
rect 386 6236 868 6266
rect 2274 6266 2306 6281
rect 2726 6266 2756 6424
rect 3164 6571 3194 6603
rect 3461 6600 3471 6634
rect 3505 6600 3515 6634
rect 3461 6584 3515 6600
rect 3557 6647 3633 6663
rect 3557 6613 3589 6647
rect 3623 6613 3633 6647
rect 3557 6597 3633 6613
rect 3856 6661 3886 6683
rect 3856 6645 3942 6661
rect 3856 6611 3892 6645
rect 3926 6611 3942 6645
rect 2890 6347 2920 6378
rect 3463 6523 3493 6584
rect 3557 6562 3587 6597
rect 3856 6595 3942 6611
rect 4114 6659 4180 6675
rect 4114 6625 4130 6659
rect 4164 6625 4180 6659
rect 4114 6609 4180 6625
rect 3856 6563 3886 6595
rect 4132 6578 4162 6609
rect 3551 6538 3587 6562
rect 3551 6523 3581 6538
rect 2872 6331 2938 6347
rect 3164 6345 3194 6371
rect 3463 6339 3493 6365
rect 3551 6339 3581 6365
rect 5351 6815 5381 6841
rect 5439 6815 5469 6841
rect 5744 6813 5774 6839
rect 6316 6838 6382 6866
rect 8204 6900 8270 6916
rect 8318 6912 8348 6938
rect 10110 6916 10140 6938
rect 8204 6866 8220 6900
rect 8254 6866 8270 6900
rect 6316 6819 6494 6838
rect 6940 6821 6970 6847
rect 4760 6659 4826 6675
rect 4760 6625 4776 6659
rect 4810 6625 4826 6659
rect 4760 6609 4826 6625
rect 5052 6669 5082 6691
rect 5052 6653 5138 6669
rect 5052 6619 5088 6653
rect 5122 6619 5138 6653
rect 5351 6650 5381 6711
rect 5439 6696 5469 6711
rect 5439 6672 5475 6696
rect 6316 6806 6444 6819
rect 6428 6785 6444 6806
rect 6478 6785 6494 6819
rect 6428 6769 6494 6785
rect 6350 6738 6380 6764
rect 6446 6738 6476 6769
rect 5445 6663 5475 6672
rect 4778 6578 4808 6609
rect 5052 6603 5138 6619
rect 5349 6634 5403 6650
rect 4462 6507 4492 6538
rect 4444 6491 4510 6507
rect 4444 6457 4460 6491
rect 4494 6457 4510 6491
rect 4444 6441 4510 6457
rect 4558 6454 4588 6538
rect 4558 6424 4644 6454
rect 3856 6337 3886 6363
rect 4132 6348 4162 6378
rect 4132 6347 4194 6348
rect 2872 6297 2888 6331
rect 2922 6297 2938 6331
rect 2872 6281 2938 6297
rect 4114 6331 4194 6347
rect 4114 6297 4130 6331
rect 4164 6297 4194 6331
rect 4114 6281 4194 6297
rect 2274 6236 2756 6266
rect 4162 6266 4194 6281
rect 4614 6266 4644 6424
rect 5052 6571 5082 6603
rect 5349 6600 5359 6634
rect 5393 6600 5403 6634
rect 5349 6584 5403 6600
rect 5445 6647 5521 6663
rect 5445 6613 5477 6647
rect 5511 6613 5521 6647
rect 5445 6597 5521 6613
rect 5744 6661 5774 6683
rect 5744 6645 5830 6661
rect 5744 6611 5780 6645
rect 5814 6611 5830 6645
rect 4778 6347 4808 6378
rect 5351 6523 5381 6584
rect 5445 6562 5475 6597
rect 5744 6595 5830 6611
rect 6002 6659 6068 6675
rect 6002 6625 6018 6659
rect 6052 6625 6068 6659
rect 6002 6609 6068 6625
rect 5744 6563 5774 6595
rect 6020 6578 6050 6609
rect 5439 6538 5475 6562
rect 5439 6523 5469 6538
rect 4760 6331 4826 6347
rect 5052 6345 5082 6371
rect 5351 6339 5381 6365
rect 5439 6339 5469 6365
rect 7239 6815 7269 6841
rect 7327 6815 7357 6841
rect 7632 6813 7662 6839
rect 8204 6838 8270 6866
rect 10092 6900 10158 6916
rect 10206 6912 10236 6938
rect 11998 6916 12028 6938
rect 10092 6866 10108 6900
rect 10142 6866 10158 6900
rect 8204 6819 8382 6838
rect 8828 6821 8858 6847
rect 6648 6659 6714 6675
rect 6648 6625 6664 6659
rect 6698 6625 6714 6659
rect 6648 6609 6714 6625
rect 6940 6669 6970 6691
rect 6940 6653 7026 6669
rect 6940 6619 6976 6653
rect 7010 6619 7026 6653
rect 7239 6650 7269 6711
rect 7327 6696 7357 6711
rect 7327 6672 7363 6696
rect 8204 6806 8332 6819
rect 8316 6785 8332 6806
rect 8366 6785 8382 6819
rect 8316 6769 8382 6785
rect 8238 6738 8268 6764
rect 8334 6738 8364 6769
rect 7333 6663 7363 6672
rect 6666 6578 6696 6609
rect 6940 6603 7026 6619
rect 7237 6634 7291 6650
rect 6350 6507 6380 6538
rect 6332 6491 6398 6507
rect 6332 6457 6348 6491
rect 6382 6457 6398 6491
rect 6332 6441 6398 6457
rect 6446 6454 6476 6538
rect 6446 6424 6532 6454
rect 5744 6337 5774 6363
rect 6020 6348 6050 6378
rect 6020 6347 6082 6348
rect 4760 6297 4776 6331
rect 4810 6297 4826 6331
rect 4760 6281 4826 6297
rect 6002 6331 6082 6347
rect 6002 6297 6018 6331
rect 6052 6297 6082 6331
rect 6002 6281 6082 6297
rect 4162 6236 4644 6266
rect 6050 6266 6082 6281
rect 6502 6266 6532 6424
rect 6940 6571 6970 6603
rect 7237 6600 7247 6634
rect 7281 6600 7291 6634
rect 7237 6584 7291 6600
rect 7333 6647 7409 6663
rect 7333 6613 7365 6647
rect 7399 6613 7409 6647
rect 7333 6597 7409 6613
rect 7632 6661 7662 6683
rect 7632 6645 7718 6661
rect 7632 6611 7668 6645
rect 7702 6611 7718 6645
rect 6666 6347 6696 6378
rect 7239 6523 7269 6584
rect 7333 6562 7363 6597
rect 7632 6595 7718 6611
rect 7890 6659 7956 6675
rect 7890 6625 7906 6659
rect 7940 6625 7956 6659
rect 7890 6609 7956 6625
rect 7632 6563 7662 6595
rect 7908 6578 7938 6609
rect 7327 6538 7363 6562
rect 7327 6523 7357 6538
rect 6648 6331 6714 6347
rect 6940 6345 6970 6371
rect 7239 6339 7269 6365
rect 7327 6339 7357 6365
rect 9127 6815 9157 6841
rect 9215 6815 9245 6841
rect 9520 6813 9550 6839
rect 10092 6838 10158 6866
rect 11980 6900 12046 6916
rect 12094 6912 12124 6938
rect 13886 6916 13916 6938
rect 11980 6866 11996 6900
rect 12030 6866 12046 6900
rect 10092 6819 10270 6838
rect 10716 6821 10746 6847
rect 8536 6659 8602 6675
rect 8536 6625 8552 6659
rect 8586 6625 8602 6659
rect 8536 6609 8602 6625
rect 8828 6669 8858 6691
rect 8828 6653 8914 6669
rect 8828 6619 8864 6653
rect 8898 6619 8914 6653
rect 9127 6650 9157 6711
rect 9215 6696 9245 6711
rect 9215 6672 9251 6696
rect 10092 6806 10220 6819
rect 10204 6785 10220 6806
rect 10254 6785 10270 6819
rect 10204 6769 10270 6785
rect 10126 6738 10156 6764
rect 10222 6738 10252 6769
rect 9221 6663 9251 6672
rect 8554 6578 8584 6609
rect 8828 6603 8914 6619
rect 9125 6634 9179 6650
rect 8238 6507 8268 6538
rect 8220 6491 8286 6507
rect 8220 6457 8236 6491
rect 8270 6457 8286 6491
rect 8220 6441 8286 6457
rect 8334 6454 8364 6538
rect 8334 6424 8420 6454
rect 7632 6337 7662 6363
rect 7908 6348 7938 6378
rect 7908 6347 7970 6348
rect 6648 6297 6664 6331
rect 6698 6297 6714 6331
rect 6648 6281 6714 6297
rect 7890 6331 7970 6347
rect 7890 6297 7906 6331
rect 7940 6297 7970 6331
rect 7890 6281 7970 6297
rect 6050 6236 6532 6266
rect 7938 6266 7970 6281
rect 8390 6266 8420 6424
rect 8828 6571 8858 6603
rect 9125 6600 9135 6634
rect 9169 6600 9179 6634
rect 9125 6584 9179 6600
rect 9221 6647 9297 6663
rect 9221 6613 9253 6647
rect 9287 6613 9297 6647
rect 9221 6597 9297 6613
rect 9520 6661 9550 6683
rect 9520 6645 9606 6661
rect 9520 6611 9556 6645
rect 9590 6611 9606 6645
rect 8554 6347 8584 6378
rect 9127 6523 9157 6584
rect 9221 6562 9251 6597
rect 9520 6595 9606 6611
rect 9778 6659 9844 6675
rect 9778 6625 9794 6659
rect 9828 6625 9844 6659
rect 9778 6609 9844 6625
rect 9520 6563 9550 6595
rect 9796 6578 9826 6609
rect 9215 6538 9251 6562
rect 9215 6523 9245 6538
rect 8536 6331 8602 6347
rect 8828 6345 8858 6371
rect 9127 6339 9157 6365
rect 9215 6339 9245 6365
rect 11015 6815 11045 6841
rect 11103 6815 11133 6841
rect 11408 6813 11438 6839
rect 11980 6838 12046 6866
rect 13868 6900 13934 6916
rect 13982 6912 14012 6938
rect 15768 6916 15798 6938
rect 13868 6866 13884 6900
rect 13918 6866 13934 6900
rect 11980 6819 12158 6838
rect 12604 6821 12634 6847
rect 10424 6659 10490 6675
rect 10424 6625 10440 6659
rect 10474 6625 10490 6659
rect 10424 6609 10490 6625
rect 10716 6669 10746 6691
rect 10716 6653 10802 6669
rect 10716 6619 10752 6653
rect 10786 6619 10802 6653
rect 11015 6650 11045 6711
rect 11103 6696 11133 6711
rect 11103 6672 11139 6696
rect 11980 6806 12108 6819
rect 12092 6785 12108 6806
rect 12142 6785 12158 6819
rect 12092 6769 12158 6785
rect 12014 6738 12044 6764
rect 12110 6738 12140 6769
rect 11109 6663 11139 6672
rect 10442 6578 10472 6609
rect 10716 6603 10802 6619
rect 11013 6634 11067 6650
rect 10126 6507 10156 6538
rect 10108 6491 10174 6507
rect 10108 6457 10124 6491
rect 10158 6457 10174 6491
rect 10108 6441 10174 6457
rect 10222 6454 10252 6538
rect 10222 6424 10308 6454
rect 9520 6337 9550 6363
rect 9796 6348 9826 6378
rect 9796 6347 9858 6348
rect 8536 6297 8552 6331
rect 8586 6297 8602 6331
rect 8536 6281 8602 6297
rect 9778 6331 9858 6347
rect 9778 6297 9794 6331
rect 9828 6297 9858 6331
rect 9778 6281 9858 6297
rect 7938 6236 8420 6266
rect 9826 6266 9858 6281
rect 10278 6266 10308 6424
rect 10716 6571 10746 6603
rect 11013 6600 11023 6634
rect 11057 6600 11067 6634
rect 11013 6584 11067 6600
rect 11109 6647 11185 6663
rect 11109 6613 11141 6647
rect 11175 6613 11185 6647
rect 11109 6597 11185 6613
rect 11408 6661 11438 6683
rect 11408 6645 11494 6661
rect 11408 6611 11444 6645
rect 11478 6611 11494 6645
rect 10442 6347 10472 6378
rect 11015 6523 11045 6584
rect 11109 6562 11139 6597
rect 11408 6595 11494 6611
rect 11666 6659 11732 6675
rect 11666 6625 11682 6659
rect 11716 6625 11732 6659
rect 11666 6609 11732 6625
rect 11408 6563 11438 6595
rect 11684 6578 11714 6609
rect 11103 6538 11139 6562
rect 11103 6523 11133 6538
rect 10424 6331 10490 6347
rect 10716 6345 10746 6371
rect 11015 6339 11045 6365
rect 11103 6339 11133 6365
rect 12903 6815 12933 6841
rect 12991 6815 13021 6841
rect 13296 6813 13326 6839
rect 13868 6838 13934 6866
rect 15750 6900 15816 6916
rect 15864 6912 15894 6938
rect 17656 6916 17686 6938
rect 15750 6866 15766 6900
rect 15800 6866 15816 6900
rect 13868 6819 14046 6838
rect 14492 6821 14522 6847
rect 12312 6659 12378 6675
rect 12312 6625 12328 6659
rect 12362 6625 12378 6659
rect 12312 6609 12378 6625
rect 12604 6669 12634 6691
rect 12604 6653 12690 6669
rect 12604 6619 12640 6653
rect 12674 6619 12690 6653
rect 12903 6650 12933 6711
rect 12991 6696 13021 6711
rect 12991 6672 13027 6696
rect 13868 6806 13996 6819
rect 13980 6785 13996 6806
rect 14030 6785 14046 6819
rect 13980 6769 14046 6785
rect 13902 6738 13932 6764
rect 13998 6738 14028 6769
rect 12997 6663 13027 6672
rect 12330 6578 12360 6609
rect 12604 6603 12690 6619
rect 12901 6634 12955 6650
rect 12014 6507 12044 6538
rect 11996 6491 12062 6507
rect 11996 6457 12012 6491
rect 12046 6457 12062 6491
rect 11996 6441 12062 6457
rect 12110 6454 12140 6538
rect 12110 6424 12196 6454
rect 11408 6337 11438 6363
rect 11684 6348 11714 6378
rect 11684 6347 11746 6348
rect 10424 6297 10440 6331
rect 10474 6297 10490 6331
rect 10424 6281 10490 6297
rect 11666 6331 11746 6347
rect 11666 6297 11682 6331
rect 11716 6297 11746 6331
rect 11666 6281 11746 6297
rect 9826 6236 10308 6266
rect 11714 6266 11746 6281
rect 12166 6266 12196 6424
rect 12604 6571 12634 6603
rect 12901 6600 12911 6634
rect 12945 6600 12955 6634
rect 12901 6584 12955 6600
rect 12997 6647 13073 6663
rect 12997 6613 13029 6647
rect 13063 6613 13073 6647
rect 12997 6597 13073 6613
rect 13296 6661 13326 6683
rect 13296 6645 13382 6661
rect 13296 6611 13332 6645
rect 13366 6611 13382 6645
rect 12330 6347 12360 6378
rect 12903 6523 12933 6584
rect 12997 6562 13027 6597
rect 13296 6595 13382 6611
rect 13554 6659 13620 6675
rect 13554 6625 13570 6659
rect 13604 6625 13620 6659
rect 13554 6609 13620 6625
rect 13296 6563 13326 6595
rect 13572 6578 13602 6609
rect 12991 6538 13027 6562
rect 12991 6523 13021 6538
rect 12312 6331 12378 6347
rect 12604 6345 12634 6371
rect 12903 6339 12933 6365
rect 12991 6339 13021 6365
rect 14785 6815 14815 6841
rect 14873 6815 14903 6841
rect 15178 6813 15208 6839
rect 15750 6838 15816 6866
rect 17638 6900 17704 6916
rect 17752 6912 17782 6938
rect 19544 6916 19574 6938
rect 17638 6866 17654 6900
rect 17688 6866 17704 6900
rect 15750 6819 15928 6838
rect 16374 6821 16404 6847
rect 14200 6659 14266 6675
rect 14200 6625 14216 6659
rect 14250 6625 14266 6659
rect 14200 6609 14266 6625
rect 14492 6669 14522 6691
rect 14492 6653 14578 6669
rect 14492 6619 14528 6653
rect 14562 6619 14578 6653
rect 14785 6650 14815 6711
rect 14873 6696 14903 6711
rect 14873 6672 14909 6696
rect 15750 6806 15878 6819
rect 15862 6785 15878 6806
rect 15912 6785 15928 6819
rect 15862 6769 15928 6785
rect 15784 6738 15814 6764
rect 15880 6738 15910 6769
rect 14879 6663 14909 6672
rect 14218 6578 14248 6609
rect 14492 6603 14578 6619
rect 14783 6634 14837 6650
rect 13902 6507 13932 6538
rect 13884 6491 13950 6507
rect 13884 6457 13900 6491
rect 13934 6457 13950 6491
rect 13884 6441 13950 6457
rect 13998 6454 14028 6538
rect 13998 6424 14084 6454
rect 13296 6337 13326 6363
rect 13572 6348 13602 6378
rect 13572 6347 13634 6348
rect 12312 6297 12328 6331
rect 12362 6297 12378 6331
rect 12312 6281 12378 6297
rect 13554 6331 13634 6347
rect 13554 6297 13570 6331
rect 13604 6297 13634 6331
rect 13554 6281 13634 6297
rect 11714 6236 12196 6266
rect 13602 6266 13634 6281
rect 14054 6266 14084 6424
rect 14492 6571 14522 6603
rect 14783 6600 14793 6634
rect 14827 6600 14837 6634
rect 14783 6584 14837 6600
rect 14879 6647 14955 6663
rect 14879 6613 14911 6647
rect 14945 6613 14955 6647
rect 14879 6597 14955 6613
rect 15178 6661 15208 6683
rect 15178 6645 15264 6661
rect 15178 6611 15214 6645
rect 15248 6611 15264 6645
rect 14218 6347 14248 6378
rect 14785 6523 14815 6584
rect 14879 6562 14909 6597
rect 15178 6595 15264 6611
rect 15436 6659 15502 6675
rect 15436 6625 15452 6659
rect 15486 6625 15502 6659
rect 15436 6609 15502 6625
rect 15178 6563 15208 6595
rect 15454 6578 15484 6609
rect 14873 6538 14909 6562
rect 14873 6523 14903 6538
rect 14200 6331 14266 6347
rect 14492 6345 14522 6371
rect 14785 6339 14815 6365
rect 14873 6339 14903 6365
rect 16673 6815 16703 6841
rect 16761 6815 16791 6841
rect 17066 6813 17096 6839
rect 17638 6838 17704 6866
rect 19526 6900 19592 6916
rect 19640 6912 19670 6938
rect 21432 6916 21462 6938
rect 19526 6866 19542 6900
rect 19576 6866 19592 6900
rect 17638 6819 17816 6838
rect 18262 6821 18292 6847
rect 16082 6659 16148 6675
rect 16082 6625 16098 6659
rect 16132 6625 16148 6659
rect 16082 6609 16148 6625
rect 16374 6669 16404 6691
rect 16374 6653 16460 6669
rect 16374 6619 16410 6653
rect 16444 6619 16460 6653
rect 16673 6650 16703 6711
rect 16761 6696 16791 6711
rect 16761 6672 16797 6696
rect 17638 6806 17766 6819
rect 17750 6785 17766 6806
rect 17800 6785 17816 6819
rect 17750 6769 17816 6785
rect 17672 6738 17702 6764
rect 17768 6738 17798 6769
rect 16767 6663 16797 6672
rect 16100 6578 16130 6609
rect 16374 6603 16460 6619
rect 16671 6634 16725 6650
rect 15784 6507 15814 6538
rect 15766 6491 15832 6507
rect 15766 6457 15782 6491
rect 15816 6457 15832 6491
rect 15766 6441 15832 6457
rect 15880 6454 15910 6538
rect 15880 6424 15966 6454
rect 15178 6337 15208 6363
rect 15454 6348 15484 6378
rect 15454 6347 15516 6348
rect 14200 6297 14216 6331
rect 14250 6297 14266 6331
rect 14200 6281 14266 6297
rect 15436 6331 15516 6347
rect 15436 6297 15452 6331
rect 15486 6297 15516 6331
rect 15436 6281 15516 6297
rect 13602 6236 14084 6266
rect 15484 6266 15516 6281
rect 15936 6266 15966 6424
rect 16374 6571 16404 6603
rect 16671 6600 16681 6634
rect 16715 6600 16725 6634
rect 16671 6584 16725 6600
rect 16767 6647 16843 6663
rect 16767 6613 16799 6647
rect 16833 6613 16843 6647
rect 16767 6597 16843 6613
rect 17066 6661 17096 6683
rect 17066 6645 17152 6661
rect 17066 6611 17102 6645
rect 17136 6611 17152 6645
rect 16100 6347 16130 6378
rect 16673 6523 16703 6584
rect 16767 6562 16797 6597
rect 17066 6595 17152 6611
rect 17324 6659 17390 6675
rect 17324 6625 17340 6659
rect 17374 6625 17390 6659
rect 17324 6609 17390 6625
rect 17066 6563 17096 6595
rect 17342 6578 17372 6609
rect 16761 6538 16797 6562
rect 16761 6523 16791 6538
rect 16082 6331 16148 6347
rect 16374 6345 16404 6371
rect 16673 6339 16703 6365
rect 16761 6339 16791 6365
rect 18561 6815 18591 6841
rect 18649 6815 18679 6841
rect 18954 6813 18984 6839
rect 19526 6838 19592 6866
rect 21414 6900 21480 6916
rect 21528 6912 21558 6938
rect 23320 6916 23350 6938
rect 21414 6866 21430 6900
rect 21464 6866 21480 6900
rect 19526 6819 19704 6838
rect 20150 6821 20180 6847
rect 17970 6659 18036 6675
rect 17970 6625 17986 6659
rect 18020 6625 18036 6659
rect 17970 6609 18036 6625
rect 18262 6669 18292 6691
rect 18262 6653 18348 6669
rect 18262 6619 18298 6653
rect 18332 6619 18348 6653
rect 18561 6650 18591 6711
rect 18649 6696 18679 6711
rect 18649 6672 18685 6696
rect 19526 6806 19654 6819
rect 19638 6785 19654 6806
rect 19688 6785 19704 6819
rect 19638 6769 19704 6785
rect 19560 6738 19590 6764
rect 19656 6738 19686 6769
rect 18655 6663 18685 6672
rect 17988 6578 18018 6609
rect 18262 6603 18348 6619
rect 18559 6634 18613 6650
rect 17672 6507 17702 6538
rect 17654 6491 17720 6507
rect 17654 6457 17670 6491
rect 17704 6457 17720 6491
rect 17654 6441 17720 6457
rect 17768 6454 17798 6538
rect 17768 6424 17854 6454
rect 17066 6337 17096 6363
rect 17342 6348 17372 6378
rect 17342 6347 17404 6348
rect 16082 6297 16098 6331
rect 16132 6297 16148 6331
rect 16082 6281 16148 6297
rect 17324 6331 17404 6347
rect 17324 6297 17340 6331
rect 17374 6297 17404 6331
rect 17324 6281 17404 6297
rect 15484 6236 15966 6266
rect 17372 6266 17404 6281
rect 17824 6266 17854 6424
rect 18262 6571 18292 6603
rect 18559 6600 18569 6634
rect 18603 6600 18613 6634
rect 18559 6584 18613 6600
rect 18655 6647 18731 6663
rect 18655 6613 18687 6647
rect 18721 6613 18731 6647
rect 18655 6597 18731 6613
rect 18954 6661 18984 6683
rect 18954 6645 19040 6661
rect 18954 6611 18990 6645
rect 19024 6611 19040 6645
rect 17988 6347 18018 6378
rect 18561 6523 18591 6584
rect 18655 6562 18685 6597
rect 18954 6595 19040 6611
rect 19212 6659 19278 6675
rect 19212 6625 19228 6659
rect 19262 6625 19278 6659
rect 19212 6609 19278 6625
rect 18954 6563 18984 6595
rect 19230 6578 19260 6609
rect 18649 6538 18685 6562
rect 18649 6523 18679 6538
rect 17970 6331 18036 6347
rect 18262 6345 18292 6371
rect 18561 6339 18591 6365
rect 18649 6339 18679 6365
rect 20449 6815 20479 6841
rect 20537 6815 20567 6841
rect 20842 6813 20872 6839
rect 21414 6838 21480 6866
rect 23302 6900 23368 6916
rect 23416 6912 23446 6938
rect 25208 6916 25238 6938
rect 23302 6866 23318 6900
rect 23352 6866 23368 6900
rect 21414 6819 21592 6838
rect 22038 6821 22068 6847
rect 19858 6659 19924 6675
rect 19858 6625 19874 6659
rect 19908 6625 19924 6659
rect 19858 6609 19924 6625
rect 20150 6669 20180 6691
rect 20150 6653 20236 6669
rect 20150 6619 20186 6653
rect 20220 6619 20236 6653
rect 20449 6650 20479 6711
rect 20537 6696 20567 6711
rect 20537 6672 20573 6696
rect 21414 6806 21542 6819
rect 21526 6785 21542 6806
rect 21576 6785 21592 6819
rect 21526 6769 21592 6785
rect 21448 6738 21478 6764
rect 21544 6738 21574 6769
rect 20543 6663 20573 6672
rect 19876 6578 19906 6609
rect 20150 6603 20236 6619
rect 20447 6634 20501 6650
rect 19560 6507 19590 6538
rect 19542 6491 19608 6507
rect 19542 6457 19558 6491
rect 19592 6457 19608 6491
rect 19542 6441 19608 6457
rect 19656 6454 19686 6538
rect 19656 6424 19742 6454
rect 18954 6337 18984 6363
rect 19230 6348 19260 6378
rect 19230 6347 19292 6348
rect 17970 6297 17986 6331
rect 18020 6297 18036 6331
rect 17970 6281 18036 6297
rect 19212 6331 19292 6347
rect 19212 6297 19228 6331
rect 19262 6297 19292 6331
rect 19212 6281 19292 6297
rect 17372 6236 17854 6266
rect 19260 6266 19292 6281
rect 19712 6266 19742 6424
rect 20150 6571 20180 6603
rect 20447 6600 20457 6634
rect 20491 6600 20501 6634
rect 20447 6584 20501 6600
rect 20543 6647 20619 6663
rect 20543 6613 20575 6647
rect 20609 6613 20619 6647
rect 20543 6597 20619 6613
rect 20842 6661 20872 6683
rect 20842 6645 20928 6661
rect 20842 6611 20878 6645
rect 20912 6611 20928 6645
rect 19876 6347 19906 6378
rect 20449 6523 20479 6584
rect 20543 6562 20573 6597
rect 20842 6595 20928 6611
rect 21100 6659 21166 6675
rect 21100 6625 21116 6659
rect 21150 6625 21166 6659
rect 21100 6609 21166 6625
rect 20842 6563 20872 6595
rect 21118 6578 21148 6609
rect 20537 6538 20573 6562
rect 20537 6523 20567 6538
rect 19858 6331 19924 6347
rect 20150 6345 20180 6371
rect 20449 6339 20479 6365
rect 20537 6339 20567 6365
rect 22337 6815 22367 6841
rect 22425 6815 22455 6841
rect 22730 6813 22760 6839
rect 23302 6838 23368 6866
rect 25190 6900 25256 6916
rect 25304 6912 25334 6938
rect 27096 6916 27126 6938
rect 25190 6866 25206 6900
rect 25240 6866 25256 6900
rect 23302 6819 23480 6838
rect 23926 6821 23956 6847
rect 21746 6659 21812 6675
rect 21746 6625 21762 6659
rect 21796 6625 21812 6659
rect 21746 6609 21812 6625
rect 22038 6669 22068 6691
rect 22038 6653 22124 6669
rect 22038 6619 22074 6653
rect 22108 6619 22124 6653
rect 22337 6650 22367 6711
rect 22425 6696 22455 6711
rect 22425 6672 22461 6696
rect 23302 6806 23430 6819
rect 23414 6785 23430 6806
rect 23464 6785 23480 6819
rect 23414 6769 23480 6785
rect 23336 6738 23366 6764
rect 23432 6738 23462 6769
rect 22431 6663 22461 6672
rect 21764 6578 21794 6609
rect 22038 6603 22124 6619
rect 22335 6634 22389 6650
rect 21448 6507 21478 6538
rect 21430 6491 21496 6507
rect 21430 6457 21446 6491
rect 21480 6457 21496 6491
rect 21430 6441 21496 6457
rect 21544 6454 21574 6538
rect 21544 6424 21630 6454
rect 20842 6337 20872 6363
rect 21118 6348 21148 6378
rect 21118 6347 21180 6348
rect 19858 6297 19874 6331
rect 19908 6297 19924 6331
rect 19858 6281 19924 6297
rect 21100 6331 21180 6347
rect 21100 6297 21116 6331
rect 21150 6297 21180 6331
rect 21100 6281 21180 6297
rect 19260 6236 19742 6266
rect 21148 6266 21180 6281
rect 21600 6266 21630 6424
rect 22038 6571 22068 6603
rect 22335 6600 22345 6634
rect 22379 6600 22389 6634
rect 22335 6584 22389 6600
rect 22431 6647 22507 6663
rect 22431 6613 22463 6647
rect 22497 6613 22507 6647
rect 22431 6597 22507 6613
rect 22730 6661 22760 6683
rect 22730 6645 22816 6661
rect 22730 6611 22766 6645
rect 22800 6611 22816 6645
rect 21764 6347 21794 6378
rect 22337 6523 22367 6584
rect 22431 6562 22461 6597
rect 22730 6595 22816 6611
rect 22988 6659 23054 6675
rect 22988 6625 23004 6659
rect 23038 6625 23054 6659
rect 22988 6609 23054 6625
rect 22730 6563 22760 6595
rect 23006 6578 23036 6609
rect 22425 6538 22461 6562
rect 22425 6523 22455 6538
rect 21746 6331 21812 6347
rect 22038 6345 22068 6371
rect 22337 6339 22367 6365
rect 22425 6339 22455 6365
rect 24225 6815 24255 6841
rect 24313 6815 24343 6841
rect 24618 6813 24648 6839
rect 25190 6838 25256 6866
rect 27078 6900 27144 6916
rect 27192 6912 27222 6938
rect 28984 6916 29014 6938
rect 27078 6866 27094 6900
rect 27128 6866 27144 6900
rect 25190 6819 25368 6838
rect 25814 6821 25844 6847
rect 23634 6659 23700 6675
rect 23634 6625 23650 6659
rect 23684 6625 23700 6659
rect 23634 6609 23700 6625
rect 23926 6669 23956 6691
rect 23926 6653 24012 6669
rect 23926 6619 23962 6653
rect 23996 6619 24012 6653
rect 24225 6650 24255 6711
rect 24313 6696 24343 6711
rect 24313 6672 24349 6696
rect 25190 6806 25318 6819
rect 25302 6785 25318 6806
rect 25352 6785 25368 6819
rect 25302 6769 25368 6785
rect 25224 6738 25254 6764
rect 25320 6738 25350 6769
rect 24319 6663 24349 6672
rect 23652 6578 23682 6609
rect 23926 6603 24012 6619
rect 24223 6634 24277 6650
rect 23336 6507 23366 6538
rect 23318 6491 23384 6507
rect 23318 6457 23334 6491
rect 23368 6457 23384 6491
rect 23318 6441 23384 6457
rect 23432 6454 23462 6538
rect 23432 6424 23518 6454
rect 22730 6337 22760 6363
rect 23006 6348 23036 6378
rect 23006 6347 23068 6348
rect 21746 6297 21762 6331
rect 21796 6297 21812 6331
rect 21746 6281 21812 6297
rect 22988 6331 23068 6347
rect 22988 6297 23004 6331
rect 23038 6297 23068 6331
rect 22988 6281 23068 6297
rect 21148 6236 21630 6266
rect 23036 6266 23068 6281
rect 23488 6266 23518 6424
rect 23926 6571 23956 6603
rect 24223 6600 24233 6634
rect 24267 6600 24277 6634
rect 24223 6584 24277 6600
rect 24319 6647 24395 6663
rect 24319 6613 24351 6647
rect 24385 6613 24395 6647
rect 24319 6597 24395 6613
rect 24618 6661 24648 6683
rect 24618 6645 24704 6661
rect 24618 6611 24654 6645
rect 24688 6611 24704 6645
rect 23652 6347 23682 6378
rect 24225 6523 24255 6584
rect 24319 6562 24349 6597
rect 24618 6595 24704 6611
rect 24876 6659 24942 6675
rect 24876 6625 24892 6659
rect 24926 6625 24942 6659
rect 24876 6609 24942 6625
rect 24618 6563 24648 6595
rect 24894 6578 24924 6609
rect 24313 6538 24349 6562
rect 24313 6523 24343 6538
rect 23634 6331 23700 6347
rect 23926 6345 23956 6371
rect 24225 6339 24255 6365
rect 24313 6339 24343 6365
rect 26113 6815 26143 6841
rect 26201 6815 26231 6841
rect 26506 6813 26536 6839
rect 27078 6838 27144 6866
rect 28966 6900 29032 6916
rect 29080 6912 29110 6938
rect 30872 6916 30902 6938
rect 28966 6866 28982 6900
rect 29016 6866 29032 6900
rect 27078 6819 27256 6838
rect 27702 6821 27732 6847
rect 25522 6659 25588 6675
rect 25522 6625 25538 6659
rect 25572 6625 25588 6659
rect 25522 6609 25588 6625
rect 25814 6669 25844 6691
rect 25814 6653 25900 6669
rect 25814 6619 25850 6653
rect 25884 6619 25900 6653
rect 26113 6650 26143 6711
rect 26201 6696 26231 6711
rect 26201 6672 26237 6696
rect 27078 6806 27206 6819
rect 27190 6785 27206 6806
rect 27240 6785 27256 6819
rect 27190 6769 27256 6785
rect 27112 6738 27142 6764
rect 27208 6738 27238 6769
rect 26207 6663 26237 6672
rect 25540 6578 25570 6609
rect 25814 6603 25900 6619
rect 26111 6634 26165 6650
rect 25224 6507 25254 6538
rect 25206 6491 25272 6507
rect 25206 6457 25222 6491
rect 25256 6457 25272 6491
rect 25206 6441 25272 6457
rect 25320 6454 25350 6538
rect 25320 6424 25406 6454
rect 24618 6337 24648 6363
rect 24894 6348 24924 6378
rect 24894 6347 24956 6348
rect 23634 6297 23650 6331
rect 23684 6297 23700 6331
rect 23634 6281 23700 6297
rect 24876 6331 24956 6347
rect 24876 6297 24892 6331
rect 24926 6297 24956 6331
rect 24876 6281 24956 6297
rect 23036 6236 23518 6266
rect 24924 6266 24956 6281
rect 25376 6266 25406 6424
rect 25814 6571 25844 6603
rect 26111 6600 26121 6634
rect 26155 6600 26165 6634
rect 26111 6584 26165 6600
rect 26207 6647 26283 6663
rect 26207 6613 26239 6647
rect 26273 6613 26283 6647
rect 26207 6597 26283 6613
rect 26506 6661 26536 6683
rect 26506 6645 26592 6661
rect 26506 6611 26542 6645
rect 26576 6611 26592 6645
rect 25540 6347 25570 6378
rect 26113 6523 26143 6584
rect 26207 6562 26237 6597
rect 26506 6595 26592 6611
rect 26764 6659 26830 6675
rect 26764 6625 26780 6659
rect 26814 6625 26830 6659
rect 26764 6609 26830 6625
rect 26506 6563 26536 6595
rect 26782 6578 26812 6609
rect 26201 6538 26237 6562
rect 26201 6523 26231 6538
rect 25522 6331 25588 6347
rect 25814 6345 25844 6371
rect 26113 6339 26143 6365
rect 26201 6339 26231 6365
rect 28001 6815 28031 6841
rect 28089 6815 28119 6841
rect 28394 6813 28424 6839
rect 28966 6838 29032 6866
rect 30854 6900 30920 6916
rect 30968 6912 30998 6938
rect 32760 6916 32790 6938
rect 30854 6866 30870 6900
rect 30904 6866 30920 6900
rect 28966 6819 29144 6838
rect 29590 6821 29620 6847
rect 27410 6659 27476 6675
rect 27410 6625 27426 6659
rect 27460 6625 27476 6659
rect 27410 6609 27476 6625
rect 27702 6669 27732 6691
rect 27702 6653 27788 6669
rect 27702 6619 27738 6653
rect 27772 6619 27788 6653
rect 28001 6650 28031 6711
rect 28089 6696 28119 6711
rect 28089 6672 28125 6696
rect 28966 6806 29094 6819
rect 29078 6785 29094 6806
rect 29128 6785 29144 6819
rect 29078 6769 29144 6785
rect 29000 6738 29030 6764
rect 29096 6738 29126 6769
rect 28095 6663 28125 6672
rect 27428 6578 27458 6609
rect 27702 6603 27788 6619
rect 27999 6634 28053 6650
rect 27112 6507 27142 6538
rect 27094 6491 27160 6507
rect 27094 6457 27110 6491
rect 27144 6457 27160 6491
rect 27094 6441 27160 6457
rect 27208 6454 27238 6538
rect 27208 6424 27294 6454
rect 26506 6337 26536 6363
rect 26782 6348 26812 6378
rect 26782 6347 26844 6348
rect 25522 6297 25538 6331
rect 25572 6297 25588 6331
rect 25522 6281 25588 6297
rect 26764 6331 26844 6347
rect 26764 6297 26780 6331
rect 26814 6297 26844 6331
rect 26764 6281 26844 6297
rect 24924 6236 25406 6266
rect 26812 6266 26844 6281
rect 27264 6266 27294 6424
rect 27702 6571 27732 6603
rect 27999 6600 28009 6634
rect 28043 6600 28053 6634
rect 27999 6584 28053 6600
rect 28095 6647 28171 6663
rect 28095 6613 28127 6647
rect 28161 6613 28171 6647
rect 28095 6597 28171 6613
rect 28394 6661 28424 6683
rect 28394 6645 28480 6661
rect 28394 6611 28430 6645
rect 28464 6611 28480 6645
rect 27428 6347 27458 6378
rect 28001 6523 28031 6584
rect 28095 6562 28125 6597
rect 28394 6595 28480 6611
rect 28652 6659 28718 6675
rect 28652 6625 28668 6659
rect 28702 6625 28718 6659
rect 28652 6609 28718 6625
rect 28394 6563 28424 6595
rect 28670 6578 28700 6609
rect 28089 6538 28125 6562
rect 28089 6523 28119 6538
rect 27410 6331 27476 6347
rect 27702 6345 27732 6371
rect 28001 6339 28031 6365
rect 28089 6339 28119 6365
rect 29889 6815 29919 6841
rect 29977 6815 30007 6841
rect 30282 6813 30312 6839
rect 30854 6838 30920 6866
rect 32742 6900 32808 6916
rect 32856 6912 32886 6938
rect 34648 6916 34678 6938
rect 32742 6866 32758 6900
rect 32792 6866 32808 6900
rect 30854 6819 31032 6838
rect 31478 6821 31508 6847
rect 29298 6659 29364 6675
rect 29298 6625 29314 6659
rect 29348 6625 29364 6659
rect 29298 6609 29364 6625
rect 29590 6669 29620 6691
rect 29590 6653 29676 6669
rect 29590 6619 29626 6653
rect 29660 6619 29676 6653
rect 29889 6650 29919 6711
rect 29977 6696 30007 6711
rect 29977 6672 30013 6696
rect 30854 6806 30982 6819
rect 30966 6785 30982 6806
rect 31016 6785 31032 6819
rect 30966 6769 31032 6785
rect 30888 6738 30918 6764
rect 30984 6738 31014 6769
rect 29983 6663 30013 6672
rect 29316 6578 29346 6609
rect 29590 6603 29676 6619
rect 29887 6634 29941 6650
rect 29000 6507 29030 6538
rect 28982 6491 29048 6507
rect 28982 6457 28998 6491
rect 29032 6457 29048 6491
rect 28982 6441 29048 6457
rect 29096 6454 29126 6538
rect 29096 6424 29182 6454
rect 28394 6337 28424 6363
rect 28670 6348 28700 6378
rect 28670 6347 28732 6348
rect 27410 6297 27426 6331
rect 27460 6297 27476 6331
rect 27410 6281 27476 6297
rect 28652 6331 28732 6347
rect 28652 6297 28668 6331
rect 28702 6297 28732 6331
rect 28652 6281 28732 6297
rect 26812 6236 27294 6266
rect 28700 6266 28732 6281
rect 29152 6266 29182 6424
rect 29590 6571 29620 6603
rect 29887 6600 29897 6634
rect 29931 6600 29941 6634
rect 29887 6584 29941 6600
rect 29983 6647 30059 6663
rect 29983 6613 30015 6647
rect 30049 6613 30059 6647
rect 29983 6597 30059 6613
rect 30282 6661 30312 6683
rect 30282 6645 30368 6661
rect 30282 6611 30318 6645
rect 30352 6611 30368 6645
rect 29316 6347 29346 6378
rect 29889 6523 29919 6584
rect 29983 6562 30013 6597
rect 30282 6595 30368 6611
rect 30540 6659 30606 6675
rect 30540 6625 30556 6659
rect 30590 6625 30606 6659
rect 30540 6609 30606 6625
rect 30282 6563 30312 6595
rect 30558 6578 30588 6609
rect 29977 6538 30013 6562
rect 29977 6523 30007 6538
rect 29298 6331 29364 6347
rect 29590 6345 29620 6371
rect 29889 6339 29919 6365
rect 29977 6339 30007 6365
rect 31777 6815 31807 6841
rect 31865 6815 31895 6841
rect 32170 6813 32200 6839
rect 32742 6838 32808 6866
rect 34630 6900 34696 6916
rect 34744 6912 34774 6938
rect 36536 6916 36566 6938
rect 34630 6866 34646 6900
rect 34680 6866 34696 6900
rect 32742 6819 32920 6838
rect 33366 6821 33396 6847
rect 31186 6659 31252 6675
rect 31186 6625 31202 6659
rect 31236 6625 31252 6659
rect 31186 6609 31252 6625
rect 31478 6669 31508 6691
rect 31478 6653 31564 6669
rect 31478 6619 31514 6653
rect 31548 6619 31564 6653
rect 31777 6650 31807 6711
rect 31865 6696 31895 6711
rect 31865 6672 31901 6696
rect 32742 6806 32870 6819
rect 32854 6785 32870 6806
rect 32904 6785 32920 6819
rect 32854 6769 32920 6785
rect 32776 6738 32806 6764
rect 32872 6738 32902 6769
rect 31871 6663 31901 6672
rect 31204 6578 31234 6609
rect 31478 6603 31564 6619
rect 31775 6634 31829 6650
rect 30888 6507 30918 6538
rect 30870 6491 30936 6507
rect 30870 6457 30886 6491
rect 30920 6457 30936 6491
rect 30870 6441 30936 6457
rect 30984 6454 31014 6538
rect 30984 6424 31070 6454
rect 30282 6337 30312 6363
rect 30558 6348 30588 6378
rect 30558 6347 30620 6348
rect 29298 6297 29314 6331
rect 29348 6297 29364 6331
rect 29298 6281 29364 6297
rect 30540 6331 30620 6347
rect 30540 6297 30556 6331
rect 30590 6297 30620 6331
rect 30540 6281 30620 6297
rect 28700 6236 29182 6266
rect 30588 6266 30620 6281
rect 31040 6266 31070 6424
rect 31478 6571 31508 6603
rect 31775 6600 31785 6634
rect 31819 6600 31829 6634
rect 31775 6584 31829 6600
rect 31871 6647 31947 6663
rect 31871 6613 31903 6647
rect 31937 6613 31947 6647
rect 31871 6597 31947 6613
rect 32170 6661 32200 6683
rect 32170 6645 32256 6661
rect 32170 6611 32206 6645
rect 32240 6611 32256 6645
rect 31204 6347 31234 6378
rect 31777 6523 31807 6584
rect 31871 6562 31901 6597
rect 32170 6595 32256 6611
rect 32428 6659 32494 6675
rect 32428 6625 32444 6659
rect 32478 6625 32494 6659
rect 32428 6609 32494 6625
rect 32170 6563 32200 6595
rect 32446 6578 32476 6609
rect 31865 6538 31901 6562
rect 31865 6523 31895 6538
rect 31186 6331 31252 6347
rect 31478 6345 31508 6371
rect 31777 6339 31807 6365
rect 31865 6339 31895 6365
rect 33665 6815 33695 6841
rect 33753 6815 33783 6841
rect 34058 6813 34088 6839
rect 34630 6838 34696 6866
rect 36518 6900 36584 6916
rect 36632 6912 36662 6938
rect 38424 6916 38454 6938
rect 36518 6866 36534 6900
rect 36568 6866 36584 6900
rect 34630 6819 34808 6838
rect 35254 6821 35284 6847
rect 33074 6659 33140 6675
rect 33074 6625 33090 6659
rect 33124 6625 33140 6659
rect 33074 6609 33140 6625
rect 33366 6669 33396 6691
rect 33366 6653 33452 6669
rect 33366 6619 33402 6653
rect 33436 6619 33452 6653
rect 33665 6650 33695 6711
rect 33753 6696 33783 6711
rect 33753 6672 33789 6696
rect 34630 6806 34758 6819
rect 34742 6785 34758 6806
rect 34792 6785 34808 6819
rect 34742 6769 34808 6785
rect 34664 6738 34694 6764
rect 34760 6738 34790 6769
rect 33759 6663 33789 6672
rect 33092 6578 33122 6609
rect 33366 6603 33452 6619
rect 33663 6634 33717 6650
rect 32776 6507 32806 6538
rect 32758 6491 32824 6507
rect 32758 6457 32774 6491
rect 32808 6457 32824 6491
rect 32758 6441 32824 6457
rect 32872 6454 32902 6538
rect 32872 6424 32958 6454
rect 32170 6337 32200 6363
rect 32446 6348 32476 6378
rect 32446 6347 32508 6348
rect 31186 6297 31202 6331
rect 31236 6297 31252 6331
rect 31186 6281 31252 6297
rect 32428 6331 32508 6347
rect 32428 6297 32444 6331
rect 32478 6297 32508 6331
rect 32428 6281 32508 6297
rect 30588 6236 31070 6266
rect 32476 6266 32508 6281
rect 32928 6266 32958 6424
rect 33366 6571 33396 6603
rect 33663 6600 33673 6634
rect 33707 6600 33717 6634
rect 33663 6584 33717 6600
rect 33759 6647 33835 6663
rect 33759 6613 33791 6647
rect 33825 6613 33835 6647
rect 33759 6597 33835 6613
rect 34058 6661 34088 6683
rect 34058 6645 34144 6661
rect 34058 6611 34094 6645
rect 34128 6611 34144 6645
rect 33092 6347 33122 6378
rect 33665 6523 33695 6584
rect 33759 6562 33789 6597
rect 34058 6595 34144 6611
rect 34316 6659 34382 6675
rect 34316 6625 34332 6659
rect 34366 6625 34382 6659
rect 34316 6609 34382 6625
rect 34058 6563 34088 6595
rect 34334 6578 34364 6609
rect 33753 6538 33789 6562
rect 33753 6523 33783 6538
rect 33074 6331 33140 6347
rect 33366 6345 33396 6371
rect 33665 6339 33695 6365
rect 33753 6339 33783 6365
rect 35553 6815 35583 6841
rect 35641 6815 35671 6841
rect 35946 6813 35976 6839
rect 36518 6838 36584 6866
rect 38406 6900 38472 6916
rect 38520 6912 38550 6938
rect 40312 6916 40342 6938
rect 38406 6866 38422 6900
rect 38456 6866 38472 6900
rect 36518 6819 36696 6838
rect 37142 6821 37172 6847
rect 34962 6659 35028 6675
rect 34962 6625 34978 6659
rect 35012 6625 35028 6659
rect 34962 6609 35028 6625
rect 35254 6669 35284 6691
rect 35254 6653 35340 6669
rect 35254 6619 35290 6653
rect 35324 6619 35340 6653
rect 35553 6650 35583 6711
rect 35641 6696 35671 6711
rect 35641 6672 35677 6696
rect 36518 6806 36646 6819
rect 36630 6785 36646 6806
rect 36680 6785 36696 6819
rect 36630 6769 36696 6785
rect 36552 6738 36582 6764
rect 36648 6738 36678 6769
rect 35647 6663 35677 6672
rect 34980 6578 35010 6609
rect 35254 6603 35340 6619
rect 35551 6634 35605 6650
rect 34664 6507 34694 6538
rect 34646 6491 34712 6507
rect 34646 6457 34662 6491
rect 34696 6457 34712 6491
rect 34646 6441 34712 6457
rect 34760 6454 34790 6538
rect 34760 6424 34846 6454
rect 34058 6337 34088 6363
rect 34334 6348 34364 6378
rect 34334 6347 34396 6348
rect 33074 6297 33090 6331
rect 33124 6297 33140 6331
rect 33074 6281 33140 6297
rect 34316 6331 34396 6347
rect 34316 6297 34332 6331
rect 34366 6297 34396 6331
rect 34316 6281 34396 6297
rect 32476 6236 32958 6266
rect 34364 6266 34396 6281
rect 34816 6266 34846 6424
rect 35254 6571 35284 6603
rect 35551 6600 35561 6634
rect 35595 6600 35605 6634
rect 35551 6584 35605 6600
rect 35647 6647 35723 6663
rect 35647 6613 35679 6647
rect 35713 6613 35723 6647
rect 35647 6597 35723 6613
rect 35946 6661 35976 6683
rect 35946 6645 36032 6661
rect 35946 6611 35982 6645
rect 36016 6611 36032 6645
rect 34980 6347 35010 6378
rect 35553 6523 35583 6584
rect 35647 6562 35677 6597
rect 35946 6595 36032 6611
rect 36204 6659 36270 6675
rect 36204 6625 36220 6659
rect 36254 6625 36270 6659
rect 36204 6609 36270 6625
rect 35946 6563 35976 6595
rect 36222 6578 36252 6609
rect 35641 6538 35677 6562
rect 35641 6523 35671 6538
rect 34962 6331 35028 6347
rect 35254 6345 35284 6371
rect 35553 6339 35583 6365
rect 35641 6339 35671 6365
rect 37441 6815 37471 6841
rect 37529 6815 37559 6841
rect 37834 6813 37864 6839
rect 38406 6838 38472 6866
rect 40294 6900 40360 6916
rect 40408 6912 40438 6938
rect 42200 6916 42230 6938
rect 40294 6866 40310 6900
rect 40344 6866 40360 6900
rect 38406 6819 38584 6838
rect 39030 6821 39060 6847
rect 36850 6659 36916 6675
rect 36850 6625 36866 6659
rect 36900 6625 36916 6659
rect 36850 6609 36916 6625
rect 37142 6669 37172 6691
rect 37142 6653 37228 6669
rect 37142 6619 37178 6653
rect 37212 6619 37228 6653
rect 37441 6650 37471 6711
rect 37529 6696 37559 6711
rect 37529 6672 37565 6696
rect 38406 6806 38534 6819
rect 38518 6785 38534 6806
rect 38568 6785 38584 6819
rect 38518 6769 38584 6785
rect 38440 6738 38470 6764
rect 38536 6738 38566 6769
rect 37535 6663 37565 6672
rect 36868 6578 36898 6609
rect 37142 6603 37228 6619
rect 37439 6634 37493 6650
rect 36552 6507 36582 6538
rect 36534 6491 36600 6507
rect 36534 6457 36550 6491
rect 36584 6457 36600 6491
rect 36534 6441 36600 6457
rect 36648 6454 36678 6538
rect 36648 6424 36734 6454
rect 35946 6337 35976 6363
rect 36222 6348 36252 6378
rect 36222 6347 36284 6348
rect 34962 6297 34978 6331
rect 35012 6297 35028 6331
rect 34962 6281 35028 6297
rect 36204 6331 36284 6347
rect 36204 6297 36220 6331
rect 36254 6297 36284 6331
rect 36204 6281 36284 6297
rect 34364 6236 34846 6266
rect 36252 6266 36284 6281
rect 36704 6266 36734 6424
rect 37142 6571 37172 6603
rect 37439 6600 37449 6634
rect 37483 6600 37493 6634
rect 37439 6584 37493 6600
rect 37535 6647 37611 6663
rect 37535 6613 37567 6647
rect 37601 6613 37611 6647
rect 37535 6597 37611 6613
rect 37834 6661 37864 6683
rect 37834 6645 37920 6661
rect 37834 6611 37870 6645
rect 37904 6611 37920 6645
rect 36868 6347 36898 6378
rect 37441 6523 37471 6584
rect 37535 6562 37565 6597
rect 37834 6595 37920 6611
rect 38092 6659 38158 6675
rect 38092 6625 38108 6659
rect 38142 6625 38158 6659
rect 38092 6609 38158 6625
rect 37834 6563 37864 6595
rect 38110 6578 38140 6609
rect 37529 6538 37565 6562
rect 37529 6523 37559 6538
rect 36850 6331 36916 6347
rect 37142 6345 37172 6371
rect 37441 6339 37471 6365
rect 37529 6339 37559 6365
rect 39329 6815 39359 6841
rect 39417 6815 39447 6841
rect 39722 6813 39752 6839
rect 40294 6838 40360 6866
rect 42182 6900 42248 6916
rect 42296 6912 42326 6938
rect 44088 6916 44118 6938
rect 42182 6866 42198 6900
rect 42232 6866 42248 6900
rect 40294 6819 40472 6838
rect 40918 6821 40948 6847
rect 38738 6659 38804 6675
rect 38738 6625 38754 6659
rect 38788 6625 38804 6659
rect 38738 6609 38804 6625
rect 39030 6669 39060 6691
rect 39030 6653 39116 6669
rect 39030 6619 39066 6653
rect 39100 6619 39116 6653
rect 39329 6650 39359 6711
rect 39417 6696 39447 6711
rect 39417 6672 39453 6696
rect 40294 6806 40422 6819
rect 40406 6785 40422 6806
rect 40456 6785 40472 6819
rect 40406 6769 40472 6785
rect 40328 6738 40358 6764
rect 40424 6738 40454 6769
rect 39423 6663 39453 6672
rect 38756 6578 38786 6609
rect 39030 6603 39116 6619
rect 39327 6634 39381 6650
rect 38440 6507 38470 6538
rect 38422 6491 38488 6507
rect 38422 6457 38438 6491
rect 38472 6457 38488 6491
rect 38422 6441 38488 6457
rect 38536 6454 38566 6538
rect 38536 6424 38622 6454
rect 37834 6337 37864 6363
rect 38110 6348 38140 6378
rect 38110 6347 38172 6348
rect 36850 6297 36866 6331
rect 36900 6297 36916 6331
rect 36850 6281 36916 6297
rect 38092 6331 38172 6347
rect 38092 6297 38108 6331
rect 38142 6297 38172 6331
rect 38092 6281 38172 6297
rect 36252 6236 36734 6266
rect 38140 6266 38172 6281
rect 38592 6266 38622 6424
rect 39030 6571 39060 6603
rect 39327 6600 39337 6634
rect 39371 6600 39381 6634
rect 39327 6584 39381 6600
rect 39423 6647 39499 6663
rect 39423 6613 39455 6647
rect 39489 6613 39499 6647
rect 39423 6597 39499 6613
rect 39722 6661 39752 6683
rect 39722 6645 39808 6661
rect 39722 6611 39758 6645
rect 39792 6611 39808 6645
rect 38756 6347 38786 6378
rect 39329 6523 39359 6584
rect 39423 6562 39453 6597
rect 39722 6595 39808 6611
rect 39980 6659 40046 6675
rect 39980 6625 39996 6659
rect 40030 6625 40046 6659
rect 39980 6609 40046 6625
rect 39722 6563 39752 6595
rect 39998 6578 40028 6609
rect 39417 6538 39453 6562
rect 39417 6523 39447 6538
rect 38738 6331 38804 6347
rect 39030 6345 39060 6371
rect 39329 6339 39359 6365
rect 39417 6339 39447 6365
rect 41217 6815 41247 6841
rect 41305 6815 41335 6841
rect 41610 6813 41640 6839
rect 42182 6838 42248 6866
rect 44070 6900 44136 6916
rect 44184 6912 44214 6938
rect 45970 6916 46000 6938
rect 44070 6866 44086 6900
rect 44120 6866 44136 6900
rect 42182 6819 42360 6838
rect 42806 6821 42836 6847
rect 40626 6659 40692 6675
rect 40626 6625 40642 6659
rect 40676 6625 40692 6659
rect 40626 6609 40692 6625
rect 40918 6669 40948 6691
rect 40918 6653 41004 6669
rect 40918 6619 40954 6653
rect 40988 6619 41004 6653
rect 41217 6650 41247 6711
rect 41305 6696 41335 6711
rect 41305 6672 41341 6696
rect 42182 6806 42310 6819
rect 42294 6785 42310 6806
rect 42344 6785 42360 6819
rect 42294 6769 42360 6785
rect 42216 6738 42246 6764
rect 42312 6738 42342 6769
rect 41311 6663 41341 6672
rect 40644 6578 40674 6609
rect 40918 6603 41004 6619
rect 41215 6634 41269 6650
rect 40328 6507 40358 6538
rect 40310 6491 40376 6507
rect 40310 6457 40326 6491
rect 40360 6457 40376 6491
rect 40310 6441 40376 6457
rect 40424 6454 40454 6538
rect 40424 6424 40510 6454
rect 39722 6337 39752 6363
rect 39998 6348 40028 6378
rect 39998 6347 40060 6348
rect 38738 6297 38754 6331
rect 38788 6297 38804 6331
rect 38738 6281 38804 6297
rect 39980 6331 40060 6347
rect 39980 6297 39996 6331
rect 40030 6297 40060 6331
rect 39980 6281 40060 6297
rect 38140 6236 38622 6266
rect 40028 6266 40060 6281
rect 40480 6266 40510 6424
rect 40918 6571 40948 6603
rect 41215 6600 41225 6634
rect 41259 6600 41269 6634
rect 41215 6584 41269 6600
rect 41311 6647 41387 6663
rect 41311 6613 41343 6647
rect 41377 6613 41387 6647
rect 41311 6597 41387 6613
rect 41610 6661 41640 6683
rect 41610 6645 41696 6661
rect 41610 6611 41646 6645
rect 41680 6611 41696 6645
rect 40644 6347 40674 6378
rect 41217 6523 41247 6584
rect 41311 6562 41341 6597
rect 41610 6595 41696 6611
rect 41868 6659 41934 6675
rect 41868 6625 41884 6659
rect 41918 6625 41934 6659
rect 41868 6609 41934 6625
rect 41610 6563 41640 6595
rect 41886 6578 41916 6609
rect 41305 6538 41341 6562
rect 41305 6523 41335 6538
rect 40626 6331 40692 6347
rect 40918 6345 40948 6371
rect 41217 6339 41247 6365
rect 41305 6339 41335 6365
rect 43105 6815 43135 6841
rect 43193 6815 43223 6841
rect 43498 6813 43528 6839
rect 44070 6838 44136 6866
rect 45952 6900 46018 6916
rect 46066 6912 46096 6938
rect 47858 6916 47888 6938
rect 45952 6866 45968 6900
rect 46002 6866 46018 6900
rect 44070 6819 44248 6838
rect 44694 6821 44724 6847
rect 42514 6659 42580 6675
rect 42514 6625 42530 6659
rect 42564 6625 42580 6659
rect 42514 6609 42580 6625
rect 42806 6669 42836 6691
rect 42806 6653 42892 6669
rect 42806 6619 42842 6653
rect 42876 6619 42892 6653
rect 43105 6650 43135 6711
rect 43193 6696 43223 6711
rect 43193 6672 43229 6696
rect 44070 6806 44198 6819
rect 44182 6785 44198 6806
rect 44232 6785 44248 6819
rect 44182 6769 44248 6785
rect 44104 6738 44134 6764
rect 44200 6738 44230 6769
rect 43199 6663 43229 6672
rect 42532 6578 42562 6609
rect 42806 6603 42892 6619
rect 43103 6634 43157 6650
rect 42216 6507 42246 6538
rect 42198 6491 42264 6507
rect 42198 6457 42214 6491
rect 42248 6457 42264 6491
rect 42198 6441 42264 6457
rect 42312 6454 42342 6538
rect 42312 6424 42398 6454
rect 41610 6337 41640 6363
rect 41886 6348 41916 6378
rect 41886 6347 41948 6348
rect 40626 6297 40642 6331
rect 40676 6297 40692 6331
rect 40626 6281 40692 6297
rect 41868 6331 41948 6347
rect 41868 6297 41884 6331
rect 41918 6297 41948 6331
rect 41868 6281 41948 6297
rect 40028 6236 40510 6266
rect 41916 6266 41948 6281
rect 42368 6266 42398 6424
rect 42806 6571 42836 6603
rect 43103 6600 43113 6634
rect 43147 6600 43157 6634
rect 43103 6584 43157 6600
rect 43199 6647 43275 6663
rect 43199 6613 43231 6647
rect 43265 6613 43275 6647
rect 43199 6597 43275 6613
rect 43498 6661 43528 6683
rect 43498 6645 43584 6661
rect 43498 6611 43534 6645
rect 43568 6611 43584 6645
rect 42532 6347 42562 6378
rect 43105 6523 43135 6584
rect 43199 6562 43229 6597
rect 43498 6595 43584 6611
rect 43756 6659 43822 6675
rect 43756 6625 43772 6659
rect 43806 6625 43822 6659
rect 43756 6609 43822 6625
rect 43498 6563 43528 6595
rect 43774 6578 43804 6609
rect 43193 6538 43229 6562
rect 43193 6523 43223 6538
rect 42514 6331 42580 6347
rect 42806 6345 42836 6371
rect 43105 6339 43135 6365
rect 43193 6339 43223 6365
rect 44987 6815 45017 6841
rect 45075 6815 45105 6841
rect 45380 6813 45410 6839
rect 45952 6838 46018 6866
rect 47840 6900 47906 6916
rect 47954 6912 47984 6938
rect 49746 6916 49776 6938
rect 47840 6866 47856 6900
rect 47890 6866 47906 6900
rect 45952 6819 46130 6838
rect 46576 6821 46606 6847
rect 44402 6659 44468 6675
rect 44402 6625 44418 6659
rect 44452 6625 44468 6659
rect 44402 6609 44468 6625
rect 44694 6669 44724 6691
rect 44694 6653 44780 6669
rect 44694 6619 44730 6653
rect 44764 6619 44780 6653
rect 44987 6650 45017 6711
rect 45075 6696 45105 6711
rect 45075 6672 45111 6696
rect 45952 6806 46080 6819
rect 46064 6785 46080 6806
rect 46114 6785 46130 6819
rect 46064 6769 46130 6785
rect 45986 6738 46016 6764
rect 46082 6738 46112 6769
rect 45081 6663 45111 6672
rect 44420 6578 44450 6609
rect 44694 6603 44780 6619
rect 44985 6634 45039 6650
rect 44104 6507 44134 6538
rect 44086 6491 44152 6507
rect 44086 6457 44102 6491
rect 44136 6457 44152 6491
rect 44086 6441 44152 6457
rect 44200 6454 44230 6538
rect 44200 6424 44286 6454
rect 43498 6337 43528 6363
rect 43774 6348 43804 6378
rect 43774 6347 43836 6348
rect 42514 6297 42530 6331
rect 42564 6297 42580 6331
rect 42514 6281 42580 6297
rect 43756 6331 43836 6347
rect 43756 6297 43772 6331
rect 43806 6297 43836 6331
rect 43756 6281 43836 6297
rect 41916 6236 42398 6266
rect 43804 6266 43836 6281
rect 44256 6266 44286 6424
rect 44694 6571 44724 6603
rect 44985 6600 44995 6634
rect 45029 6600 45039 6634
rect 44985 6584 45039 6600
rect 45081 6647 45157 6663
rect 45081 6613 45113 6647
rect 45147 6613 45157 6647
rect 45081 6597 45157 6613
rect 45380 6661 45410 6683
rect 45380 6645 45466 6661
rect 45380 6611 45416 6645
rect 45450 6611 45466 6645
rect 44420 6347 44450 6378
rect 44987 6523 45017 6584
rect 45081 6562 45111 6597
rect 45380 6595 45466 6611
rect 45638 6659 45704 6675
rect 45638 6625 45654 6659
rect 45688 6625 45704 6659
rect 45638 6609 45704 6625
rect 45380 6563 45410 6595
rect 45656 6578 45686 6609
rect 45075 6538 45111 6562
rect 45075 6523 45105 6538
rect 44402 6331 44468 6347
rect 44694 6345 44724 6371
rect 44987 6339 45017 6365
rect 45075 6339 45105 6365
rect 46875 6815 46905 6841
rect 46963 6815 46993 6841
rect 47268 6813 47298 6839
rect 47840 6838 47906 6866
rect 49728 6900 49794 6916
rect 49842 6912 49872 6938
rect 51634 6916 51664 6938
rect 49728 6866 49744 6900
rect 49778 6866 49794 6900
rect 47840 6819 48018 6838
rect 48464 6821 48494 6847
rect 46284 6659 46350 6675
rect 46284 6625 46300 6659
rect 46334 6625 46350 6659
rect 46284 6609 46350 6625
rect 46576 6669 46606 6691
rect 46576 6653 46662 6669
rect 46576 6619 46612 6653
rect 46646 6619 46662 6653
rect 46875 6650 46905 6711
rect 46963 6696 46993 6711
rect 46963 6672 46999 6696
rect 47840 6806 47968 6819
rect 47952 6785 47968 6806
rect 48002 6785 48018 6819
rect 47952 6769 48018 6785
rect 47874 6738 47904 6764
rect 47970 6738 48000 6769
rect 46969 6663 46999 6672
rect 46302 6578 46332 6609
rect 46576 6603 46662 6619
rect 46873 6634 46927 6650
rect 45986 6507 46016 6538
rect 45968 6491 46034 6507
rect 45968 6457 45984 6491
rect 46018 6457 46034 6491
rect 45968 6441 46034 6457
rect 46082 6454 46112 6538
rect 46082 6424 46168 6454
rect 45380 6337 45410 6363
rect 45656 6348 45686 6378
rect 45656 6347 45718 6348
rect 44402 6297 44418 6331
rect 44452 6297 44468 6331
rect 44402 6281 44468 6297
rect 45638 6331 45718 6347
rect 45638 6297 45654 6331
rect 45688 6297 45718 6331
rect 45638 6281 45718 6297
rect 43804 6236 44286 6266
rect 45686 6266 45718 6281
rect 46138 6266 46168 6424
rect 46576 6571 46606 6603
rect 46873 6600 46883 6634
rect 46917 6600 46927 6634
rect 46873 6584 46927 6600
rect 46969 6647 47045 6663
rect 46969 6613 47001 6647
rect 47035 6613 47045 6647
rect 46969 6597 47045 6613
rect 47268 6661 47298 6683
rect 47268 6645 47354 6661
rect 47268 6611 47304 6645
rect 47338 6611 47354 6645
rect 46302 6347 46332 6378
rect 46875 6523 46905 6584
rect 46969 6562 46999 6597
rect 47268 6595 47354 6611
rect 47526 6659 47592 6675
rect 47526 6625 47542 6659
rect 47576 6625 47592 6659
rect 47526 6609 47592 6625
rect 47268 6563 47298 6595
rect 47544 6578 47574 6609
rect 46963 6538 46999 6562
rect 46963 6523 46993 6538
rect 46284 6331 46350 6347
rect 46576 6345 46606 6371
rect 46875 6339 46905 6365
rect 46963 6339 46993 6365
rect 48763 6815 48793 6841
rect 48851 6815 48881 6841
rect 49156 6813 49186 6839
rect 49728 6838 49794 6866
rect 51616 6900 51682 6916
rect 51730 6912 51760 6938
rect 53522 6916 53552 6938
rect 51616 6866 51632 6900
rect 51666 6866 51682 6900
rect 49728 6819 49906 6838
rect 50352 6821 50382 6847
rect 48172 6659 48238 6675
rect 48172 6625 48188 6659
rect 48222 6625 48238 6659
rect 48172 6609 48238 6625
rect 48464 6669 48494 6691
rect 48464 6653 48550 6669
rect 48464 6619 48500 6653
rect 48534 6619 48550 6653
rect 48763 6650 48793 6711
rect 48851 6696 48881 6711
rect 48851 6672 48887 6696
rect 49728 6806 49856 6819
rect 49840 6785 49856 6806
rect 49890 6785 49906 6819
rect 49840 6769 49906 6785
rect 49762 6738 49792 6764
rect 49858 6738 49888 6769
rect 48857 6663 48887 6672
rect 48190 6578 48220 6609
rect 48464 6603 48550 6619
rect 48761 6634 48815 6650
rect 47874 6507 47904 6538
rect 47856 6491 47922 6507
rect 47856 6457 47872 6491
rect 47906 6457 47922 6491
rect 47856 6441 47922 6457
rect 47970 6454 48000 6538
rect 47970 6424 48056 6454
rect 47268 6337 47298 6363
rect 47544 6348 47574 6378
rect 47544 6347 47606 6348
rect 46284 6297 46300 6331
rect 46334 6297 46350 6331
rect 46284 6281 46350 6297
rect 47526 6331 47606 6347
rect 47526 6297 47542 6331
rect 47576 6297 47606 6331
rect 47526 6281 47606 6297
rect 45686 6236 46168 6266
rect 47574 6266 47606 6281
rect 48026 6266 48056 6424
rect 48464 6571 48494 6603
rect 48761 6600 48771 6634
rect 48805 6600 48815 6634
rect 48761 6584 48815 6600
rect 48857 6647 48933 6663
rect 48857 6613 48889 6647
rect 48923 6613 48933 6647
rect 48857 6597 48933 6613
rect 49156 6661 49186 6683
rect 49156 6645 49242 6661
rect 49156 6611 49192 6645
rect 49226 6611 49242 6645
rect 48190 6347 48220 6378
rect 48763 6523 48793 6584
rect 48857 6562 48887 6597
rect 49156 6595 49242 6611
rect 49414 6659 49480 6675
rect 49414 6625 49430 6659
rect 49464 6625 49480 6659
rect 49414 6609 49480 6625
rect 49156 6563 49186 6595
rect 49432 6578 49462 6609
rect 48851 6538 48887 6562
rect 48851 6523 48881 6538
rect 48172 6331 48238 6347
rect 48464 6345 48494 6371
rect 48763 6339 48793 6365
rect 48851 6339 48881 6365
rect 50651 6815 50681 6841
rect 50739 6815 50769 6841
rect 51044 6813 51074 6839
rect 51616 6838 51682 6866
rect 53504 6900 53570 6916
rect 53618 6912 53648 6938
rect 55410 6916 55440 6938
rect 53504 6866 53520 6900
rect 53554 6866 53570 6900
rect 51616 6819 51794 6838
rect 52240 6821 52270 6847
rect 50060 6659 50126 6675
rect 50060 6625 50076 6659
rect 50110 6625 50126 6659
rect 50060 6609 50126 6625
rect 50352 6669 50382 6691
rect 50352 6653 50438 6669
rect 50352 6619 50388 6653
rect 50422 6619 50438 6653
rect 50651 6650 50681 6711
rect 50739 6696 50769 6711
rect 50739 6672 50775 6696
rect 51616 6806 51744 6819
rect 51728 6785 51744 6806
rect 51778 6785 51794 6819
rect 51728 6769 51794 6785
rect 51650 6738 51680 6764
rect 51746 6738 51776 6769
rect 50745 6663 50775 6672
rect 50078 6578 50108 6609
rect 50352 6603 50438 6619
rect 50649 6634 50703 6650
rect 49762 6507 49792 6538
rect 49744 6491 49810 6507
rect 49744 6457 49760 6491
rect 49794 6457 49810 6491
rect 49744 6441 49810 6457
rect 49858 6454 49888 6538
rect 49858 6424 49944 6454
rect 49156 6337 49186 6363
rect 49432 6348 49462 6378
rect 49432 6347 49494 6348
rect 48172 6297 48188 6331
rect 48222 6297 48238 6331
rect 48172 6281 48238 6297
rect 49414 6331 49494 6347
rect 49414 6297 49430 6331
rect 49464 6297 49494 6331
rect 49414 6281 49494 6297
rect 47574 6236 48056 6266
rect 49462 6266 49494 6281
rect 49914 6266 49944 6424
rect 50352 6571 50382 6603
rect 50649 6600 50659 6634
rect 50693 6600 50703 6634
rect 50649 6584 50703 6600
rect 50745 6647 50821 6663
rect 50745 6613 50777 6647
rect 50811 6613 50821 6647
rect 50745 6597 50821 6613
rect 51044 6661 51074 6683
rect 51044 6645 51130 6661
rect 51044 6611 51080 6645
rect 51114 6611 51130 6645
rect 50078 6347 50108 6378
rect 50651 6523 50681 6584
rect 50745 6562 50775 6597
rect 51044 6595 51130 6611
rect 51302 6659 51368 6675
rect 51302 6625 51318 6659
rect 51352 6625 51368 6659
rect 51302 6609 51368 6625
rect 51044 6563 51074 6595
rect 51320 6578 51350 6609
rect 50739 6538 50775 6562
rect 50739 6523 50769 6538
rect 50060 6331 50126 6347
rect 50352 6345 50382 6371
rect 50651 6339 50681 6365
rect 50739 6339 50769 6365
rect 52539 6815 52569 6841
rect 52627 6815 52657 6841
rect 52932 6813 52962 6839
rect 53504 6838 53570 6866
rect 55392 6900 55458 6916
rect 55506 6912 55536 6938
rect 57298 6916 57328 6938
rect 55392 6866 55408 6900
rect 55442 6866 55458 6900
rect 53504 6819 53682 6838
rect 54128 6821 54158 6847
rect 51948 6659 52014 6675
rect 51948 6625 51964 6659
rect 51998 6625 52014 6659
rect 51948 6609 52014 6625
rect 52240 6669 52270 6691
rect 52240 6653 52326 6669
rect 52240 6619 52276 6653
rect 52310 6619 52326 6653
rect 52539 6650 52569 6711
rect 52627 6696 52657 6711
rect 52627 6672 52663 6696
rect 53504 6806 53632 6819
rect 53616 6785 53632 6806
rect 53666 6785 53682 6819
rect 53616 6769 53682 6785
rect 53538 6738 53568 6764
rect 53634 6738 53664 6769
rect 52633 6663 52663 6672
rect 51966 6578 51996 6609
rect 52240 6603 52326 6619
rect 52537 6634 52591 6650
rect 51650 6507 51680 6538
rect 51632 6491 51698 6507
rect 51632 6457 51648 6491
rect 51682 6457 51698 6491
rect 51632 6441 51698 6457
rect 51746 6454 51776 6538
rect 51746 6424 51832 6454
rect 51044 6337 51074 6363
rect 51320 6348 51350 6378
rect 51320 6347 51382 6348
rect 50060 6297 50076 6331
rect 50110 6297 50126 6331
rect 50060 6281 50126 6297
rect 51302 6331 51382 6347
rect 51302 6297 51318 6331
rect 51352 6297 51382 6331
rect 51302 6281 51382 6297
rect 49462 6236 49944 6266
rect 51350 6266 51382 6281
rect 51802 6266 51832 6424
rect 52240 6571 52270 6603
rect 52537 6600 52547 6634
rect 52581 6600 52591 6634
rect 52537 6584 52591 6600
rect 52633 6647 52709 6663
rect 52633 6613 52665 6647
rect 52699 6613 52709 6647
rect 52633 6597 52709 6613
rect 52932 6661 52962 6683
rect 52932 6645 53018 6661
rect 52932 6611 52968 6645
rect 53002 6611 53018 6645
rect 51966 6347 51996 6378
rect 52539 6523 52569 6584
rect 52633 6562 52663 6597
rect 52932 6595 53018 6611
rect 53190 6659 53256 6675
rect 53190 6625 53206 6659
rect 53240 6625 53256 6659
rect 53190 6609 53256 6625
rect 52932 6563 52962 6595
rect 53208 6578 53238 6609
rect 52627 6538 52663 6562
rect 52627 6523 52657 6538
rect 51948 6331 52014 6347
rect 52240 6345 52270 6371
rect 52539 6339 52569 6365
rect 52627 6339 52657 6365
rect 54427 6815 54457 6841
rect 54515 6815 54545 6841
rect 54820 6813 54850 6839
rect 55392 6838 55458 6866
rect 57280 6900 57346 6916
rect 57394 6912 57424 6938
rect 59186 6916 59216 6938
rect 57280 6866 57296 6900
rect 57330 6866 57346 6900
rect 55392 6819 55570 6838
rect 56016 6821 56046 6847
rect 53836 6659 53902 6675
rect 53836 6625 53852 6659
rect 53886 6625 53902 6659
rect 53836 6609 53902 6625
rect 54128 6669 54158 6691
rect 54128 6653 54214 6669
rect 54128 6619 54164 6653
rect 54198 6619 54214 6653
rect 54427 6650 54457 6711
rect 54515 6696 54545 6711
rect 54515 6672 54551 6696
rect 55392 6806 55520 6819
rect 55504 6785 55520 6806
rect 55554 6785 55570 6819
rect 55504 6769 55570 6785
rect 55426 6738 55456 6764
rect 55522 6738 55552 6769
rect 54521 6663 54551 6672
rect 53854 6578 53884 6609
rect 54128 6603 54214 6619
rect 54425 6634 54479 6650
rect 53538 6507 53568 6538
rect 53520 6491 53586 6507
rect 53520 6457 53536 6491
rect 53570 6457 53586 6491
rect 53520 6441 53586 6457
rect 53634 6454 53664 6538
rect 53634 6424 53720 6454
rect 52932 6337 52962 6363
rect 53208 6348 53238 6378
rect 53208 6347 53270 6348
rect 51948 6297 51964 6331
rect 51998 6297 52014 6331
rect 51948 6281 52014 6297
rect 53190 6331 53270 6347
rect 53190 6297 53206 6331
rect 53240 6297 53270 6331
rect 53190 6281 53270 6297
rect 51350 6236 51832 6266
rect 53238 6266 53270 6281
rect 53690 6266 53720 6424
rect 54128 6571 54158 6603
rect 54425 6600 54435 6634
rect 54469 6600 54479 6634
rect 54425 6584 54479 6600
rect 54521 6647 54597 6663
rect 54521 6613 54553 6647
rect 54587 6613 54597 6647
rect 54521 6597 54597 6613
rect 54820 6661 54850 6683
rect 54820 6645 54906 6661
rect 54820 6611 54856 6645
rect 54890 6611 54906 6645
rect 53854 6347 53884 6378
rect 54427 6523 54457 6584
rect 54521 6562 54551 6597
rect 54820 6595 54906 6611
rect 55078 6659 55144 6675
rect 55078 6625 55094 6659
rect 55128 6625 55144 6659
rect 55078 6609 55144 6625
rect 54820 6563 54850 6595
rect 55096 6578 55126 6609
rect 54515 6538 54551 6562
rect 54515 6523 54545 6538
rect 53836 6331 53902 6347
rect 54128 6345 54158 6371
rect 54427 6339 54457 6365
rect 54515 6339 54545 6365
rect 56315 6815 56345 6841
rect 56403 6815 56433 6841
rect 56708 6813 56738 6839
rect 57280 6838 57346 6866
rect 59168 6900 59234 6916
rect 59282 6912 59312 6938
rect 59168 6866 59184 6900
rect 59218 6866 59234 6900
rect 57280 6819 57458 6838
rect 57904 6821 57934 6847
rect 55724 6659 55790 6675
rect 55724 6625 55740 6659
rect 55774 6625 55790 6659
rect 55724 6609 55790 6625
rect 56016 6669 56046 6691
rect 56016 6653 56102 6669
rect 56016 6619 56052 6653
rect 56086 6619 56102 6653
rect 56315 6650 56345 6711
rect 56403 6696 56433 6711
rect 56403 6672 56439 6696
rect 57280 6806 57408 6819
rect 57392 6785 57408 6806
rect 57442 6785 57458 6819
rect 57392 6769 57458 6785
rect 57314 6738 57344 6764
rect 57410 6738 57440 6769
rect 56409 6663 56439 6672
rect 55742 6578 55772 6609
rect 56016 6603 56102 6619
rect 56313 6634 56367 6650
rect 55426 6507 55456 6538
rect 55408 6491 55474 6507
rect 55408 6457 55424 6491
rect 55458 6457 55474 6491
rect 55408 6441 55474 6457
rect 55522 6454 55552 6538
rect 55522 6424 55608 6454
rect 54820 6337 54850 6363
rect 55096 6348 55126 6378
rect 55096 6347 55158 6348
rect 53836 6297 53852 6331
rect 53886 6297 53902 6331
rect 53836 6281 53902 6297
rect 55078 6331 55158 6347
rect 55078 6297 55094 6331
rect 55128 6297 55158 6331
rect 55078 6281 55158 6297
rect 53238 6236 53720 6266
rect 55126 6266 55158 6281
rect 55578 6266 55608 6424
rect 56016 6571 56046 6603
rect 56313 6600 56323 6634
rect 56357 6600 56367 6634
rect 56313 6584 56367 6600
rect 56409 6647 56485 6663
rect 56409 6613 56441 6647
rect 56475 6613 56485 6647
rect 56409 6597 56485 6613
rect 56708 6661 56738 6683
rect 56708 6645 56794 6661
rect 56708 6611 56744 6645
rect 56778 6611 56794 6645
rect 55742 6347 55772 6378
rect 56315 6523 56345 6584
rect 56409 6562 56439 6597
rect 56708 6595 56794 6611
rect 56966 6659 57032 6675
rect 56966 6625 56982 6659
rect 57016 6625 57032 6659
rect 56966 6609 57032 6625
rect 56708 6563 56738 6595
rect 56984 6578 57014 6609
rect 56403 6538 56439 6562
rect 56403 6523 56433 6538
rect 55724 6331 55790 6347
rect 56016 6345 56046 6371
rect 56315 6339 56345 6365
rect 56403 6339 56433 6365
rect 58203 6815 58233 6841
rect 58291 6815 58321 6841
rect 58596 6813 58626 6839
rect 59168 6838 59234 6866
rect 59168 6819 59346 6838
rect 59792 6821 59822 6847
rect 57612 6659 57678 6675
rect 57612 6625 57628 6659
rect 57662 6625 57678 6659
rect 57612 6609 57678 6625
rect 57904 6669 57934 6691
rect 57904 6653 57990 6669
rect 57904 6619 57940 6653
rect 57974 6619 57990 6653
rect 58203 6650 58233 6711
rect 58291 6696 58321 6711
rect 58291 6672 58327 6696
rect 59168 6806 59296 6819
rect 59280 6785 59296 6806
rect 59330 6785 59346 6819
rect 59280 6769 59346 6785
rect 59202 6738 59232 6764
rect 59298 6738 59328 6769
rect 58297 6663 58327 6672
rect 57630 6578 57660 6609
rect 57904 6603 57990 6619
rect 58201 6634 58255 6650
rect 57314 6507 57344 6538
rect 57296 6491 57362 6507
rect 57296 6457 57312 6491
rect 57346 6457 57362 6491
rect 57296 6441 57362 6457
rect 57410 6454 57440 6538
rect 57410 6424 57496 6454
rect 56708 6337 56738 6363
rect 56984 6348 57014 6378
rect 56984 6347 57046 6348
rect 55724 6297 55740 6331
rect 55774 6297 55790 6331
rect 55724 6281 55790 6297
rect 56966 6331 57046 6347
rect 56966 6297 56982 6331
rect 57016 6297 57046 6331
rect 56966 6281 57046 6297
rect 55126 6236 55608 6266
rect 57014 6266 57046 6281
rect 57466 6266 57496 6424
rect 57904 6571 57934 6603
rect 58201 6600 58211 6634
rect 58245 6600 58255 6634
rect 58201 6584 58255 6600
rect 58297 6647 58373 6663
rect 58297 6613 58329 6647
rect 58363 6613 58373 6647
rect 58297 6597 58373 6613
rect 58596 6661 58626 6683
rect 58596 6645 58682 6661
rect 58596 6611 58632 6645
rect 58666 6611 58682 6645
rect 57630 6347 57660 6378
rect 58203 6523 58233 6584
rect 58297 6562 58327 6597
rect 58596 6595 58682 6611
rect 58854 6659 58920 6675
rect 58854 6625 58870 6659
rect 58904 6625 58920 6659
rect 58854 6609 58920 6625
rect 58596 6563 58626 6595
rect 58872 6578 58902 6609
rect 58291 6538 58327 6562
rect 58291 6523 58321 6538
rect 57612 6331 57678 6347
rect 57904 6345 57934 6371
rect 58203 6339 58233 6365
rect 58291 6339 58321 6365
rect 59500 6659 59566 6675
rect 59500 6625 59516 6659
rect 59550 6625 59566 6659
rect 59500 6609 59566 6625
rect 59792 6669 59822 6691
rect 59792 6653 59878 6669
rect 59792 6619 59828 6653
rect 59862 6619 59878 6653
rect 59518 6578 59548 6609
rect 59792 6603 59878 6619
rect 59202 6507 59232 6538
rect 59184 6491 59250 6507
rect 59184 6457 59200 6491
rect 59234 6457 59250 6491
rect 59184 6441 59250 6457
rect 59298 6454 59328 6538
rect 59298 6424 59384 6454
rect 58596 6337 58626 6363
rect 58872 6348 58902 6378
rect 58872 6347 58934 6348
rect 57612 6297 57628 6331
rect 57662 6297 57678 6331
rect 57612 6281 57678 6297
rect 58854 6331 58934 6347
rect 58854 6297 58870 6331
rect 58904 6297 58934 6331
rect 58854 6281 58934 6297
rect 57014 6236 57496 6266
rect 58902 6266 58934 6281
rect 59354 6266 59384 6424
rect 59792 6571 59822 6603
rect 59518 6347 59548 6378
rect 59500 6331 59566 6347
rect 59792 6345 59822 6371
rect 59500 6297 59516 6331
rect 59550 6297 59566 6331
rect 59500 6281 59566 6297
rect 58902 6236 59384 6266
rect 564 6068 594 6236
rect 746 6084 812 6100
rect 564 6038 698 6068
rect 668 6012 698 6038
rect 746 6050 762 6084
rect 796 6050 812 6084
rect 746 6034 812 6050
rect 2452 6068 2482 6236
rect 2634 6084 2700 6100
rect 2452 6038 2586 6068
rect 764 6012 794 6034
rect 2556 6012 2586 6038
rect 2634 6050 2650 6084
rect 2684 6050 2700 6084
rect 2634 6034 2700 6050
rect 4340 6068 4370 6236
rect 4522 6084 4588 6100
rect 4340 6038 4474 6068
rect 2652 6012 2682 6034
rect 4444 6012 4474 6038
rect 4522 6050 4538 6084
rect 4572 6050 4588 6084
rect 4522 6034 4588 6050
rect 6228 6068 6258 6236
rect 6410 6084 6476 6100
rect 6228 6038 6362 6068
rect 4540 6012 4570 6034
rect 6332 6012 6362 6038
rect 6410 6050 6426 6084
rect 6460 6050 6476 6084
rect 6410 6034 6476 6050
rect 8116 6068 8146 6236
rect 8298 6084 8364 6100
rect 8116 6038 8250 6068
rect 6428 6012 6458 6034
rect 8220 6012 8250 6038
rect 8298 6050 8314 6084
rect 8348 6050 8364 6084
rect 8298 6034 8364 6050
rect 10004 6068 10034 6236
rect 10186 6084 10252 6100
rect 10004 6038 10138 6068
rect 8316 6012 8346 6034
rect 10108 6012 10138 6038
rect 10186 6050 10202 6084
rect 10236 6050 10252 6084
rect 10186 6034 10252 6050
rect 11892 6068 11922 6236
rect 12074 6084 12140 6100
rect 11892 6038 12026 6068
rect 10204 6012 10234 6034
rect 11996 6012 12026 6038
rect 12074 6050 12090 6084
rect 12124 6050 12140 6084
rect 12074 6034 12140 6050
rect 13780 6068 13810 6236
rect 13962 6084 14028 6100
rect 13780 6038 13914 6068
rect 12092 6012 12122 6034
rect 13884 6012 13914 6038
rect 13962 6050 13978 6084
rect 14012 6050 14028 6084
rect 13962 6034 14028 6050
rect 15662 6068 15692 6236
rect 15844 6084 15910 6100
rect 15662 6038 15796 6068
rect 13980 6012 14010 6034
rect 15766 6012 15796 6038
rect 15844 6050 15860 6084
rect 15894 6050 15910 6084
rect 15844 6034 15910 6050
rect 17550 6068 17580 6236
rect 17732 6084 17798 6100
rect 17550 6038 17684 6068
rect 15862 6012 15892 6034
rect 17654 6012 17684 6038
rect 17732 6050 17748 6084
rect 17782 6050 17798 6084
rect 17732 6034 17798 6050
rect 19438 6068 19468 6236
rect 19620 6084 19686 6100
rect 19438 6038 19572 6068
rect 17750 6012 17780 6034
rect 19542 6012 19572 6038
rect 19620 6050 19636 6084
rect 19670 6050 19686 6084
rect 19620 6034 19686 6050
rect 21326 6068 21356 6236
rect 21508 6084 21574 6100
rect 21326 6038 21460 6068
rect 19638 6012 19668 6034
rect 21430 6012 21460 6038
rect 21508 6050 21524 6084
rect 21558 6050 21574 6084
rect 21508 6034 21574 6050
rect 23214 6068 23244 6236
rect 23396 6084 23462 6100
rect 23214 6038 23348 6068
rect 21526 6012 21556 6034
rect 23318 6012 23348 6038
rect 23396 6050 23412 6084
rect 23446 6050 23462 6084
rect 23396 6034 23462 6050
rect 25102 6068 25132 6236
rect 25284 6084 25350 6100
rect 25102 6038 25236 6068
rect 23414 6012 23444 6034
rect 25206 6012 25236 6038
rect 25284 6050 25300 6084
rect 25334 6050 25350 6084
rect 25284 6034 25350 6050
rect 26990 6068 27020 6236
rect 27172 6084 27238 6100
rect 26990 6038 27124 6068
rect 25302 6012 25332 6034
rect 27094 6012 27124 6038
rect 27172 6050 27188 6084
rect 27222 6050 27238 6084
rect 27172 6034 27238 6050
rect 28878 6068 28908 6236
rect 29060 6084 29126 6100
rect 28878 6038 29012 6068
rect 27190 6012 27220 6034
rect 28982 6012 29012 6038
rect 29060 6050 29076 6084
rect 29110 6050 29126 6084
rect 29060 6034 29126 6050
rect 30766 6068 30796 6236
rect 30948 6084 31014 6100
rect 30766 6038 30900 6068
rect 29078 6012 29108 6034
rect 30870 6012 30900 6038
rect 30948 6050 30964 6084
rect 30998 6050 31014 6084
rect 30948 6034 31014 6050
rect 32654 6068 32684 6236
rect 32836 6084 32902 6100
rect 32654 6038 32788 6068
rect 30966 6012 30996 6034
rect 32758 6012 32788 6038
rect 32836 6050 32852 6084
rect 32886 6050 32902 6084
rect 32836 6034 32902 6050
rect 34542 6068 34572 6236
rect 34724 6084 34790 6100
rect 34542 6038 34676 6068
rect 32854 6012 32884 6034
rect 34646 6012 34676 6038
rect 34724 6050 34740 6084
rect 34774 6050 34790 6084
rect 34724 6034 34790 6050
rect 36430 6068 36460 6236
rect 36612 6084 36678 6100
rect 36430 6038 36564 6068
rect 34742 6012 34772 6034
rect 36534 6012 36564 6038
rect 36612 6050 36628 6084
rect 36662 6050 36678 6084
rect 36612 6034 36678 6050
rect 38318 6068 38348 6236
rect 38500 6084 38566 6100
rect 38318 6038 38452 6068
rect 36630 6012 36660 6034
rect 38422 6012 38452 6038
rect 38500 6050 38516 6084
rect 38550 6050 38566 6084
rect 38500 6034 38566 6050
rect 40206 6068 40236 6236
rect 40388 6084 40454 6100
rect 40206 6038 40340 6068
rect 38518 6012 38548 6034
rect 40310 6012 40340 6038
rect 40388 6050 40404 6084
rect 40438 6050 40454 6084
rect 40388 6034 40454 6050
rect 42094 6068 42124 6236
rect 42276 6084 42342 6100
rect 42094 6038 42228 6068
rect 40406 6012 40436 6034
rect 42198 6012 42228 6038
rect 42276 6050 42292 6084
rect 42326 6050 42342 6084
rect 42276 6034 42342 6050
rect 43982 6068 44012 6236
rect 44164 6084 44230 6100
rect 43982 6038 44116 6068
rect 42294 6012 42324 6034
rect 44086 6012 44116 6038
rect 44164 6050 44180 6084
rect 44214 6050 44230 6084
rect 44164 6034 44230 6050
rect 45864 6068 45894 6236
rect 46046 6084 46112 6100
rect 45864 6038 45998 6068
rect 44182 6012 44212 6034
rect 45968 6012 45998 6038
rect 46046 6050 46062 6084
rect 46096 6050 46112 6084
rect 46046 6034 46112 6050
rect 47752 6068 47782 6236
rect 47934 6084 48000 6100
rect 47752 6038 47886 6068
rect 46064 6012 46094 6034
rect 47856 6012 47886 6038
rect 47934 6050 47950 6084
rect 47984 6050 48000 6084
rect 47934 6034 48000 6050
rect 49640 6068 49670 6236
rect 49822 6084 49888 6100
rect 49640 6038 49774 6068
rect 47952 6012 47982 6034
rect 49744 6012 49774 6038
rect 49822 6050 49838 6084
rect 49872 6050 49888 6084
rect 49822 6034 49888 6050
rect 51528 6068 51558 6236
rect 51710 6084 51776 6100
rect 51528 6038 51662 6068
rect 49840 6012 49870 6034
rect 51632 6012 51662 6038
rect 51710 6050 51726 6084
rect 51760 6050 51776 6084
rect 51710 6034 51776 6050
rect 53416 6068 53446 6236
rect 53598 6084 53664 6100
rect 53416 6038 53550 6068
rect 51728 6012 51758 6034
rect 53520 6012 53550 6038
rect 53598 6050 53614 6084
rect 53648 6050 53664 6084
rect 53598 6034 53664 6050
rect 55304 6068 55334 6236
rect 55486 6084 55552 6100
rect 55304 6038 55438 6068
rect 53616 6012 53646 6034
rect 55408 6012 55438 6038
rect 55486 6050 55502 6084
rect 55536 6050 55552 6084
rect 55486 6034 55552 6050
rect 57192 6068 57222 6236
rect 57374 6084 57440 6100
rect 57192 6038 57326 6068
rect 55504 6012 55534 6034
rect 57296 6012 57326 6038
rect 57374 6050 57390 6084
rect 57424 6050 57440 6084
rect 57374 6034 57440 6050
rect 59080 6068 59110 6236
rect 59262 6084 59328 6100
rect 59080 6038 59214 6068
rect 57392 6012 57422 6034
rect 59184 6012 59214 6038
rect 59262 6050 59278 6084
rect 59312 6050 59328 6084
rect 59262 6034 59328 6050
rect 59280 6012 59310 6034
rect 668 5860 698 5882
rect 650 5844 716 5860
rect 764 5856 794 5882
rect 2556 5860 2586 5882
rect 650 5810 666 5844
rect 700 5810 716 5844
rect 241 5767 271 5793
rect 325 5767 355 5793
rect 650 5782 716 5810
rect 2538 5844 2604 5860
rect 2652 5856 2682 5882
rect 4444 5860 4474 5882
rect 2538 5810 2554 5844
rect 2588 5810 2604 5844
rect 650 5763 828 5782
rect 1055 5767 1085 5793
rect 1139 5767 1169 5793
rect 2129 5767 2159 5793
rect 2213 5767 2243 5793
rect 2538 5782 2604 5810
rect 4426 5844 4492 5860
rect 4540 5856 4570 5882
rect 6332 5860 6362 5882
rect 4426 5810 4442 5844
rect 4476 5810 4492 5844
rect 650 5750 778 5763
rect 762 5729 778 5750
rect 812 5729 828 5763
rect 762 5713 828 5729
rect 684 5682 714 5708
rect 780 5682 810 5713
rect 241 5615 271 5637
rect 179 5599 271 5615
rect 179 5565 195 5599
rect 229 5579 271 5599
rect 325 5615 355 5637
rect 325 5599 412 5615
rect 229 5565 283 5579
rect 179 5549 283 5565
rect 253 5517 283 5549
rect 325 5565 363 5599
rect 397 5565 412 5599
rect 325 5549 412 5565
rect 325 5517 355 5549
rect 2538 5763 2716 5782
rect 2943 5767 2973 5793
rect 3027 5767 3057 5793
rect 4017 5767 4047 5793
rect 4101 5767 4131 5793
rect 4426 5782 4492 5810
rect 6314 5844 6380 5860
rect 6428 5856 6458 5882
rect 8220 5860 8250 5882
rect 6314 5810 6330 5844
rect 6364 5810 6380 5844
rect 2538 5750 2666 5763
rect 2650 5729 2666 5750
rect 2700 5729 2716 5763
rect 2650 5713 2716 5729
rect 2572 5682 2602 5708
rect 2668 5682 2698 5713
rect 1055 5615 1085 5637
rect 993 5599 1085 5615
rect 993 5565 1009 5599
rect 1043 5579 1085 5599
rect 1139 5615 1169 5637
rect 2129 5615 2159 5637
rect 1139 5599 1226 5615
rect 1043 5565 1097 5579
rect 993 5549 1097 5565
rect 1067 5517 1097 5549
rect 1139 5565 1177 5599
rect 1211 5565 1226 5599
rect 1139 5549 1226 5565
rect 2067 5599 2159 5615
rect 2067 5565 2083 5599
rect 2117 5579 2159 5599
rect 2213 5615 2243 5637
rect 2213 5599 2300 5615
rect 2117 5565 2171 5579
rect 2067 5549 2171 5565
rect 1139 5517 1169 5549
rect 2141 5517 2171 5549
rect 2213 5565 2251 5599
rect 2285 5565 2300 5599
rect 2213 5549 2300 5565
rect 2213 5517 2243 5549
rect 684 5451 714 5482
rect 780 5456 810 5482
rect 666 5435 732 5451
rect 666 5401 682 5435
rect 716 5401 732 5435
rect 666 5385 732 5401
rect 253 5291 283 5317
rect 325 5291 355 5317
rect 4426 5763 4604 5782
rect 4831 5767 4861 5793
rect 4915 5767 4945 5793
rect 5905 5767 5935 5793
rect 5989 5767 6019 5793
rect 6314 5782 6380 5810
rect 8202 5844 8268 5860
rect 8316 5856 8346 5882
rect 10108 5860 10138 5882
rect 8202 5810 8218 5844
rect 8252 5810 8268 5844
rect 4426 5750 4554 5763
rect 4538 5729 4554 5750
rect 4588 5729 4604 5763
rect 4538 5713 4604 5729
rect 4460 5682 4490 5708
rect 4556 5682 4586 5713
rect 2943 5615 2973 5637
rect 2881 5599 2973 5615
rect 2881 5565 2897 5599
rect 2931 5579 2973 5599
rect 3027 5615 3057 5637
rect 4017 5615 4047 5637
rect 3027 5599 3114 5615
rect 2931 5565 2985 5579
rect 2881 5549 2985 5565
rect 2955 5517 2985 5549
rect 3027 5565 3065 5599
rect 3099 5565 3114 5599
rect 3027 5549 3114 5565
rect 3955 5599 4047 5615
rect 3955 5565 3971 5599
rect 4005 5579 4047 5599
rect 4101 5615 4131 5637
rect 4101 5599 4188 5615
rect 4005 5565 4059 5579
rect 3955 5549 4059 5565
rect 3027 5517 3057 5549
rect 4029 5517 4059 5549
rect 4101 5565 4139 5599
rect 4173 5565 4188 5599
rect 4101 5549 4188 5565
rect 4101 5517 4131 5549
rect 2572 5451 2602 5482
rect 2668 5456 2698 5482
rect 2554 5435 2620 5451
rect 2554 5401 2570 5435
rect 2604 5401 2620 5435
rect 2554 5385 2620 5401
rect 1067 5291 1097 5317
rect 1139 5291 1169 5317
rect 2141 5291 2171 5317
rect 2213 5291 2243 5317
rect 6314 5763 6492 5782
rect 6719 5767 6749 5793
rect 6803 5767 6833 5793
rect 7793 5767 7823 5793
rect 7877 5767 7907 5793
rect 8202 5782 8268 5810
rect 10090 5844 10156 5860
rect 10204 5856 10234 5882
rect 11996 5860 12026 5882
rect 10090 5810 10106 5844
rect 10140 5810 10156 5844
rect 6314 5750 6442 5763
rect 6426 5729 6442 5750
rect 6476 5729 6492 5763
rect 6426 5713 6492 5729
rect 6348 5682 6378 5708
rect 6444 5682 6474 5713
rect 4831 5615 4861 5637
rect 4769 5599 4861 5615
rect 4769 5565 4785 5599
rect 4819 5579 4861 5599
rect 4915 5615 4945 5637
rect 5905 5615 5935 5637
rect 4915 5599 5002 5615
rect 4819 5565 4873 5579
rect 4769 5549 4873 5565
rect 4843 5517 4873 5549
rect 4915 5565 4953 5599
rect 4987 5565 5002 5599
rect 4915 5549 5002 5565
rect 5843 5599 5935 5615
rect 5843 5565 5859 5599
rect 5893 5579 5935 5599
rect 5989 5615 6019 5637
rect 5989 5599 6076 5615
rect 5893 5565 5947 5579
rect 5843 5549 5947 5565
rect 4915 5517 4945 5549
rect 5917 5517 5947 5549
rect 5989 5565 6027 5599
rect 6061 5565 6076 5599
rect 5989 5549 6076 5565
rect 5989 5517 6019 5549
rect 4460 5451 4490 5482
rect 4556 5456 4586 5482
rect 4442 5435 4508 5451
rect 4442 5401 4458 5435
rect 4492 5401 4508 5435
rect 4442 5385 4508 5401
rect 2955 5291 2985 5317
rect 3027 5291 3057 5317
rect 4029 5291 4059 5317
rect 4101 5291 4131 5317
rect 8202 5763 8380 5782
rect 8607 5767 8637 5793
rect 8691 5767 8721 5793
rect 9681 5767 9711 5793
rect 9765 5767 9795 5793
rect 10090 5782 10156 5810
rect 11978 5844 12044 5860
rect 12092 5856 12122 5882
rect 13884 5860 13914 5882
rect 11978 5810 11994 5844
rect 12028 5810 12044 5844
rect 8202 5750 8330 5763
rect 8314 5729 8330 5750
rect 8364 5729 8380 5763
rect 8314 5713 8380 5729
rect 8236 5682 8266 5708
rect 8332 5682 8362 5713
rect 6719 5615 6749 5637
rect 6657 5599 6749 5615
rect 6657 5565 6673 5599
rect 6707 5579 6749 5599
rect 6803 5615 6833 5637
rect 7793 5615 7823 5637
rect 6803 5599 6890 5615
rect 6707 5565 6761 5579
rect 6657 5549 6761 5565
rect 6731 5517 6761 5549
rect 6803 5565 6841 5599
rect 6875 5565 6890 5599
rect 6803 5549 6890 5565
rect 7731 5599 7823 5615
rect 7731 5565 7747 5599
rect 7781 5579 7823 5599
rect 7877 5615 7907 5637
rect 7877 5599 7964 5615
rect 7781 5565 7835 5579
rect 7731 5549 7835 5565
rect 6803 5517 6833 5549
rect 7805 5517 7835 5549
rect 7877 5565 7915 5599
rect 7949 5565 7964 5599
rect 7877 5549 7964 5565
rect 7877 5517 7907 5549
rect 6348 5451 6378 5482
rect 6444 5456 6474 5482
rect 6330 5435 6396 5451
rect 6330 5401 6346 5435
rect 6380 5401 6396 5435
rect 6330 5385 6396 5401
rect 4843 5291 4873 5317
rect 4915 5291 4945 5317
rect 5917 5291 5947 5317
rect 5989 5291 6019 5317
rect 10090 5763 10268 5782
rect 10495 5767 10525 5793
rect 10579 5767 10609 5793
rect 11569 5767 11599 5793
rect 11653 5767 11683 5793
rect 11978 5782 12044 5810
rect 13866 5844 13932 5860
rect 13980 5856 14010 5882
rect 15766 5860 15796 5882
rect 13866 5810 13882 5844
rect 13916 5810 13932 5844
rect 10090 5750 10218 5763
rect 10202 5729 10218 5750
rect 10252 5729 10268 5763
rect 10202 5713 10268 5729
rect 10124 5682 10154 5708
rect 10220 5682 10250 5713
rect 8607 5615 8637 5637
rect 8545 5599 8637 5615
rect 8545 5565 8561 5599
rect 8595 5579 8637 5599
rect 8691 5615 8721 5637
rect 9681 5615 9711 5637
rect 8691 5599 8778 5615
rect 8595 5565 8649 5579
rect 8545 5549 8649 5565
rect 8619 5517 8649 5549
rect 8691 5565 8729 5599
rect 8763 5565 8778 5599
rect 8691 5549 8778 5565
rect 9619 5599 9711 5615
rect 9619 5565 9635 5599
rect 9669 5579 9711 5599
rect 9765 5615 9795 5637
rect 9765 5599 9852 5615
rect 9669 5565 9723 5579
rect 9619 5549 9723 5565
rect 8691 5517 8721 5549
rect 9693 5517 9723 5549
rect 9765 5565 9803 5599
rect 9837 5565 9852 5599
rect 9765 5549 9852 5565
rect 9765 5517 9795 5549
rect 8236 5451 8266 5482
rect 8332 5456 8362 5482
rect 8218 5435 8284 5451
rect 8218 5401 8234 5435
rect 8268 5401 8284 5435
rect 8218 5385 8284 5401
rect 6731 5291 6761 5317
rect 6803 5291 6833 5317
rect 7805 5291 7835 5317
rect 7877 5291 7907 5317
rect 11978 5763 12156 5782
rect 12383 5767 12413 5793
rect 12467 5767 12497 5793
rect 13457 5767 13487 5793
rect 13541 5767 13571 5793
rect 13866 5782 13932 5810
rect 15748 5844 15814 5860
rect 15862 5856 15892 5882
rect 17654 5860 17684 5882
rect 15748 5810 15764 5844
rect 15798 5810 15814 5844
rect 11978 5750 12106 5763
rect 12090 5729 12106 5750
rect 12140 5729 12156 5763
rect 12090 5713 12156 5729
rect 12012 5682 12042 5708
rect 12108 5682 12138 5713
rect 10495 5615 10525 5637
rect 10433 5599 10525 5615
rect 10433 5565 10449 5599
rect 10483 5579 10525 5599
rect 10579 5615 10609 5637
rect 11569 5615 11599 5637
rect 10579 5599 10666 5615
rect 10483 5565 10537 5579
rect 10433 5549 10537 5565
rect 10507 5517 10537 5549
rect 10579 5565 10617 5599
rect 10651 5565 10666 5599
rect 10579 5549 10666 5565
rect 11507 5599 11599 5615
rect 11507 5565 11523 5599
rect 11557 5579 11599 5599
rect 11653 5615 11683 5637
rect 11653 5599 11740 5615
rect 11557 5565 11611 5579
rect 11507 5549 11611 5565
rect 10579 5517 10609 5549
rect 11581 5517 11611 5549
rect 11653 5565 11691 5599
rect 11725 5565 11740 5599
rect 11653 5549 11740 5565
rect 11653 5517 11683 5549
rect 10124 5451 10154 5482
rect 10220 5456 10250 5482
rect 10106 5435 10172 5451
rect 10106 5401 10122 5435
rect 10156 5401 10172 5435
rect 10106 5385 10172 5401
rect 8619 5291 8649 5317
rect 8691 5291 8721 5317
rect 9693 5291 9723 5317
rect 9765 5291 9795 5317
rect 13866 5763 14044 5782
rect 14271 5767 14301 5793
rect 14355 5767 14385 5793
rect 15339 5767 15369 5793
rect 15423 5767 15453 5793
rect 15748 5782 15814 5810
rect 17636 5844 17702 5860
rect 17750 5856 17780 5882
rect 19542 5860 19572 5882
rect 17636 5810 17652 5844
rect 17686 5810 17702 5844
rect 13866 5750 13994 5763
rect 13978 5729 13994 5750
rect 14028 5729 14044 5763
rect 13978 5713 14044 5729
rect 13900 5682 13930 5708
rect 13996 5682 14026 5713
rect 12383 5615 12413 5637
rect 12321 5599 12413 5615
rect 12321 5565 12337 5599
rect 12371 5579 12413 5599
rect 12467 5615 12497 5637
rect 13457 5615 13487 5637
rect 12467 5599 12554 5615
rect 12371 5565 12425 5579
rect 12321 5549 12425 5565
rect 12395 5517 12425 5549
rect 12467 5565 12505 5599
rect 12539 5565 12554 5599
rect 12467 5549 12554 5565
rect 13395 5599 13487 5615
rect 13395 5565 13411 5599
rect 13445 5579 13487 5599
rect 13541 5615 13571 5637
rect 13541 5599 13628 5615
rect 13445 5565 13499 5579
rect 13395 5549 13499 5565
rect 12467 5517 12497 5549
rect 13469 5517 13499 5549
rect 13541 5565 13579 5599
rect 13613 5565 13628 5599
rect 13541 5549 13628 5565
rect 13541 5517 13571 5549
rect 12012 5451 12042 5482
rect 12108 5456 12138 5482
rect 11994 5435 12060 5451
rect 11994 5401 12010 5435
rect 12044 5401 12060 5435
rect 11994 5385 12060 5401
rect 10507 5291 10537 5317
rect 10579 5291 10609 5317
rect 11581 5291 11611 5317
rect 11653 5291 11683 5317
rect 15748 5763 15926 5782
rect 16153 5767 16183 5793
rect 16237 5767 16267 5793
rect 17227 5767 17257 5793
rect 17311 5767 17341 5793
rect 17636 5782 17702 5810
rect 19524 5844 19590 5860
rect 19638 5856 19668 5882
rect 21430 5860 21460 5882
rect 19524 5810 19540 5844
rect 19574 5810 19590 5844
rect 15748 5750 15876 5763
rect 15860 5729 15876 5750
rect 15910 5729 15926 5763
rect 15860 5713 15926 5729
rect 15782 5682 15812 5708
rect 15878 5682 15908 5713
rect 14271 5615 14301 5637
rect 14209 5599 14301 5615
rect 14209 5565 14225 5599
rect 14259 5579 14301 5599
rect 14355 5615 14385 5637
rect 15339 5615 15369 5637
rect 14355 5599 14442 5615
rect 14259 5565 14313 5579
rect 14209 5549 14313 5565
rect 14283 5517 14313 5549
rect 14355 5565 14393 5599
rect 14427 5565 14442 5599
rect 14355 5549 14442 5565
rect 15277 5599 15369 5615
rect 15277 5565 15293 5599
rect 15327 5579 15369 5599
rect 15423 5615 15453 5637
rect 15423 5599 15510 5615
rect 15327 5565 15381 5579
rect 15277 5549 15381 5565
rect 14355 5517 14385 5549
rect 15351 5517 15381 5549
rect 15423 5565 15461 5599
rect 15495 5565 15510 5599
rect 15423 5549 15510 5565
rect 15423 5517 15453 5549
rect 13900 5451 13930 5482
rect 13996 5456 14026 5482
rect 13882 5435 13948 5451
rect 13882 5401 13898 5435
rect 13932 5401 13948 5435
rect 13882 5385 13948 5401
rect 12395 5291 12425 5317
rect 12467 5291 12497 5317
rect 13469 5291 13499 5317
rect 13541 5291 13571 5317
rect 17636 5763 17814 5782
rect 18041 5767 18071 5793
rect 18125 5767 18155 5793
rect 19115 5767 19145 5793
rect 19199 5767 19229 5793
rect 19524 5782 19590 5810
rect 21412 5844 21478 5860
rect 21526 5856 21556 5882
rect 23318 5860 23348 5882
rect 21412 5810 21428 5844
rect 21462 5810 21478 5844
rect 17636 5750 17764 5763
rect 17748 5729 17764 5750
rect 17798 5729 17814 5763
rect 17748 5713 17814 5729
rect 17670 5682 17700 5708
rect 17766 5682 17796 5713
rect 16153 5615 16183 5637
rect 16091 5599 16183 5615
rect 16091 5565 16107 5599
rect 16141 5579 16183 5599
rect 16237 5615 16267 5637
rect 17227 5615 17257 5637
rect 16237 5599 16324 5615
rect 16141 5565 16195 5579
rect 16091 5549 16195 5565
rect 16165 5517 16195 5549
rect 16237 5565 16275 5599
rect 16309 5565 16324 5599
rect 16237 5549 16324 5565
rect 17165 5599 17257 5615
rect 17165 5565 17181 5599
rect 17215 5579 17257 5599
rect 17311 5615 17341 5637
rect 17311 5599 17398 5615
rect 17215 5565 17269 5579
rect 17165 5549 17269 5565
rect 16237 5517 16267 5549
rect 17239 5517 17269 5549
rect 17311 5565 17349 5599
rect 17383 5565 17398 5599
rect 17311 5549 17398 5565
rect 17311 5517 17341 5549
rect 15782 5451 15812 5482
rect 15878 5456 15908 5482
rect 15764 5435 15830 5451
rect 15764 5401 15780 5435
rect 15814 5401 15830 5435
rect 15764 5385 15830 5401
rect 14283 5291 14313 5317
rect 14355 5291 14385 5317
rect 15351 5291 15381 5317
rect 15423 5291 15453 5317
rect 19524 5763 19702 5782
rect 19929 5767 19959 5793
rect 20013 5767 20043 5793
rect 21003 5767 21033 5793
rect 21087 5767 21117 5793
rect 21412 5782 21478 5810
rect 23300 5844 23366 5860
rect 23414 5856 23444 5882
rect 25206 5860 25236 5882
rect 23300 5810 23316 5844
rect 23350 5810 23366 5844
rect 19524 5750 19652 5763
rect 19636 5729 19652 5750
rect 19686 5729 19702 5763
rect 19636 5713 19702 5729
rect 19558 5682 19588 5708
rect 19654 5682 19684 5713
rect 18041 5615 18071 5637
rect 17979 5599 18071 5615
rect 17979 5565 17995 5599
rect 18029 5579 18071 5599
rect 18125 5615 18155 5637
rect 19115 5615 19145 5637
rect 18125 5599 18212 5615
rect 18029 5565 18083 5579
rect 17979 5549 18083 5565
rect 18053 5517 18083 5549
rect 18125 5565 18163 5599
rect 18197 5565 18212 5599
rect 18125 5549 18212 5565
rect 19053 5599 19145 5615
rect 19053 5565 19069 5599
rect 19103 5579 19145 5599
rect 19199 5615 19229 5637
rect 19199 5599 19286 5615
rect 19103 5565 19157 5579
rect 19053 5549 19157 5565
rect 18125 5517 18155 5549
rect 19127 5517 19157 5549
rect 19199 5565 19237 5599
rect 19271 5565 19286 5599
rect 19199 5549 19286 5565
rect 19199 5517 19229 5549
rect 17670 5451 17700 5482
rect 17766 5456 17796 5482
rect 17652 5435 17718 5451
rect 17652 5401 17668 5435
rect 17702 5401 17718 5435
rect 17652 5385 17718 5401
rect 16165 5291 16195 5317
rect 16237 5291 16267 5317
rect 17239 5291 17269 5317
rect 17311 5291 17341 5317
rect 21412 5763 21590 5782
rect 21817 5767 21847 5793
rect 21901 5767 21931 5793
rect 22891 5767 22921 5793
rect 22975 5767 23005 5793
rect 23300 5782 23366 5810
rect 25188 5844 25254 5860
rect 25302 5856 25332 5882
rect 27094 5860 27124 5882
rect 25188 5810 25204 5844
rect 25238 5810 25254 5844
rect 21412 5750 21540 5763
rect 21524 5729 21540 5750
rect 21574 5729 21590 5763
rect 21524 5713 21590 5729
rect 21446 5682 21476 5708
rect 21542 5682 21572 5713
rect 19929 5615 19959 5637
rect 19867 5599 19959 5615
rect 19867 5565 19883 5599
rect 19917 5579 19959 5599
rect 20013 5615 20043 5637
rect 21003 5615 21033 5637
rect 20013 5599 20100 5615
rect 19917 5565 19971 5579
rect 19867 5549 19971 5565
rect 19941 5517 19971 5549
rect 20013 5565 20051 5599
rect 20085 5565 20100 5599
rect 20013 5549 20100 5565
rect 20941 5599 21033 5615
rect 20941 5565 20957 5599
rect 20991 5579 21033 5599
rect 21087 5615 21117 5637
rect 21087 5599 21174 5615
rect 20991 5565 21045 5579
rect 20941 5549 21045 5565
rect 20013 5517 20043 5549
rect 21015 5517 21045 5549
rect 21087 5565 21125 5599
rect 21159 5565 21174 5599
rect 21087 5549 21174 5565
rect 21087 5517 21117 5549
rect 19558 5451 19588 5482
rect 19654 5456 19684 5482
rect 19540 5435 19606 5451
rect 19540 5401 19556 5435
rect 19590 5401 19606 5435
rect 19540 5385 19606 5401
rect 18053 5291 18083 5317
rect 18125 5291 18155 5317
rect 19127 5291 19157 5317
rect 19199 5291 19229 5317
rect 23300 5763 23478 5782
rect 23705 5767 23735 5793
rect 23789 5767 23819 5793
rect 24779 5767 24809 5793
rect 24863 5767 24893 5793
rect 25188 5782 25254 5810
rect 27076 5844 27142 5860
rect 27190 5856 27220 5882
rect 28982 5860 29012 5882
rect 27076 5810 27092 5844
rect 27126 5810 27142 5844
rect 23300 5750 23428 5763
rect 23412 5729 23428 5750
rect 23462 5729 23478 5763
rect 23412 5713 23478 5729
rect 23334 5682 23364 5708
rect 23430 5682 23460 5713
rect 21817 5615 21847 5637
rect 21755 5599 21847 5615
rect 21755 5565 21771 5599
rect 21805 5579 21847 5599
rect 21901 5615 21931 5637
rect 22891 5615 22921 5637
rect 21901 5599 21988 5615
rect 21805 5565 21859 5579
rect 21755 5549 21859 5565
rect 21829 5517 21859 5549
rect 21901 5565 21939 5599
rect 21973 5565 21988 5599
rect 21901 5549 21988 5565
rect 22829 5599 22921 5615
rect 22829 5565 22845 5599
rect 22879 5579 22921 5599
rect 22975 5615 23005 5637
rect 22975 5599 23062 5615
rect 22879 5565 22933 5579
rect 22829 5549 22933 5565
rect 21901 5517 21931 5549
rect 22903 5517 22933 5549
rect 22975 5565 23013 5599
rect 23047 5565 23062 5599
rect 22975 5549 23062 5565
rect 22975 5517 23005 5549
rect 21446 5451 21476 5482
rect 21542 5456 21572 5482
rect 21428 5435 21494 5451
rect 21428 5401 21444 5435
rect 21478 5401 21494 5435
rect 21428 5385 21494 5401
rect 19941 5291 19971 5317
rect 20013 5291 20043 5317
rect 21015 5291 21045 5317
rect 21087 5291 21117 5317
rect 25188 5763 25366 5782
rect 25593 5767 25623 5793
rect 25677 5767 25707 5793
rect 26667 5767 26697 5793
rect 26751 5767 26781 5793
rect 27076 5782 27142 5810
rect 28964 5844 29030 5860
rect 29078 5856 29108 5882
rect 30870 5860 30900 5882
rect 28964 5810 28980 5844
rect 29014 5810 29030 5844
rect 25188 5750 25316 5763
rect 25300 5729 25316 5750
rect 25350 5729 25366 5763
rect 25300 5713 25366 5729
rect 25222 5682 25252 5708
rect 25318 5682 25348 5713
rect 23705 5615 23735 5637
rect 23643 5599 23735 5615
rect 23643 5565 23659 5599
rect 23693 5579 23735 5599
rect 23789 5615 23819 5637
rect 24779 5615 24809 5637
rect 23789 5599 23876 5615
rect 23693 5565 23747 5579
rect 23643 5549 23747 5565
rect 23717 5517 23747 5549
rect 23789 5565 23827 5599
rect 23861 5565 23876 5599
rect 23789 5549 23876 5565
rect 24717 5599 24809 5615
rect 24717 5565 24733 5599
rect 24767 5579 24809 5599
rect 24863 5615 24893 5637
rect 24863 5599 24950 5615
rect 24767 5565 24821 5579
rect 24717 5549 24821 5565
rect 23789 5517 23819 5549
rect 24791 5517 24821 5549
rect 24863 5565 24901 5599
rect 24935 5565 24950 5599
rect 24863 5549 24950 5565
rect 24863 5517 24893 5549
rect 23334 5451 23364 5482
rect 23430 5456 23460 5482
rect 23316 5435 23382 5451
rect 23316 5401 23332 5435
rect 23366 5401 23382 5435
rect 23316 5385 23382 5401
rect 21829 5291 21859 5317
rect 21901 5291 21931 5317
rect 22903 5291 22933 5317
rect 22975 5291 23005 5317
rect 27076 5763 27254 5782
rect 27481 5767 27511 5793
rect 27565 5767 27595 5793
rect 28555 5767 28585 5793
rect 28639 5767 28669 5793
rect 28964 5782 29030 5810
rect 30852 5844 30918 5860
rect 30966 5856 30996 5882
rect 32758 5860 32788 5882
rect 30852 5810 30868 5844
rect 30902 5810 30918 5844
rect 27076 5750 27204 5763
rect 27188 5729 27204 5750
rect 27238 5729 27254 5763
rect 27188 5713 27254 5729
rect 27110 5682 27140 5708
rect 27206 5682 27236 5713
rect 25593 5615 25623 5637
rect 25531 5599 25623 5615
rect 25531 5565 25547 5599
rect 25581 5579 25623 5599
rect 25677 5615 25707 5637
rect 26667 5615 26697 5637
rect 25677 5599 25764 5615
rect 25581 5565 25635 5579
rect 25531 5549 25635 5565
rect 25605 5517 25635 5549
rect 25677 5565 25715 5599
rect 25749 5565 25764 5599
rect 25677 5549 25764 5565
rect 26605 5599 26697 5615
rect 26605 5565 26621 5599
rect 26655 5579 26697 5599
rect 26751 5615 26781 5637
rect 26751 5599 26838 5615
rect 26655 5565 26709 5579
rect 26605 5549 26709 5565
rect 25677 5517 25707 5549
rect 26679 5517 26709 5549
rect 26751 5565 26789 5599
rect 26823 5565 26838 5599
rect 26751 5549 26838 5565
rect 26751 5517 26781 5549
rect 25222 5451 25252 5482
rect 25318 5456 25348 5482
rect 25204 5435 25270 5451
rect 25204 5401 25220 5435
rect 25254 5401 25270 5435
rect 25204 5385 25270 5401
rect 23717 5291 23747 5317
rect 23789 5291 23819 5317
rect 24791 5291 24821 5317
rect 24863 5291 24893 5317
rect 28964 5763 29142 5782
rect 29369 5767 29399 5793
rect 29453 5767 29483 5793
rect 30443 5767 30473 5793
rect 30527 5767 30557 5793
rect 30852 5782 30918 5810
rect 32740 5844 32806 5860
rect 32854 5856 32884 5882
rect 34646 5860 34676 5882
rect 32740 5810 32756 5844
rect 32790 5810 32806 5844
rect 28964 5750 29092 5763
rect 29076 5729 29092 5750
rect 29126 5729 29142 5763
rect 29076 5713 29142 5729
rect 28998 5682 29028 5708
rect 29094 5682 29124 5713
rect 27481 5615 27511 5637
rect 27419 5599 27511 5615
rect 27419 5565 27435 5599
rect 27469 5579 27511 5599
rect 27565 5615 27595 5637
rect 28555 5615 28585 5637
rect 27565 5599 27652 5615
rect 27469 5565 27523 5579
rect 27419 5549 27523 5565
rect 27493 5517 27523 5549
rect 27565 5565 27603 5599
rect 27637 5565 27652 5599
rect 27565 5549 27652 5565
rect 28493 5599 28585 5615
rect 28493 5565 28509 5599
rect 28543 5579 28585 5599
rect 28639 5615 28669 5637
rect 28639 5599 28726 5615
rect 28543 5565 28597 5579
rect 28493 5549 28597 5565
rect 27565 5517 27595 5549
rect 28567 5517 28597 5549
rect 28639 5565 28677 5599
rect 28711 5565 28726 5599
rect 28639 5549 28726 5565
rect 28639 5517 28669 5549
rect 27110 5451 27140 5482
rect 27206 5456 27236 5482
rect 27092 5435 27158 5451
rect 27092 5401 27108 5435
rect 27142 5401 27158 5435
rect 27092 5385 27158 5401
rect 25605 5291 25635 5317
rect 25677 5291 25707 5317
rect 26679 5291 26709 5317
rect 26751 5291 26781 5317
rect 30852 5763 31030 5782
rect 31257 5767 31287 5793
rect 31341 5767 31371 5793
rect 32331 5767 32361 5793
rect 32415 5767 32445 5793
rect 32740 5782 32806 5810
rect 34628 5844 34694 5860
rect 34742 5856 34772 5882
rect 36534 5860 36564 5882
rect 34628 5810 34644 5844
rect 34678 5810 34694 5844
rect 30852 5750 30980 5763
rect 30964 5729 30980 5750
rect 31014 5729 31030 5763
rect 30964 5713 31030 5729
rect 30886 5682 30916 5708
rect 30982 5682 31012 5713
rect 29369 5615 29399 5637
rect 29307 5599 29399 5615
rect 29307 5565 29323 5599
rect 29357 5579 29399 5599
rect 29453 5615 29483 5637
rect 30443 5615 30473 5637
rect 29453 5599 29540 5615
rect 29357 5565 29411 5579
rect 29307 5549 29411 5565
rect 29381 5517 29411 5549
rect 29453 5565 29491 5599
rect 29525 5565 29540 5599
rect 29453 5549 29540 5565
rect 30381 5599 30473 5615
rect 30381 5565 30397 5599
rect 30431 5579 30473 5599
rect 30527 5615 30557 5637
rect 30527 5599 30614 5615
rect 30431 5565 30485 5579
rect 30381 5549 30485 5565
rect 29453 5517 29483 5549
rect 30455 5517 30485 5549
rect 30527 5565 30565 5599
rect 30599 5565 30614 5599
rect 30527 5549 30614 5565
rect 30527 5517 30557 5549
rect 28998 5451 29028 5482
rect 29094 5456 29124 5482
rect 28980 5435 29046 5451
rect 28980 5401 28996 5435
rect 29030 5401 29046 5435
rect 28980 5385 29046 5401
rect 27493 5291 27523 5317
rect 27565 5291 27595 5317
rect 28567 5291 28597 5317
rect 28639 5291 28669 5317
rect 32740 5763 32918 5782
rect 33145 5767 33175 5793
rect 33229 5767 33259 5793
rect 34219 5767 34249 5793
rect 34303 5767 34333 5793
rect 34628 5782 34694 5810
rect 36516 5844 36582 5860
rect 36630 5856 36660 5882
rect 38422 5860 38452 5882
rect 36516 5810 36532 5844
rect 36566 5810 36582 5844
rect 32740 5750 32868 5763
rect 32852 5729 32868 5750
rect 32902 5729 32918 5763
rect 32852 5713 32918 5729
rect 32774 5682 32804 5708
rect 32870 5682 32900 5713
rect 31257 5615 31287 5637
rect 31195 5599 31287 5615
rect 31195 5565 31211 5599
rect 31245 5579 31287 5599
rect 31341 5615 31371 5637
rect 32331 5615 32361 5637
rect 31341 5599 31428 5615
rect 31245 5565 31299 5579
rect 31195 5549 31299 5565
rect 31269 5517 31299 5549
rect 31341 5565 31379 5599
rect 31413 5565 31428 5599
rect 31341 5549 31428 5565
rect 32269 5599 32361 5615
rect 32269 5565 32285 5599
rect 32319 5579 32361 5599
rect 32415 5615 32445 5637
rect 32415 5599 32502 5615
rect 32319 5565 32373 5579
rect 32269 5549 32373 5565
rect 31341 5517 31371 5549
rect 32343 5517 32373 5549
rect 32415 5565 32453 5599
rect 32487 5565 32502 5599
rect 32415 5549 32502 5565
rect 32415 5517 32445 5549
rect 30886 5451 30916 5482
rect 30982 5456 31012 5482
rect 30868 5435 30934 5451
rect 30868 5401 30884 5435
rect 30918 5401 30934 5435
rect 30868 5385 30934 5401
rect 29381 5291 29411 5317
rect 29453 5291 29483 5317
rect 30455 5291 30485 5317
rect 30527 5291 30557 5317
rect 34628 5763 34806 5782
rect 35033 5767 35063 5793
rect 35117 5767 35147 5793
rect 36107 5767 36137 5793
rect 36191 5767 36221 5793
rect 36516 5782 36582 5810
rect 38404 5844 38470 5860
rect 38518 5856 38548 5882
rect 40310 5860 40340 5882
rect 38404 5810 38420 5844
rect 38454 5810 38470 5844
rect 34628 5750 34756 5763
rect 34740 5729 34756 5750
rect 34790 5729 34806 5763
rect 34740 5713 34806 5729
rect 34662 5682 34692 5708
rect 34758 5682 34788 5713
rect 33145 5615 33175 5637
rect 33083 5599 33175 5615
rect 33083 5565 33099 5599
rect 33133 5579 33175 5599
rect 33229 5615 33259 5637
rect 34219 5615 34249 5637
rect 33229 5599 33316 5615
rect 33133 5565 33187 5579
rect 33083 5549 33187 5565
rect 33157 5517 33187 5549
rect 33229 5565 33267 5599
rect 33301 5565 33316 5599
rect 33229 5549 33316 5565
rect 34157 5599 34249 5615
rect 34157 5565 34173 5599
rect 34207 5579 34249 5599
rect 34303 5615 34333 5637
rect 34303 5599 34390 5615
rect 34207 5565 34261 5579
rect 34157 5549 34261 5565
rect 33229 5517 33259 5549
rect 34231 5517 34261 5549
rect 34303 5565 34341 5599
rect 34375 5565 34390 5599
rect 34303 5549 34390 5565
rect 34303 5517 34333 5549
rect 32774 5451 32804 5482
rect 32870 5456 32900 5482
rect 32756 5435 32822 5451
rect 32756 5401 32772 5435
rect 32806 5401 32822 5435
rect 32756 5385 32822 5401
rect 31269 5291 31299 5317
rect 31341 5291 31371 5317
rect 32343 5291 32373 5317
rect 32415 5291 32445 5317
rect 36516 5763 36694 5782
rect 36921 5767 36951 5793
rect 37005 5767 37035 5793
rect 37995 5767 38025 5793
rect 38079 5767 38109 5793
rect 38404 5782 38470 5810
rect 40292 5844 40358 5860
rect 40406 5856 40436 5882
rect 42198 5860 42228 5882
rect 40292 5810 40308 5844
rect 40342 5810 40358 5844
rect 36516 5750 36644 5763
rect 36628 5729 36644 5750
rect 36678 5729 36694 5763
rect 36628 5713 36694 5729
rect 36550 5682 36580 5708
rect 36646 5682 36676 5713
rect 35033 5615 35063 5637
rect 34971 5599 35063 5615
rect 34971 5565 34987 5599
rect 35021 5579 35063 5599
rect 35117 5615 35147 5637
rect 36107 5615 36137 5637
rect 35117 5599 35204 5615
rect 35021 5565 35075 5579
rect 34971 5549 35075 5565
rect 35045 5517 35075 5549
rect 35117 5565 35155 5599
rect 35189 5565 35204 5599
rect 35117 5549 35204 5565
rect 36045 5599 36137 5615
rect 36045 5565 36061 5599
rect 36095 5579 36137 5599
rect 36191 5615 36221 5637
rect 36191 5599 36278 5615
rect 36095 5565 36149 5579
rect 36045 5549 36149 5565
rect 35117 5517 35147 5549
rect 36119 5517 36149 5549
rect 36191 5565 36229 5599
rect 36263 5565 36278 5599
rect 36191 5549 36278 5565
rect 36191 5517 36221 5549
rect 34662 5451 34692 5482
rect 34758 5456 34788 5482
rect 34644 5435 34710 5451
rect 34644 5401 34660 5435
rect 34694 5401 34710 5435
rect 34644 5385 34710 5401
rect 33157 5291 33187 5317
rect 33229 5291 33259 5317
rect 34231 5291 34261 5317
rect 34303 5291 34333 5317
rect 38404 5763 38582 5782
rect 38809 5767 38839 5793
rect 38893 5767 38923 5793
rect 39883 5767 39913 5793
rect 39967 5767 39997 5793
rect 40292 5782 40358 5810
rect 42180 5844 42246 5860
rect 42294 5856 42324 5882
rect 44086 5860 44116 5882
rect 42180 5810 42196 5844
rect 42230 5810 42246 5844
rect 38404 5750 38532 5763
rect 38516 5729 38532 5750
rect 38566 5729 38582 5763
rect 38516 5713 38582 5729
rect 38438 5682 38468 5708
rect 38534 5682 38564 5713
rect 36921 5615 36951 5637
rect 36859 5599 36951 5615
rect 36859 5565 36875 5599
rect 36909 5579 36951 5599
rect 37005 5615 37035 5637
rect 37995 5615 38025 5637
rect 37005 5599 37092 5615
rect 36909 5565 36963 5579
rect 36859 5549 36963 5565
rect 36933 5517 36963 5549
rect 37005 5565 37043 5599
rect 37077 5565 37092 5599
rect 37005 5549 37092 5565
rect 37933 5599 38025 5615
rect 37933 5565 37949 5599
rect 37983 5579 38025 5599
rect 38079 5615 38109 5637
rect 38079 5599 38166 5615
rect 37983 5565 38037 5579
rect 37933 5549 38037 5565
rect 37005 5517 37035 5549
rect 38007 5517 38037 5549
rect 38079 5565 38117 5599
rect 38151 5565 38166 5599
rect 38079 5549 38166 5565
rect 38079 5517 38109 5549
rect 36550 5451 36580 5482
rect 36646 5456 36676 5482
rect 36532 5435 36598 5451
rect 36532 5401 36548 5435
rect 36582 5401 36598 5435
rect 36532 5385 36598 5401
rect 35045 5291 35075 5317
rect 35117 5291 35147 5317
rect 36119 5291 36149 5317
rect 36191 5291 36221 5317
rect 40292 5763 40470 5782
rect 40697 5767 40727 5793
rect 40781 5767 40811 5793
rect 41771 5767 41801 5793
rect 41855 5767 41885 5793
rect 42180 5782 42246 5810
rect 44068 5844 44134 5860
rect 44182 5856 44212 5882
rect 45968 5860 45998 5882
rect 44068 5810 44084 5844
rect 44118 5810 44134 5844
rect 40292 5750 40420 5763
rect 40404 5729 40420 5750
rect 40454 5729 40470 5763
rect 40404 5713 40470 5729
rect 40326 5682 40356 5708
rect 40422 5682 40452 5713
rect 38809 5615 38839 5637
rect 38747 5599 38839 5615
rect 38747 5565 38763 5599
rect 38797 5579 38839 5599
rect 38893 5615 38923 5637
rect 39883 5615 39913 5637
rect 38893 5599 38980 5615
rect 38797 5565 38851 5579
rect 38747 5549 38851 5565
rect 38821 5517 38851 5549
rect 38893 5565 38931 5599
rect 38965 5565 38980 5599
rect 38893 5549 38980 5565
rect 39821 5599 39913 5615
rect 39821 5565 39837 5599
rect 39871 5579 39913 5599
rect 39967 5615 39997 5637
rect 39967 5599 40054 5615
rect 39871 5565 39925 5579
rect 39821 5549 39925 5565
rect 38893 5517 38923 5549
rect 39895 5517 39925 5549
rect 39967 5565 40005 5599
rect 40039 5565 40054 5599
rect 39967 5549 40054 5565
rect 39967 5517 39997 5549
rect 38438 5451 38468 5482
rect 38534 5456 38564 5482
rect 38420 5435 38486 5451
rect 38420 5401 38436 5435
rect 38470 5401 38486 5435
rect 38420 5385 38486 5401
rect 36933 5291 36963 5317
rect 37005 5291 37035 5317
rect 38007 5291 38037 5317
rect 38079 5291 38109 5317
rect 42180 5763 42358 5782
rect 42585 5767 42615 5793
rect 42669 5767 42699 5793
rect 43659 5767 43689 5793
rect 43743 5767 43773 5793
rect 44068 5782 44134 5810
rect 45950 5844 46016 5860
rect 46064 5856 46094 5882
rect 47856 5860 47886 5882
rect 45950 5810 45966 5844
rect 46000 5810 46016 5844
rect 42180 5750 42308 5763
rect 42292 5729 42308 5750
rect 42342 5729 42358 5763
rect 42292 5713 42358 5729
rect 42214 5682 42244 5708
rect 42310 5682 42340 5713
rect 40697 5615 40727 5637
rect 40635 5599 40727 5615
rect 40635 5565 40651 5599
rect 40685 5579 40727 5599
rect 40781 5615 40811 5637
rect 41771 5615 41801 5637
rect 40781 5599 40868 5615
rect 40685 5565 40739 5579
rect 40635 5549 40739 5565
rect 40709 5517 40739 5549
rect 40781 5565 40819 5599
rect 40853 5565 40868 5599
rect 40781 5549 40868 5565
rect 41709 5599 41801 5615
rect 41709 5565 41725 5599
rect 41759 5579 41801 5599
rect 41855 5615 41885 5637
rect 41855 5599 41942 5615
rect 41759 5565 41813 5579
rect 41709 5549 41813 5565
rect 40781 5517 40811 5549
rect 41783 5517 41813 5549
rect 41855 5565 41893 5599
rect 41927 5565 41942 5599
rect 41855 5549 41942 5565
rect 41855 5517 41885 5549
rect 40326 5451 40356 5482
rect 40422 5456 40452 5482
rect 40308 5435 40374 5451
rect 40308 5401 40324 5435
rect 40358 5401 40374 5435
rect 40308 5385 40374 5401
rect 38821 5291 38851 5317
rect 38893 5291 38923 5317
rect 39895 5291 39925 5317
rect 39967 5291 39997 5317
rect 44068 5763 44246 5782
rect 44473 5767 44503 5793
rect 44557 5767 44587 5793
rect 45541 5767 45571 5793
rect 45625 5767 45655 5793
rect 45950 5782 46016 5810
rect 47838 5844 47904 5860
rect 47952 5856 47982 5882
rect 49744 5860 49774 5882
rect 47838 5810 47854 5844
rect 47888 5810 47904 5844
rect 44068 5750 44196 5763
rect 44180 5729 44196 5750
rect 44230 5729 44246 5763
rect 44180 5713 44246 5729
rect 44102 5682 44132 5708
rect 44198 5682 44228 5713
rect 42585 5615 42615 5637
rect 42523 5599 42615 5615
rect 42523 5565 42539 5599
rect 42573 5579 42615 5599
rect 42669 5615 42699 5637
rect 43659 5615 43689 5637
rect 42669 5599 42756 5615
rect 42573 5565 42627 5579
rect 42523 5549 42627 5565
rect 42597 5517 42627 5549
rect 42669 5565 42707 5599
rect 42741 5565 42756 5599
rect 42669 5549 42756 5565
rect 43597 5599 43689 5615
rect 43597 5565 43613 5599
rect 43647 5579 43689 5599
rect 43743 5615 43773 5637
rect 43743 5599 43830 5615
rect 43647 5565 43701 5579
rect 43597 5549 43701 5565
rect 42669 5517 42699 5549
rect 43671 5517 43701 5549
rect 43743 5565 43781 5599
rect 43815 5565 43830 5599
rect 43743 5549 43830 5565
rect 43743 5517 43773 5549
rect 42214 5451 42244 5482
rect 42310 5456 42340 5482
rect 42196 5435 42262 5451
rect 42196 5401 42212 5435
rect 42246 5401 42262 5435
rect 42196 5385 42262 5401
rect 40709 5291 40739 5317
rect 40781 5291 40811 5317
rect 41783 5291 41813 5317
rect 41855 5291 41885 5317
rect 45950 5763 46128 5782
rect 46355 5767 46385 5793
rect 46439 5767 46469 5793
rect 47429 5767 47459 5793
rect 47513 5767 47543 5793
rect 47838 5782 47904 5810
rect 49726 5844 49792 5860
rect 49840 5856 49870 5882
rect 51632 5860 51662 5882
rect 49726 5810 49742 5844
rect 49776 5810 49792 5844
rect 45950 5750 46078 5763
rect 46062 5729 46078 5750
rect 46112 5729 46128 5763
rect 46062 5713 46128 5729
rect 45984 5682 46014 5708
rect 46080 5682 46110 5713
rect 44473 5615 44503 5637
rect 44411 5599 44503 5615
rect 44411 5565 44427 5599
rect 44461 5579 44503 5599
rect 44557 5615 44587 5637
rect 45541 5615 45571 5637
rect 44557 5599 44644 5615
rect 44461 5565 44515 5579
rect 44411 5549 44515 5565
rect 44485 5517 44515 5549
rect 44557 5565 44595 5599
rect 44629 5565 44644 5599
rect 44557 5549 44644 5565
rect 45479 5599 45571 5615
rect 45479 5565 45495 5599
rect 45529 5579 45571 5599
rect 45625 5615 45655 5637
rect 45625 5599 45712 5615
rect 45529 5565 45583 5579
rect 45479 5549 45583 5565
rect 44557 5517 44587 5549
rect 45553 5517 45583 5549
rect 45625 5565 45663 5599
rect 45697 5565 45712 5599
rect 45625 5549 45712 5565
rect 45625 5517 45655 5549
rect 44102 5451 44132 5482
rect 44198 5456 44228 5482
rect 44084 5435 44150 5451
rect 44084 5401 44100 5435
rect 44134 5401 44150 5435
rect 44084 5385 44150 5401
rect 42597 5291 42627 5317
rect 42669 5291 42699 5317
rect 43671 5291 43701 5317
rect 43743 5291 43773 5317
rect 47838 5763 48016 5782
rect 48243 5767 48273 5793
rect 48327 5767 48357 5793
rect 49317 5767 49347 5793
rect 49401 5767 49431 5793
rect 49726 5782 49792 5810
rect 51614 5844 51680 5860
rect 51728 5856 51758 5882
rect 53520 5860 53550 5882
rect 51614 5810 51630 5844
rect 51664 5810 51680 5844
rect 47838 5750 47966 5763
rect 47950 5729 47966 5750
rect 48000 5729 48016 5763
rect 47950 5713 48016 5729
rect 47872 5682 47902 5708
rect 47968 5682 47998 5713
rect 46355 5615 46385 5637
rect 46293 5599 46385 5615
rect 46293 5565 46309 5599
rect 46343 5579 46385 5599
rect 46439 5615 46469 5637
rect 47429 5615 47459 5637
rect 46439 5599 46526 5615
rect 46343 5565 46397 5579
rect 46293 5549 46397 5565
rect 46367 5517 46397 5549
rect 46439 5565 46477 5599
rect 46511 5565 46526 5599
rect 46439 5549 46526 5565
rect 47367 5599 47459 5615
rect 47367 5565 47383 5599
rect 47417 5579 47459 5599
rect 47513 5615 47543 5637
rect 47513 5599 47600 5615
rect 47417 5565 47471 5579
rect 47367 5549 47471 5565
rect 46439 5517 46469 5549
rect 47441 5517 47471 5549
rect 47513 5565 47551 5599
rect 47585 5565 47600 5599
rect 47513 5549 47600 5565
rect 47513 5517 47543 5549
rect 45984 5451 46014 5482
rect 46080 5456 46110 5482
rect 45966 5435 46032 5451
rect 45966 5401 45982 5435
rect 46016 5401 46032 5435
rect 45966 5385 46032 5401
rect 44485 5291 44515 5317
rect 44557 5291 44587 5317
rect 45553 5291 45583 5317
rect 45625 5291 45655 5317
rect 49726 5763 49904 5782
rect 50131 5767 50161 5793
rect 50215 5767 50245 5793
rect 51205 5767 51235 5793
rect 51289 5767 51319 5793
rect 51614 5782 51680 5810
rect 53502 5844 53568 5860
rect 53616 5856 53646 5882
rect 55408 5860 55438 5882
rect 53502 5810 53518 5844
rect 53552 5810 53568 5844
rect 49726 5750 49854 5763
rect 49838 5729 49854 5750
rect 49888 5729 49904 5763
rect 49838 5713 49904 5729
rect 49760 5682 49790 5708
rect 49856 5682 49886 5713
rect 48243 5615 48273 5637
rect 48181 5599 48273 5615
rect 48181 5565 48197 5599
rect 48231 5579 48273 5599
rect 48327 5615 48357 5637
rect 49317 5615 49347 5637
rect 48327 5599 48414 5615
rect 48231 5565 48285 5579
rect 48181 5549 48285 5565
rect 48255 5517 48285 5549
rect 48327 5565 48365 5599
rect 48399 5565 48414 5599
rect 48327 5549 48414 5565
rect 49255 5599 49347 5615
rect 49255 5565 49271 5599
rect 49305 5579 49347 5599
rect 49401 5615 49431 5637
rect 49401 5599 49488 5615
rect 49305 5565 49359 5579
rect 49255 5549 49359 5565
rect 48327 5517 48357 5549
rect 49329 5517 49359 5549
rect 49401 5565 49439 5599
rect 49473 5565 49488 5599
rect 49401 5549 49488 5565
rect 49401 5517 49431 5549
rect 47872 5451 47902 5482
rect 47968 5456 47998 5482
rect 47854 5435 47920 5451
rect 47854 5401 47870 5435
rect 47904 5401 47920 5435
rect 47854 5385 47920 5401
rect 46367 5291 46397 5317
rect 46439 5291 46469 5317
rect 47441 5291 47471 5317
rect 47513 5291 47543 5317
rect 51614 5763 51792 5782
rect 52019 5767 52049 5793
rect 52103 5767 52133 5793
rect 53093 5767 53123 5793
rect 53177 5767 53207 5793
rect 53502 5782 53568 5810
rect 55390 5844 55456 5860
rect 55504 5856 55534 5882
rect 57296 5860 57326 5882
rect 55390 5810 55406 5844
rect 55440 5810 55456 5844
rect 51614 5750 51742 5763
rect 51726 5729 51742 5750
rect 51776 5729 51792 5763
rect 51726 5713 51792 5729
rect 51648 5682 51678 5708
rect 51744 5682 51774 5713
rect 50131 5615 50161 5637
rect 50069 5599 50161 5615
rect 50069 5565 50085 5599
rect 50119 5579 50161 5599
rect 50215 5615 50245 5637
rect 51205 5615 51235 5637
rect 50215 5599 50302 5615
rect 50119 5565 50173 5579
rect 50069 5549 50173 5565
rect 50143 5517 50173 5549
rect 50215 5565 50253 5599
rect 50287 5565 50302 5599
rect 50215 5549 50302 5565
rect 51143 5599 51235 5615
rect 51143 5565 51159 5599
rect 51193 5579 51235 5599
rect 51289 5615 51319 5637
rect 51289 5599 51376 5615
rect 51193 5565 51247 5579
rect 51143 5549 51247 5565
rect 50215 5517 50245 5549
rect 51217 5517 51247 5549
rect 51289 5565 51327 5599
rect 51361 5565 51376 5599
rect 51289 5549 51376 5565
rect 51289 5517 51319 5549
rect 49760 5451 49790 5482
rect 49856 5456 49886 5482
rect 49742 5435 49808 5451
rect 49742 5401 49758 5435
rect 49792 5401 49808 5435
rect 49742 5385 49808 5401
rect 48255 5291 48285 5317
rect 48327 5291 48357 5317
rect 49329 5291 49359 5317
rect 49401 5291 49431 5317
rect 53502 5763 53680 5782
rect 53907 5767 53937 5793
rect 53991 5767 54021 5793
rect 54981 5767 55011 5793
rect 55065 5767 55095 5793
rect 55390 5782 55456 5810
rect 57278 5844 57344 5860
rect 57392 5856 57422 5882
rect 59184 5860 59214 5882
rect 57278 5810 57294 5844
rect 57328 5810 57344 5844
rect 53502 5750 53630 5763
rect 53614 5729 53630 5750
rect 53664 5729 53680 5763
rect 53614 5713 53680 5729
rect 53536 5682 53566 5708
rect 53632 5682 53662 5713
rect 52019 5615 52049 5637
rect 51957 5599 52049 5615
rect 51957 5565 51973 5599
rect 52007 5579 52049 5599
rect 52103 5615 52133 5637
rect 53093 5615 53123 5637
rect 52103 5599 52190 5615
rect 52007 5565 52061 5579
rect 51957 5549 52061 5565
rect 52031 5517 52061 5549
rect 52103 5565 52141 5599
rect 52175 5565 52190 5599
rect 52103 5549 52190 5565
rect 53031 5599 53123 5615
rect 53031 5565 53047 5599
rect 53081 5579 53123 5599
rect 53177 5615 53207 5637
rect 53177 5599 53264 5615
rect 53081 5565 53135 5579
rect 53031 5549 53135 5565
rect 52103 5517 52133 5549
rect 53105 5517 53135 5549
rect 53177 5565 53215 5599
rect 53249 5565 53264 5599
rect 53177 5549 53264 5565
rect 53177 5517 53207 5549
rect 51648 5451 51678 5482
rect 51744 5456 51774 5482
rect 51630 5435 51696 5451
rect 51630 5401 51646 5435
rect 51680 5401 51696 5435
rect 51630 5385 51696 5401
rect 50143 5291 50173 5317
rect 50215 5291 50245 5317
rect 51217 5291 51247 5317
rect 51289 5291 51319 5317
rect 55390 5763 55568 5782
rect 55795 5767 55825 5793
rect 55879 5767 55909 5793
rect 56869 5767 56899 5793
rect 56953 5767 56983 5793
rect 57278 5782 57344 5810
rect 59166 5844 59232 5860
rect 59280 5856 59310 5882
rect 59166 5810 59182 5844
rect 59216 5810 59232 5844
rect 55390 5750 55518 5763
rect 55502 5729 55518 5750
rect 55552 5729 55568 5763
rect 55502 5713 55568 5729
rect 55424 5682 55454 5708
rect 55520 5682 55550 5713
rect 53907 5615 53937 5637
rect 53845 5599 53937 5615
rect 53845 5565 53861 5599
rect 53895 5579 53937 5599
rect 53991 5615 54021 5637
rect 54981 5615 55011 5637
rect 53991 5599 54078 5615
rect 53895 5565 53949 5579
rect 53845 5549 53949 5565
rect 53919 5517 53949 5549
rect 53991 5565 54029 5599
rect 54063 5565 54078 5599
rect 53991 5549 54078 5565
rect 54919 5599 55011 5615
rect 54919 5565 54935 5599
rect 54969 5579 55011 5599
rect 55065 5615 55095 5637
rect 55065 5599 55152 5615
rect 54969 5565 55023 5579
rect 54919 5549 55023 5565
rect 53991 5517 54021 5549
rect 54993 5517 55023 5549
rect 55065 5565 55103 5599
rect 55137 5565 55152 5599
rect 55065 5549 55152 5565
rect 55065 5517 55095 5549
rect 53536 5451 53566 5482
rect 53632 5456 53662 5482
rect 53518 5435 53584 5451
rect 53518 5401 53534 5435
rect 53568 5401 53584 5435
rect 53518 5385 53584 5401
rect 52031 5291 52061 5317
rect 52103 5291 52133 5317
rect 53105 5291 53135 5317
rect 53177 5291 53207 5317
rect 57278 5763 57456 5782
rect 57683 5767 57713 5793
rect 57767 5767 57797 5793
rect 58757 5767 58787 5793
rect 58841 5767 58871 5793
rect 59166 5782 59232 5810
rect 57278 5750 57406 5763
rect 57390 5729 57406 5750
rect 57440 5729 57456 5763
rect 57390 5713 57456 5729
rect 57312 5682 57342 5708
rect 57408 5682 57438 5713
rect 55795 5615 55825 5637
rect 55733 5599 55825 5615
rect 55733 5565 55749 5599
rect 55783 5579 55825 5599
rect 55879 5615 55909 5637
rect 56869 5615 56899 5637
rect 55879 5599 55966 5615
rect 55783 5565 55837 5579
rect 55733 5549 55837 5565
rect 55807 5517 55837 5549
rect 55879 5565 55917 5599
rect 55951 5565 55966 5599
rect 55879 5549 55966 5565
rect 56807 5599 56899 5615
rect 56807 5565 56823 5599
rect 56857 5579 56899 5599
rect 56953 5615 56983 5637
rect 56953 5599 57040 5615
rect 56857 5565 56911 5579
rect 56807 5549 56911 5565
rect 55879 5517 55909 5549
rect 56881 5517 56911 5549
rect 56953 5565 56991 5599
rect 57025 5565 57040 5599
rect 56953 5549 57040 5565
rect 56953 5517 56983 5549
rect 55424 5451 55454 5482
rect 55520 5456 55550 5482
rect 55406 5435 55472 5451
rect 55406 5401 55422 5435
rect 55456 5401 55472 5435
rect 55406 5385 55472 5401
rect 53919 5291 53949 5317
rect 53991 5291 54021 5317
rect 54993 5291 55023 5317
rect 55065 5291 55095 5317
rect 59166 5763 59344 5782
rect 59571 5767 59601 5793
rect 59655 5767 59685 5793
rect 59166 5750 59294 5763
rect 59278 5729 59294 5750
rect 59328 5729 59344 5763
rect 59278 5713 59344 5729
rect 59200 5682 59230 5708
rect 59296 5682 59326 5713
rect 57683 5615 57713 5637
rect 57621 5599 57713 5615
rect 57621 5565 57637 5599
rect 57671 5579 57713 5599
rect 57767 5615 57797 5637
rect 58757 5615 58787 5637
rect 57767 5599 57854 5615
rect 57671 5565 57725 5579
rect 57621 5549 57725 5565
rect 57695 5517 57725 5549
rect 57767 5565 57805 5599
rect 57839 5565 57854 5599
rect 57767 5549 57854 5565
rect 58695 5599 58787 5615
rect 58695 5565 58711 5599
rect 58745 5579 58787 5599
rect 58841 5615 58871 5637
rect 58841 5599 58928 5615
rect 58745 5565 58799 5579
rect 58695 5549 58799 5565
rect 57767 5517 57797 5549
rect 58769 5517 58799 5549
rect 58841 5565 58879 5599
rect 58913 5565 58928 5599
rect 58841 5549 58928 5565
rect 58841 5517 58871 5549
rect 57312 5451 57342 5482
rect 57408 5456 57438 5482
rect 57294 5435 57360 5451
rect 57294 5401 57310 5435
rect 57344 5401 57360 5435
rect 57294 5385 57360 5401
rect 55807 5291 55837 5317
rect 55879 5291 55909 5317
rect 56881 5291 56911 5317
rect 56953 5291 56983 5317
rect 59571 5615 59601 5637
rect 59509 5599 59601 5615
rect 59509 5565 59525 5599
rect 59559 5579 59601 5599
rect 59655 5615 59685 5637
rect 59655 5599 59742 5615
rect 59559 5565 59613 5579
rect 59509 5549 59613 5565
rect 59583 5517 59613 5549
rect 59655 5565 59693 5599
rect 59727 5565 59742 5599
rect 59655 5549 59742 5565
rect 59655 5517 59685 5549
rect 59200 5451 59230 5482
rect 59296 5456 59326 5482
rect 59182 5435 59248 5451
rect 59182 5401 59198 5435
rect 59232 5401 59248 5435
rect 59182 5385 59248 5401
rect 57695 5291 57725 5317
rect 57767 5291 57797 5317
rect 58769 5291 58799 5317
rect 58841 5291 58871 5317
rect 59583 5291 59613 5317
rect 59655 5291 59685 5317
rect 5754 5145 5784 5171
rect 5838 5145 5868 5171
rect 5922 5145 5952 5171
rect 6006 5145 6036 5171
rect 6090 5145 6120 5171
rect 6174 5145 6204 5171
rect 6258 5145 6288 5171
rect 6342 5145 6372 5171
rect 6426 5145 6456 5171
rect 6510 5145 6540 5171
rect 6594 5145 6624 5171
rect 6678 5145 6708 5171
rect 6762 5145 6792 5171
rect 6846 5145 6876 5171
rect 6930 5145 6960 5171
rect 7014 5145 7044 5171
rect 7636 5143 7666 5169
rect 7720 5143 7750 5169
rect 7804 5143 7834 5169
rect 7888 5143 7918 5169
rect 7972 5143 8002 5169
rect 8056 5143 8086 5169
rect 8140 5143 8170 5169
rect 8224 5143 8254 5169
rect 8308 5143 8338 5169
rect 8392 5143 8422 5169
rect 8476 5143 8506 5169
rect 8560 5143 8590 5169
rect 8644 5143 8674 5169
rect 8728 5143 8758 5169
rect 8812 5143 8842 5169
rect 8896 5143 8926 5169
rect 20852 5145 20882 5171
rect 20936 5145 20966 5171
rect 21020 5145 21050 5171
rect 21104 5145 21134 5171
rect 21188 5145 21218 5171
rect 21272 5145 21302 5171
rect 21356 5145 21386 5171
rect 21440 5145 21470 5171
rect 21524 5145 21554 5171
rect 21608 5145 21638 5171
rect 21692 5145 21722 5171
rect 21776 5145 21806 5171
rect 21860 5145 21890 5171
rect 21944 5145 21974 5171
rect 22028 5145 22058 5171
rect 22112 5145 22142 5171
rect 5754 4913 5784 4945
rect 5838 4913 5868 4945
rect 5922 4913 5952 4945
rect 6006 4913 6036 4945
rect 6090 4913 6120 4945
rect 6174 4913 6204 4945
rect 6258 4913 6288 4945
rect 6342 4913 6372 4945
rect 6426 4913 6456 4945
rect 6510 4913 6540 4945
rect 6594 4913 6624 4945
rect 6678 4913 6708 4945
rect 6762 4913 6792 4945
rect 6846 4913 6876 4945
rect 6930 4913 6960 4945
rect 7014 4913 7044 4945
rect 22734 5143 22764 5169
rect 22818 5143 22848 5169
rect 22902 5143 22932 5169
rect 22986 5143 23016 5169
rect 23070 5143 23100 5169
rect 23154 5143 23184 5169
rect 23238 5143 23268 5169
rect 23322 5143 23352 5169
rect 23406 5143 23436 5169
rect 23490 5143 23520 5169
rect 23574 5143 23604 5169
rect 23658 5143 23688 5169
rect 23742 5143 23772 5169
rect 23826 5143 23856 5169
rect 23910 5143 23940 5169
rect 23994 5143 24024 5169
rect 35956 5145 35986 5171
rect 36040 5145 36070 5171
rect 36124 5145 36154 5171
rect 36208 5145 36238 5171
rect 36292 5145 36322 5171
rect 36376 5145 36406 5171
rect 36460 5145 36490 5171
rect 36544 5145 36574 5171
rect 36628 5145 36658 5171
rect 36712 5145 36742 5171
rect 36796 5145 36826 5171
rect 36880 5145 36910 5171
rect 36964 5145 36994 5171
rect 37048 5145 37078 5171
rect 37132 5145 37162 5171
rect 37216 5145 37246 5171
rect 5754 4897 7110 4913
rect 5754 4863 6047 4897
rect 6081 4863 6214 4897
rect 6248 4863 6382 4897
rect 6416 4863 6549 4897
rect 6583 4863 6718 4897
rect 6752 4863 6886 4897
rect 6920 4863 7060 4897
rect 7094 4863 7110 4897
rect 5754 4847 7110 4863
rect 7636 4911 7666 4943
rect 7720 4911 7750 4943
rect 7804 4911 7834 4943
rect 7888 4911 7918 4943
rect 7972 4911 8002 4943
rect 8056 4911 8086 4943
rect 8140 4911 8170 4943
rect 8224 4911 8254 4943
rect 8308 4911 8338 4943
rect 8392 4911 8422 4943
rect 8476 4911 8506 4943
rect 8560 4911 8590 4943
rect 8644 4911 8674 4943
rect 8728 4911 8758 4943
rect 8812 4911 8842 4943
rect 8896 4911 8926 4943
rect 20852 4913 20882 4945
rect 20936 4913 20966 4945
rect 21020 4913 21050 4945
rect 21104 4913 21134 4945
rect 21188 4913 21218 4945
rect 21272 4913 21302 4945
rect 21356 4913 21386 4945
rect 21440 4913 21470 4945
rect 21524 4913 21554 4945
rect 21608 4913 21638 4945
rect 21692 4913 21722 4945
rect 21776 4913 21806 4945
rect 21860 4913 21890 4945
rect 21944 4913 21974 4945
rect 22028 4913 22058 4945
rect 22112 4913 22142 4945
rect 37838 5143 37868 5169
rect 37922 5143 37952 5169
rect 38006 5143 38036 5169
rect 38090 5143 38120 5169
rect 38174 5143 38204 5169
rect 38258 5143 38288 5169
rect 38342 5143 38372 5169
rect 38426 5143 38456 5169
rect 38510 5143 38540 5169
rect 38594 5143 38624 5169
rect 38678 5143 38708 5169
rect 38762 5143 38792 5169
rect 38846 5143 38876 5169
rect 38930 5143 38960 5169
rect 39014 5143 39044 5169
rect 39098 5143 39128 5169
rect 51054 5145 51084 5171
rect 51138 5145 51168 5171
rect 51222 5145 51252 5171
rect 51306 5145 51336 5171
rect 51390 5145 51420 5171
rect 51474 5145 51504 5171
rect 51558 5145 51588 5171
rect 51642 5145 51672 5171
rect 51726 5145 51756 5171
rect 51810 5145 51840 5171
rect 51894 5145 51924 5171
rect 51978 5145 52008 5171
rect 52062 5145 52092 5171
rect 52146 5145 52176 5171
rect 52230 5145 52260 5171
rect 52314 5145 52344 5171
rect 7636 4895 8992 4911
rect 7636 4861 7929 4895
rect 7963 4861 8096 4895
rect 8130 4861 8264 4895
rect 8298 4861 8431 4895
rect 8465 4861 8600 4895
rect 8634 4861 8768 4895
rect 8802 4861 8942 4895
rect 8976 4861 8992 4895
rect 5754 4825 5784 4847
rect 5838 4825 5868 4847
rect 5922 4825 5952 4847
rect 6006 4825 6036 4847
rect 6090 4825 6120 4847
rect 6174 4825 6204 4847
rect 6258 4825 6288 4847
rect 6342 4825 6372 4847
rect 6426 4825 6456 4847
rect 6510 4825 6540 4847
rect 6594 4825 6624 4847
rect 6678 4825 6708 4847
rect 6762 4825 6792 4847
rect 6846 4825 6876 4847
rect 6930 4825 6960 4847
rect 7014 4825 7044 4847
rect 7636 4845 8992 4861
rect 20852 4897 22208 4913
rect 20852 4863 21145 4897
rect 21179 4863 21312 4897
rect 21346 4863 21480 4897
rect 21514 4863 21647 4897
rect 21681 4863 21816 4897
rect 21850 4863 21984 4897
rect 22018 4863 22158 4897
rect 22192 4863 22208 4897
rect 20852 4847 22208 4863
rect 22734 4911 22764 4943
rect 22818 4911 22848 4943
rect 22902 4911 22932 4943
rect 22986 4911 23016 4943
rect 23070 4911 23100 4943
rect 23154 4911 23184 4943
rect 23238 4911 23268 4943
rect 23322 4911 23352 4943
rect 23406 4911 23436 4943
rect 23490 4911 23520 4943
rect 23574 4911 23604 4943
rect 23658 4911 23688 4943
rect 23742 4911 23772 4943
rect 23826 4911 23856 4943
rect 23910 4911 23940 4943
rect 23994 4911 24024 4943
rect 35956 4913 35986 4945
rect 36040 4913 36070 4945
rect 36124 4913 36154 4945
rect 36208 4913 36238 4945
rect 36292 4913 36322 4945
rect 36376 4913 36406 4945
rect 36460 4913 36490 4945
rect 36544 4913 36574 4945
rect 36628 4913 36658 4945
rect 36712 4913 36742 4945
rect 36796 4913 36826 4945
rect 36880 4913 36910 4945
rect 36964 4913 36994 4945
rect 37048 4913 37078 4945
rect 37132 4913 37162 4945
rect 37216 4913 37246 4945
rect 52936 5143 52966 5169
rect 53020 5143 53050 5169
rect 53104 5143 53134 5169
rect 53188 5143 53218 5169
rect 53272 5143 53302 5169
rect 53356 5143 53386 5169
rect 53440 5143 53470 5169
rect 53524 5143 53554 5169
rect 53608 5143 53638 5169
rect 53692 5143 53722 5169
rect 53776 5143 53806 5169
rect 53860 5143 53890 5169
rect 53944 5143 53974 5169
rect 54028 5143 54058 5169
rect 54112 5143 54142 5169
rect 54196 5143 54226 5169
rect 22734 4895 24090 4911
rect 22734 4861 23027 4895
rect 23061 4861 23194 4895
rect 23228 4861 23362 4895
rect 23396 4861 23529 4895
rect 23563 4861 23698 4895
rect 23732 4861 23866 4895
rect 23900 4861 24040 4895
rect 24074 4861 24090 4895
rect 7636 4823 7666 4845
rect 7720 4823 7750 4845
rect 7804 4823 7834 4845
rect 7888 4823 7918 4845
rect 7972 4823 8002 4845
rect 8056 4823 8086 4845
rect 8140 4823 8170 4845
rect 8224 4823 8254 4845
rect 8308 4823 8338 4845
rect 8392 4823 8422 4845
rect 8476 4823 8506 4845
rect 8560 4823 8590 4845
rect 8644 4823 8674 4845
rect 8728 4823 8758 4845
rect 8812 4823 8842 4845
rect 8896 4823 8926 4845
rect 20852 4825 20882 4847
rect 20936 4825 20966 4847
rect 21020 4825 21050 4847
rect 21104 4825 21134 4847
rect 21188 4825 21218 4847
rect 21272 4825 21302 4847
rect 21356 4825 21386 4847
rect 21440 4825 21470 4847
rect 21524 4825 21554 4847
rect 21608 4825 21638 4847
rect 21692 4825 21722 4847
rect 21776 4825 21806 4847
rect 21860 4825 21890 4847
rect 21944 4825 21974 4847
rect 22028 4825 22058 4847
rect 22112 4825 22142 4847
rect 22734 4845 24090 4861
rect 35956 4897 37312 4913
rect 35956 4863 36249 4897
rect 36283 4863 36416 4897
rect 36450 4863 36584 4897
rect 36618 4863 36751 4897
rect 36785 4863 36920 4897
rect 36954 4863 37088 4897
rect 37122 4863 37262 4897
rect 37296 4863 37312 4897
rect 35956 4847 37312 4863
rect 37838 4911 37868 4943
rect 37922 4911 37952 4943
rect 38006 4911 38036 4943
rect 38090 4911 38120 4943
rect 38174 4911 38204 4943
rect 38258 4911 38288 4943
rect 38342 4911 38372 4943
rect 38426 4911 38456 4943
rect 38510 4911 38540 4943
rect 38594 4911 38624 4943
rect 38678 4911 38708 4943
rect 38762 4911 38792 4943
rect 38846 4911 38876 4943
rect 38930 4911 38960 4943
rect 39014 4911 39044 4943
rect 39098 4911 39128 4943
rect 51054 4913 51084 4945
rect 51138 4913 51168 4945
rect 51222 4913 51252 4945
rect 51306 4913 51336 4945
rect 51390 4913 51420 4945
rect 51474 4913 51504 4945
rect 51558 4913 51588 4945
rect 51642 4913 51672 4945
rect 51726 4913 51756 4945
rect 51810 4913 51840 4945
rect 51894 4913 51924 4945
rect 51978 4913 52008 4945
rect 52062 4913 52092 4945
rect 52146 4913 52176 4945
rect 52230 4913 52260 4945
rect 52314 4913 52344 4945
rect 37838 4895 39194 4911
rect 37838 4861 38131 4895
rect 38165 4861 38298 4895
rect 38332 4861 38466 4895
rect 38500 4861 38633 4895
rect 38667 4861 38802 4895
rect 38836 4861 38970 4895
rect 39004 4861 39144 4895
rect 39178 4861 39194 4895
rect 5754 4669 5784 4695
rect 5838 4669 5868 4695
rect 5922 4669 5952 4695
rect 6006 4669 6036 4695
rect 6090 4669 6120 4695
rect 6174 4669 6204 4695
rect 6258 4669 6288 4695
rect 6342 4669 6372 4695
rect 6426 4669 6456 4695
rect 6510 4669 6540 4695
rect 6594 4669 6624 4695
rect 6678 4669 6708 4695
rect 6762 4669 6792 4695
rect 6846 4669 6876 4695
rect 6930 4669 6960 4695
rect 7014 4669 7044 4695
rect 22734 4823 22764 4845
rect 22818 4823 22848 4845
rect 22902 4823 22932 4845
rect 22986 4823 23016 4845
rect 23070 4823 23100 4845
rect 23154 4823 23184 4845
rect 23238 4823 23268 4845
rect 23322 4823 23352 4845
rect 23406 4823 23436 4845
rect 23490 4823 23520 4845
rect 23574 4823 23604 4845
rect 23658 4823 23688 4845
rect 23742 4823 23772 4845
rect 23826 4823 23856 4845
rect 23910 4823 23940 4845
rect 23994 4823 24024 4845
rect 35956 4825 35986 4847
rect 36040 4825 36070 4847
rect 36124 4825 36154 4847
rect 36208 4825 36238 4847
rect 36292 4825 36322 4847
rect 36376 4825 36406 4847
rect 36460 4825 36490 4847
rect 36544 4825 36574 4847
rect 36628 4825 36658 4847
rect 36712 4825 36742 4847
rect 36796 4825 36826 4847
rect 36880 4825 36910 4847
rect 36964 4825 36994 4847
rect 37048 4825 37078 4847
rect 37132 4825 37162 4847
rect 37216 4825 37246 4847
rect 37838 4845 39194 4861
rect 51054 4897 52410 4913
rect 51054 4863 51347 4897
rect 51381 4863 51514 4897
rect 51548 4863 51682 4897
rect 51716 4863 51849 4897
rect 51883 4863 52018 4897
rect 52052 4863 52186 4897
rect 52220 4863 52360 4897
rect 52394 4863 52410 4897
rect 51054 4847 52410 4863
rect 52936 4911 52966 4943
rect 53020 4911 53050 4943
rect 53104 4911 53134 4943
rect 53188 4911 53218 4943
rect 53272 4911 53302 4943
rect 53356 4911 53386 4943
rect 53440 4911 53470 4943
rect 53524 4911 53554 4943
rect 53608 4911 53638 4943
rect 53692 4911 53722 4943
rect 53776 4911 53806 4943
rect 53860 4911 53890 4943
rect 53944 4911 53974 4943
rect 54028 4911 54058 4943
rect 54112 4911 54142 4943
rect 54196 4911 54226 4943
rect 52936 4895 54292 4911
rect 52936 4861 53229 4895
rect 53263 4861 53396 4895
rect 53430 4861 53564 4895
rect 53598 4861 53731 4895
rect 53765 4861 53900 4895
rect 53934 4861 54068 4895
rect 54102 4861 54242 4895
rect 54276 4861 54292 4895
rect 7636 4667 7666 4693
rect 7720 4667 7750 4693
rect 7804 4667 7834 4693
rect 7888 4667 7918 4693
rect 7972 4667 8002 4693
rect 8056 4667 8086 4693
rect 8140 4667 8170 4693
rect 8224 4667 8254 4693
rect 8308 4667 8338 4693
rect 8392 4667 8422 4693
rect 8476 4667 8506 4693
rect 8560 4667 8590 4693
rect 8644 4667 8674 4693
rect 8728 4667 8758 4693
rect 8812 4667 8842 4693
rect 8896 4667 8926 4693
rect 20852 4669 20882 4695
rect 20936 4669 20966 4695
rect 21020 4669 21050 4695
rect 21104 4669 21134 4695
rect 21188 4669 21218 4695
rect 21272 4669 21302 4695
rect 21356 4669 21386 4695
rect 21440 4669 21470 4695
rect 21524 4669 21554 4695
rect 21608 4669 21638 4695
rect 21692 4669 21722 4695
rect 21776 4669 21806 4695
rect 21860 4669 21890 4695
rect 21944 4669 21974 4695
rect 22028 4669 22058 4695
rect 22112 4669 22142 4695
rect 37838 4823 37868 4845
rect 37922 4823 37952 4845
rect 38006 4823 38036 4845
rect 38090 4823 38120 4845
rect 38174 4823 38204 4845
rect 38258 4823 38288 4845
rect 38342 4823 38372 4845
rect 38426 4823 38456 4845
rect 38510 4823 38540 4845
rect 38594 4823 38624 4845
rect 38678 4823 38708 4845
rect 38762 4823 38792 4845
rect 38846 4823 38876 4845
rect 38930 4823 38960 4845
rect 39014 4823 39044 4845
rect 39098 4823 39128 4845
rect 51054 4825 51084 4847
rect 51138 4825 51168 4847
rect 51222 4825 51252 4847
rect 51306 4825 51336 4847
rect 51390 4825 51420 4847
rect 51474 4825 51504 4847
rect 51558 4825 51588 4847
rect 51642 4825 51672 4847
rect 51726 4825 51756 4847
rect 51810 4825 51840 4847
rect 51894 4825 51924 4847
rect 51978 4825 52008 4847
rect 52062 4825 52092 4847
rect 52146 4825 52176 4847
rect 52230 4825 52260 4847
rect 52314 4825 52344 4847
rect 52936 4845 54292 4861
rect 22734 4667 22764 4693
rect 22818 4667 22848 4693
rect 22902 4667 22932 4693
rect 22986 4667 23016 4693
rect 23070 4667 23100 4693
rect 23154 4667 23184 4693
rect 23238 4667 23268 4693
rect 23322 4667 23352 4693
rect 23406 4667 23436 4693
rect 23490 4667 23520 4693
rect 23574 4667 23604 4693
rect 23658 4667 23688 4693
rect 23742 4667 23772 4693
rect 23826 4667 23856 4693
rect 23910 4667 23940 4693
rect 23994 4667 24024 4693
rect 35956 4669 35986 4695
rect 36040 4669 36070 4695
rect 36124 4669 36154 4695
rect 36208 4669 36238 4695
rect 36292 4669 36322 4695
rect 36376 4669 36406 4695
rect 36460 4669 36490 4695
rect 36544 4669 36574 4695
rect 36628 4669 36658 4695
rect 36712 4669 36742 4695
rect 36796 4669 36826 4695
rect 36880 4669 36910 4695
rect 36964 4669 36994 4695
rect 37048 4669 37078 4695
rect 37132 4669 37162 4695
rect 37216 4669 37246 4695
rect 52936 4823 52966 4845
rect 53020 4823 53050 4845
rect 53104 4823 53134 4845
rect 53188 4823 53218 4845
rect 53272 4823 53302 4845
rect 53356 4823 53386 4845
rect 53440 4823 53470 4845
rect 53524 4823 53554 4845
rect 53608 4823 53638 4845
rect 53692 4823 53722 4845
rect 53776 4823 53806 4845
rect 53860 4823 53890 4845
rect 53944 4823 53974 4845
rect 54028 4823 54058 4845
rect 54112 4823 54142 4845
rect 54196 4823 54226 4845
rect 37838 4667 37868 4693
rect 37922 4667 37952 4693
rect 38006 4667 38036 4693
rect 38090 4667 38120 4693
rect 38174 4667 38204 4693
rect 38258 4667 38288 4693
rect 38342 4667 38372 4693
rect 38426 4667 38456 4693
rect 38510 4667 38540 4693
rect 38594 4667 38624 4693
rect 38678 4667 38708 4693
rect 38762 4667 38792 4693
rect 38846 4667 38876 4693
rect 38930 4667 38960 4693
rect 39014 4667 39044 4693
rect 39098 4667 39128 4693
rect 51054 4669 51084 4695
rect 51138 4669 51168 4695
rect 51222 4669 51252 4695
rect 51306 4669 51336 4695
rect 51390 4669 51420 4695
rect 51474 4669 51504 4695
rect 51558 4669 51588 4695
rect 51642 4669 51672 4695
rect 51726 4669 51756 4695
rect 51810 4669 51840 4695
rect 51894 4669 51924 4695
rect 51978 4669 52008 4695
rect 52062 4669 52092 4695
rect 52146 4669 52176 4695
rect 52230 4669 52260 4695
rect 52314 4669 52344 4695
rect 52936 4667 52966 4693
rect 53020 4667 53050 4693
rect 53104 4667 53134 4693
rect 53188 4667 53218 4693
rect 53272 4667 53302 4693
rect 53356 4667 53386 4693
rect 53440 4667 53470 4693
rect 53524 4667 53554 4693
rect 53608 4667 53638 4693
rect 53692 4667 53722 4693
rect 53776 4667 53806 4693
rect 53860 4667 53890 4693
rect 53944 4667 53974 4693
rect 54028 4667 54058 4693
rect 54112 4667 54142 4693
rect 54196 4667 54226 4693
rect 30116 4068 30146 4094
rect 30200 4068 30230 4094
rect 30284 4068 30314 4094
rect 30368 4068 30398 4094
rect 30647 4068 30677 4094
rect 30731 4068 30761 4094
rect 30815 4068 30845 4094
rect 30899 4068 30929 4094
rect 30983 4068 31013 4094
rect 31067 4068 31097 4094
rect 31151 4068 31181 4094
rect 31235 4068 31265 4094
rect 31319 4068 31349 4094
rect 31403 4068 31433 4094
rect 31487 4068 31517 4094
rect 31571 4068 31601 4094
rect 31655 4068 31685 4094
rect 31739 4068 31769 4094
rect 31823 4068 31853 4094
rect 31907 4068 31937 4094
rect 30116 3836 30146 3868
rect 30200 3836 30230 3868
rect 30284 3836 30314 3868
rect 30368 3836 30398 3868
rect 30647 3836 30677 3868
rect 30731 3836 30761 3868
rect 30815 3836 30845 3868
rect 30899 3836 30929 3868
rect 30983 3836 31013 3868
rect 31067 3836 31097 3868
rect 31151 3836 31181 3868
rect 31235 3836 31265 3868
rect 31319 3836 31349 3868
rect 31403 3836 31433 3868
rect 31487 3836 31517 3868
rect 31571 3836 31601 3868
rect 31655 3836 31685 3868
rect 31739 3836 31769 3868
rect 31823 3836 31853 3868
rect 31907 3836 31937 3868
rect 43473 3852 43503 3878
rect 43557 3852 43587 3878
rect 43641 3852 43671 3878
rect 43725 3852 43755 3878
rect 43809 3852 43839 3878
rect 43893 3852 43923 3878
rect 43977 3852 44007 3878
rect 44061 3852 44091 3878
rect 44145 3852 44175 3878
rect 44229 3852 44259 3878
rect 44313 3852 44343 3878
rect 44397 3852 44427 3878
rect 44481 3852 44511 3878
rect 44565 3852 44595 3878
rect 44649 3852 44679 3878
rect 44733 3852 44763 3878
rect 45403 3852 45433 3878
rect 45487 3852 45517 3878
rect 45571 3852 45601 3878
rect 45655 3852 45685 3878
rect 45739 3852 45769 3878
rect 45823 3852 45853 3878
rect 45907 3852 45937 3878
rect 45991 3852 46021 3878
rect 46075 3852 46105 3878
rect 46159 3852 46189 3878
rect 46243 3852 46273 3878
rect 46327 3852 46357 3878
rect 46411 3852 46441 3878
rect 46495 3852 46525 3878
rect 46579 3852 46609 3878
rect 46663 3852 46693 3878
rect 30048 3820 30398 3836
rect 30048 3786 30064 3820
rect 30098 3786 30156 3820
rect 30190 3786 30240 3820
rect 30274 3786 30324 3820
rect 30358 3786 30398 3820
rect 30048 3770 30398 3786
rect 30581 3820 31937 3836
rect 30581 3786 30597 3820
rect 30631 3786 30771 3820
rect 30805 3786 30939 3820
rect 30973 3786 31108 3820
rect 31142 3786 31275 3820
rect 31309 3786 31443 3820
rect 31477 3786 31610 3820
rect 31644 3786 31937 3820
rect 30581 3770 31937 3786
rect 30116 3748 30146 3770
rect 30200 3748 30230 3770
rect 30284 3748 30314 3770
rect 30368 3748 30398 3770
rect 30647 3748 30677 3770
rect 30731 3748 30761 3770
rect 30815 3748 30845 3770
rect 30899 3748 30929 3770
rect 30983 3748 31013 3770
rect 31067 3748 31097 3770
rect 31151 3748 31181 3770
rect 31235 3748 31265 3770
rect 31319 3748 31349 3770
rect 31403 3748 31433 3770
rect 31487 3748 31517 3770
rect 31571 3748 31601 3770
rect 31655 3748 31685 3770
rect 31739 3748 31769 3770
rect 31823 3748 31853 3770
rect 31907 3748 31937 3770
rect 13331 3692 13361 3718
rect 13415 3692 13445 3718
rect 13499 3692 13529 3718
rect 13583 3692 13613 3718
rect 13667 3692 13697 3718
rect 13751 3692 13781 3718
rect 13835 3692 13865 3718
rect 13919 3692 13949 3718
rect 14003 3692 14033 3718
rect 14087 3692 14117 3718
rect 14171 3692 14201 3718
rect 14255 3692 14285 3718
rect 14339 3692 14369 3718
rect 14423 3692 14453 3718
rect 14507 3692 14537 3718
rect 14591 3692 14621 3718
rect 15261 3692 15291 3718
rect 15345 3692 15375 3718
rect 15429 3692 15459 3718
rect 15513 3692 15543 3718
rect 15597 3692 15627 3718
rect 15681 3692 15711 3718
rect 15765 3692 15795 3718
rect 15849 3692 15879 3718
rect 15933 3692 15963 3718
rect 16017 3692 16047 3718
rect 16101 3692 16131 3718
rect 16185 3692 16215 3718
rect 16269 3692 16299 3718
rect 16353 3692 16383 3718
rect 16437 3692 16467 3718
rect 16521 3692 16551 3718
rect 43473 3620 43503 3652
rect 43557 3620 43587 3652
rect 43641 3620 43671 3652
rect 43725 3620 43755 3652
rect 43809 3620 43839 3652
rect 43893 3620 43923 3652
rect 43977 3620 44007 3652
rect 44061 3620 44091 3652
rect 44145 3620 44175 3652
rect 44229 3620 44259 3652
rect 44313 3620 44343 3652
rect 44397 3620 44427 3652
rect 44481 3620 44511 3652
rect 44565 3620 44595 3652
rect 44649 3620 44679 3652
rect 44733 3620 44763 3652
rect 45403 3620 45433 3652
rect 45487 3620 45517 3652
rect 45571 3620 45601 3652
rect 45655 3620 45685 3652
rect 45739 3620 45769 3652
rect 45823 3620 45853 3652
rect 45907 3620 45937 3652
rect 45991 3620 46021 3652
rect 46075 3620 46105 3652
rect 46159 3620 46189 3652
rect 46243 3620 46273 3652
rect 46327 3620 46357 3652
rect 46411 3620 46441 3652
rect 46495 3620 46525 3652
rect 46579 3620 46609 3652
rect 46663 3620 46693 3652
rect 30116 3592 30146 3618
rect 30200 3592 30230 3618
rect 30284 3592 30314 3618
rect 30368 3592 30398 3618
rect 30647 3592 30677 3618
rect 30731 3592 30761 3618
rect 30815 3592 30845 3618
rect 30899 3592 30929 3618
rect 30983 3592 31013 3618
rect 31067 3592 31097 3618
rect 31151 3592 31181 3618
rect 31235 3592 31265 3618
rect 31319 3592 31349 3618
rect 31403 3592 31433 3618
rect 31487 3592 31517 3618
rect 31571 3592 31601 3618
rect 31655 3592 31685 3618
rect 31739 3592 31769 3618
rect 31823 3592 31853 3618
rect 31907 3592 31937 3618
rect 43407 3604 44763 3620
rect 43407 3570 43423 3604
rect 43457 3570 43597 3604
rect 43631 3570 43765 3604
rect 43799 3570 43934 3604
rect 43968 3570 44101 3604
rect 44135 3570 44269 3604
rect 44303 3570 44436 3604
rect 44470 3570 44763 3604
rect 43407 3554 44763 3570
rect 45337 3604 46693 3620
rect 45337 3570 45353 3604
rect 45387 3570 45527 3604
rect 45561 3570 45695 3604
rect 45729 3570 45864 3604
rect 45898 3570 46031 3604
rect 46065 3570 46199 3604
rect 46233 3570 46366 3604
rect 46400 3570 46693 3604
rect 45337 3554 46693 3570
rect 43473 3532 43503 3554
rect 43557 3532 43587 3554
rect 43641 3532 43671 3554
rect 43725 3532 43755 3554
rect 43809 3532 43839 3554
rect 43893 3532 43923 3554
rect 43977 3532 44007 3554
rect 44061 3532 44091 3554
rect 44145 3532 44175 3554
rect 44229 3532 44259 3554
rect 44313 3532 44343 3554
rect 44397 3532 44427 3554
rect 44481 3532 44511 3554
rect 44565 3532 44595 3554
rect 44649 3532 44679 3554
rect 44733 3532 44763 3554
rect 45403 3532 45433 3554
rect 45487 3532 45517 3554
rect 45571 3532 45601 3554
rect 45655 3532 45685 3554
rect 45739 3532 45769 3554
rect 45823 3532 45853 3554
rect 45907 3532 45937 3554
rect 45991 3532 46021 3554
rect 46075 3532 46105 3554
rect 46159 3532 46189 3554
rect 46243 3532 46273 3554
rect 46327 3532 46357 3554
rect 46411 3532 46441 3554
rect 46495 3532 46525 3554
rect 46579 3532 46609 3554
rect 46663 3532 46693 3554
rect 13331 3460 13361 3492
rect 13415 3460 13445 3492
rect 13499 3460 13529 3492
rect 13583 3460 13613 3492
rect 13667 3460 13697 3492
rect 13751 3460 13781 3492
rect 13835 3460 13865 3492
rect 13919 3460 13949 3492
rect 14003 3460 14033 3492
rect 14087 3460 14117 3492
rect 14171 3460 14201 3492
rect 14255 3460 14285 3492
rect 14339 3460 14369 3492
rect 14423 3460 14453 3492
rect 14507 3460 14537 3492
rect 14591 3460 14621 3492
rect 15261 3460 15291 3492
rect 15345 3460 15375 3492
rect 15429 3460 15459 3492
rect 15513 3460 15543 3492
rect 15597 3460 15627 3492
rect 15681 3460 15711 3492
rect 15765 3460 15795 3492
rect 15849 3460 15879 3492
rect 15933 3460 15963 3492
rect 16017 3460 16047 3492
rect 16101 3460 16131 3492
rect 16185 3460 16215 3492
rect 16269 3460 16299 3492
rect 16353 3460 16383 3492
rect 16437 3460 16467 3492
rect 16521 3460 16551 3492
rect 13265 3444 14621 3460
rect 13265 3410 13281 3444
rect 13315 3410 13455 3444
rect 13489 3410 13623 3444
rect 13657 3410 13792 3444
rect 13826 3410 13959 3444
rect 13993 3410 14127 3444
rect 14161 3410 14294 3444
rect 14328 3410 14621 3444
rect 13265 3394 14621 3410
rect 15195 3444 16551 3460
rect 15195 3410 15211 3444
rect 15245 3410 15385 3444
rect 15419 3410 15553 3444
rect 15587 3410 15722 3444
rect 15756 3410 15889 3444
rect 15923 3410 16057 3444
rect 16091 3410 16224 3444
rect 16258 3410 16551 3444
rect 15195 3394 16551 3410
rect 13331 3372 13361 3394
rect 13415 3372 13445 3394
rect 13499 3372 13529 3394
rect 13583 3372 13613 3394
rect 13667 3372 13697 3394
rect 13751 3372 13781 3394
rect 13835 3372 13865 3394
rect 13919 3372 13949 3394
rect 14003 3372 14033 3394
rect 14087 3372 14117 3394
rect 14171 3372 14201 3394
rect 14255 3372 14285 3394
rect 14339 3372 14369 3394
rect 14423 3372 14453 3394
rect 14507 3372 14537 3394
rect 14591 3372 14621 3394
rect 15261 3372 15291 3394
rect 15345 3372 15375 3394
rect 15429 3372 15459 3394
rect 15513 3372 15543 3394
rect 15597 3372 15627 3394
rect 15681 3372 15711 3394
rect 15765 3372 15795 3394
rect 15849 3372 15879 3394
rect 15933 3372 15963 3394
rect 16017 3372 16047 3394
rect 16101 3372 16131 3394
rect 16185 3372 16215 3394
rect 16269 3372 16299 3394
rect 16353 3372 16383 3394
rect 16437 3372 16467 3394
rect 16521 3372 16551 3394
rect 43473 3376 43503 3402
rect 43557 3376 43587 3402
rect 43641 3376 43671 3402
rect 43725 3376 43755 3402
rect 43809 3376 43839 3402
rect 43893 3376 43923 3402
rect 43977 3376 44007 3402
rect 44061 3376 44091 3402
rect 44145 3376 44175 3402
rect 44229 3376 44259 3402
rect 44313 3376 44343 3402
rect 44397 3376 44427 3402
rect 44481 3376 44511 3402
rect 44565 3376 44595 3402
rect 44649 3376 44679 3402
rect 44733 3376 44763 3402
rect 45403 3376 45433 3402
rect 45487 3376 45517 3402
rect 45571 3376 45601 3402
rect 45655 3376 45685 3402
rect 45739 3376 45769 3402
rect 45823 3376 45853 3402
rect 45907 3376 45937 3402
rect 45991 3376 46021 3402
rect 46075 3376 46105 3402
rect 46159 3376 46189 3402
rect 46243 3376 46273 3402
rect 46327 3376 46357 3402
rect 46411 3376 46441 3402
rect 46495 3376 46525 3402
rect 46579 3376 46609 3402
rect 46663 3376 46693 3402
rect 13331 3216 13361 3242
rect 13415 3216 13445 3242
rect 13499 3216 13529 3242
rect 13583 3216 13613 3242
rect 13667 3216 13697 3242
rect 13751 3216 13781 3242
rect 13835 3216 13865 3242
rect 13919 3216 13949 3242
rect 14003 3216 14033 3242
rect 14087 3216 14117 3242
rect 14171 3216 14201 3242
rect 14255 3216 14285 3242
rect 14339 3216 14369 3242
rect 14423 3216 14453 3242
rect 14507 3216 14537 3242
rect 14591 3216 14621 3242
rect 15261 3216 15291 3242
rect 15345 3216 15375 3242
rect 15429 3216 15459 3242
rect 15513 3216 15543 3242
rect 15597 3216 15627 3242
rect 15681 3216 15711 3242
rect 15765 3216 15795 3242
rect 15849 3216 15879 3242
rect 15933 3216 15963 3242
rect 16017 3216 16047 3242
rect 16101 3216 16131 3242
rect 16185 3216 16215 3242
rect 16269 3216 16299 3242
rect 16353 3216 16383 3242
rect 16437 3216 16467 3242
rect 16521 3216 16551 3242
rect 5756 2747 5786 2773
rect 5840 2747 5870 2773
rect 5924 2747 5954 2773
rect 6008 2747 6038 2773
rect 6092 2747 6122 2773
rect 6176 2747 6206 2773
rect 6260 2747 6290 2773
rect 6344 2747 6374 2773
rect 6428 2747 6458 2773
rect 6512 2747 6542 2773
rect 6596 2747 6626 2773
rect 6680 2747 6710 2773
rect 6764 2747 6794 2773
rect 6848 2747 6878 2773
rect 6932 2747 6962 2773
rect 7016 2747 7046 2773
rect 7638 2745 7668 2771
rect 7722 2745 7752 2771
rect 7806 2745 7836 2771
rect 7890 2745 7920 2771
rect 7974 2745 8004 2771
rect 8058 2745 8088 2771
rect 8142 2745 8172 2771
rect 8226 2745 8256 2771
rect 8310 2745 8340 2771
rect 8394 2745 8424 2771
rect 8478 2745 8508 2771
rect 8562 2745 8592 2771
rect 8646 2745 8676 2771
rect 8730 2745 8760 2771
rect 8814 2745 8844 2771
rect 8898 2745 8928 2771
rect 20854 2747 20884 2773
rect 20938 2747 20968 2773
rect 21022 2747 21052 2773
rect 21106 2747 21136 2773
rect 21190 2747 21220 2773
rect 21274 2747 21304 2773
rect 21358 2747 21388 2773
rect 21442 2747 21472 2773
rect 21526 2747 21556 2773
rect 21610 2747 21640 2773
rect 21694 2747 21724 2773
rect 21778 2747 21808 2773
rect 21862 2747 21892 2773
rect 21946 2747 21976 2773
rect 22030 2747 22060 2773
rect 22114 2747 22144 2773
rect 5756 2595 5786 2617
rect 5840 2595 5870 2617
rect 5924 2595 5954 2617
rect 6008 2595 6038 2617
rect 6092 2595 6122 2617
rect 6176 2595 6206 2617
rect 6260 2595 6290 2617
rect 6344 2595 6374 2617
rect 6428 2595 6458 2617
rect 6512 2595 6542 2617
rect 6596 2595 6626 2617
rect 6680 2595 6710 2617
rect 6764 2595 6794 2617
rect 6848 2595 6878 2617
rect 6932 2595 6962 2617
rect 7016 2595 7046 2617
rect 22736 2745 22766 2771
rect 22820 2745 22850 2771
rect 22904 2745 22934 2771
rect 22988 2745 23018 2771
rect 23072 2745 23102 2771
rect 23156 2745 23186 2771
rect 23240 2745 23270 2771
rect 23324 2745 23354 2771
rect 23408 2745 23438 2771
rect 23492 2745 23522 2771
rect 23576 2745 23606 2771
rect 23660 2745 23690 2771
rect 23744 2745 23774 2771
rect 23828 2745 23858 2771
rect 23912 2745 23942 2771
rect 23996 2745 24026 2771
rect 35958 2747 35988 2773
rect 36042 2747 36072 2773
rect 36126 2747 36156 2773
rect 36210 2747 36240 2773
rect 36294 2747 36324 2773
rect 36378 2747 36408 2773
rect 36462 2747 36492 2773
rect 36546 2747 36576 2773
rect 36630 2747 36660 2773
rect 36714 2747 36744 2773
rect 36798 2747 36828 2773
rect 36882 2747 36912 2773
rect 36966 2747 36996 2773
rect 37050 2747 37080 2773
rect 37134 2747 37164 2773
rect 37218 2747 37248 2773
rect 5690 2579 7046 2595
rect 7638 2593 7668 2615
rect 7722 2593 7752 2615
rect 7806 2593 7836 2615
rect 7890 2593 7920 2615
rect 7974 2593 8004 2615
rect 8058 2593 8088 2615
rect 8142 2593 8172 2615
rect 8226 2593 8256 2615
rect 8310 2593 8340 2615
rect 8394 2593 8424 2615
rect 8478 2593 8508 2615
rect 8562 2593 8592 2615
rect 8646 2593 8676 2615
rect 8730 2593 8760 2615
rect 8814 2593 8844 2615
rect 8898 2593 8928 2615
rect 20854 2595 20884 2617
rect 20938 2595 20968 2617
rect 21022 2595 21052 2617
rect 21106 2595 21136 2617
rect 21190 2595 21220 2617
rect 21274 2595 21304 2617
rect 21358 2595 21388 2617
rect 21442 2595 21472 2617
rect 21526 2595 21556 2617
rect 21610 2595 21640 2617
rect 21694 2595 21724 2617
rect 21778 2595 21808 2617
rect 21862 2595 21892 2617
rect 21946 2595 21976 2617
rect 22030 2595 22060 2617
rect 22114 2595 22144 2617
rect 37840 2745 37870 2771
rect 37924 2745 37954 2771
rect 38008 2745 38038 2771
rect 38092 2745 38122 2771
rect 38176 2745 38206 2771
rect 38260 2745 38290 2771
rect 38344 2745 38374 2771
rect 38428 2745 38458 2771
rect 38512 2745 38542 2771
rect 38596 2745 38626 2771
rect 38680 2745 38710 2771
rect 38764 2745 38794 2771
rect 38848 2745 38878 2771
rect 38932 2745 38962 2771
rect 39016 2745 39046 2771
rect 39100 2745 39130 2771
rect 51056 2747 51086 2773
rect 51140 2747 51170 2773
rect 51224 2747 51254 2773
rect 51308 2747 51338 2773
rect 51392 2747 51422 2773
rect 51476 2747 51506 2773
rect 51560 2747 51590 2773
rect 51644 2747 51674 2773
rect 51728 2747 51758 2773
rect 51812 2747 51842 2773
rect 51896 2747 51926 2773
rect 51980 2747 52010 2773
rect 52064 2747 52094 2773
rect 52148 2747 52178 2773
rect 52232 2747 52262 2773
rect 52316 2747 52346 2773
rect 5690 2545 5706 2579
rect 5740 2545 5880 2579
rect 5914 2545 6048 2579
rect 6082 2545 6217 2579
rect 6251 2545 6384 2579
rect 6418 2545 6552 2579
rect 6586 2545 6719 2579
rect 6753 2545 7046 2579
rect 5690 2529 7046 2545
rect 5756 2497 5786 2529
rect 5840 2497 5870 2529
rect 5924 2497 5954 2529
rect 6008 2497 6038 2529
rect 6092 2497 6122 2529
rect 6176 2497 6206 2529
rect 6260 2497 6290 2529
rect 6344 2497 6374 2529
rect 6428 2497 6458 2529
rect 6512 2497 6542 2529
rect 6596 2497 6626 2529
rect 6680 2497 6710 2529
rect 6764 2497 6794 2529
rect 6848 2497 6878 2529
rect 6932 2497 6962 2529
rect 7016 2497 7046 2529
rect 7572 2577 8928 2593
rect 7572 2543 7588 2577
rect 7622 2543 7762 2577
rect 7796 2543 7930 2577
rect 7964 2543 8099 2577
rect 8133 2543 8266 2577
rect 8300 2543 8434 2577
rect 8468 2543 8601 2577
rect 8635 2543 8928 2577
rect 7572 2527 8928 2543
rect 20788 2579 22144 2595
rect 22736 2593 22766 2615
rect 22820 2593 22850 2615
rect 22904 2593 22934 2615
rect 22988 2593 23018 2615
rect 23072 2593 23102 2615
rect 23156 2593 23186 2615
rect 23240 2593 23270 2615
rect 23324 2593 23354 2615
rect 23408 2593 23438 2615
rect 23492 2593 23522 2615
rect 23576 2593 23606 2615
rect 23660 2593 23690 2615
rect 23744 2593 23774 2615
rect 23828 2593 23858 2615
rect 23912 2593 23942 2615
rect 23996 2593 24026 2615
rect 35958 2595 35988 2617
rect 36042 2595 36072 2617
rect 36126 2595 36156 2617
rect 36210 2595 36240 2617
rect 36294 2595 36324 2617
rect 36378 2595 36408 2617
rect 36462 2595 36492 2617
rect 36546 2595 36576 2617
rect 36630 2595 36660 2617
rect 36714 2595 36744 2617
rect 36798 2595 36828 2617
rect 36882 2595 36912 2617
rect 36966 2595 36996 2617
rect 37050 2595 37080 2617
rect 37134 2595 37164 2617
rect 37218 2595 37248 2617
rect 52938 2745 52968 2771
rect 53022 2745 53052 2771
rect 53106 2745 53136 2771
rect 53190 2745 53220 2771
rect 53274 2745 53304 2771
rect 53358 2745 53388 2771
rect 53442 2745 53472 2771
rect 53526 2745 53556 2771
rect 53610 2745 53640 2771
rect 53694 2745 53724 2771
rect 53778 2745 53808 2771
rect 53862 2745 53892 2771
rect 53946 2745 53976 2771
rect 54030 2745 54060 2771
rect 54114 2745 54144 2771
rect 54198 2745 54228 2771
rect 20788 2545 20804 2579
rect 20838 2545 20978 2579
rect 21012 2545 21146 2579
rect 21180 2545 21315 2579
rect 21349 2545 21482 2579
rect 21516 2545 21650 2579
rect 21684 2545 21817 2579
rect 21851 2545 22144 2579
rect 20788 2529 22144 2545
rect 7638 2495 7668 2527
rect 7722 2495 7752 2527
rect 7806 2495 7836 2527
rect 7890 2495 7920 2527
rect 7974 2495 8004 2527
rect 8058 2495 8088 2527
rect 8142 2495 8172 2527
rect 8226 2495 8256 2527
rect 8310 2495 8340 2527
rect 8394 2495 8424 2527
rect 8478 2495 8508 2527
rect 8562 2495 8592 2527
rect 8646 2495 8676 2527
rect 8730 2495 8760 2527
rect 8814 2495 8844 2527
rect 8898 2495 8928 2527
rect 20854 2497 20884 2529
rect 20938 2497 20968 2529
rect 21022 2497 21052 2529
rect 21106 2497 21136 2529
rect 21190 2497 21220 2529
rect 21274 2497 21304 2529
rect 21358 2497 21388 2529
rect 21442 2497 21472 2529
rect 21526 2497 21556 2529
rect 21610 2497 21640 2529
rect 21694 2497 21724 2529
rect 21778 2497 21808 2529
rect 21862 2497 21892 2529
rect 21946 2497 21976 2529
rect 22030 2497 22060 2529
rect 22114 2497 22144 2529
rect 22670 2577 24026 2593
rect 22670 2543 22686 2577
rect 22720 2543 22860 2577
rect 22894 2543 23028 2577
rect 23062 2543 23197 2577
rect 23231 2543 23364 2577
rect 23398 2543 23532 2577
rect 23566 2543 23699 2577
rect 23733 2543 24026 2577
rect 22670 2527 24026 2543
rect 35892 2579 37248 2595
rect 37840 2593 37870 2615
rect 37924 2593 37954 2615
rect 38008 2593 38038 2615
rect 38092 2593 38122 2615
rect 38176 2593 38206 2615
rect 38260 2593 38290 2615
rect 38344 2593 38374 2615
rect 38428 2593 38458 2615
rect 38512 2593 38542 2615
rect 38596 2593 38626 2615
rect 38680 2593 38710 2615
rect 38764 2593 38794 2615
rect 38848 2593 38878 2615
rect 38932 2593 38962 2615
rect 39016 2593 39046 2615
rect 39100 2593 39130 2615
rect 51056 2595 51086 2617
rect 51140 2595 51170 2617
rect 51224 2595 51254 2617
rect 51308 2595 51338 2617
rect 51392 2595 51422 2617
rect 51476 2595 51506 2617
rect 51560 2595 51590 2617
rect 51644 2595 51674 2617
rect 51728 2595 51758 2617
rect 51812 2595 51842 2617
rect 51896 2595 51926 2617
rect 51980 2595 52010 2617
rect 52064 2595 52094 2617
rect 52148 2595 52178 2617
rect 52232 2595 52262 2617
rect 52316 2595 52346 2617
rect 35892 2545 35908 2579
rect 35942 2545 36082 2579
rect 36116 2545 36250 2579
rect 36284 2545 36419 2579
rect 36453 2545 36586 2579
rect 36620 2545 36754 2579
rect 36788 2545 36921 2579
rect 36955 2545 37248 2579
rect 35892 2529 37248 2545
rect 5756 2271 5786 2297
rect 5840 2271 5870 2297
rect 5924 2271 5954 2297
rect 6008 2271 6038 2297
rect 6092 2271 6122 2297
rect 6176 2271 6206 2297
rect 6260 2271 6290 2297
rect 6344 2271 6374 2297
rect 6428 2271 6458 2297
rect 6512 2271 6542 2297
rect 6596 2271 6626 2297
rect 6680 2271 6710 2297
rect 6764 2271 6794 2297
rect 6848 2271 6878 2297
rect 6932 2271 6962 2297
rect 7016 2271 7046 2297
rect 22736 2495 22766 2527
rect 22820 2495 22850 2527
rect 22904 2495 22934 2527
rect 22988 2495 23018 2527
rect 23072 2495 23102 2527
rect 23156 2495 23186 2527
rect 23240 2495 23270 2527
rect 23324 2495 23354 2527
rect 23408 2495 23438 2527
rect 23492 2495 23522 2527
rect 23576 2495 23606 2527
rect 23660 2495 23690 2527
rect 23744 2495 23774 2527
rect 23828 2495 23858 2527
rect 23912 2495 23942 2527
rect 23996 2495 24026 2527
rect 35958 2497 35988 2529
rect 36042 2497 36072 2529
rect 36126 2497 36156 2529
rect 36210 2497 36240 2529
rect 36294 2497 36324 2529
rect 36378 2497 36408 2529
rect 36462 2497 36492 2529
rect 36546 2497 36576 2529
rect 36630 2497 36660 2529
rect 36714 2497 36744 2529
rect 36798 2497 36828 2529
rect 36882 2497 36912 2529
rect 36966 2497 36996 2529
rect 37050 2497 37080 2529
rect 37134 2497 37164 2529
rect 37218 2497 37248 2529
rect 37774 2577 39130 2593
rect 37774 2543 37790 2577
rect 37824 2543 37964 2577
rect 37998 2543 38132 2577
rect 38166 2543 38301 2577
rect 38335 2543 38468 2577
rect 38502 2543 38636 2577
rect 38670 2543 38803 2577
rect 38837 2543 39130 2577
rect 37774 2527 39130 2543
rect 50990 2579 52346 2595
rect 52938 2593 52968 2615
rect 53022 2593 53052 2615
rect 53106 2593 53136 2615
rect 53190 2593 53220 2615
rect 53274 2593 53304 2615
rect 53358 2593 53388 2615
rect 53442 2593 53472 2615
rect 53526 2593 53556 2615
rect 53610 2593 53640 2615
rect 53694 2593 53724 2615
rect 53778 2593 53808 2615
rect 53862 2593 53892 2615
rect 53946 2593 53976 2615
rect 54030 2593 54060 2615
rect 54114 2593 54144 2615
rect 54198 2593 54228 2615
rect 50990 2545 51006 2579
rect 51040 2545 51180 2579
rect 51214 2545 51348 2579
rect 51382 2545 51517 2579
rect 51551 2545 51684 2579
rect 51718 2545 51852 2579
rect 51886 2545 52019 2579
rect 52053 2545 52346 2579
rect 50990 2529 52346 2545
rect 7638 2269 7668 2295
rect 7722 2269 7752 2295
rect 7806 2269 7836 2295
rect 7890 2269 7920 2295
rect 7974 2269 8004 2295
rect 8058 2269 8088 2295
rect 8142 2269 8172 2295
rect 8226 2269 8256 2295
rect 8310 2269 8340 2295
rect 8394 2269 8424 2295
rect 8478 2269 8508 2295
rect 8562 2269 8592 2295
rect 8646 2269 8676 2295
rect 8730 2269 8760 2295
rect 8814 2269 8844 2295
rect 8898 2269 8928 2295
rect 20854 2271 20884 2297
rect 20938 2271 20968 2297
rect 21022 2271 21052 2297
rect 21106 2271 21136 2297
rect 21190 2271 21220 2297
rect 21274 2271 21304 2297
rect 21358 2271 21388 2297
rect 21442 2271 21472 2297
rect 21526 2271 21556 2297
rect 21610 2271 21640 2297
rect 21694 2271 21724 2297
rect 21778 2271 21808 2297
rect 21862 2271 21892 2297
rect 21946 2271 21976 2297
rect 22030 2271 22060 2297
rect 22114 2271 22144 2297
rect 37840 2495 37870 2527
rect 37924 2495 37954 2527
rect 38008 2495 38038 2527
rect 38092 2495 38122 2527
rect 38176 2495 38206 2527
rect 38260 2495 38290 2527
rect 38344 2495 38374 2527
rect 38428 2495 38458 2527
rect 38512 2495 38542 2527
rect 38596 2495 38626 2527
rect 38680 2495 38710 2527
rect 38764 2495 38794 2527
rect 38848 2495 38878 2527
rect 38932 2495 38962 2527
rect 39016 2495 39046 2527
rect 39100 2495 39130 2527
rect 51056 2497 51086 2529
rect 51140 2497 51170 2529
rect 51224 2497 51254 2529
rect 51308 2497 51338 2529
rect 51392 2497 51422 2529
rect 51476 2497 51506 2529
rect 51560 2497 51590 2529
rect 51644 2497 51674 2529
rect 51728 2497 51758 2529
rect 51812 2497 51842 2529
rect 51896 2497 51926 2529
rect 51980 2497 52010 2529
rect 52064 2497 52094 2529
rect 52148 2497 52178 2529
rect 52232 2497 52262 2529
rect 52316 2497 52346 2529
rect 52872 2577 54228 2593
rect 52872 2543 52888 2577
rect 52922 2543 53062 2577
rect 53096 2543 53230 2577
rect 53264 2543 53399 2577
rect 53433 2543 53566 2577
rect 53600 2543 53734 2577
rect 53768 2543 53901 2577
rect 53935 2543 54228 2577
rect 52872 2527 54228 2543
rect 22736 2269 22766 2295
rect 22820 2269 22850 2295
rect 22904 2269 22934 2295
rect 22988 2269 23018 2295
rect 23072 2269 23102 2295
rect 23156 2269 23186 2295
rect 23240 2269 23270 2295
rect 23324 2269 23354 2295
rect 23408 2269 23438 2295
rect 23492 2269 23522 2295
rect 23576 2269 23606 2295
rect 23660 2269 23690 2295
rect 23744 2269 23774 2295
rect 23828 2269 23858 2295
rect 23912 2269 23942 2295
rect 23996 2269 24026 2295
rect 35958 2271 35988 2297
rect 36042 2271 36072 2297
rect 36126 2271 36156 2297
rect 36210 2271 36240 2297
rect 36294 2271 36324 2297
rect 36378 2271 36408 2297
rect 36462 2271 36492 2297
rect 36546 2271 36576 2297
rect 36630 2271 36660 2297
rect 36714 2271 36744 2297
rect 36798 2271 36828 2297
rect 36882 2271 36912 2297
rect 36966 2271 36996 2297
rect 37050 2271 37080 2297
rect 37134 2271 37164 2297
rect 37218 2271 37248 2297
rect 52938 2495 52968 2527
rect 53022 2495 53052 2527
rect 53106 2495 53136 2527
rect 53190 2495 53220 2527
rect 53274 2495 53304 2527
rect 53358 2495 53388 2527
rect 53442 2495 53472 2527
rect 53526 2495 53556 2527
rect 53610 2495 53640 2527
rect 53694 2495 53724 2527
rect 53778 2495 53808 2527
rect 53862 2495 53892 2527
rect 53946 2495 53976 2527
rect 54030 2495 54060 2527
rect 54114 2495 54144 2527
rect 54198 2495 54228 2527
rect 37840 2269 37870 2295
rect 37924 2269 37954 2295
rect 38008 2269 38038 2295
rect 38092 2269 38122 2295
rect 38176 2269 38206 2295
rect 38260 2269 38290 2295
rect 38344 2269 38374 2295
rect 38428 2269 38458 2295
rect 38512 2269 38542 2295
rect 38596 2269 38626 2295
rect 38680 2269 38710 2295
rect 38764 2269 38794 2295
rect 38848 2269 38878 2295
rect 38932 2269 38962 2295
rect 39016 2269 39046 2295
rect 39100 2269 39130 2295
rect 51056 2271 51086 2297
rect 51140 2271 51170 2297
rect 51224 2271 51254 2297
rect 51308 2271 51338 2297
rect 51392 2271 51422 2297
rect 51476 2271 51506 2297
rect 51560 2271 51590 2297
rect 51644 2271 51674 2297
rect 51728 2271 51758 2297
rect 51812 2271 51842 2297
rect 51896 2271 51926 2297
rect 51980 2271 52010 2297
rect 52064 2271 52094 2297
rect 52148 2271 52178 2297
rect 52232 2271 52262 2297
rect 52316 2271 52346 2297
rect 52938 2269 52968 2295
rect 53022 2269 53052 2295
rect 53106 2269 53136 2295
rect 53190 2269 53220 2295
rect 53274 2269 53304 2295
rect 53358 2269 53388 2295
rect 53442 2269 53472 2295
rect 53526 2269 53556 2295
rect 53610 2269 53640 2295
rect 53694 2269 53724 2295
rect 53778 2269 53808 2295
rect 53862 2269 53892 2295
rect 53946 2269 53976 2295
rect 54030 2269 54060 2295
rect 54114 2269 54144 2295
rect 54198 2269 54228 2295
rect 297 2123 327 2149
rect 369 2123 399 2149
rect 1111 2123 1141 2149
rect 1183 2123 1213 2149
rect 2185 2123 2215 2149
rect 2257 2123 2287 2149
rect 734 2039 800 2055
rect 734 2005 750 2039
rect 784 2005 800 2039
rect 734 1989 800 2005
rect 656 1958 686 1984
rect 752 1958 782 1989
rect 297 1891 327 1923
rect 240 1875 327 1891
rect 240 1841 255 1875
rect 289 1841 327 1875
rect 369 1891 399 1923
rect 369 1875 473 1891
rect 369 1861 423 1875
rect 240 1825 327 1841
rect 297 1803 327 1825
rect 381 1841 423 1861
rect 457 1841 473 1875
rect 381 1825 473 1841
rect 381 1803 411 1825
rect 2999 2123 3029 2149
rect 3071 2123 3101 2149
rect 4073 2123 4103 2149
rect 4145 2123 4175 2149
rect 2622 2039 2688 2055
rect 2622 2005 2638 2039
rect 2672 2005 2688 2039
rect 2622 1989 2688 2005
rect 2544 1958 2574 1984
rect 2640 1958 2670 1989
rect 1111 1891 1141 1923
rect 1054 1875 1141 1891
rect 1054 1841 1069 1875
rect 1103 1841 1141 1875
rect 1183 1891 1213 1923
rect 2185 1891 2215 1923
rect 1183 1875 1287 1891
rect 1183 1861 1237 1875
rect 1054 1825 1141 1841
rect 1111 1803 1141 1825
rect 1195 1841 1237 1861
rect 1271 1841 1287 1875
rect 1195 1825 1287 1841
rect 2128 1875 2215 1891
rect 2128 1841 2143 1875
rect 2177 1841 2215 1875
rect 2257 1891 2287 1923
rect 2257 1875 2361 1891
rect 2257 1861 2311 1875
rect 2128 1825 2215 1841
rect 1195 1803 1225 1825
rect 2185 1803 2215 1825
rect 2269 1841 2311 1861
rect 2345 1841 2361 1875
rect 2269 1825 2361 1841
rect 2269 1803 2299 1825
rect 656 1727 686 1758
rect 752 1732 782 1758
rect 638 1711 704 1727
rect 638 1677 654 1711
rect 688 1690 704 1711
rect 688 1677 816 1690
rect 297 1647 327 1673
rect 381 1647 411 1673
rect 638 1658 816 1677
rect 4887 2123 4917 2149
rect 4959 2123 4989 2149
rect 5961 2123 5991 2149
rect 6033 2123 6063 2149
rect 4510 2039 4576 2055
rect 4510 2005 4526 2039
rect 4560 2005 4576 2039
rect 4510 1989 4576 2005
rect 4432 1958 4462 1984
rect 4528 1958 4558 1989
rect 2999 1891 3029 1923
rect 2942 1875 3029 1891
rect 2942 1841 2957 1875
rect 2991 1841 3029 1875
rect 3071 1891 3101 1923
rect 4073 1891 4103 1923
rect 3071 1875 3175 1891
rect 3071 1861 3125 1875
rect 2942 1825 3029 1841
rect 2999 1803 3029 1825
rect 3083 1841 3125 1861
rect 3159 1841 3175 1875
rect 3083 1825 3175 1841
rect 4016 1875 4103 1891
rect 4016 1841 4031 1875
rect 4065 1841 4103 1875
rect 4145 1891 4175 1923
rect 4145 1875 4249 1891
rect 4145 1861 4199 1875
rect 4016 1825 4103 1841
rect 3083 1803 3113 1825
rect 4073 1803 4103 1825
rect 4157 1841 4199 1861
rect 4233 1841 4249 1875
rect 4157 1825 4249 1841
rect 4157 1803 4187 1825
rect 2544 1727 2574 1758
rect 2640 1732 2670 1758
rect 2526 1711 2592 1727
rect 2526 1677 2542 1711
rect 2576 1690 2592 1711
rect 2576 1677 2704 1690
rect 750 1630 816 1658
rect 1111 1647 1141 1673
rect 1195 1647 1225 1673
rect 2185 1647 2215 1673
rect 2269 1647 2299 1673
rect 2526 1658 2704 1677
rect 6775 2123 6805 2149
rect 6847 2123 6877 2149
rect 7849 2123 7879 2149
rect 7921 2123 7951 2149
rect 6398 2039 6464 2055
rect 6398 2005 6414 2039
rect 6448 2005 6464 2039
rect 6398 1989 6464 2005
rect 6320 1958 6350 1984
rect 6416 1958 6446 1989
rect 4887 1891 4917 1923
rect 4830 1875 4917 1891
rect 4830 1841 4845 1875
rect 4879 1841 4917 1875
rect 4959 1891 4989 1923
rect 5961 1891 5991 1923
rect 4959 1875 5063 1891
rect 4959 1861 5013 1875
rect 4830 1825 4917 1841
rect 4887 1803 4917 1825
rect 4971 1841 5013 1861
rect 5047 1841 5063 1875
rect 4971 1825 5063 1841
rect 5904 1875 5991 1891
rect 5904 1841 5919 1875
rect 5953 1841 5991 1875
rect 6033 1891 6063 1923
rect 6033 1875 6137 1891
rect 6033 1861 6087 1875
rect 5904 1825 5991 1841
rect 4971 1803 5001 1825
rect 5961 1803 5991 1825
rect 6045 1841 6087 1861
rect 6121 1841 6137 1875
rect 6045 1825 6137 1841
rect 6045 1803 6075 1825
rect 4432 1727 4462 1758
rect 4528 1732 4558 1758
rect 4414 1711 4480 1727
rect 4414 1677 4430 1711
rect 4464 1690 4480 1711
rect 4464 1677 4592 1690
rect 750 1596 766 1630
rect 800 1596 816 1630
rect 672 1558 702 1584
rect 750 1580 816 1596
rect 2638 1630 2704 1658
rect 2999 1647 3029 1673
rect 3083 1647 3113 1673
rect 4073 1647 4103 1673
rect 4157 1647 4187 1673
rect 4414 1658 4592 1677
rect 8663 2123 8693 2149
rect 8735 2123 8765 2149
rect 9737 2123 9767 2149
rect 9809 2123 9839 2149
rect 8286 2039 8352 2055
rect 8286 2005 8302 2039
rect 8336 2005 8352 2039
rect 8286 1989 8352 2005
rect 8208 1958 8238 1984
rect 8304 1958 8334 1989
rect 6775 1891 6805 1923
rect 6718 1875 6805 1891
rect 6718 1841 6733 1875
rect 6767 1841 6805 1875
rect 6847 1891 6877 1923
rect 7849 1891 7879 1923
rect 6847 1875 6951 1891
rect 6847 1861 6901 1875
rect 6718 1825 6805 1841
rect 6775 1803 6805 1825
rect 6859 1841 6901 1861
rect 6935 1841 6951 1875
rect 6859 1825 6951 1841
rect 7792 1875 7879 1891
rect 7792 1841 7807 1875
rect 7841 1841 7879 1875
rect 7921 1891 7951 1923
rect 7921 1875 8025 1891
rect 7921 1861 7975 1875
rect 7792 1825 7879 1841
rect 6859 1803 6889 1825
rect 7849 1803 7879 1825
rect 7933 1841 7975 1861
rect 8009 1841 8025 1875
rect 7933 1825 8025 1841
rect 7933 1803 7963 1825
rect 6320 1727 6350 1758
rect 6416 1732 6446 1758
rect 6302 1711 6368 1727
rect 6302 1677 6318 1711
rect 6352 1690 6368 1711
rect 6352 1677 6480 1690
rect 2638 1596 2654 1630
rect 2688 1596 2704 1630
rect 768 1558 798 1580
rect 2560 1558 2590 1584
rect 2638 1580 2704 1596
rect 4526 1630 4592 1658
rect 4887 1647 4917 1673
rect 4971 1647 5001 1673
rect 5961 1647 5991 1673
rect 6045 1647 6075 1673
rect 6302 1658 6480 1677
rect 10551 2123 10581 2149
rect 10623 2123 10653 2149
rect 11625 2123 11655 2149
rect 11697 2123 11727 2149
rect 10174 2039 10240 2055
rect 10174 2005 10190 2039
rect 10224 2005 10240 2039
rect 10174 1989 10240 2005
rect 10096 1958 10126 1984
rect 10192 1958 10222 1989
rect 8663 1891 8693 1923
rect 8606 1875 8693 1891
rect 8606 1841 8621 1875
rect 8655 1841 8693 1875
rect 8735 1891 8765 1923
rect 9737 1891 9767 1923
rect 8735 1875 8839 1891
rect 8735 1861 8789 1875
rect 8606 1825 8693 1841
rect 8663 1803 8693 1825
rect 8747 1841 8789 1861
rect 8823 1841 8839 1875
rect 8747 1825 8839 1841
rect 9680 1875 9767 1891
rect 9680 1841 9695 1875
rect 9729 1841 9767 1875
rect 9809 1891 9839 1923
rect 9809 1875 9913 1891
rect 9809 1861 9863 1875
rect 9680 1825 9767 1841
rect 8747 1803 8777 1825
rect 9737 1803 9767 1825
rect 9821 1841 9863 1861
rect 9897 1841 9913 1875
rect 9821 1825 9913 1841
rect 9821 1803 9851 1825
rect 8208 1727 8238 1758
rect 8304 1732 8334 1758
rect 8190 1711 8256 1727
rect 8190 1677 8206 1711
rect 8240 1690 8256 1711
rect 8240 1677 8368 1690
rect 4526 1596 4542 1630
rect 4576 1596 4592 1630
rect 2656 1558 2686 1580
rect 4448 1558 4478 1584
rect 4526 1580 4592 1596
rect 6414 1630 6480 1658
rect 6775 1647 6805 1673
rect 6859 1647 6889 1673
rect 7849 1647 7879 1673
rect 7933 1647 7963 1673
rect 8190 1658 8368 1677
rect 12439 2123 12469 2149
rect 12511 2123 12541 2149
rect 13513 2123 13543 2149
rect 13585 2123 13615 2149
rect 12062 2039 12128 2055
rect 12062 2005 12078 2039
rect 12112 2005 12128 2039
rect 12062 1989 12128 2005
rect 11984 1958 12014 1984
rect 12080 1958 12110 1989
rect 10551 1891 10581 1923
rect 10494 1875 10581 1891
rect 10494 1841 10509 1875
rect 10543 1841 10581 1875
rect 10623 1891 10653 1923
rect 11625 1891 11655 1923
rect 10623 1875 10727 1891
rect 10623 1861 10677 1875
rect 10494 1825 10581 1841
rect 10551 1803 10581 1825
rect 10635 1841 10677 1861
rect 10711 1841 10727 1875
rect 10635 1825 10727 1841
rect 11568 1875 11655 1891
rect 11568 1841 11583 1875
rect 11617 1841 11655 1875
rect 11697 1891 11727 1923
rect 11697 1875 11801 1891
rect 11697 1861 11751 1875
rect 11568 1825 11655 1841
rect 10635 1803 10665 1825
rect 11625 1803 11655 1825
rect 11709 1841 11751 1861
rect 11785 1841 11801 1875
rect 11709 1825 11801 1841
rect 11709 1803 11739 1825
rect 10096 1727 10126 1758
rect 10192 1732 10222 1758
rect 10078 1711 10144 1727
rect 10078 1677 10094 1711
rect 10128 1690 10144 1711
rect 10128 1677 10256 1690
rect 6414 1596 6430 1630
rect 6464 1596 6480 1630
rect 4544 1558 4574 1580
rect 6336 1558 6366 1584
rect 6414 1580 6480 1596
rect 8302 1630 8368 1658
rect 8663 1647 8693 1673
rect 8747 1647 8777 1673
rect 9737 1647 9767 1673
rect 9821 1647 9851 1673
rect 10078 1658 10256 1677
rect 14327 2123 14357 2149
rect 14399 2123 14429 2149
rect 15395 2123 15425 2149
rect 15467 2123 15497 2149
rect 13950 2039 14016 2055
rect 13950 2005 13966 2039
rect 14000 2005 14016 2039
rect 13950 1989 14016 2005
rect 13872 1958 13902 1984
rect 13968 1958 13998 1989
rect 12439 1891 12469 1923
rect 12382 1875 12469 1891
rect 12382 1841 12397 1875
rect 12431 1841 12469 1875
rect 12511 1891 12541 1923
rect 13513 1891 13543 1923
rect 12511 1875 12615 1891
rect 12511 1861 12565 1875
rect 12382 1825 12469 1841
rect 12439 1803 12469 1825
rect 12523 1841 12565 1861
rect 12599 1841 12615 1875
rect 12523 1825 12615 1841
rect 13456 1875 13543 1891
rect 13456 1841 13471 1875
rect 13505 1841 13543 1875
rect 13585 1891 13615 1923
rect 13585 1875 13689 1891
rect 13585 1861 13639 1875
rect 13456 1825 13543 1841
rect 12523 1803 12553 1825
rect 13513 1803 13543 1825
rect 13597 1841 13639 1861
rect 13673 1841 13689 1875
rect 13597 1825 13689 1841
rect 13597 1803 13627 1825
rect 11984 1727 12014 1758
rect 12080 1732 12110 1758
rect 11966 1711 12032 1727
rect 11966 1677 11982 1711
rect 12016 1690 12032 1711
rect 12016 1677 12144 1690
rect 8302 1596 8318 1630
rect 8352 1596 8368 1630
rect 6432 1558 6462 1580
rect 8224 1558 8254 1584
rect 8302 1580 8368 1596
rect 10190 1630 10256 1658
rect 10551 1647 10581 1673
rect 10635 1647 10665 1673
rect 11625 1647 11655 1673
rect 11709 1647 11739 1673
rect 11966 1658 12144 1677
rect 16209 2123 16239 2149
rect 16281 2123 16311 2149
rect 17283 2123 17313 2149
rect 17355 2123 17385 2149
rect 15832 2039 15898 2055
rect 15832 2005 15848 2039
rect 15882 2005 15898 2039
rect 15832 1989 15898 2005
rect 15754 1958 15784 1984
rect 15850 1958 15880 1989
rect 14327 1891 14357 1923
rect 14270 1875 14357 1891
rect 14270 1841 14285 1875
rect 14319 1841 14357 1875
rect 14399 1891 14429 1923
rect 15395 1891 15425 1923
rect 14399 1875 14503 1891
rect 14399 1861 14453 1875
rect 14270 1825 14357 1841
rect 14327 1803 14357 1825
rect 14411 1841 14453 1861
rect 14487 1841 14503 1875
rect 14411 1825 14503 1841
rect 15338 1875 15425 1891
rect 15338 1841 15353 1875
rect 15387 1841 15425 1875
rect 15467 1891 15497 1923
rect 15467 1875 15571 1891
rect 15467 1861 15521 1875
rect 15338 1825 15425 1841
rect 14411 1803 14441 1825
rect 15395 1803 15425 1825
rect 15479 1841 15521 1861
rect 15555 1841 15571 1875
rect 15479 1825 15571 1841
rect 15479 1803 15509 1825
rect 13872 1727 13902 1758
rect 13968 1732 13998 1758
rect 13854 1711 13920 1727
rect 13854 1677 13870 1711
rect 13904 1690 13920 1711
rect 13904 1677 14032 1690
rect 10190 1596 10206 1630
rect 10240 1596 10256 1630
rect 8320 1558 8350 1580
rect 10112 1558 10142 1584
rect 10190 1580 10256 1596
rect 12078 1630 12144 1658
rect 12439 1647 12469 1673
rect 12523 1647 12553 1673
rect 13513 1647 13543 1673
rect 13597 1647 13627 1673
rect 13854 1658 14032 1677
rect 18097 2123 18127 2149
rect 18169 2123 18199 2149
rect 19171 2123 19201 2149
rect 19243 2123 19273 2149
rect 17720 2039 17786 2055
rect 17720 2005 17736 2039
rect 17770 2005 17786 2039
rect 17720 1989 17786 2005
rect 17642 1958 17672 1984
rect 17738 1958 17768 1989
rect 16209 1891 16239 1923
rect 16152 1875 16239 1891
rect 16152 1841 16167 1875
rect 16201 1841 16239 1875
rect 16281 1891 16311 1923
rect 17283 1891 17313 1923
rect 16281 1875 16385 1891
rect 16281 1861 16335 1875
rect 16152 1825 16239 1841
rect 16209 1803 16239 1825
rect 16293 1841 16335 1861
rect 16369 1841 16385 1875
rect 16293 1825 16385 1841
rect 17226 1875 17313 1891
rect 17226 1841 17241 1875
rect 17275 1841 17313 1875
rect 17355 1891 17385 1923
rect 17355 1875 17459 1891
rect 17355 1861 17409 1875
rect 17226 1825 17313 1841
rect 16293 1803 16323 1825
rect 17283 1803 17313 1825
rect 17367 1841 17409 1861
rect 17443 1841 17459 1875
rect 17367 1825 17459 1841
rect 17367 1803 17397 1825
rect 15754 1727 15784 1758
rect 15850 1732 15880 1758
rect 15736 1711 15802 1727
rect 15736 1677 15752 1711
rect 15786 1690 15802 1711
rect 15786 1677 15914 1690
rect 12078 1596 12094 1630
rect 12128 1596 12144 1630
rect 10208 1558 10238 1580
rect 12000 1558 12030 1584
rect 12078 1580 12144 1596
rect 13966 1630 14032 1658
rect 14327 1647 14357 1673
rect 14411 1647 14441 1673
rect 15395 1647 15425 1673
rect 15479 1647 15509 1673
rect 15736 1658 15914 1677
rect 19985 2123 20015 2149
rect 20057 2123 20087 2149
rect 21059 2123 21089 2149
rect 21131 2123 21161 2149
rect 19608 2039 19674 2055
rect 19608 2005 19624 2039
rect 19658 2005 19674 2039
rect 19608 1989 19674 2005
rect 19530 1958 19560 1984
rect 19626 1958 19656 1989
rect 18097 1891 18127 1923
rect 18040 1875 18127 1891
rect 18040 1841 18055 1875
rect 18089 1841 18127 1875
rect 18169 1891 18199 1923
rect 19171 1891 19201 1923
rect 18169 1875 18273 1891
rect 18169 1861 18223 1875
rect 18040 1825 18127 1841
rect 18097 1803 18127 1825
rect 18181 1841 18223 1861
rect 18257 1841 18273 1875
rect 18181 1825 18273 1841
rect 19114 1875 19201 1891
rect 19114 1841 19129 1875
rect 19163 1841 19201 1875
rect 19243 1891 19273 1923
rect 19243 1875 19347 1891
rect 19243 1861 19297 1875
rect 19114 1825 19201 1841
rect 18181 1803 18211 1825
rect 19171 1803 19201 1825
rect 19255 1841 19297 1861
rect 19331 1841 19347 1875
rect 19255 1825 19347 1841
rect 19255 1803 19285 1825
rect 17642 1727 17672 1758
rect 17738 1732 17768 1758
rect 17624 1711 17690 1727
rect 17624 1677 17640 1711
rect 17674 1690 17690 1711
rect 17674 1677 17802 1690
rect 13966 1596 13982 1630
rect 14016 1596 14032 1630
rect 12096 1558 12126 1580
rect 13888 1558 13918 1584
rect 13966 1580 14032 1596
rect 15848 1630 15914 1658
rect 16209 1647 16239 1673
rect 16293 1647 16323 1673
rect 17283 1647 17313 1673
rect 17367 1647 17397 1673
rect 17624 1658 17802 1677
rect 21873 2123 21903 2149
rect 21945 2123 21975 2149
rect 22947 2123 22977 2149
rect 23019 2123 23049 2149
rect 21496 2039 21562 2055
rect 21496 2005 21512 2039
rect 21546 2005 21562 2039
rect 21496 1989 21562 2005
rect 21418 1958 21448 1984
rect 21514 1958 21544 1989
rect 19985 1891 20015 1923
rect 19928 1875 20015 1891
rect 19928 1841 19943 1875
rect 19977 1841 20015 1875
rect 20057 1891 20087 1923
rect 21059 1891 21089 1923
rect 20057 1875 20161 1891
rect 20057 1861 20111 1875
rect 19928 1825 20015 1841
rect 19985 1803 20015 1825
rect 20069 1841 20111 1861
rect 20145 1841 20161 1875
rect 20069 1825 20161 1841
rect 21002 1875 21089 1891
rect 21002 1841 21017 1875
rect 21051 1841 21089 1875
rect 21131 1891 21161 1923
rect 21131 1875 21235 1891
rect 21131 1861 21185 1875
rect 21002 1825 21089 1841
rect 20069 1803 20099 1825
rect 21059 1803 21089 1825
rect 21143 1841 21185 1861
rect 21219 1841 21235 1875
rect 21143 1825 21235 1841
rect 21143 1803 21173 1825
rect 19530 1727 19560 1758
rect 19626 1732 19656 1758
rect 19512 1711 19578 1727
rect 19512 1677 19528 1711
rect 19562 1690 19578 1711
rect 19562 1677 19690 1690
rect 15848 1596 15864 1630
rect 15898 1596 15914 1630
rect 13984 1558 14014 1580
rect 15770 1558 15800 1584
rect 15848 1580 15914 1596
rect 17736 1630 17802 1658
rect 18097 1647 18127 1673
rect 18181 1647 18211 1673
rect 19171 1647 19201 1673
rect 19255 1647 19285 1673
rect 19512 1658 19690 1677
rect 23761 2123 23791 2149
rect 23833 2123 23863 2149
rect 24835 2123 24865 2149
rect 24907 2123 24937 2149
rect 23384 2039 23450 2055
rect 23384 2005 23400 2039
rect 23434 2005 23450 2039
rect 23384 1989 23450 2005
rect 23306 1958 23336 1984
rect 23402 1958 23432 1989
rect 21873 1891 21903 1923
rect 21816 1875 21903 1891
rect 21816 1841 21831 1875
rect 21865 1841 21903 1875
rect 21945 1891 21975 1923
rect 22947 1891 22977 1923
rect 21945 1875 22049 1891
rect 21945 1861 21999 1875
rect 21816 1825 21903 1841
rect 21873 1803 21903 1825
rect 21957 1841 21999 1861
rect 22033 1841 22049 1875
rect 21957 1825 22049 1841
rect 22890 1875 22977 1891
rect 22890 1841 22905 1875
rect 22939 1841 22977 1875
rect 23019 1891 23049 1923
rect 23019 1875 23123 1891
rect 23019 1861 23073 1875
rect 22890 1825 22977 1841
rect 21957 1803 21987 1825
rect 22947 1803 22977 1825
rect 23031 1841 23073 1861
rect 23107 1841 23123 1875
rect 23031 1825 23123 1841
rect 23031 1803 23061 1825
rect 21418 1727 21448 1758
rect 21514 1732 21544 1758
rect 21400 1711 21466 1727
rect 21400 1677 21416 1711
rect 21450 1690 21466 1711
rect 21450 1677 21578 1690
rect 17736 1596 17752 1630
rect 17786 1596 17802 1630
rect 15866 1558 15896 1580
rect 17658 1558 17688 1584
rect 17736 1580 17802 1596
rect 19624 1630 19690 1658
rect 19985 1647 20015 1673
rect 20069 1647 20099 1673
rect 21059 1647 21089 1673
rect 21143 1647 21173 1673
rect 21400 1658 21578 1677
rect 25649 2123 25679 2149
rect 25721 2123 25751 2149
rect 26723 2123 26753 2149
rect 26795 2123 26825 2149
rect 25272 2039 25338 2055
rect 25272 2005 25288 2039
rect 25322 2005 25338 2039
rect 25272 1989 25338 2005
rect 25194 1958 25224 1984
rect 25290 1958 25320 1989
rect 23761 1891 23791 1923
rect 23704 1875 23791 1891
rect 23704 1841 23719 1875
rect 23753 1841 23791 1875
rect 23833 1891 23863 1923
rect 24835 1891 24865 1923
rect 23833 1875 23937 1891
rect 23833 1861 23887 1875
rect 23704 1825 23791 1841
rect 23761 1803 23791 1825
rect 23845 1841 23887 1861
rect 23921 1841 23937 1875
rect 23845 1825 23937 1841
rect 24778 1875 24865 1891
rect 24778 1841 24793 1875
rect 24827 1841 24865 1875
rect 24907 1891 24937 1923
rect 24907 1875 25011 1891
rect 24907 1861 24961 1875
rect 24778 1825 24865 1841
rect 23845 1803 23875 1825
rect 24835 1803 24865 1825
rect 24919 1841 24961 1861
rect 24995 1841 25011 1875
rect 24919 1825 25011 1841
rect 24919 1803 24949 1825
rect 23306 1727 23336 1758
rect 23402 1732 23432 1758
rect 23288 1711 23354 1727
rect 23288 1677 23304 1711
rect 23338 1690 23354 1711
rect 23338 1677 23466 1690
rect 19624 1596 19640 1630
rect 19674 1596 19690 1630
rect 17754 1558 17784 1580
rect 19546 1558 19576 1584
rect 19624 1580 19690 1596
rect 21512 1630 21578 1658
rect 21873 1647 21903 1673
rect 21957 1647 21987 1673
rect 22947 1647 22977 1673
rect 23031 1647 23061 1673
rect 23288 1658 23466 1677
rect 27537 2123 27567 2149
rect 27609 2123 27639 2149
rect 28611 2123 28641 2149
rect 28683 2123 28713 2149
rect 27160 2039 27226 2055
rect 27160 2005 27176 2039
rect 27210 2005 27226 2039
rect 27160 1989 27226 2005
rect 27082 1958 27112 1984
rect 27178 1958 27208 1989
rect 25649 1891 25679 1923
rect 25592 1875 25679 1891
rect 25592 1841 25607 1875
rect 25641 1841 25679 1875
rect 25721 1891 25751 1923
rect 26723 1891 26753 1923
rect 25721 1875 25825 1891
rect 25721 1861 25775 1875
rect 25592 1825 25679 1841
rect 25649 1803 25679 1825
rect 25733 1841 25775 1861
rect 25809 1841 25825 1875
rect 25733 1825 25825 1841
rect 26666 1875 26753 1891
rect 26666 1841 26681 1875
rect 26715 1841 26753 1875
rect 26795 1891 26825 1923
rect 26795 1875 26899 1891
rect 26795 1861 26849 1875
rect 26666 1825 26753 1841
rect 25733 1803 25763 1825
rect 26723 1803 26753 1825
rect 26807 1841 26849 1861
rect 26883 1841 26899 1875
rect 26807 1825 26899 1841
rect 26807 1803 26837 1825
rect 25194 1727 25224 1758
rect 25290 1732 25320 1758
rect 25176 1711 25242 1727
rect 25176 1677 25192 1711
rect 25226 1690 25242 1711
rect 25226 1677 25354 1690
rect 21512 1596 21528 1630
rect 21562 1596 21578 1630
rect 19642 1558 19672 1580
rect 21434 1558 21464 1584
rect 21512 1580 21578 1596
rect 23400 1630 23466 1658
rect 23761 1647 23791 1673
rect 23845 1647 23875 1673
rect 24835 1647 24865 1673
rect 24919 1647 24949 1673
rect 25176 1658 25354 1677
rect 29425 2123 29455 2149
rect 29497 2123 29527 2149
rect 30499 2123 30529 2149
rect 30571 2123 30601 2149
rect 29048 2039 29114 2055
rect 29048 2005 29064 2039
rect 29098 2005 29114 2039
rect 29048 1989 29114 2005
rect 28970 1958 29000 1984
rect 29066 1958 29096 1989
rect 27537 1891 27567 1923
rect 27480 1875 27567 1891
rect 27480 1841 27495 1875
rect 27529 1841 27567 1875
rect 27609 1891 27639 1923
rect 28611 1891 28641 1923
rect 27609 1875 27713 1891
rect 27609 1861 27663 1875
rect 27480 1825 27567 1841
rect 27537 1803 27567 1825
rect 27621 1841 27663 1861
rect 27697 1841 27713 1875
rect 27621 1825 27713 1841
rect 28554 1875 28641 1891
rect 28554 1841 28569 1875
rect 28603 1841 28641 1875
rect 28683 1891 28713 1923
rect 28683 1875 28787 1891
rect 28683 1861 28737 1875
rect 28554 1825 28641 1841
rect 27621 1803 27651 1825
rect 28611 1803 28641 1825
rect 28695 1841 28737 1861
rect 28771 1841 28787 1875
rect 28695 1825 28787 1841
rect 28695 1803 28725 1825
rect 27082 1727 27112 1758
rect 27178 1732 27208 1758
rect 27064 1711 27130 1727
rect 27064 1677 27080 1711
rect 27114 1690 27130 1711
rect 27114 1677 27242 1690
rect 23400 1596 23416 1630
rect 23450 1596 23466 1630
rect 21530 1558 21560 1580
rect 23322 1558 23352 1584
rect 23400 1580 23466 1596
rect 25288 1630 25354 1658
rect 25649 1647 25679 1673
rect 25733 1647 25763 1673
rect 26723 1647 26753 1673
rect 26807 1647 26837 1673
rect 27064 1658 27242 1677
rect 31313 2123 31343 2149
rect 31385 2123 31415 2149
rect 32387 2123 32417 2149
rect 32459 2123 32489 2149
rect 30936 2039 31002 2055
rect 30936 2005 30952 2039
rect 30986 2005 31002 2039
rect 30936 1989 31002 2005
rect 30858 1958 30888 1984
rect 30954 1958 30984 1989
rect 29425 1891 29455 1923
rect 29368 1875 29455 1891
rect 29368 1841 29383 1875
rect 29417 1841 29455 1875
rect 29497 1891 29527 1923
rect 30499 1891 30529 1923
rect 29497 1875 29601 1891
rect 29497 1861 29551 1875
rect 29368 1825 29455 1841
rect 29425 1803 29455 1825
rect 29509 1841 29551 1861
rect 29585 1841 29601 1875
rect 29509 1825 29601 1841
rect 30442 1875 30529 1891
rect 30442 1841 30457 1875
rect 30491 1841 30529 1875
rect 30571 1891 30601 1923
rect 30571 1875 30675 1891
rect 30571 1861 30625 1875
rect 30442 1825 30529 1841
rect 29509 1803 29539 1825
rect 30499 1803 30529 1825
rect 30583 1841 30625 1861
rect 30659 1841 30675 1875
rect 30583 1825 30675 1841
rect 30583 1803 30613 1825
rect 28970 1727 29000 1758
rect 29066 1732 29096 1758
rect 28952 1711 29018 1727
rect 28952 1677 28968 1711
rect 29002 1690 29018 1711
rect 29002 1677 29130 1690
rect 25288 1596 25304 1630
rect 25338 1596 25354 1630
rect 23418 1558 23448 1580
rect 25210 1558 25240 1584
rect 25288 1580 25354 1596
rect 27176 1630 27242 1658
rect 27537 1647 27567 1673
rect 27621 1647 27651 1673
rect 28611 1647 28641 1673
rect 28695 1647 28725 1673
rect 28952 1658 29130 1677
rect 33201 2123 33231 2149
rect 33273 2123 33303 2149
rect 34275 2123 34305 2149
rect 34347 2123 34377 2149
rect 32824 2039 32890 2055
rect 32824 2005 32840 2039
rect 32874 2005 32890 2039
rect 32824 1989 32890 2005
rect 32746 1958 32776 1984
rect 32842 1958 32872 1989
rect 31313 1891 31343 1923
rect 31256 1875 31343 1891
rect 31256 1841 31271 1875
rect 31305 1841 31343 1875
rect 31385 1891 31415 1923
rect 32387 1891 32417 1923
rect 31385 1875 31489 1891
rect 31385 1861 31439 1875
rect 31256 1825 31343 1841
rect 31313 1803 31343 1825
rect 31397 1841 31439 1861
rect 31473 1841 31489 1875
rect 31397 1825 31489 1841
rect 32330 1875 32417 1891
rect 32330 1841 32345 1875
rect 32379 1841 32417 1875
rect 32459 1891 32489 1923
rect 32459 1875 32563 1891
rect 32459 1861 32513 1875
rect 32330 1825 32417 1841
rect 31397 1803 31427 1825
rect 32387 1803 32417 1825
rect 32471 1841 32513 1861
rect 32547 1841 32563 1875
rect 32471 1825 32563 1841
rect 32471 1803 32501 1825
rect 30858 1727 30888 1758
rect 30954 1732 30984 1758
rect 30840 1711 30906 1727
rect 30840 1677 30856 1711
rect 30890 1690 30906 1711
rect 30890 1677 31018 1690
rect 27176 1596 27192 1630
rect 27226 1596 27242 1630
rect 25306 1558 25336 1580
rect 27098 1558 27128 1584
rect 27176 1580 27242 1596
rect 29064 1630 29130 1658
rect 29425 1647 29455 1673
rect 29509 1647 29539 1673
rect 30499 1647 30529 1673
rect 30583 1647 30613 1673
rect 30840 1658 31018 1677
rect 35089 2123 35119 2149
rect 35161 2123 35191 2149
rect 36163 2123 36193 2149
rect 36235 2123 36265 2149
rect 34712 2039 34778 2055
rect 34712 2005 34728 2039
rect 34762 2005 34778 2039
rect 34712 1989 34778 2005
rect 34634 1958 34664 1984
rect 34730 1958 34760 1989
rect 33201 1891 33231 1923
rect 33144 1875 33231 1891
rect 33144 1841 33159 1875
rect 33193 1841 33231 1875
rect 33273 1891 33303 1923
rect 34275 1891 34305 1923
rect 33273 1875 33377 1891
rect 33273 1861 33327 1875
rect 33144 1825 33231 1841
rect 33201 1803 33231 1825
rect 33285 1841 33327 1861
rect 33361 1841 33377 1875
rect 33285 1825 33377 1841
rect 34218 1875 34305 1891
rect 34218 1841 34233 1875
rect 34267 1841 34305 1875
rect 34347 1891 34377 1923
rect 34347 1875 34451 1891
rect 34347 1861 34401 1875
rect 34218 1825 34305 1841
rect 33285 1803 33315 1825
rect 34275 1803 34305 1825
rect 34359 1841 34401 1861
rect 34435 1841 34451 1875
rect 34359 1825 34451 1841
rect 34359 1803 34389 1825
rect 32746 1727 32776 1758
rect 32842 1732 32872 1758
rect 32728 1711 32794 1727
rect 32728 1677 32744 1711
rect 32778 1690 32794 1711
rect 32778 1677 32906 1690
rect 29064 1596 29080 1630
rect 29114 1596 29130 1630
rect 27194 1558 27224 1580
rect 28986 1558 29016 1584
rect 29064 1580 29130 1596
rect 30952 1630 31018 1658
rect 31313 1647 31343 1673
rect 31397 1647 31427 1673
rect 32387 1647 32417 1673
rect 32471 1647 32501 1673
rect 32728 1658 32906 1677
rect 36977 2123 37007 2149
rect 37049 2123 37079 2149
rect 38051 2123 38081 2149
rect 38123 2123 38153 2149
rect 36600 2039 36666 2055
rect 36600 2005 36616 2039
rect 36650 2005 36666 2039
rect 36600 1989 36666 2005
rect 36522 1958 36552 1984
rect 36618 1958 36648 1989
rect 35089 1891 35119 1923
rect 35032 1875 35119 1891
rect 35032 1841 35047 1875
rect 35081 1841 35119 1875
rect 35161 1891 35191 1923
rect 36163 1891 36193 1923
rect 35161 1875 35265 1891
rect 35161 1861 35215 1875
rect 35032 1825 35119 1841
rect 35089 1803 35119 1825
rect 35173 1841 35215 1861
rect 35249 1841 35265 1875
rect 35173 1825 35265 1841
rect 36106 1875 36193 1891
rect 36106 1841 36121 1875
rect 36155 1841 36193 1875
rect 36235 1891 36265 1923
rect 36235 1875 36339 1891
rect 36235 1861 36289 1875
rect 36106 1825 36193 1841
rect 35173 1803 35203 1825
rect 36163 1803 36193 1825
rect 36247 1841 36289 1861
rect 36323 1841 36339 1875
rect 36247 1825 36339 1841
rect 36247 1803 36277 1825
rect 34634 1727 34664 1758
rect 34730 1732 34760 1758
rect 34616 1711 34682 1727
rect 34616 1677 34632 1711
rect 34666 1690 34682 1711
rect 34666 1677 34794 1690
rect 30952 1596 30968 1630
rect 31002 1596 31018 1630
rect 29082 1558 29112 1580
rect 30874 1558 30904 1584
rect 30952 1580 31018 1596
rect 32840 1630 32906 1658
rect 33201 1647 33231 1673
rect 33285 1647 33315 1673
rect 34275 1647 34305 1673
rect 34359 1647 34389 1673
rect 34616 1658 34794 1677
rect 38865 2123 38895 2149
rect 38937 2123 38967 2149
rect 39939 2123 39969 2149
rect 40011 2123 40041 2149
rect 38488 2039 38554 2055
rect 38488 2005 38504 2039
rect 38538 2005 38554 2039
rect 38488 1989 38554 2005
rect 38410 1958 38440 1984
rect 38506 1958 38536 1989
rect 36977 1891 37007 1923
rect 36920 1875 37007 1891
rect 36920 1841 36935 1875
rect 36969 1841 37007 1875
rect 37049 1891 37079 1923
rect 38051 1891 38081 1923
rect 37049 1875 37153 1891
rect 37049 1861 37103 1875
rect 36920 1825 37007 1841
rect 36977 1803 37007 1825
rect 37061 1841 37103 1861
rect 37137 1841 37153 1875
rect 37061 1825 37153 1841
rect 37994 1875 38081 1891
rect 37994 1841 38009 1875
rect 38043 1841 38081 1875
rect 38123 1891 38153 1923
rect 38123 1875 38227 1891
rect 38123 1861 38177 1875
rect 37994 1825 38081 1841
rect 37061 1803 37091 1825
rect 38051 1803 38081 1825
rect 38135 1841 38177 1861
rect 38211 1841 38227 1875
rect 38135 1825 38227 1841
rect 38135 1803 38165 1825
rect 36522 1727 36552 1758
rect 36618 1732 36648 1758
rect 36504 1711 36570 1727
rect 36504 1677 36520 1711
rect 36554 1690 36570 1711
rect 36554 1677 36682 1690
rect 32840 1596 32856 1630
rect 32890 1596 32906 1630
rect 30970 1558 31000 1580
rect 32762 1558 32792 1584
rect 32840 1580 32906 1596
rect 34728 1630 34794 1658
rect 35089 1647 35119 1673
rect 35173 1647 35203 1673
rect 36163 1647 36193 1673
rect 36247 1647 36277 1673
rect 36504 1658 36682 1677
rect 40753 2123 40783 2149
rect 40825 2123 40855 2149
rect 41827 2123 41857 2149
rect 41899 2123 41929 2149
rect 40376 2039 40442 2055
rect 40376 2005 40392 2039
rect 40426 2005 40442 2039
rect 40376 1989 40442 2005
rect 40298 1958 40328 1984
rect 40394 1958 40424 1989
rect 38865 1891 38895 1923
rect 38808 1875 38895 1891
rect 38808 1841 38823 1875
rect 38857 1841 38895 1875
rect 38937 1891 38967 1923
rect 39939 1891 39969 1923
rect 38937 1875 39041 1891
rect 38937 1861 38991 1875
rect 38808 1825 38895 1841
rect 38865 1803 38895 1825
rect 38949 1841 38991 1861
rect 39025 1841 39041 1875
rect 38949 1825 39041 1841
rect 39882 1875 39969 1891
rect 39882 1841 39897 1875
rect 39931 1841 39969 1875
rect 40011 1891 40041 1923
rect 40011 1875 40115 1891
rect 40011 1861 40065 1875
rect 39882 1825 39969 1841
rect 38949 1803 38979 1825
rect 39939 1803 39969 1825
rect 40023 1841 40065 1861
rect 40099 1841 40115 1875
rect 40023 1825 40115 1841
rect 40023 1803 40053 1825
rect 38410 1727 38440 1758
rect 38506 1732 38536 1758
rect 38392 1711 38458 1727
rect 38392 1677 38408 1711
rect 38442 1690 38458 1711
rect 38442 1677 38570 1690
rect 34728 1596 34744 1630
rect 34778 1596 34794 1630
rect 32858 1558 32888 1580
rect 34650 1558 34680 1584
rect 34728 1580 34794 1596
rect 36616 1630 36682 1658
rect 36977 1647 37007 1673
rect 37061 1647 37091 1673
rect 38051 1647 38081 1673
rect 38135 1647 38165 1673
rect 38392 1658 38570 1677
rect 42641 2123 42671 2149
rect 42713 2123 42743 2149
rect 43715 2123 43745 2149
rect 43787 2123 43817 2149
rect 42264 2039 42330 2055
rect 42264 2005 42280 2039
rect 42314 2005 42330 2039
rect 42264 1989 42330 2005
rect 42186 1958 42216 1984
rect 42282 1958 42312 1989
rect 40753 1891 40783 1923
rect 40696 1875 40783 1891
rect 40696 1841 40711 1875
rect 40745 1841 40783 1875
rect 40825 1891 40855 1923
rect 41827 1891 41857 1923
rect 40825 1875 40929 1891
rect 40825 1861 40879 1875
rect 40696 1825 40783 1841
rect 40753 1803 40783 1825
rect 40837 1841 40879 1861
rect 40913 1841 40929 1875
rect 40837 1825 40929 1841
rect 41770 1875 41857 1891
rect 41770 1841 41785 1875
rect 41819 1841 41857 1875
rect 41899 1891 41929 1923
rect 41899 1875 42003 1891
rect 41899 1861 41953 1875
rect 41770 1825 41857 1841
rect 40837 1803 40867 1825
rect 41827 1803 41857 1825
rect 41911 1841 41953 1861
rect 41987 1841 42003 1875
rect 41911 1825 42003 1841
rect 41911 1803 41941 1825
rect 40298 1727 40328 1758
rect 40394 1732 40424 1758
rect 40280 1711 40346 1727
rect 40280 1677 40296 1711
rect 40330 1690 40346 1711
rect 40330 1677 40458 1690
rect 36616 1596 36632 1630
rect 36666 1596 36682 1630
rect 34746 1558 34776 1580
rect 36538 1558 36568 1584
rect 36616 1580 36682 1596
rect 38504 1630 38570 1658
rect 38865 1647 38895 1673
rect 38949 1647 38979 1673
rect 39939 1647 39969 1673
rect 40023 1647 40053 1673
rect 40280 1658 40458 1677
rect 44529 2123 44559 2149
rect 44601 2123 44631 2149
rect 45597 2123 45627 2149
rect 45669 2123 45699 2149
rect 44152 2039 44218 2055
rect 44152 2005 44168 2039
rect 44202 2005 44218 2039
rect 44152 1989 44218 2005
rect 44074 1958 44104 1984
rect 44170 1958 44200 1989
rect 42641 1891 42671 1923
rect 42584 1875 42671 1891
rect 42584 1841 42599 1875
rect 42633 1841 42671 1875
rect 42713 1891 42743 1923
rect 43715 1891 43745 1923
rect 42713 1875 42817 1891
rect 42713 1861 42767 1875
rect 42584 1825 42671 1841
rect 42641 1803 42671 1825
rect 42725 1841 42767 1861
rect 42801 1841 42817 1875
rect 42725 1825 42817 1841
rect 43658 1875 43745 1891
rect 43658 1841 43673 1875
rect 43707 1841 43745 1875
rect 43787 1891 43817 1923
rect 43787 1875 43891 1891
rect 43787 1861 43841 1875
rect 43658 1825 43745 1841
rect 42725 1803 42755 1825
rect 43715 1803 43745 1825
rect 43799 1841 43841 1861
rect 43875 1841 43891 1875
rect 43799 1825 43891 1841
rect 43799 1803 43829 1825
rect 42186 1727 42216 1758
rect 42282 1732 42312 1758
rect 42168 1711 42234 1727
rect 42168 1677 42184 1711
rect 42218 1690 42234 1711
rect 42218 1677 42346 1690
rect 38504 1596 38520 1630
rect 38554 1596 38570 1630
rect 36634 1558 36664 1580
rect 38426 1558 38456 1584
rect 38504 1580 38570 1596
rect 40392 1630 40458 1658
rect 40753 1647 40783 1673
rect 40837 1647 40867 1673
rect 41827 1647 41857 1673
rect 41911 1647 41941 1673
rect 42168 1658 42346 1677
rect 46411 2123 46441 2149
rect 46483 2123 46513 2149
rect 47485 2123 47515 2149
rect 47557 2123 47587 2149
rect 46034 2039 46100 2055
rect 46034 2005 46050 2039
rect 46084 2005 46100 2039
rect 46034 1989 46100 2005
rect 45956 1958 45986 1984
rect 46052 1958 46082 1989
rect 44529 1891 44559 1923
rect 44472 1875 44559 1891
rect 44472 1841 44487 1875
rect 44521 1841 44559 1875
rect 44601 1891 44631 1923
rect 45597 1891 45627 1923
rect 44601 1875 44705 1891
rect 44601 1861 44655 1875
rect 44472 1825 44559 1841
rect 44529 1803 44559 1825
rect 44613 1841 44655 1861
rect 44689 1841 44705 1875
rect 44613 1825 44705 1841
rect 45540 1875 45627 1891
rect 45540 1841 45555 1875
rect 45589 1841 45627 1875
rect 45669 1891 45699 1923
rect 45669 1875 45773 1891
rect 45669 1861 45723 1875
rect 45540 1825 45627 1841
rect 44613 1803 44643 1825
rect 45597 1803 45627 1825
rect 45681 1841 45723 1861
rect 45757 1841 45773 1875
rect 45681 1825 45773 1841
rect 45681 1803 45711 1825
rect 44074 1727 44104 1758
rect 44170 1732 44200 1758
rect 44056 1711 44122 1727
rect 44056 1677 44072 1711
rect 44106 1690 44122 1711
rect 44106 1677 44234 1690
rect 40392 1596 40408 1630
rect 40442 1596 40458 1630
rect 38522 1558 38552 1580
rect 40314 1558 40344 1584
rect 40392 1580 40458 1596
rect 42280 1630 42346 1658
rect 42641 1647 42671 1673
rect 42725 1647 42755 1673
rect 43715 1647 43745 1673
rect 43799 1647 43829 1673
rect 44056 1658 44234 1677
rect 48299 2123 48329 2149
rect 48371 2123 48401 2149
rect 49373 2123 49403 2149
rect 49445 2123 49475 2149
rect 47922 2039 47988 2055
rect 47922 2005 47938 2039
rect 47972 2005 47988 2039
rect 47922 1989 47988 2005
rect 47844 1958 47874 1984
rect 47940 1958 47970 1989
rect 46411 1891 46441 1923
rect 46354 1875 46441 1891
rect 46354 1841 46369 1875
rect 46403 1841 46441 1875
rect 46483 1891 46513 1923
rect 47485 1891 47515 1923
rect 46483 1875 46587 1891
rect 46483 1861 46537 1875
rect 46354 1825 46441 1841
rect 46411 1803 46441 1825
rect 46495 1841 46537 1861
rect 46571 1841 46587 1875
rect 46495 1825 46587 1841
rect 47428 1875 47515 1891
rect 47428 1841 47443 1875
rect 47477 1841 47515 1875
rect 47557 1891 47587 1923
rect 47557 1875 47661 1891
rect 47557 1861 47611 1875
rect 47428 1825 47515 1841
rect 46495 1803 46525 1825
rect 47485 1803 47515 1825
rect 47569 1841 47611 1861
rect 47645 1841 47661 1875
rect 47569 1825 47661 1841
rect 47569 1803 47599 1825
rect 45956 1727 45986 1758
rect 46052 1732 46082 1758
rect 45938 1711 46004 1727
rect 45938 1677 45954 1711
rect 45988 1690 46004 1711
rect 45988 1677 46116 1690
rect 42280 1596 42296 1630
rect 42330 1596 42346 1630
rect 40410 1558 40440 1580
rect 42202 1558 42232 1584
rect 42280 1580 42346 1596
rect 44168 1630 44234 1658
rect 44529 1647 44559 1673
rect 44613 1647 44643 1673
rect 45597 1647 45627 1673
rect 45681 1647 45711 1673
rect 45938 1658 46116 1677
rect 50187 2123 50217 2149
rect 50259 2123 50289 2149
rect 51261 2123 51291 2149
rect 51333 2123 51363 2149
rect 49810 2039 49876 2055
rect 49810 2005 49826 2039
rect 49860 2005 49876 2039
rect 49810 1989 49876 2005
rect 49732 1958 49762 1984
rect 49828 1958 49858 1989
rect 48299 1891 48329 1923
rect 48242 1875 48329 1891
rect 48242 1841 48257 1875
rect 48291 1841 48329 1875
rect 48371 1891 48401 1923
rect 49373 1891 49403 1923
rect 48371 1875 48475 1891
rect 48371 1861 48425 1875
rect 48242 1825 48329 1841
rect 48299 1803 48329 1825
rect 48383 1841 48425 1861
rect 48459 1841 48475 1875
rect 48383 1825 48475 1841
rect 49316 1875 49403 1891
rect 49316 1841 49331 1875
rect 49365 1841 49403 1875
rect 49445 1891 49475 1923
rect 49445 1875 49549 1891
rect 49445 1861 49499 1875
rect 49316 1825 49403 1841
rect 48383 1803 48413 1825
rect 49373 1803 49403 1825
rect 49457 1841 49499 1861
rect 49533 1841 49549 1875
rect 49457 1825 49549 1841
rect 49457 1803 49487 1825
rect 47844 1727 47874 1758
rect 47940 1732 47970 1758
rect 47826 1711 47892 1727
rect 47826 1677 47842 1711
rect 47876 1690 47892 1711
rect 47876 1677 48004 1690
rect 44168 1596 44184 1630
rect 44218 1596 44234 1630
rect 42298 1558 42328 1580
rect 44090 1558 44120 1584
rect 44168 1580 44234 1596
rect 46050 1630 46116 1658
rect 46411 1647 46441 1673
rect 46495 1647 46525 1673
rect 47485 1647 47515 1673
rect 47569 1647 47599 1673
rect 47826 1658 48004 1677
rect 52075 2123 52105 2149
rect 52147 2123 52177 2149
rect 53149 2123 53179 2149
rect 53221 2123 53251 2149
rect 51698 2039 51764 2055
rect 51698 2005 51714 2039
rect 51748 2005 51764 2039
rect 51698 1989 51764 2005
rect 51620 1958 51650 1984
rect 51716 1958 51746 1989
rect 50187 1891 50217 1923
rect 50130 1875 50217 1891
rect 50130 1841 50145 1875
rect 50179 1841 50217 1875
rect 50259 1891 50289 1923
rect 51261 1891 51291 1923
rect 50259 1875 50363 1891
rect 50259 1861 50313 1875
rect 50130 1825 50217 1841
rect 50187 1803 50217 1825
rect 50271 1841 50313 1861
rect 50347 1841 50363 1875
rect 50271 1825 50363 1841
rect 51204 1875 51291 1891
rect 51204 1841 51219 1875
rect 51253 1841 51291 1875
rect 51333 1891 51363 1923
rect 51333 1875 51437 1891
rect 51333 1861 51387 1875
rect 51204 1825 51291 1841
rect 50271 1803 50301 1825
rect 51261 1803 51291 1825
rect 51345 1841 51387 1861
rect 51421 1841 51437 1875
rect 51345 1825 51437 1841
rect 51345 1803 51375 1825
rect 49732 1727 49762 1758
rect 49828 1732 49858 1758
rect 49714 1711 49780 1727
rect 49714 1677 49730 1711
rect 49764 1690 49780 1711
rect 49764 1677 49892 1690
rect 46050 1596 46066 1630
rect 46100 1596 46116 1630
rect 44186 1558 44216 1580
rect 45972 1558 46002 1584
rect 46050 1580 46116 1596
rect 47938 1630 48004 1658
rect 48299 1647 48329 1673
rect 48383 1647 48413 1673
rect 49373 1647 49403 1673
rect 49457 1647 49487 1673
rect 49714 1658 49892 1677
rect 53963 2123 53993 2149
rect 54035 2123 54065 2149
rect 55037 2123 55067 2149
rect 55109 2123 55139 2149
rect 53586 2039 53652 2055
rect 53586 2005 53602 2039
rect 53636 2005 53652 2039
rect 53586 1989 53652 2005
rect 53508 1958 53538 1984
rect 53604 1958 53634 1989
rect 52075 1891 52105 1923
rect 52018 1875 52105 1891
rect 52018 1841 52033 1875
rect 52067 1841 52105 1875
rect 52147 1891 52177 1923
rect 53149 1891 53179 1923
rect 52147 1875 52251 1891
rect 52147 1861 52201 1875
rect 52018 1825 52105 1841
rect 52075 1803 52105 1825
rect 52159 1841 52201 1861
rect 52235 1841 52251 1875
rect 52159 1825 52251 1841
rect 53092 1875 53179 1891
rect 53092 1841 53107 1875
rect 53141 1841 53179 1875
rect 53221 1891 53251 1923
rect 53221 1875 53325 1891
rect 53221 1861 53275 1875
rect 53092 1825 53179 1841
rect 52159 1803 52189 1825
rect 53149 1803 53179 1825
rect 53233 1841 53275 1861
rect 53309 1841 53325 1875
rect 53233 1825 53325 1841
rect 53233 1803 53263 1825
rect 51620 1727 51650 1758
rect 51716 1732 51746 1758
rect 51602 1711 51668 1727
rect 51602 1677 51618 1711
rect 51652 1690 51668 1711
rect 51652 1677 51780 1690
rect 47938 1596 47954 1630
rect 47988 1596 48004 1630
rect 46068 1558 46098 1580
rect 47860 1558 47890 1584
rect 47938 1580 48004 1596
rect 49826 1630 49892 1658
rect 50187 1647 50217 1673
rect 50271 1647 50301 1673
rect 51261 1647 51291 1673
rect 51345 1647 51375 1673
rect 51602 1658 51780 1677
rect 55851 2123 55881 2149
rect 55923 2123 55953 2149
rect 56925 2123 56955 2149
rect 56997 2123 57027 2149
rect 55474 2039 55540 2055
rect 55474 2005 55490 2039
rect 55524 2005 55540 2039
rect 55474 1989 55540 2005
rect 55396 1958 55426 1984
rect 55492 1958 55522 1989
rect 53963 1891 53993 1923
rect 53906 1875 53993 1891
rect 53906 1841 53921 1875
rect 53955 1841 53993 1875
rect 54035 1891 54065 1923
rect 55037 1891 55067 1923
rect 54035 1875 54139 1891
rect 54035 1861 54089 1875
rect 53906 1825 53993 1841
rect 53963 1803 53993 1825
rect 54047 1841 54089 1861
rect 54123 1841 54139 1875
rect 54047 1825 54139 1841
rect 54980 1875 55067 1891
rect 54980 1841 54995 1875
rect 55029 1841 55067 1875
rect 55109 1891 55139 1923
rect 55109 1875 55213 1891
rect 55109 1861 55163 1875
rect 54980 1825 55067 1841
rect 54047 1803 54077 1825
rect 55037 1803 55067 1825
rect 55121 1841 55163 1861
rect 55197 1841 55213 1875
rect 55121 1825 55213 1841
rect 55121 1803 55151 1825
rect 53508 1727 53538 1758
rect 53604 1732 53634 1758
rect 53490 1711 53556 1727
rect 53490 1677 53506 1711
rect 53540 1690 53556 1711
rect 53540 1677 53668 1690
rect 49826 1596 49842 1630
rect 49876 1596 49892 1630
rect 47956 1558 47986 1580
rect 49748 1558 49778 1584
rect 49826 1580 49892 1596
rect 51714 1630 51780 1658
rect 52075 1647 52105 1673
rect 52159 1647 52189 1673
rect 53149 1647 53179 1673
rect 53233 1647 53263 1673
rect 53490 1658 53668 1677
rect 57739 2123 57769 2149
rect 57811 2123 57841 2149
rect 58813 2123 58843 2149
rect 58885 2123 58915 2149
rect 57362 2039 57428 2055
rect 57362 2005 57378 2039
rect 57412 2005 57428 2039
rect 57362 1989 57428 2005
rect 57284 1958 57314 1984
rect 57380 1958 57410 1989
rect 55851 1891 55881 1923
rect 55794 1875 55881 1891
rect 55794 1841 55809 1875
rect 55843 1841 55881 1875
rect 55923 1891 55953 1923
rect 56925 1891 56955 1923
rect 55923 1875 56027 1891
rect 55923 1861 55977 1875
rect 55794 1825 55881 1841
rect 55851 1803 55881 1825
rect 55935 1841 55977 1861
rect 56011 1841 56027 1875
rect 55935 1825 56027 1841
rect 56868 1875 56955 1891
rect 56868 1841 56883 1875
rect 56917 1841 56955 1875
rect 56997 1891 57027 1923
rect 56997 1875 57101 1891
rect 56997 1861 57051 1875
rect 56868 1825 56955 1841
rect 55935 1803 55965 1825
rect 56925 1803 56955 1825
rect 57009 1841 57051 1861
rect 57085 1841 57101 1875
rect 57009 1825 57101 1841
rect 57009 1803 57039 1825
rect 55396 1727 55426 1758
rect 55492 1732 55522 1758
rect 55378 1711 55444 1727
rect 55378 1677 55394 1711
rect 55428 1690 55444 1711
rect 55428 1677 55556 1690
rect 51714 1596 51730 1630
rect 51764 1596 51780 1630
rect 49844 1558 49874 1580
rect 51636 1558 51666 1584
rect 51714 1580 51780 1596
rect 53602 1630 53668 1658
rect 53963 1647 53993 1673
rect 54047 1647 54077 1673
rect 55037 1647 55067 1673
rect 55121 1647 55151 1673
rect 55378 1658 55556 1677
rect 59627 2123 59657 2149
rect 59699 2123 59729 2149
rect 59250 2039 59316 2055
rect 59250 2005 59266 2039
rect 59300 2005 59316 2039
rect 59250 1989 59316 2005
rect 59172 1958 59202 1984
rect 59268 1958 59298 1989
rect 57739 1891 57769 1923
rect 57682 1875 57769 1891
rect 57682 1841 57697 1875
rect 57731 1841 57769 1875
rect 57811 1891 57841 1923
rect 58813 1891 58843 1923
rect 57811 1875 57915 1891
rect 57811 1861 57865 1875
rect 57682 1825 57769 1841
rect 57739 1803 57769 1825
rect 57823 1841 57865 1861
rect 57899 1841 57915 1875
rect 57823 1825 57915 1841
rect 58756 1875 58843 1891
rect 58756 1841 58771 1875
rect 58805 1841 58843 1875
rect 58885 1891 58915 1923
rect 58885 1875 58989 1891
rect 58885 1861 58939 1875
rect 58756 1825 58843 1841
rect 57823 1803 57853 1825
rect 58813 1803 58843 1825
rect 58897 1841 58939 1861
rect 58973 1841 58989 1875
rect 58897 1825 58989 1841
rect 58897 1803 58927 1825
rect 57284 1727 57314 1758
rect 57380 1732 57410 1758
rect 57266 1711 57332 1727
rect 57266 1677 57282 1711
rect 57316 1690 57332 1711
rect 57316 1677 57444 1690
rect 53602 1596 53618 1630
rect 53652 1596 53668 1630
rect 51732 1558 51762 1580
rect 53524 1558 53554 1584
rect 53602 1580 53668 1596
rect 55490 1630 55556 1658
rect 55851 1647 55881 1673
rect 55935 1647 55965 1673
rect 56925 1647 56955 1673
rect 57009 1647 57039 1673
rect 57266 1658 57444 1677
rect 59627 1891 59657 1923
rect 59570 1875 59657 1891
rect 59570 1841 59585 1875
rect 59619 1841 59657 1875
rect 59699 1891 59729 1923
rect 59699 1875 59803 1891
rect 59699 1861 59753 1875
rect 59570 1825 59657 1841
rect 59627 1803 59657 1825
rect 59711 1841 59753 1861
rect 59787 1841 59803 1875
rect 59711 1825 59803 1841
rect 59711 1803 59741 1825
rect 59172 1727 59202 1758
rect 59268 1732 59298 1758
rect 59154 1711 59220 1727
rect 59154 1677 59170 1711
rect 59204 1690 59220 1711
rect 59204 1677 59332 1690
rect 55490 1596 55506 1630
rect 55540 1596 55556 1630
rect 53620 1558 53650 1580
rect 55412 1558 55442 1584
rect 55490 1580 55556 1596
rect 57378 1630 57444 1658
rect 57739 1647 57769 1673
rect 57823 1647 57853 1673
rect 58813 1647 58843 1673
rect 58897 1647 58927 1673
rect 59154 1658 59332 1677
rect 57378 1596 57394 1630
rect 57428 1596 57444 1630
rect 55508 1558 55538 1580
rect 57300 1558 57330 1584
rect 57378 1580 57444 1596
rect 59266 1630 59332 1658
rect 59627 1647 59657 1673
rect 59711 1647 59741 1673
rect 59266 1596 59282 1630
rect 59316 1596 59332 1630
rect 57396 1558 57426 1580
rect 59188 1558 59218 1584
rect 59266 1580 59332 1596
rect 59284 1558 59314 1580
rect 672 1406 702 1428
rect 654 1390 720 1406
rect 654 1356 670 1390
rect 704 1356 720 1390
rect 768 1402 798 1428
rect 2560 1406 2590 1428
rect 768 1372 902 1402
rect 654 1340 720 1356
rect 872 1204 902 1372
rect 2542 1390 2608 1406
rect 2542 1356 2558 1390
rect 2592 1356 2608 1390
rect 2656 1402 2686 1428
rect 4448 1406 4478 1428
rect 2656 1372 2790 1402
rect 2542 1340 2608 1356
rect 2760 1204 2790 1372
rect 4430 1390 4496 1406
rect 4430 1356 4446 1390
rect 4480 1356 4496 1390
rect 4544 1402 4574 1428
rect 6336 1406 6366 1428
rect 4544 1372 4678 1402
rect 4430 1340 4496 1356
rect 4648 1204 4678 1372
rect 6318 1390 6384 1406
rect 6318 1356 6334 1390
rect 6368 1356 6384 1390
rect 6432 1402 6462 1428
rect 8224 1406 8254 1428
rect 6432 1372 6566 1402
rect 6318 1340 6384 1356
rect 6536 1204 6566 1372
rect 8206 1390 8272 1406
rect 8206 1356 8222 1390
rect 8256 1356 8272 1390
rect 8320 1402 8350 1428
rect 10112 1406 10142 1428
rect 8320 1372 8454 1402
rect 8206 1340 8272 1356
rect 8424 1204 8454 1372
rect 10094 1390 10160 1406
rect 10094 1356 10110 1390
rect 10144 1356 10160 1390
rect 10208 1402 10238 1428
rect 12000 1406 12030 1428
rect 10208 1372 10342 1402
rect 10094 1340 10160 1356
rect 10312 1204 10342 1372
rect 11982 1390 12048 1406
rect 11982 1356 11998 1390
rect 12032 1356 12048 1390
rect 12096 1402 12126 1428
rect 13888 1406 13918 1428
rect 12096 1372 12230 1402
rect 11982 1340 12048 1356
rect 12200 1204 12230 1372
rect 13870 1390 13936 1406
rect 13870 1356 13886 1390
rect 13920 1356 13936 1390
rect 13984 1402 14014 1428
rect 15770 1406 15800 1428
rect 13984 1372 14118 1402
rect 13870 1340 13936 1356
rect 14088 1204 14118 1372
rect 15752 1390 15818 1406
rect 15752 1356 15768 1390
rect 15802 1356 15818 1390
rect 15866 1402 15896 1428
rect 17658 1406 17688 1428
rect 15866 1372 16000 1402
rect 15752 1340 15818 1356
rect 15970 1204 16000 1372
rect 17640 1390 17706 1406
rect 17640 1356 17656 1390
rect 17690 1356 17706 1390
rect 17754 1402 17784 1428
rect 19546 1406 19576 1428
rect 17754 1372 17888 1402
rect 17640 1340 17706 1356
rect 17858 1204 17888 1372
rect 19528 1390 19594 1406
rect 19528 1356 19544 1390
rect 19578 1356 19594 1390
rect 19642 1402 19672 1428
rect 21434 1406 21464 1428
rect 19642 1372 19776 1402
rect 19528 1340 19594 1356
rect 19746 1204 19776 1372
rect 21416 1390 21482 1406
rect 21416 1356 21432 1390
rect 21466 1356 21482 1390
rect 21530 1402 21560 1428
rect 23322 1406 23352 1428
rect 21530 1372 21664 1402
rect 21416 1340 21482 1356
rect 21634 1204 21664 1372
rect 23304 1390 23370 1406
rect 23304 1356 23320 1390
rect 23354 1356 23370 1390
rect 23418 1402 23448 1428
rect 25210 1406 25240 1428
rect 23418 1372 23552 1402
rect 23304 1340 23370 1356
rect 23522 1204 23552 1372
rect 25192 1390 25258 1406
rect 25192 1356 25208 1390
rect 25242 1356 25258 1390
rect 25306 1402 25336 1428
rect 27098 1406 27128 1428
rect 25306 1372 25440 1402
rect 25192 1340 25258 1356
rect 25410 1204 25440 1372
rect 27080 1390 27146 1406
rect 27080 1356 27096 1390
rect 27130 1356 27146 1390
rect 27194 1402 27224 1428
rect 28986 1406 29016 1428
rect 27194 1372 27328 1402
rect 27080 1340 27146 1356
rect 27298 1204 27328 1372
rect 28968 1390 29034 1406
rect 28968 1356 28984 1390
rect 29018 1356 29034 1390
rect 29082 1402 29112 1428
rect 30874 1406 30904 1428
rect 29082 1372 29216 1402
rect 28968 1340 29034 1356
rect 29186 1204 29216 1372
rect 30856 1390 30922 1406
rect 30856 1356 30872 1390
rect 30906 1356 30922 1390
rect 30970 1402 31000 1428
rect 32762 1406 32792 1428
rect 30970 1372 31104 1402
rect 30856 1340 30922 1356
rect 31074 1204 31104 1372
rect 32744 1390 32810 1406
rect 32744 1356 32760 1390
rect 32794 1356 32810 1390
rect 32858 1402 32888 1428
rect 34650 1406 34680 1428
rect 32858 1372 32992 1402
rect 32744 1340 32810 1356
rect 32962 1204 32992 1372
rect 34632 1390 34698 1406
rect 34632 1356 34648 1390
rect 34682 1356 34698 1390
rect 34746 1402 34776 1428
rect 36538 1406 36568 1428
rect 34746 1372 34880 1402
rect 34632 1340 34698 1356
rect 34850 1204 34880 1372
rect 36520 1390 36586 1406
rect 36520 1356 36536 1390
rect 36570 1356 36586 1390
rect 36634 1402 36664 1428
rect 38426 1406 38456 1428
rect 36634 1372 36768 1402
rect 36520 1340 36586 1356
rect 36738 1204 36768 1372
rect 38408 1390 38474 1406
rect 38408 1356 38424 1390
rect 38458 1356 38474 1390
rect 38522 1402 38552 1428
rect 40314 1406 40344 1428
rect 38522 1372 38656 1402
rect 38408 1340 38474 1356
rect 38626 1204 38656 1372
rect 40296 1390 40362 1406
rect 40296 1356 40312 1390
rect 40346 1356 40362 1390
rect 40410 1402 40440 1428
rect 42202 1406 42232 1428
rect 40410 1372 40544 1402
rect 40296 1340 40362 1356
rect 40514 1204 40544 1372
rect 42184 1390 42250 1406
rect 42184 1356 42200 1390
rect 42234 1356 42250 1390
rect 42298 1402 42328 1428
rect 44090 1406 44120 1428
rect 42298 1372 42432 1402
rect 42184 1340 42250 1356
rect 42402 1204 42432 1372
rect 44072 1390 44138 1406
rect 44072 1356 44088 1390
rect 44122 1356 44138 1390
rect 44186 1402 44216 1428
rect 45972 1406 46002 1428
rect 44186 1372 44320 1402
rect 44072 1340 44138 1356
rect 44290 1204 44320 1372
rect 45954 1390 46020 1406
rect 45954 1356 45970 1390
rect 46004 1356 46020 1390
rect 46068 1402 46098 1428
rect 47860 1406 47890 1428
rect 46068 1372 46202 1402
rect 45954 1340 46020 1356
rect 46172 1204 46202 1372
rect 47842 1390 47908 1406
rect 47842 1356 47858 1390
rect 47892 1356 47908 1390
rect 47956 1402 47986 1428
rect 49748 1406 49778 1428
rect 47956 1372 48090 1402
rect 47842 1340 47908 1356
rect 48060 1204 48090 1372
rect 49730 1390 49796 1406
rect 49730 1356 49746 1390
rect 49780 1356 49796 1390
rect 49844 1402 49874 1428
rect 51636 1406 51666 1428
rect 49844 1372 49978 1402
rect 49730 1340 49796 1356
rect 49948 1204 49978 1372
rect 51618 1390 51684 1406
rect 51618 1356 51634 1390
rect 51668 1356 51684 1390
rect 51732 1402 51762 1428
rect 53524 1406 53554 1428
rect 51732 1372 51866 1402
rect 51618 1340 51684 1356
rect 51836 1204 51866 1372
rect 53506 1390 53572 1406
rect 53506 1356 53522 1390
rect 53556 1356 53572 1390
rect 53620 1402 53650 1428
rect 55412 1406 55442 1428
rect 53620 1372 53754 1402
rect 53506 1340 53572 1356
rect 53724 1204 53754 1372
rect 55394 1390 55460 1406
rect 55394 1356 55410 1390
rect 55444 1356 55460 1390
rect 55508 1402 55538 1428
rect 57300 1406 57330 1428
rect 55508 1372 55642 1402
rect 55394 1340 55460 1356
rect 55612 1204 55642 1372
rect 57282 1390 57348 1406
rect 57282 1356 57298 1390
rect 57332 1356 57348 1390
rect 57396 1402 57426 1428
rect 59188 1406 59218 1428
rect 57396 1372 57530 1402
rect 57282 1340 57348 1356
rect 57500 1204 57530 1372
rect 59170 1390 59236 1406
rect 59170 1356 59186 1390
rect 59220 1356 59236 1390
rect 59284 1402 59314 1428
rect 59284 1372 59418 1402
rect 59170 1340 59236 1356
rect 59388 1204 59418 1372
rect 598 1174 1080 1204
rect 416 1143 482 1159
rect 416 1109 432 1143
rect 466 1109 482 1143
rect 160 1069 190 1095
rect 416 1093 482 1109
rect 434 1062 464 1093
rect 160 837 190 869
rect 598 1016 628 1174
rect 1048 1159 1080 1174
rect 2486 1174 2968 1204
rect 1048 1143 1128 1159
rect 1048 1109 1078 1143
rect 1112 1109 1128 1143
rect 1048 1093 1128 1109
rect 2304 1143 2370 1159
rect 2304 1109 2320 1143
rect 2354 1109 2370 1143
rect 1048 1092 1110 1093
rect 1080 1062 1110 1092
rect 1356 1077 1386 1103
rect 598 986 684 1016
rect 654 902 684 986
rect 732 983 798 999
rect 732 949 748 983
rect 782 949 798 983
rect 732 933 798 949
rect 750 902 780 933
rect 104 821 190 837
rect 434 831 464 862
rect 104 787 120 821
rect 154 787 190 821
rect 104 771 190 787
rect 160 749 190 771
rect 416 815 482 831
rect 416 781 432 815
rect 466 781 482 815
rect 416 765 482 781
rect 1661 1075 1691 1101
rect 1749 1075 1779 1101
rect 2048 1069 2078 1095
rect 2304 1093 2370 1109
rect 1661 902 1691 917
rect 1655 878 1691 902
rect 1080 831 1110 862
rect 1356 845 1386 877
rect 1062 815 1128 831
rect 1062 781 1078 815
rect 1112 781 1128 815
rect 1062 765 1128 781
rect 1300 829 1386 845
rect 1655 843 1685 878
rect 1749 856 1779 917
rect 2322 1062 2352 1093
rect 1300 795 1316 829
rect 1350 795 1386 829
rect 1300 779 1386 795
rect 1356 757 1386 779
rect 1609 827 1685 843
rect 1609 793 1619 827
rect 1653 793 1685 827
rect 1609 777 1685 793
rect 1727 840 1781 856
rect 1727 806 1737 840
rect 1771 806 1781 840
rect 2048 837 2078 869
rect 2486 1016 2516 1174
rect 2936 1159 2968 1174
rect 4374 1174 4856 1204
rect 2936 1143 3016 1159
rect 2936 1109 2966 1143
rect 3000 1109 3016 1143
rect 2936 1093 3016 1109
rect 4192 1143 4258 1159
rect 4192 1109 4208 1143
rect 4242 1109 4258 1143
rect 2936 1092 2998 1093
rect 2968 1062 2998 1092
rect 3244 1077 3274 1103
rect 2486 986 2572 1016
rect 2542 902 2572 986
rect 2620 983 2686 999
rect 2620 949 2636 983
rect 2670 949 2686 983
rect 2620 933 2686 949
rect 2638 902 2668 933
rect 1727 790 1781 806
rect 1992 821 2078 837
rect 2322 831 2352 862
rect 1655 768 1685 777
rect 654 671 684 702
rect 750 676 780 702
rect 636 655 702 671
rect 636 621 652 655
rect 686 634 702 655
rect 686 621 814 634
rect 1655 744 1691 768
rect 1661 729 1691 744
rect 1749 729 1779 790
rect 1992 787 2008 821
rect 2042 787 2078 821
rect 1992 771 2078 787
rect 2048 749 2078 771
rect 2304 815 2370 831
rect 2304 781 2320 815
rect 2354 781 2370 815
rect 2304 765 2370 781
rect 160 593 190 619
rect 636 602 814 621
rect 748 574 814 602
rect 1356 601 1386 627
rect 1661 599 1691 625
rect 1749 599 1779 625
rect 3549 1075 3579 1101
rect 3637 1075 3667 1101
rect 3936 1069 3966 1095
rect 4192 1093 4258 1109
rect 3549 902 3579 917
rect 3543 878 3579 902
rect 2968 831 2998 862
rect 3244 845 3274 877
rect 2950 815 3016 831
rect 2950 781 2966 815
rect 3000 781 3016 815
rect 2950 765 3016 781
rect 3188 829 3274 845
rect 3543 843 3573 878
rect 3637 856 3667 917
rect 4210 1062 4240 1093
rect 3188 795 3204 829
rect 3238 795 3274 829
rect 3188 779 3274 795
rect 3244 757 3274 779
rect 3497 827 3573 843
rect 3497 793 3507 827
rect 3541 793 3573 827
rect 3497 777 3573 793
rect 3615 840 3669 856
rect 3615 806 3625 840
rect 3659 806 3669 840
rect 3936 837 3966 869
rect 4374 1016 4404 1174
rect 4824 1159 4856 1174
rect 6262 1174 6744 1204
rect 4824 1143 4904 1159
rect 4824 1109 4854 1143
rect 4888 1109 4904 1143
rect 4824 1093 4904 1109
rect 6080 1143 6146 1159
rect 6080 1109 6096 1143
rect 6130 1109 6146 1143
rect 4824 1092 4886 1093
rect 4856 1062 4886 1092
rect 5132 1077 5162 1103
rect 4374 986 4460 1016
rect 4430 902 4460 986
rect 4508 983 4574 999
rect 4508 949 4524 983
rect 4558 949 4574 983
rect 4508 933 4574 949
rect 4526 902 4556 933
rect 3615 790 3669 806
rect 3880 821 3966 837
rect 4210 831 4240 862
rect 3543 768 3573 777
rect 2542 671 2572 702
rect 2638 676 2668 702
rect 2524 655 2590 671
rect 2524 621 2540 655
rect 2574 634 2590 655
rect 2574 621 2702 634
rect 3543 744 3579 768
rect 3549 729 3579 744
rect 3637 729 3667 790
rect 3880 787 3896 821
rect 3930 787 3966 821
rect 3880 771 3966 787
rect 3936 749 3966 771
rect 4192 815 4258 831
rect 4192 781 4208 815
rect 4242 781 4258 815
rect 4192 765 4258 781
rect 2048 593 2078 619
rect 2524 602 2702 621
rect 748 540 764 574
rect 798 540 814 574
rect 670 502 700 528
rect 748 524 814 540
rect 2636 574 2702 602
rect 3244 601 3274 627
rect 3549 599 3579 625
rect 3637 599 3667 625
rect 5437 1075 5467 1101
rect 5525 1075 5555 1101
rect 5824 1069 5854 1095
rect 6080 1093 6146 1109
rect 5437 902 5467 917
rect 5431 878 5467 902
rect 4856 831 4886 862
rect 5132 845 5162 877
rect 4838 815 4904 831
rect 4838 781 4854 815
rect 4888 781 4904 815
rect 4838 765 4904 781
rect 5076 829 5162 845
rect 5431 843 5461 878
rect 5525 856 5555 917
rect 6098 1062 6128 1093
rect 5076 795 5092 829
rect 5126 795 5162 829
rect 5076 779 5162 795
rect 5132 757 5162 779
rect 5385 827 5461 843
rect 5385 793 5395 827
rect 5429 793 5461 827
rect 5385 777 5461 793
rect 5503 840 5557 856
rect 5503 806 5513 840
rect 5547 806 5557 840
rect 5824 837 5854 869
rect 6262 1016 6292 1174
rect 6712 1159 6744 1174
rect 8150 1174 8632 1204
rect 6712 1143 6792 1159
rect 6712 1109 6742 1143
rect 6776 1109 6792 1143
rect 6712 1093 6792 1109
rect 7968 1143 8034 1159
rect 7968 1109 7984 1143
rect 8018 1109 8034 1143
rect 6712 1092 6774 1093
rect 6744 1062 6774 1092
rect 7020 1077 7050 1103
rect 6262 986 6348 1016
rect 6318 902 6348 986
rect 6396 983 6462 999
rect 6396 949 6412 983
rect 6446 949 6462 983
rect 6396 933 6462 949
rect 6414 902 6444 933
rect 5503 790 5557 806
rect 5768 821 5854 837
rect 6098 831 6128 862
rect 5431 768 5461 777
rect 4430 671 4460 702
rect 4526 676 4556 702
rect 4412 655 4478 671
rect 4412 621 4428 655
rect 4462 634 4478 655
rect 4462 621 4590 634
rect 5431 744 5467 768
rect 5437 729 5467 744
rect 5525 729 5555 790
rect 5768 787 5784 821
rect 5818 787 5854 821
rect 5768 771 5854 787
rect 5824 749 5854 771
rect 6080 815 6146 831
rect 6080 781 6096 815
rect 6130 781 6146 815
rect 6080 765 6146 781
rect 3936 593 3966 619
rect 4412 602 4590 621
rect 2636 540 2652 574
rect 2686 540 2702 574
rect 766 502 796 524
rect 2558 502 2588 528
rect 2636 524 2702 540
rect 4524 574 4590 602
rect 5132 601 5162 627
rect 5437 599 5467 625
rect 5525 599 5555 625
rect 7325 1075 7355 1101
rect 7413 1075 7443 1101
rect 7712 1069 7742 1095
rect 7968 1093 8034 1109
rect 7325 902 7355 917
rect 7319 878 7355 902
rect 6744 831 6774 862
rect 7020 845 7050 877
rect 6726 815 6792 831
rect 6726 781 6742 815
rect 6776 781 6792 815
rect 6726 765 6792 781
rect 6964 829 7050 845
rect 7319 843 7349 878
rect 7413 856 7443 917
rect 7986 1062 8016 1093
rect 6964 795 6980 829
rect 7014 795 7050 829
rect 6964 779 7050 795
rect 7020 757 7050 779
rect 7273 827 7349 843
rect 7273 793 7283 827
rect 7317 793 7349 827
rect 7273 777 7349 793
rect 7391 840 7445 856
rect 7391 806 7401 840
rect 7435 806 7445 840
rect 7712 837 7742 869
rect 8150 1016 8180 1174
rect 8600 1159 8632 1174
rect 10038 1174 10520 1204
rect 8600 1143 8680 1159
rect 8600 1109 8630 1143
rect 8664 1109 8680 1143
rect 8600 1093 8680 1109
rect 9856 1143 9922 1159
rect 9856 1109 9872 1143
rect 9906 1109 9922 1143
rect 8600 1092 8662 1093
rect 8632 1062 8662 1092
rect 8908 1077 8938 1103
rect 8150 986 8236 1016
rect 8206 902 8236 986
rect 8284 983 8350 999
rect 8284 949 8300 983
rect 8334 949 8350 983
rect 8284 933 8350 949
rect 8302 902 8332 933
rect 7391 790 7445 806
rect 7656 821 7742 837
rect 7986 831 8016 862
rect 7319 768 7349 777
rect 6318 671 6348 702
rect 6414 676 6444 702
rect 6300 655 6366 671
rect 6300 621 6316 655
rect 6350 634 6366 655
rect 6350 621 6478 634
rect 7319 744 7355 768
rect 7325 729 7355 744
rect 7413 729 7443 790
rect 7656 787 7672 821
rect 7706 787 7742 821
rect 7656 771 7742 787
rect 7712 749 7742 771
rect 7968 815 8034 831
rect 7968 781 7984 815
rect 8018 781 8034 815
rect 7968 765 8034 781
rect 5824 593 5854 619
rect 6300 602 6478 621
rect 4524 540 4540 574
rect 4574 540 4590 574
rect 2654 502 2684 524
rect 4446 502 4476 528
rect 4524 524 4590 540
rect 6412 574 6478 602
rect 7020 601 7050 627
rect 7325 599 7355 625
rect 7413 599 7443 625
rect 9213 1075 9243 1101
rect 9301 1075 9331 1101
rect 9600 1069 9630 1095
rect 9856 1093 9922 1109
rect 9213 902 9243 917
rect 9207 878 9243 902
rect 8632 831 8662 862
rect 8908 845 8938 877
rect 8614 815 8680 831
rect 8614 781 8630 815
rect 8664 781 8680 815
rect 8614 765 8680 781
rect 8852 829 8938 845
rect 9207 843 9237 878
rect 9301 856 9331 917
rect 9874 1062 9904 1093
rect 8852 795 8868 829
rect 8902 795 8938 829
rect 8852 779 8938 795
rect 8908 757 8938 779
rect 9161 827 9237 843
rect 9161 793 9171 827
rect 9205 793 9237 827
rect 9161 777 9237 793
rect 9279 840 9333 856
rect 9279 806 9289 840
rect 9323 806 9333 840
rect 9600 837 9630 869
rect 10038 1016 10068 1174
rect 10488 1159 10520 1174
rect 11926 1174 12408 1204
rect 10488 1143 10568 1159
rect 10488 1109 10518 1143
rect 10552 1109 10568 1143
rect 10488 1093 10568 1109
rect 11744 1143 11810 1159
rect 11744 1109 11760 1143
rect 11794 1109 11810 1143
rect 10488 1092 10550 1093
rect 10520 1062 10550 1092
rect 10796 1077 10826 1103
rect 10038 986 10124 1016
rect 10094 902 10124 986
rect 10172 983 10238 999
rect 10172 949 10188 983
rect 10222 949 10238 983
rect 10172 933 10238 949
rect 10190 902 10220 933
rect 9279 790 9333 806
rect 9544 821 9630 837
rect 9874 831 9904 862
rect 9207 768 9237 777
rect 8206 671 8236 702
rect 8302 676 8332 702
rect 8188 655 8254 671
rect 8188 621 8204 655
rect 8238 634 8254 655
rect 8238 621 8366 634
rect 9207 744 9243 768
rect 9213 729 9243 744
rect 9301 729 9331 790
rect 9544 787 9560 821
rect 9594 787 9630 821
rect 9544 771 9630 787
rect 9600 749 9630 771
rect 9856 815 9922 831
rect 9856 781 9872 815
rect 9906 781 9922 815
rect 9856 765 9922 781
rect 7712 593 7742 619
rect 8188 602 8366 621
rect 6412 540 6428 574
rect 6462 540 6478 574
rect 4542 502 4572 524
rect 6334 502 6364 528
rect 6412 524 6478 540
rect 8300 574 8366 602
rect 8908 601 8938 627
rect 9213 599 9243 625
rect 9301 599 9331 625
rect 11101 1075 11131 1101
rect 11189 1075 11219 1101
rect 11488 1069 11518 1095
rect 11744 1093 11810 1109
rect 11101 902 11131 917
rect 11095 878 11131 902
rect 10520 831 10550 862
rect 10796 845 10826 877
rect 10502 815 10568 831
rect 10502 781 10518 815
rect 10552 781 10568 815
rect 10502 765 10568 781
rect 10740 829 10826 845
rect 11095 843 11125 878
rect 11189 856 11219 917
rect 11762 1062 11792 1093
rect 10740 795 10756 829
rect 10790 795 10826 829
rect 10740 779 10826 795
rect 10796 757 10826 779
rect 11049 827 11125 843
rect 11049 793 11059 827
rect 11093 793 11125 827
rect 11049 777 11125 793
rect 11167 840 11221 856
rect 11167 806 11177 840
rect 11211 806 11221 840
rect 11488 837 11518 869
rect 11926 1016 11956 1174
rect 12376 1159 12408 1174
rect 13814 1174 14296 1204
rect 12376 1143 12456 1159
rect 12376 1109 12406 1143
rect 12440 1109 12456 1143
rect 12376 1093 12456 1109
rect 13632 1143 13698 1159
rect 13632 1109 13648 1143
rect 13682 1109 13698 1143
rect 12376 1092 12438 1093
rect 12408 1062 12438 1092
rect 12684 1077 12714 1103
rect 11926 986 12012 1016
rect 11982 902 12012 986
rect 12060 983 12126 999
rect 12060 949 12076 983
rect 12110 949 12126 983
rect 12060 933 12126 949
rect 12078 902 12108 933
rect 11167 790 11221 806
rect 11432 821 11518 837
rect 11762 831 11792 862
rect 11095 768 11125 777
rect 10094 671 10124 702
rect 10190 676 10220 702
rect 10076 655 10142 671
rect 10076 621 10092 655
rect 10126 634 10142 655
rect 10126 621 10254 634
rect 11095 744 11131 768
rect 11101 729 11131 744
rect 11189 729 11219 790
rect 11432 787 11448 821
rect 11482 787 11518 821
rect 11432 771 11518 787
rect 11488 749 11518 771
rect 11744 815 11810 831
rect 11744 781 11760 815
rect 11794 781 11810 815
rect 11744 765 11810 781
rect 9600 593 9630 619
rect 10076 602 10254 621
rect 8300 540 8316 574
rect 8350 540 8366 574
rect 6430 502 6460 524
rect 8222 502 8252 528
rect 8300 524 8366 540
rect 10188 574 10254 602
rect 10796 601 10826 627
rect 11101 599 11131 625
rect 11189 599 11219 625
rect 12989 1075 13019 1101
rect 13077 1075 13107 1101
rect 13376 1069 13406 1095
rect 13632 1093 13698 1109
rect 12989 902 13019 917
rect 12983 878 13019 902
rect 12408 831 12438 862
rect 12684 845 12714 877
rect 12390 815 12456 831
rect 12390 781 12406 815
rect 12440 781 12456 815
rect 12390 765 12456 781
rect 12628 829 12714 845
rect 12983 843 13013 878
rect 13077 856 13107 917
rect 13650 1062 13680 1093
rect 12628 795 12644 829
rect 12678 795 12714 829
rect 12628 779 12714 795
rect 12684 757 12714 779
rect 12937 827 13013 843
rect 12937 793 12947 827
rect 12981 793 13013 827
rect 12937 777 13013 793
rect 13055 840 13109 856
rect 13055 806 13065 840
rect 13099 806 13109 840
rect 13376 837 13406 869
rect 13814 1016 13844 1174
rect 14264 1159 14296 1174
rect 15696 1174 16178 1204
rect 14264 1143 14344 1159
rect 14264 1109 14294 1143
rect 14328 1109 14344 1143
rect 14264 1093 14344 1109
rect 15514 1143 15580 1159
rect 15514 1109 15530 1143
rect 15564 1109 15580 1143
rect 14264 1092 14326 1093
rect 14296 1062 14326 1092
rect 14572 1077 14602 1103
rect 13814 986 13900 1016
rect 13870 902 13900 986
rect 13948 983 14014 999
rect 13948 949 13964 983
rect 13998 949 14014 983
rect 13948 933 14014 949
rect 13966 902 13996 933
rect 13055 790 13109 806
rect 13320 821 13406 837
rect 13650 831 13680 862
rect 12983 768 13013 777
rect 11982 671 12012 702
rect 12078 676 12108 702
rect 11964 655 12030 671
rect 11964 621 11980 655
rect 12014 634 12030 655
rect 12014 621 12142 634
rect 12983 744 13019 768
rect 12989 729 13019 744
rect 13077 729 13107 790
rect 13320 787 13336 821
rect 13370 787 13406 821
rect 13320 771 13406 787
rect 13376 749 13406 771
rect 13632 815 13698 831
rect 13632 781 13648 815
rect 13682 781 13698 815
rect 13632 765 13698 781
rect 11488 593 11518 619
rect 11964 602 12142 621
rect 10188 540 10204 574
rect 10238 540 10254 574
rect 8318 502 8348 524
rect 10110 502 10140 528
rect 10188 524 10254 540
rect 12076 574 12142 602
rect 12684 601 12714 627
rect 12989 599 13019 625
rect 13077 599 13107 625
rect 14877 1075 14907 1101
rect 14965 1075 14995 1101
rect 15258 1069 15288 1095
rect 15514 1093 15580 1109
rect 14877 902 14907 917
rect 14871 878 14907 902
rect 14296 831 14326 862
rect 14572 845 14602 877
rect 14278 815 14344 831
rect 14278 781 14294 815
rect 14328 781 14344 815
rect 14278 765 14344 781
rect 14516 829 14602 845
rect 14871 843 14901 878
rect 14965 856 14995 917
rect 15532 1062 15562 1093
rect 14516 795 14532 829
rect 14566 795 14602 829
rect 14516 779 14602 795
rect 14572 757 14602 779
rect 14825 827 14901 843
rect 14825 793 14835 827
rect 14869 793 14901 827
rect 14825 777 14901 793
rect 14943 840 14997 856
rect 14943 806 14953 840
rect 14987 806 14997 840
rect 15258 837 15288 869
rect 15696 1016 15726 1174
rect 16146 1159 16178 1174
rect 17584 1174 18066 1204
rect 16146 1143 16226 1159
rect 16146 1109 16176 1143
rect 16210 1109 16226 1143
rect 16146 1093 16226 1109
rect 17402 1143 17468 1159
rect 17402 1109 17418 1143
rect 17452 1109 17468 1143
rect 16146 1092 16208 1093
rect 16178 1062 16208 1092
rect 16454 1077 16484 1103
rect 15696 986 15782 1016
rect 15752 902 15782 986
rect 15830 983 15896 999
rect 15830 949 15846 983
rect 15880 949 15896 983
rect 15830 933 15896 949
rect 15848 902 15878 933
rect 14943 790 14997 806
rect 15202 821 15288 837
rect 15532 831 15562 862
rect 14871 768 14901 777
rect 13870 671 13900 702
rect 13966 676 13996 702
rect 13852 655 13918 671
rect 13852 621 13868 655
rect 13902 634 13918 655
rect 13902 621 14030 634
rect 14871 744 14907 768
rect 14877 729 14907 744
rect 14965 729 14995 790
rect 15202 787 15218 821
rect 15252 787 15288 821
rect 15202 771 15288 787
rect 15258 749 15288 771
rect 15514 815 15580 831
rect 15514 781 15530 815
rect 15564 781 15580 815
rect 15514 765 15580 781
rect 13376 593 13406 619
rect 13852 602 14030 621
rect 12076 540 12092 574
rect 12126 540 12142 574
rect 10206 502 10236 524
rect 11998 502 12028 528
rect 12076 524 12142 540
rect 13964 574 14030 602
rect 14572 601 14602 627
rect 14877 599 14907 625
rect 14965 599 14995 625
rect 16759 1075 16789 1101
rect 16847 1075 16877 1101
rect 17146 1069 17176 1095
rect 17402 1093 17468 1109
rect 16759 902 16789 917
rect 16753 878 16789 902
rect 16178 831 16208 862
rect 16454 845 16484 877
rect 16160 815 16226 831
rect 16160 781 16176 815
rect 16210 781 16226 815
rect 16160 765 16226 781
rect 16398 829 16484 845
rect 16753 843 16783 878
rect 16847 856 16877 917
rect 17420 1062 17450 1093
rect 16398 795 16414 829
rect 16448 795 16484 829
rect 16398 779 16484 795
rect 16454 757 16484 779
rect 16707 827 16783 843
rect 16707 793 16717 827
rect 16751 793 16783 827
rect 16707 777 16783 793
rect 16825 840 16879 856
rect 16825 806 16835 840
rect 16869 806 16879 840
rect 17146 837 17176 869
rect 17584 1016 17614 1174
rect 18034 1159 18066 1174
rect 19472 1174 19954 1204
rect 18034 1143 18114 1159
rect 18034 1109 18064 1143
rect 18098 1109 18114 1143
rect 18034 1093 18114 1109
rect 19290 1143 19356 1159
rect 19290 1109 19306 1143
rect 19340 1109 19356 1143
rect 18034 1092 18096 1093
rect 18066 1062 18096 1092
rect 18342 1077 18372 1103
rect 17584 986 17670 1016
rect 17640 902 17670 986
rect 17718 983 17784 999
rect 17718 949 17734 983
rect 17768 949 17784 983
rect 17718 933 17784 949
rect 17736 902 17766 933
rect 16825 790 16879 806
rect 17090 821 17176 837
rect 17420 831 17450 862
rect 16753 768 16783 777
rect 15752 671 15782 702
rect 15848 676 15878 702
rect 15734 655 15800 671
rect 15734 621 15750 655
rect 15784 634 15800 655
rect 15784 621 15912 634
rect 16753 744 16789 768
rect 16759 729 16789 744
rect 16847 729 16877 790
rect 17090 787 17106 821
rect 17140 787 17176 821
rect 17090 771 17176 787
rect 17146 749 17176 771
rect 17402 815 17468 831
rect 17402 781 17418 815
rect 17452 781 17468 815
rect 17402 765 17468 781
rect 15258 593 15288 619
rect 15734 602 15912 621
rect 13964 540 13980 574
rect 14014 540 14030 574
rect 12094 502 12124 524
rect 13886 502 13916 528
rect 13964 524 14030 540
rect 15846 574 15912 602
rect 16454 601 16484 627
rect 16759 599 16789 625
rect 16847 599 16877 625
rect 18647 1075 18677 1101
rect 18735 1075 18765 1101
rect 19034 1069 19064 1095
rect 19290 1093 19356 1109
rect 18647 902 18677 917
rect 18641 878 18677 902
rect 18066 831 18096 862
rect 18342 845 18372 877
rect 18048 815 18114 831
rect 18048 781 18064 815
rect 18098 781 18114 815
rect 18048 765 18114 781
rect 18286 829 18372 845
rect 18641 843 18671 878
rect 18735 856 18765 917
rect 19308 1062 19338 1093
rect 18286 795 18302 829
rect 18336 795 18372 829
rect 18286 779 18372 795
rect 18342 757 18372 779
rect 18595 827 18671 843
rect 18595 793 18605 827
rect 18639 793 18671 827
rect 18595 777 18671 793
rect 18713 840 18767 856
rect 18713 806 18723 840
rect 18757 806 18767 840
rect 19034 837 19064 869
rect 19472 1016 19502 1174
rect 19922 1159 19954 1174
rect 21360 1174 21842 1204
rect 19922 1143 20002 1159
rect 19922 1109 19952 1143
rect 19986 1109 20002 1143
rect 19922 1093 20002 1109
rect 21178 1143 21244 1159
rect 21178 1109 21194 1143
rect 21228 1109 21244 1143
rect 19922 1092 19984 1093
rect 19954 1062 19984 1092
rect 20230 1077 20260 1103
rect 19472 986 19558 1016
rect 19528 902 19558 986
rect 19606 983 19672 999
rect 19606 949 19622 983
rect 19656 949 19672 983
rect 19606 933 19672 949
rect 19624 902 19654 933
rect 18713 790 18767 806
rect 18978 821 19064 837
rect 19308 831 19338 862
rect 18641 768 18671 777
rect 17640 671 17670 702
rect 17736 676 17766 702
rect 17622 655 17688 671
rect 17622 621 17638 655
rect 17672 634 17688 655
rect 17672 621 17800 634
rect 18641 744 18677 768
rect 18647 729 18677 744
rect 18735 729 18765 790
rect 18978 787 18994 821
rect 19028 787 19064 821
rect 18978 771 19064 787
rect 19034 749 19064 771
rect 19290 815 19356 831
rect 19290 781 19306 815
rect 19340 781 19356 815
rect 19290 765 19356 781
rect 17146 593 17176 619
rect 17622 602 17800 621
rect 15846 540 15862 574
rect 15896 540 15912 574
rect 13982 502 14012 524
rect 15768 502 15798 528
rect 15846 524 15912 540
rect 17734 574 17800 602
rect 18342 601 18372 627
rect 18647 599 18677 625
rect 18735 599 18765 625
rect 20535 1075 20565 1101
rect 20623 1075 20653 1101
rect 20922 1069 20952 1095
rect 21178 1093 21244 1109
rect 20535 902 20565 917
rect 20529 878 20565 902
rect 19954 831 19984 862
rect 20230 845 20260 877
rect 19936 815 20002 831
rect 19936 781 19952 815
rect 19986 781 20002 815
rect 19936 765 20002 781
rect 20174 829 20260 845
rect 20529 843 20559 878
rect 20623 856 20653 917
rect 21196 1062 21226 1093
rect 20174 795 20190 829
rect 20224 795 20260 829
rect 20174 779 20260 795
rect 20230 757 20260 779
rect 20483 827 20559 843
rect 20483 793 20493 827
rect 20527 793 20559 827
rect 20483 777 20559 793
rect 20601 840 20655 856
rect 20601 806 20611 840
rect 20645 806 20655 840
rect 20922 837 20952 869
rect 21360 1016 21390 1174
rect 21810 1159 21842 1174
rect 23248 1174 23730 1204
rect 21810 1143 21890 1159
rect 21810 1109 21840 1143
rect 21874 1109 21890 1143
rect 21810 1093 21890 1109
rect 23066 1143 23132 1159
rect 23066 1109 23082 1143
rect 23116 1109 23132 1143
rect 21810 1092 21872 1093
rect 21842 1062 21872 1092
rect 22118 1077 22148 1103
rect 21360 986 21446 1016
rect 21416 902 21446 986
rect 21494 983 21560 999
rect 21494 949 21510 983
rect 21544 949 21560 983
rect 21494 933 21560 949
rect 21512 902 21542 933
rect 20601 790 20655 806
rect 20866 821 20952 837
rect 21196 831 21226 862
rect 20529 768 20559 777
rect 19528 671 19558 702
rect 19624 676 19654 702
rect 19510 655 19576 671
rect 19510 621 19526 655
rect 19560 634 19576 655
rect 19560 621 19688 634
rect 20529 744 20565 768
rect 20535 729 20565 744
rect 20623 729 20653 790
rect 20866 787 20882 821
rect 20916 787 20952 821
rect 20866 771 20952 787
rect 20922 749 20952 771
rect 21178 815 21244 831
rect 21178 781 21194 815
rect 21228 781 21244 815
rect 21178 765 21244 781
rect 19034 593 19064 619
rect 19510 602 19688 621
rect 17734 540 17750 574
rect 17784 540 17800 574
rect 15864 502 15894 524
rect 17656 502 17686 528
rect 17734 524 17800 540
rect 19622 574 19688 602
rect 20230 601 20260 627
rect 20535 599 20565 625
rect 20623 599 20653 625
rect 22423 1075 22453 1101
rect 22511 1075 22541 1101
rect 22810 1069 22840 1095
rect 23066 1093 23132 1109
rect 22423 902 22453 917
rect 22417 878 22453 902
rect 21842 831 21872 862
rect 22118 845 22148 877
rect 21824 815 21890 831
rect 21824 781 21840 815
rect 21874 781 21890 815
rect 21824 765 21890 781
rect 22062 829 22148 845
rect 22417 843 22447 878
rect 22511 856 22541 917
rect 23084 1062 23114 1093
rect 22062 795 22078 829
rect 22112 795 22148 829
rect 22062 779 22148 795
rect 22118 757 22148 779
rect 22371 827 22447 843
rect 22371 793 22381 827
rect 22415 793 22447 827
rect 22371 777 22447 793
rect 22489 840 22543 856
rect 22489 806 22499 840
rect 22533 806 22543 840
rect 22810 837 22840 869
rect 23248 1016 23278 1174
rect 23698 1159 23730 1174
rect 25136 1174 25618 1204
rect 23698 1143 23778 1159
rect 23698 1109 23728 1143
rect 23762 1109 23778 1143
rect 23698 1093 23778 1109
rect 24954 1143 25020 1159
rect 24954 1109 24970 1143
rect 25004 1109 25020 1143
rect 23698 1092 23760 1093
rect 23730 1062 23760 1092
rect 24006 1077 24036 1103
rect 23248 986 23334 1016
rect 23304 902 23334 986
rect 23382 983 23448 999
rect 23382 949 23398 983
rect 23432 949 23448 983
rect 23382 933 23448 949
rect 23400 902 23430 933
rect 22489 790 22543 806
rect 22754 821 22840 837
rect 23084 831 23114 862
rect 22417 768 22447 777
rect 21416 671 21446 702
rect 21512 676 21542 702
rect 21398 655 21464 671
rect 21398 621 21414 655
rect 21448 634 21464 655
rect 21448 621 21576 634
rect 22417 744 22453 768
rect 22423 729 22453 744
rect 22511 729 22541 790
rect 22754 787 22770 821
rect 22804 787 22840 821
rect 22754 771 22840 787
rect 22810 749 22840 771
rect 23066 815 23132 831
rect 23066 781 23082 815
rect 23116 781 23132 815
rect 23066 765 23132 781
rect 20922 593 20952 619
rect 21398 602 21576 621
rect 19622 540 19638 574
rect 19672 540 19688 574
rect 17752 502 17782 524
rect 19544 502 19574 528
rect 19622 524 19688 540
rect 21510 574 21576 602
rect 22118 601 22148 627
rect 22423 599 22453 625
rect 22511 599 22541 625
rect 24311 1075 24341 1101
rect 24399 1075 24429 1101
rect 24698 1069 24728 1095
rect 24954 1093 25020 1109
rect 24311 902 24341 917
rect 24305 878 24341 902
rect 23730 831 23760 862
rect 24006 845 24036 877
rect 23712 815 23778 831
rect 23712 781 23728 815
rect 23762 781 23778 815
rect 23712 765 23778 781
rect 23950 829 24036 845
rect 24305 843 24335 878
rect 24399 856 24429 917
rect 24972 1062 25002 1093
rect 23950 795 23966 829
rect 24000 795 24036 829
rect 23950 779 24036 795
rect 24006 757 24036 779
rect 24259 827 24335 843
rect 24259 793 24269 827
rect 24303 793 24335 827
rect 24259 777 24335 793
rect 24377 840 24431 856
rect 24377 806 24387 840
rect 24421 806 24431 840
rect 24698 837 24728 869
rect 25136 1016 25166 1174
rect 25586 1159 25618 1174
rect 27024 1174 27506 1204
rect 25586 1143 25666 1159
rect 25586 1109 25616 1143
rect 25650 1109 25666 1143
rect 25586 1093 25666 1109
rect 26842 1143 26908 1159
rect 26842 1109 26858 1143
rect 26892 1109 26908 1143
rect 25586 1092 25648 1093
rect 25618 1062 25648 1092
rect 25894 1077 25924 1103
rect 25136 986 25222 1016
rect 25192 902 25222 986
rect 25270 983 25336 999
rect 25270 949 25286 983
rect 25320 949 25336 983
rect 25270 933 25336 949
rect 25288 902 25318 933
rect 24377 790 24431 806
rect 24642 821 24728 837
rect 24972 831 25002 862
rect 24305 768 24335 777
rect 23304 671 23334 702
rect 23400 676 23430 702
rect 23286 655 23352 671
rect 23286 621 23302 655
rect 23336 634 23352 655
rect 23336 621 23464 634
rect 24305 744 24341 768
rect 24311 729 24341 744
rect 24399 729 24429 790
rect 24642 787 24658 821
rect 24692 787 24728 821
rect 24642 771 24728 787
rect 24698 749 24728 771
rect 24954 815 25020 831
rect 24954 781 24970 815
rect 25004 781 25020 815
rect 24954 765 25020 781
rect 22810 593 22840 619
rect 23286 602 23464 621
rect 21510 540 21526 574
rect 21560 540 21576 574
rect 19640 502 19670 524
rect 21432 502 21462 528
rect 21510 524 21576 540
rect 23398 574 23464 602
rect 24006 601 24036 627
rect 24311 599 24341 625
rect 24399 599 24429 625
rect 26199 1075 26229 1101
rect 26287 1075 26317 1101
rect 26586 1069 26616 1095
rect 26842 1093 26908 1109
rect 26199 902 26229 917
rect 26193 878 26229 902
rect 25618 831 25648 862
rect 25894 845 25924 877
rect 25600 815 25666 831
rect 25600 781 25616 815
rect 25650 781 25666 815
rect 25600 765 25666 781
rect 25838 829 25924 845
rect 26193 843 26223 878
rect 26287 856 26317 917
rect 26860 1062 26890 1093
rect 25838 795 25854 829
rect 25888 795 25924 829
rect 25838 779 25924 795
rect 25894 757 25924 779
rect 26147 827 26223 843
rect 26147 793 26157 827
rect 26191 793 26223 827
rect 26147 777 26223 793
rect 26265 840 26319 856
rect 26265 806 26275 840
rect 26309 806 26319 840
rect 26586 837 26616 869
rect 27024 1016 27054 1174
rect 27474 1159 27506 1174
rect 28912 1174 29394 1204
rect 27474 1143 27554 1159
rect 27474 1109 27504 1143
rect 27538 1109 27554 1143
rect 27474 1093 27554 1109
rect 28730 1143 28796 1159
rect 28730 1109 28746 1143
rect 28780 1109 28796 1143
rect 27474 1092 27536 1093
rect 27506 1062 27536 1092
rect 27782 1077 27812 1103
rect 27024 986 27110 1016
rect 27080 902 27110 986
rect 27158 983 27224 999
rect 27158 949 27174 983
rect 27208 949 27224 983
rect 27158 933 27224 949
rect 27176 902 27206 933
rect 26265 790 26319 806
rect 26530 821 26616 837
rect 26860 831 26890 862
rect 26193 768 26223 777
rect 25192 671 25222 702
rect 25288 676 25318 702
rect 25174 655 25240 671
rect 25174 621 25190 655
rect 25224 634 25240 655
rect 25224 621 25352 634
rect 26193 744 26229 768
rect 26199 729 26229 744
rect 26287 729 26317 790
rect 26530 787 26546 821
rect 26580 787 26616 821
rect 26530 771 26616 787
rect 26586 749 26616 771
rect 26842 815 26908 831
rect 26842 781 26858 815
rect 26892 781 26908 815
rect 26842 765 26908 781
rect 24698 593 24728 619
rect 25174 602 25352 621
rect 23398 540 23414 574
rect 23448 540 23464 574
rect 21528 502 21558 524
rect 23320 502 23350 528
rect 23398 524 23464 540
rect 25286 574 25352 602
rect 25894 601 25924 627
rect 26199 599 26229 625
rect 26287 599 26317 625
rect 28087 1075 28117 1101
rect 28175 1075 28205 1101
rect 28474 1069 28504 1095
rect 28730 1093 28796 1109
rect 28087 902 28117 917
rect 28081 878 28117 902
rect 27506 831 27536 862
rect 27782 845 27812 877
rect 27488 815 27554 831
rect 27488 781 27504 815
rect 27538 781 27554 815
rect 27488 765 27554 781
rect 27726 829 27812 845
rect 28081 843 28111 878
rect 28175 856 28205 917
rect 28748 1062 28778 1093
rect 27726 795 27742 829
rect 27776 795 27812 829
rect 27726 779 27812 795
rect 27782 757 27812 779
rect 28035 827 28111 843
rect 28035 793 28045 827
rect 28079 793 28111 827
rect 28035 777 28111 793
rect 28153 840 28207 856
rect 28153 806 28163 840
rect 28197 806 28207 840
rect 28474 837 28504 869
rect 28912 1016 28942 1174
rect 29362 1159 29394 1174
rect 30800 1174 31282 1204
rect 29362 1143 29442 1159
rect 29362 1109 29392 1143
rect 29426 1109 29442 1143
rect 29362 1093 29442 1109
rect 30618 1143 30684 1159
rect 30618 1109 30634 1143
rect 30668 1109 30684 1143
rect 29362 1092 29424 1093
rect 29394 1062 29424 1092
rect 29670 1077 29700 1103
rect 28912 986 28998 1016
rect 28968 902 28998 986
rect 29046 983 29112 999
rect 29046 949 29062 983
rect 29096 949 29112 983
rect 29046 933 29112 949
rect 29064 902 29094 933
rect 28153 790 28207 806
rect 28418 821 28504 837
rect 28748 831 28778 862
rect 28081 768 28111 777
rect 27080 671 27110 702
rect 27176 676 27206 702
rect 27062 655 27128 671
rect 27062 621 27078 655
rect 27112 634 27128 655
rect 27112 621 27240 634
rect 28081 744 28117 768
rect 28087 729 28117 744
rect 28175 729 28205 790
rect 28418 787 28434 821
rect 28468 787 28504 821
rect 28418 771 28504 787
rect 28474 749 28504 771
rect 28730 815 28796 831
rect 28730 781 28746 815
rect 28780 781 28796 815
rect 28730 765 28796 781
rect 26586 593 26616 619
rect 27062 602 27240 621
rect 25286 540 25302 574
rect 25336 540 25352 574
rect 23416 502 23446 524
rect 25208 502 25238 528
rect 25286 524 25352 540
rect 27174 574 27240 602
rect 27782 601 27812 627
rect 28087 599 28117 625
rect 28175 599 28205 625
rect 29975 1075 30005 1101
rect 30063 1075 30093 1101
rect 30362 1069 30392 1095
rect 30618 1093 30684 1109
rect 29975 902 30005 917
rect 29969 878 30005 902
rect 29394 831 29424 862
rect 29670 845 29700 877
rect 29376 815 29442 831
rect 29376 781 29392 815
rect 29426 781 29442 815
rect 29376 765 29442 781
rect 29614 829 29700 845
rect 29969 843 29999 878
rect 30063 856 30093 917
rect 30636 1062 30666 1093
rect 29614 795 29630 829
rect 29664 795 29700 829
rect 29614 779 29700 795
rect 29670 757 29700 779
rect 29923 827 29999 843
rect 29923 793 29933 827
rect 29967 793 29999 827
rect 29923 777 29999 793
rect 30041 840 30095 856
rect 30041 806 30051 840
rect 30085 806 30095 840
rect 30362 837 30392 869
rect 30800 1016 30830 1174
rect 31250 1159 31282 1174
rect 32688 1174 33170 1204
rect 31250 1143 31330 1159
rect 31250 1109 31280 1143
rect 31314 1109 31330 1143
rect 31250 1093 31330 1109
rect 32506 1143 32572 1159
rect 32506 1109 32522 1143
rect 32556 1109 32572 1143
rect 31250 1092 31312 1093
rect 31282 1062 31312 1092
rect 31558 1077 31588 1103
rect 30800 986 30886 1016
rect 30856 902 30886 986
rect 30934 983 31000 999
rect 30934 949 30950 983
rect 30984 949 31000 983
rect 30934 933 31000 949
rect 30952 902 30982 933
rect 30041 790 30095 806
rect 30306 821 30392 837
rect 30636 831 30666 862
rect 29969 768 29999 777
rect 28968 671 28998 702
rect 29064 676 29094 702
rect 28950 655 29016 671
rect 28950 621 28966 655
rect 29000 634 29016 655
rect 29000 621 29128 634
rect 29969 744 30005 768
rect 29975 729 30005 744
rect 30063 729 30093 790
rect 30306 787 30322 821
rect 30356 787 30392 821
rect 30306 771 30392 787
rect 30362 749 30392 771
rect 30618 815 30684 831
rect 30618 781 30634 815
rect 30668 781 30684 815
rect 30618 765 30684 781
rect 28474 593 28504 619
rect 28950 602 29128 621
rect 27174 540 27190 574
rect 27224 540 27240 574
rect 25304 502 25334 524
rect 27096 502 27126 528
rect 27174 524 27240 540
rect 29062 574 29128 602
rect 29670 601 29700 627
rect 29975 599 30005 625
rect 30063 599 30093 625
rect 31863 1075 31893 1101
rect 31951 1075 31981 1101
rect 32250 1069 32280 1095
rect 32506 1093 32572 1109
rect 31863 902 31893 917
rect 31857 878 31893 902
rect 31282 831 31312 862
rect 31558 845 31588 877
rect 31264 815 31330 831
rect 31264 781 31280 815
rect 31314 781 31330 815
rect 31264 765 31330 781
rect 31502 829 31588 845
rect 31857 843 31887 878
rect 31951 856 31981 917
rect 32524 1062 32554 1093
rect 31502 795 31518 829
rect 31552 795 31588 829
rect 31502 779 31588 795
rect 31558 757 31588 779
rect 31811 827 31887 843
rect 31811 793 31821 827
rect 31855 793 31887 827
rect 31811 777 31887 793
rect 31929 840 31983 856
rect 31929 806 31939 840
rect 31973 806 31983 840
rect 32250 837 32280 869
rect 32688 1016 32718 1174
rect 33138 1159 33170 1174
rect 34576 1174 35058 1204
rect 33138 1143 33218 1159
rect 33138 1109 33168 1143
rect 33202 1109 33218 1143
rect 33138 1093 33218 1109
rect 34394 1143 34460 1159
rect 34394 1109 34410 1143
rect 34444 1109 34460 1143
rect 33138 1092 33200 1093
rect 33170 1062 33200 1092
rect 33446 1077 33476 1103
rect 32688 986 32774 1016
rect 32744 902 32774 986
rect 32822 983 32888 999
rect 32822 949 32838 983
rect 32872 949 32888 983
rect 32822 933 32888 949
rect 32840 902 32870 933
rect 31929 790 31983 806
rect 32194 821 32280 837
rect 32524 831 32554 862
rect 31857 768 31887 777
rect 30856 671 30886 702
rect 30952 676 30982 702
rect 30838 655 30904 671
rect 30838 621 30854 655
rect 30888 634 30904 655
rect 30888 621 31016 634
rect 31857 744 31893 768
rect 31863 729 31893 744
rect 31951 729 31981 790
rect 32194 787 32210 821
rect 32244 787 32280 821
rect 32194 771 32280 787
rect 32250 749 32280 771
rect 32506 815 32572 831
rect 32506 781 32522 815
rect 32556 781 32572 815
rect 32506 765 32572 781
rect 30362 593 30392 619
rect 30838 602 31016 621
rect 29062 540 29078 574
rect 29112 540 29128 574
rect 27192 502 27222 524
rect 28984 502 29014 528
rect 29062 524 29128 540
rect 30950 574 31016 602
rect 31558 601 31588 627
rect 31863 599 31893 625
rect 31951 599 31981 625
rect 33751 1075 33781 1101
rect 33839 1075 33869 1101
rect 34138 1069 34168 1095
rect 34394 1093 34460 1109
rect 33751 902 33781 917
rect 33745 878 33781 902
rect 33170 831 33200 862
rect 33446 845 33476 877
rect 33152 815 33218 831
rect 33152 781 33168 815
rect 33202 781 33218 815
rect 33152 765 33218 781
rect 33390 829 33476 845
rect 33745 843 33775 878
rect 33839 856 33869 917
rect 34412 1062 34442 1093
rect 33390 795 33406 829
rect 33440 795 33476 829
rect 33390 779 33476 795
rect 33446 757 33476 779
rect 33699 827 33775 843
rect 33699 793 33709 827
rect 33743 793 33775 827
rect 33699 777 33775 793
rect 33817 840 33871 856
rect 33817 806 33827 840
rect 33861 806 33871 840
rect 34138 837 34168 869
rect 34576 1016 34606 1174
rect 35026 1159 35058 1174
rect 36464 1174 36946 1204
rect 35026 1143 35106 1159
rect 35026 1109 35056 1143
rect 35090 1109 35106 1143
rect 35026 1093 35106 1109
rect 36282 1143 36348 1159
rect 36282 1109 36298 1143
rect 36332 1109 36348 1143
rect 35026 1092 35088 1093
rect 35058 1062 35088 1092
rect 35334 1077 35364 1103
rect 34576 986 34662 1016
rect 34632 902 34662 986
rect 34710 983 34776 999
rect 34710 949 34726 983
rect 34760 949 34776 983
rect 34710 933 34776 949
rect 34728 902 34758 933
rect 33817 790 33871 806
rect 34082 821 34168 837
rect 34412 831 34442 862
rect 33745 768 33775 777
rect 32744 671 32774 702
rect 32840 676 32870 702
rect 32726 655 32792 671
rect 32726 621 32742 655
rect 32776 634 32792 655
rect 32776 621 32904 634
rect 33745 744 33781 768
rect 33751 729 33781 744
rect 33839 729 33869 790
rect 34082 787 34098 821
rect 34132 787 34168 821
rect 34082 771 34168 787
rect 34138 749 34168 771
rect 34394 815 34460 831
rect 34394 781 34410 815
rect 34444 781 34460 815
rect 34394 765 34460 781
rect 32250 593 32280 619
rect 32726 602 32904 621
rect 30950 540 30966 574
rect 31000 540 31016 574
rect 29080 502 29110 524
rect 30872 502 30902 528
rect 30950 524 31016 540
rect 32838 574 32904 602
rect 33446 601 33476 627
rect 33751 599 33781 625
rect 33839 599 33869 625
rect 35639 1075 35669 1101
rect 35727 1075 35757 1101
rect 36026 1069 36056 1095
rect 36282 1093 36348 1109
rect 35639 902 35669 917
rect 35633 878 35669 902
rect 35058 831 35088 862
rect 35334 845 35364 877
rect 35040 815 35106 831
rect 35040 781 35056 815
rect 35090 781 35106 815
rect 35040 765 35106 781
rect 35278 829 35364 845
rect 35633 843 35663 878
rect 35727 856 35757 917
rect 36300 1062 36330 1093
rect 35278 795 35294 829
rect 35328 795 35364 829
rect 35278 779 35364 795
rect 35334 757 35364 779
rect 35587 827 35663 843
rect 35587 793 35597 827
rect 35631 793 35663 827
rect 35587 777 35663 793
rect 35705 840 35759 856
rect 35705 806 35715 840
rect 35749 806 35759 840
rect 36026 837 36056 869
rect 36464 1016 36494 1174
rect 36914 1159 36946 1174
rect 38352 1174 38834 1204
rect 36914 1143 36994 1159
rect 36914 1109 36944 1143
rect 36978 1109 36994 1143
rect 36914 1093 36994 1109
rect 38170 1143 38236 1159
rect 38170 1109 38186 1143
rect 38220 1109 38236 1143
rect 36914 1092 36976 1093
rect 36946 1062 36976 1092
rect 37222 1077 37252 1103
rect 36464 986 36550 1016
rect 36520 902 36550 986
rect 36598 983 36664 999
rect 36598 949 36614 983
rect 36648 949 36664 983
rect 36598 933 36664 949
rect 36616 902 36646 933
rect 35705 790 35759 806
rect 35970 821 36056 837
rect 36300 831 36330 862
rect 35633 768 35663 777
rect 34632 671 34662 702
rect 34728 676 34758 702
rect 34614 655 34680 671
rect 34614 621 34630 655
rect 34664 634 34680 655
rect 34664 621 34792 634
rect 35633 744 35669 768
rect 35639 729 35669 744
rect 35727 729 35757 790
rect 35970 787 35986 821
rect 36020 787 36056 821
rect 35970 771 36056 787
rect 36026 749 36056 771
rect 36282 815 36348 831
rect 36282 781 36298 815
rect 36332 781 36348 815
rect 36282 765 36348 781
rect 34138 593 34168 619
rect 34614 602 34792 621
rect 32838 540 32854 574
rect 32888 540 32904 574
rect 30968 502 30998 524
rect 32760 502 32790 528
rect 32838 524 32904 540
rect 34726 574 34792 602
rect 35334 601 35364 627
rect 35639 599 35669 625
rect 35727 599 35757 625
rect 37527 1075 37557 1101
rect 37615 1075 37645 1101
rect 37914 1069 37944 1095
rect 38170 1093 38236 1109
rect 37527 902 37557 917
rect 37521 878 37557 902
rect 36946 831 36976 862
rect 37222 845 37252 877
rect 36928 815 36994 831
rect 36928 781 36944 815
rect 36978 781 36994 815
rect 36928 765 36994 781
rect 37166 829 37252 845
rect 37521 843 37551 878
rect 37615 856 37645 917
rect 38188 1062 38218 1093
rect 37166 795 37182 829
rect 37216 795 37252 829
rect 37166 779 37252 795
rect 37222 757 37252 779
rect 37475 827 37551 843
rect 37475 793 37485 827
rect 37519 793 37551 827
rect 37475 777 37551 793
rect 37593 840 37647 856
rect 37593 806 37603 840
rect 37637 806 37647 840
rect 37914 837 37944 869
rect 38352 1016 38382 1174
rect 38802 1159 38834 1174
rect 40240 1174 40722 1204
rect 38802 1143 38882 1159
rect 38802 1109 38832 1143
rect 38866 1109 38882 1143
rect 38802 1093 38882 1109
rect 40058 1143 40124 1159
rect 40058 1109 40074 1143
rect 40108 1109 40124 1143
rect 38802 1092 38864 1093
rect 38834 1062 38864 1092
rect 39110 1077 39140 1103
rect 38352 986 38438 1016
rect 38408 902 38438 986
rect 38486 983 38552 999
rect 38486 949 38502 983
rect 38536 949 38552 983
rect 38486 933 38552 949
rect 38504 902 38534 933
rect 37593 790 37647 806
rect 37858 821 37944 837
rect 38188 831 38218 862
rect 37521 768 37551 777
rect 36520 671 36550 702
rect 36616 676 36646 702
rect 36502 655 36568 671
rect 36502 621 36518 655
rect 36552 634 36568 655
rect 36552 621 36680 634
rect 37521 744 37557 768
rect 37527 729 37557 744
rect 37615 729 37645 790
rect 37858 787 37874 821
rect 37908 787 37944 821
rect 37858 771 37944 787
rect 37914 749 37944 771
rect 38170 815 38236 831
rect 38170 781 38186 815
rect 38220 781 38236 815
rect 38170 765 38236 781
rect 36026 593 36056 619
rect 36502 602 36680 621
rect 34726 540 34742 574
rect 34776 540 34792 574
rect 32856 502 32886 524
rect 34648 502 34678 528
rect 34726 524 34792 540
rect 36614 574 36680 602
rect 37222 601 37252 627
rect 37527 599 37557 625
rect 37615 599 37645 625
rect 39415 1075 39445 1101
rect 39503 1075 39533 1101
rect 39802 1069 39832 1095
rect 40058 1093 40124 1109
rect 39415 902 39445 917
rect 39409 878 39445 902
rect 38834 831 38864 862
rect 39110 845 39140 877
rect 38816 815 38882 831
rect 38816 781 38832 815
rect 38866 781 38882 815
rect 38816 765 38882 781
rect 39054 829 39140 845
rect 39409 843 39439 878
rect 39503 856 39533 917
rect 40076 1062 40106 1093
rect 39054 795 39070 829
rect 39104 795 39140 829
rect 39054 779 39140 795
rect 39110 757 39140 779
rect 39363 827 39439 843
rect 39363 793 39373 827
rect 39407 793 39439 827
rect 39363 777 39439 793
rect 39481 840 39535 856
rect 39481 806 39491 840
rect 39525 806 39535 840
rect 39802 837 39832 869
rect 40240 1016 40270 1174
rect 40690 1159 40722 1174
rect 42128 1174 42610 1204
rect 40690 1143 40770 1159
rect 40690 1109 40720 1143
rect 40754 1109 40770 1143
rect 40690 1093 40770 1109
rect 41946 1143 42012 1159
rect 41946 1109 41962 1143
rect 41996 1109 42012 1143
rect 40690 1092 40752 1093
rect 40722 1062 40752 1092
rect 40998 1077 41028 1103
rect 40240 986 40326 1016
rect 40296 902 40326 986
rect 40374 983 40440 999
rect 40374 949 40390 983
rect 40424 949 40440 983
rect 40374 933 40440 949
rect 40392 902 40422 933
rect 39481 790 39535 806
rect 39746 821 39832 837
rect 40076 831 40106 862
rect 39409 768 39439 777
rect 38408 671 38438 702
rect 38504 676 38534 702
rect 38390 655 38456 671
rect 38390 621 38406 655
rect 38440 634 38456 655
rect 38440 621 38568 634
rect 39409 744 39445 768
rect 39415 729 39445 744
rect 39503 729 39533 790
rect 39746 787 39762 821
rect 39796 787 39832 821
rect 39746 771 39832 787
rect 39802 749 39832 771
rect 40058 815 40124 831
rect 40058 781 40074 815
rect 40108 781 40124 815
rect 40058 765 40124 781
rect 37914 593 37944 619
rect 38390 602 38568 621
rect 36614 540 36630 574
rect 36664 540 36680 574
rect 34744 502 34774 524
rect 36536 502 36566 528
rect 36614 524 36680 540
rect 38502 574 38568 602
rect 39110 601 39140 627
rect 39415 599 39445 625
rect 39503 599 39533 625
rect 41303 1075 41333 1101
rect 41391 1075 41421 1101
rect 41690 1069 41720 1095
rect 41946 1093 42012 1109
rect 41303 902 41333 917
rect 41297 878 41333 902
rect 40722 831 40752 862
rect 40998 845 41028 877
rect 40704 815 40770 831
rect 40704 781 40720 815
rect 40754 781 40770 815
rect 40704 765 40770 781
rect 40942 829 41028 845
rect 41297 843 41327 878
rect 41391 856 41421 917
rect 41964 1062 41994 1093
rect 40942 795 40958 829
rect 40992 795 41028 829
rect 40942 779 41028 795
rect 40998 757 41028 779
rect 41251 827 41327 843
rect 41251 793 41261 827
rect 41295 793 41327 827
rect 41251 777 41327 793
rect 41369 840 41423 856
rect 41369 806 41379 840
rect 41413 806 41423 840
rect 41690 837 41720 869
rect 42128 1016 42158 1174
rect 42578 1159 42610 1174
rect 44016 1174 44498 1204
rect 42578 1143 42658 1159
rect 42578 1109 42608 1143
rect 42642 1109 42658 1143
rect 42578 1093 42658 1109
rect 43834 1143 43900 1159
rect 43834 1109 43850 1143
rect 43884 1109 43900 1143
rect 42578 1092 42640 1093
rect 42610 1062 42640 1092
rect 42886 1077 42916 1103
rect 42128 986 42214 1016
rect 42184 902 42214 986
rect 42262 983 42328 999
rect 42262 949 42278 983
rect 42312 949 42328 983
rect 42262 933 42328 949
rect 42280 902 42310 933
rect 41369 790 41423 806
rect 41634 821 41720 837
rect 41964 831 41994 862
rect 41297 768 41327 777
rect 40296 671 40326 702
rect 40392 676 40422 702
rect 40278 655 40344 671
rect 40278 621 40294 655
rect 40328 634 40344 655
rect 40328 621 40456 634
rect 41297 744 41333 768
rect 41303 729 41333 744
rect 41391 729 41421 790
rect 41634 787 41650 821
rect 41684 787 41720 821
rect 41634 771 41720 787
rect 41690 749 41720 771
rect 41946 815 42012 831
rect 41946 781 41962 815
rect 41996 781 42012 815
rect 41946 765 42012 781
rect 39802 593 39832 619
rect 40278 602 40456 621
rect 38502 540 38518 574
rect 38552 540 38568 574
rect 36632 502 36662 524
rect 38424 502 38454 528
rect 38502 524 38568 540
rect 40390 574 40456 602
rect 40998 601 41028 627
rect 41303 599 41333 625
rect 41391 599 41421 625
rect 43191 1075 43221 1101
rect 43279 1075 43309 1101
rect 43578 1069 43608 1095
rect 43834 1093 43900 1109
rect 43191 902 43221 917
rect 43185 878 43221 902
rect 42610 831 42640 862
rect 42886 845 42916 877
rect 42592 815 42658 831
rect 42592 781 42608 815
rect 42642 781 42658 815
rect 42592 765 42658 781
rect 42830 829 42916 845
rect 43185 843 43215 878
rect 43279 856 43309 917
rect 43852 1062 43882 1093
rect 42830 795 42846 829
rect 42880 795 42916 829
rect 42830 779 42916 795
rect 42886 757 42916 779
rect 43139 827 43215 843
rect 43139 793 43149 827
rect 43183 793 43215 827
rect 43139 777 43215 793
rect 43257 840 43311 856
rect 43257 806 43267 840
rect 43301 806 43311 840
rect 43578 837 43608 869
rect 44016 1016 44046 1174
rect 44466 1159 44498 1174
rect 45898 1174 46380 1204
rect 44466 1143 44546 1159
rect 44466 1109 44496 1143
rect 44530 1109 44546 1143
rect 44466 1093 44546 1109
rect 45716 1143 45782 1159
rect 45716 1109 45732 1143
rect 45766 1109 45782 1143
rect 44466 1092 44528 1093
rect 44498 1062 44528 1092
rect 44774 1077 44804 1103
rect 44016 986 44102 1016
rect 44072 902 44102 986
rect 44150 983 44216 999
rect 44150 949 44166 983
rect 44200 949 44216 983
rect 44150 933 44216 949
rect 44168 902 44198 933
rect 43257 790 43311 806
rect 43522 821 43608 837
rect 43852 831 43882 862
rect 43185 768 43215 777
rect 42184 671 42214 702
rect 42280 676 42310 702
rect 42166 655 42232 671
rect 42166 621 42182 655
rect 42216 634 42232 655
rect 42216 621 42344 634
rect 43185 744 43221 768
rect 43191 729 43221 744
rect 43279 729 43309 790
rect 43522 787 43538 821
rect 43572 787 43608 821
rect 43522 771 43608 787
rect 43578 749 43608 771
rect 43834 815 43900 831
rect 43834 781 43850 815
rect 43884 781 43900 815
rect 43834 765 43900 781
rect 41690 593 41720 619
rect 42166 602 42344 621
rect 40390 540 40406 574
rect 40440 540 40456 574
rect 38520 502 38550 524
rect 40312 502 40342 528
rect 40390 524 40456 540
rect 42278 574 42344 602
rect 42886 601 42916 627
rect 43191 599 43221 625
rect 43279 599 43309 625
rect 45079 1075 45109 1101
rect 45167 1075 45197 1101
rect 45460 1069 45490 1095
rect 45716 1093 45782 1109
rect 45079 902 45109 917
rect 45073 878 45109 902
rect 44498 831 44528 862
rect 44774 845 44804 877
rect 44480 815 44546 831
rect 44480 781 44496 815
rect 44530 781 44546 815
rect 44480 765 44546 781
rect 44718 829 44804 845
rect 45073 843 45103 878
rect 45167 856 45197 917
rect 45734 1062 45764 1093
rect 44718 795 44734 829
rect 44768 795 44804 829
rect 44718 779 44804 795
rect 44774 757 44804 779
rect 45027 827 45103 843
rect 45027 793 45037 827
rect 45071 793 45103 827
rect 45027 777 45103 793
rect 45145 840 45199 856
rect 45145 806 45155 840
rect 45189 806 45199 840
rect 45460 837 45490 869
rect 45898 1016 45928 1174
rect 46348 1159 46380 1174
rect 47786 1174 48268 1204
rect 46348 1143 46428 1159
rect 46348 1109 46378 1143
rect 46412 1109 46428 1143
rect 46348 1093 46428 1109
rect 47604 1143 47670 1159
rect 47604 1109 47620 1143
rect 47654 1109 47670 1143
rect 46348 1092 46410 1093
rect 46380 1062 46410 1092
rect 46656 1077 46686 1103
rect 45898 986 45984 1016
rect 45954 902 45984 986
rect 46032 983 46098 999
rect 46032 949 46048 983
rect 46082 949 46098 983
rect 46032 933 46098 949
rect 46050 902 46080 933
rect 45145 790 45199 806
rect 45404 821 45490 837
rect 45734 831 45764 862
rect 45073 768 45103 777
rect 44072 671 44102 702
rect 44168 676 44198 702
rect 44054 655 44120 671
rect 44054 621 44070 655
rect 44104 634 44120 655
rect 44104 621 44232 634
rect 45073 744 45109 768
rect 45079 729 45109 744
rect 45167 729 45197 790
rect 45404 787 45420 821
rect 45454 787 45490 821
rect 45404 771 45490 787
rect 45460 749 45490 771
rect 45716 815 45782 831
rect 45716 781 45732 815
rect 45766 781 45782 815
rect 45716 765 45782 781
rect 43578 593 43608 619
rect 44054 602 44232 621
rect 42278 540 42294 574
rect 42328 540 42344 574
rect 40408 502 40438 524
rect 42200 502 42230 528
rect 42278 524 42344 540
rect 44166 574 44232 602
rect 44774 601 44804 627
rect 45079 599 45109 625
rect 45167 599 45197 625
rect 46961 1075 46991 1101
rect 47049 1075 47079 1101
rect 47348 1069 47378 1095
rect 47604 1093 47670 1109
rect 46961 902 46991 917
rect 46955 878 46991 902
rect 46380 831 46410 862
rect 46656 845 46686 877
rect 46362 815 46428 831
rect 46362 781 46378 815
rect 46412 781 46428 815
rect 46362 765 46428 781
rect 46600 829 46686 845
rect 46955 843 46985 878
rect 47049 856 47079 917
rect 47622 1062 47652 1093
rect 46600 795 46616 829
rect 46650 795 46686 829
rect 46600 779 46686 795
rect 46656 757 46686 779
rect 46909 827 46985 843
rect 46909 793 46919 827
rect 46953 793 46985 827
rect 46909 777 46985 793
rect 47027 840 47081 856
rect 47027 806 47037 840
rect 47071 806 47081 840
rect 47348 837 47378 869
rect 47786 1016 47816 1174
rect 48236 1159 48268 1174
rect 49674 1174 50156 1204
rect 48236 1143 48316 1159
rect 48236 1109 48266 1143
rect 48300 1109 48316 1143
rect 48236 1093 48316 1109
rect 49492 1143 49558 1159
rect 49492 1109 49508 1143
rect 49542 1109 49558 1143
rect 48236 1092 48298 1093
rect 48268 1062 48298 1092
rect 48544 1077 48574 1103
rect 47786 986 47872 1016
rect 47842 902 47872 986
rect 47920 983 47986 999
rect 47920 949 47936 983
rect 47970 949 47986 983
rect 47920 933 47986 949
rect 47938 902 47968 933
rect 47027 790 47081 806
rect 47292 821 47378 837
rect 47622 831 47652 862
rect 46955 768 46985 777
rect 45954 671 45984 702
rect 46050 676 46080 702
rect 45936 655 46002 671
rect 45936 621 45952 655
rect 45986 634 46002 655
rect 45986 621 46114 634
rect 46955 744 46991 768
rect 46961 729 46991 744
rect 47049 729 47079 790
rect 47292 787 47308 821
rect 47342 787 47378 821
rect 47292 771 47378 787
rect 47348 749 47378 771
rect 47604 815 47670 831
rect 47604 781 47620 815
rect 47654 781 47670 815
rect 47604 765 47670 781
rect 45460 593 45490 619
rect 45936 602 46114 621
rect 44166 540 44182 574
rect 44216 540 44232 574
rect 42296 502 42326 524
rect 44088 502 44118 528
rect 44166 524 44232 540
rect 46048 574 46114 602
rect 46656 601 46686 627
rect 46961 599 46991 625
rect 47049 599 47079 625
rect 48849 1075 48879 1101
rect 48937 1075 48967 1101
rect 49236 1069 49266 1095
rect 49492 1093 49558 1109
rect 48849 902 48879 917
rect 48843 878 48879 902
rect 48268 831 48298 862
rect 48544 845 48574 877
rect 48250 815 48316 831
rect 48250 781 48266 815
rect 48300 781 48316 815
rect 48250 765 48316 781
rect 48488 829 48574 845
rect 48843 843 48873 878
rect 48937 856 48967 917
rect 49510 1062 49540 1093
rect 48488 795 48504 829
rect 48538 795 48574 829
rect 48488 779 48574 795
rect 48544 757 48574 779
rect 48797 827 48873 843
rect 48797 793 48807 827
rect 48841 793 48873 827
rect 48797 777 48873 793
rect 48915 840 48969 856
rect 48915 806 48925 840
rect 48959 806 48969 840
rect 49236 837 49266 869
rect 49674 1016 49704 1174
rect 50124 1159 50156 1174
rect 51562 1174 52044 1204
rect 50124 1143 50204 1159
rect 50124 1109 50154 1143
rect 50188 1109 50204 1143
rect 50124 1093 50204 1109
rect 51380 1143 51446 1159
rect 51380 1109 51396 1143
rect 51430 1109 51446 1143
rect 50124 1092 50186 1093
rect 50156 1062 50186 1092
rect 50432 1077 50462 1103
rect 49674 986 49760 1016
rect 49730 902 49760 986
rect 49808 983 49874 999
rect 49808 949 49824 983
rect 49858 949 49874 983
rect 49808 933 49874 949
rect 49826 902 49856 933
rect 48915 790 48969 806
rect 49180 821 49266 837
rect 49510 831 49540 862
rect 48843 768 48873 777
rect 47842 671 47872 702
rect 47938 676 47968 702
rect 47824 655 47890 671
rect 47824 621 47840 655
rect 47874 634 47890 655
rect 47874 621 48002 634
rect 48843 744 48879 768
rect 48849 729 48879 744
rect 48937 729 48967 790
rect 49180 787 49196 821
rect 49230 787 49266 821
rect 49180 771 49266 787
rect 49236 749 49266 771
rect 49492 815 49558 831
rect 49492 781 49508 815
rect 49542 781 49558 815
rect 49492 765 49558 781
rect 47348 593 47378 619
rect 47824 602 48002 621
rect 46048 540 46064 574
rect 46098 540 46114 574
rect 44184 502 44214 524
rect 45970 502 46000 528
rect 46048 524 46114 540
rect 47936 574 48002 602
rect 48544 601 48574 627
rect 48849 599 48879 625
rect 48937 599 48967 625
rect 50737 1075 50767 1101
rect 50825 1075 50855 1101
rect 51124 1069 51154 1095
rect 51380 1093 51446 1109
rect 50737 902 50767 917
rect 50731 878 50767 902
rect 50156 831 50186 862
rect 50432 845 50462 877
rect 50138 815 50204 831
rect 50138 781 50154 815
rect 50188 781 50204 815
rect 50138 765 50204 781
rect 50376 829 50462 845
rect 50731 843 50761 878
rect 50825 856 50855 917
rect 51398 1062 51428 1093
rect 50376 795 50392 829
rect 50426 795 50462 829
rect 50376 779 50462 795
rect 50432 757 50462 779
rect 50685 827 50761 843
rect 50685 793 50695 827
rect 50729 793 50761 827
rect 50685 777 50761 793
rect 50803 840 50857 856
rect 50803 806 50813 840
rect 50847 806 50857 840
rect 51124 837 51154 869
rect 51562 1016 51592 1174
rect 52012 1159 52044 1174
rect 53450 1174 53932 1204
rect 52012 1143 52092 1159
rect 52012 1109 52042 1143
rect 52076 1109 52092 1143
rect 52012 1093 52092 1109
rect 53268 1143 53334 1159
rect 53268 1109 53284 1143
rect 53318 1109 53334 1143
rect 52012 1092 52074 1093
rect 52044 1062 52074 1092
rect 52320 1077 52350 1103
rect 51562 986 51648 1016
rect 51618 902 51648 986
rect 51696 983 51762 999
rect 51696 949 51712 983
rect 51746 949 51762 983
rect 51696 933 51762 949
rect 51714 902 51744 933
rect 50803 790 50857 806
rect 51068 821 51154 837
rect 51398 831 51428 862
rect 50731 768 50761 777
rect 49730 671 49760 702
rect 49826 676 49856 702
rect 49712 655 49778 671
rect 49712 621 49728 655
rect 49762 634 49778 655
rect 49762 621 49890 634
rect 50731 744 50767 768
rect 50737 729 50767 744
rect 50825 729 50855 790
rect 51068 787 51084 821
rect 51118 787 51154 821
rect 51068 771 51154 787
rect 51124 749 51154 771
rect 51380 815 51446 831
rect 51380 781 51396 815
rect 51430 781 51446 815
rect 51380 765 51446 781
rect 49236 593 49266 619
rect 49712 602 49890 621
rect 47936 540 47952 574
rect 47986 540 48002 574
rect 46066 502 46096 524
rect 47858 502 47888 528
rect 47936 524 48002 540
rect 49824 574 49890 602
rect 50432 601 50462 627
rect 50737 599 50767 625
rect 50825 599 50855 625
rect 52625 1075 52655 1101
rect 52713 1075 52743 1101
rect 53012 1069 53042 1095
rect 53268 1093 53334 1109
rect 52625 902 52655 917
rect 52619 878 52655 902
rect 52044 831 52074 862
rect 52320 845 52350 877
rect 52026 815 52092 831
rect 52026 781 52042 815
rect 52076 781 52092 815
rect 52026 765 52092 781
rect 52264 829 52350 845
rect 52619 843 52649 878
rect 52713 856 52743 917
rect 53286 1062 53316 1093
rect 52264 795 52280 829
rect 52314 795 52350 829
rect 52264 779 52350 795
rect 52320 757 52350 779
rect 52573 827 52649 843
rect 52573 793 52583 827
rect 52617 793 52649 827
rect 52573 777 52649 793
rect 52691 840 52745 856
rect 52691 806 52701 840
rect 52735 806 52745 840
rect 53012 837 53042 869
rect 53450 1016 53480 1174
rect 53900 1159 53932 1174
rect 55338 1174 55820 1204
rect 53900 1143 53980 1159
rect 53900 1109 53930 1143
rect 53964 1109 53980 1143
rect 53900 1093 53980 1109
rect 55156 1143 55222 1159
rect 55156 1109 55172 1143
rect 55206 1109 55222 1143
rect 53900 1092 53962 1093
rect 53932 1062 53962 1092
rect 54208 1077 54238 1103
rect 53450 986 53536 1016
rect 53506 902 53536 986
rect 53584 983 53650 999
rect 53584 949 53600 983
rect 53634 949 53650 983
rect 53584 933 53650 949
rect 53602 902 53632 933
rect 52691 790 52745 806
rect 52956 821 53042 837
rect 53286 831 53316 862
rect 52619 768 52649 777
rect 51618 671 51648 702
rect 51714 676 51744 702
rect 51600 655 51666 671
rect 51600 621 51616 655
rect 51650 634 51666 655
rect 51650 621 51778 634
rect 52619 744 52655 768
rect 52625 729 52655 744
rect 52713 729 52743 790
rect 52956 787 52972 821
rect 53006 787 53042 821
rect 52956 771 53042 787
rect 53012 749 53042 771
rect 53268 815 53334 831
rect 53268 781 53284 815
rect 53318 781 53334 815
rect 53268 765 53334 781
rect 51124 593 51154 619
rect 51600 602 51778 621
rect 49824 540 49840 574
rect 49874 540 49890 574
rect 47954 502 47984 524
rect 49746 502 49776 528
rect 49824 524 49890 540
rect 51712 574 51778 602
rect 52320 601 52350 627
rect 52625 599 52655 625
rect 52713 599 52743 625
rect 54513 1075 54543 1101
rect 54601 1075 54631 1101
rect 54900 1069 54930 1095
rect 55156 1093 55222 1109
rect 54513 902 54543 917
rect 54507 878 54543 902
rect 53932 831 53962 862
rect 54208 845 54238 877
rect 53914 815 53980 831
rect 53914 781 53930 815
rect 53964 781 53980 815
rect 53914 765 53980 781
rect 54152 829 54238 845
rect 54507 843 54537 878
rect 54601 856 54631 917
rect 55174 1062 55204 1093
rect 54152 795 54168 829
rect 54202 795 54238 829
rect 54152 779 54238 795
rect 54208 757 54238 779
rect 54461 827 54537 843
rect 54461 793 54471 827
rect 54505 793 54537 827
rect 54461 777 54537 793
rect 54579 840 54633 856
rect 54579 806 54589 840
rect 54623 806 54633 840
rect 54900 837 54930 869
rect 55338 1016 55368 1174
rect 55788 1159 55820 1174
rect 57226 1174 57708 1204
rect 55788 1143 55868 1159
rect 55788 1109 55818 1143
rect 55852 1109 55868 1143
rect 55788 1093 55868 1109
rect 57044 1143 57110 1159
rect 57044 1109 57060 1143
rect 57094 1109 57110 1143
rect 55788 1092 55850 1093
rect 55820 1062 55850 1092
rect 56096 1077 56126 1103
rect 55338 986 55424 1016
rect 55394 902 55424 986
rect 55472 983 55538 999
rect 55472 949 55488 983
rect 55522 949 55538 983
rect 55472 933 55538 949
rect 55490 902 55520 933
rect 54579 790 54633 806
rect 54844 821 54930 837
rect 55174 831 55204 862
rect 54507 768 54537 777
rect 53506 671 53536 702
rect 53602 676 53632 702
rect 53488 655 53554 671
rect 53488 621 53504 655
rect 53538 634 53554 655
rect 53538 621 53666 634
rect 54507 744 54543 768
rect 54513 729 54543 744
rect 54601 729 54631 790
rect 54844 787 54860 821
rect 54894 787 54930 821
rect 54844 771 54930 787
rect 54900 749 54930 771
rect 55156 815 55222 831
rect 55156 781 55172 815
rect 55206 781 55222 815
rect 55156 765 55222 781
rect 53012 593 53042 619
rect 53488 602 53666 621
rect 51712 540 51728 574
rect 51762 540 51778 574
rect 49842 502 49872 524
rect 51634 502 51664 528
rect 51712 524 51778 540
rect 53600 574 53666 602
rect 54208 601 54238 627
rect 54513 599 54543 625
rect 54601 599 54631 625
rect 56401 1075 56431 1101
rect 56489 1075 56519 1101
rect 56788 1069 56818 1095
rect 57044 1093 57110 1109
rect 56401 902 56431 917
rect 56395 878 56431 902
rect 55820 831 55850 862
rect 56096 845 56126 877
rect 55802 815 55868 831
rect 55802 781 55818 815
rect 55852 781 55868 815
rect 55802 765 55868 781
rect 56040 829 56126 845
rect 56395 843 56425 878
rect 56489 856 56519 917
rect 57062 1062 57092 1093
rect 56040 795 56056 829
rect 56090 795 56126 829
rect 56040 779 56126 795
rect 56096 757 56126 779
rect 56349 827 56425 843
rect 56349 793 56359 827
rect 56393 793 56425 827
rect 56349 777 56425 793
rect 56467 840 56521 856
rect 56467 806 56477 840
rect 56511 806 56521 840
rect 56788 837 56818 869
rect 57226 1016 57256 1174
rect 57676 1159 57708 1174
rect 59114 1174 59596 1204
rect 57676 1143 57756 1159
rect 57676 1109 57706 1143
rect 57740 1109 57756 1143
rect 57676 1093 57756 1109
rect 58932 1143 58998 1159
rect 58932 1109 58948 1143
rect 58982 1109 58998 1143
rect 57676 1092 57738 1093
rect 57708 1062 57738 1092
rect 57984 1077 58014 1103
rect 57226 986 57312 1016
rect 57282 902 57312 986
rect 57360 983 57426 999
rect 57360 949 57376 983
rect 57410 949 57426 983
rect 57360 933 57426 949
rect 57378 902 57408 933
rect 56467 790 56521 806
rect 56732 821 56818 837
rect 57062 831 57092 862
rect 56395 768 56425 777
rect 55394 671 55424 702
rect 55490 676 55520 702
rect 55376 655 55442 671
rect 55376 621 55392 655
rect 55426 634 55442 655
rect 55426 621 55554 634
rect 56395 744 56431 768
rect 56401 729 56431 744
rect 56489 729 56519 790
rect 56732 787 56748 821
rect 56782 787 56818 821
rect 56732 771 56818 787
rect 56788 749 56818 771
rect 57044 815 57110 831
rect 57044 781 57060 815
rect 57094 781 57110 815
rect 57044 765 57110 781
rect 54900 593 54930 619
rect 55376 602 55554 621
rect 53600 540 53616 574
rect 53650 540 53666 574
rect 51730 502 51760 524
rect 53522 502 53552 528
rect 53600 524 53666 540
rect 55488 574 55554 602
rect 56096 601 56126 627
rect 56401 599 56431 625
rect 56489 599 56519 625
rect 58289 1075 58319 1101
rect 58377 1075 58407 1101
rect 58676 1069 58706 1095
rect 58932 1093 58998 1109
rect 58289 902 58319 917
rect 58283 878 58319 902
rect 57708 831 57738 862
rect 57984 845 58014 877
rect 57690 815 57756 831
rect 57690 781 57706 815
rect 57740 781 57756 815
rect 57690 765 57756 781
rect 57928 829 58014 845
rect 58283 843 58313 878
rect 58377 856 58407 917
rect 58950 1062 58980 1093
rect 57928 795 57944 829
rect 57978 795 58014 829
rect 57928 779 58014 795
rect 57984 757 58014 779
rect 58237 827 58313 843
rect 58237 793 58247 827
rect 58281 793 58313 827
rect 58237 777 58313 793
rect 58355 840 58409 856
rect 58355 806 58365 840
rect 58399 806 58409 840
rect 58676 837 58706 869
rect 59114 1016 59144 1174
rect 59564 1159 59596 1174
rect 59564 1143 59644 1159
rect 59564 1109 59594 1143
rect 59628 1109 59644 1143
rect 59564 1093 59644 1109
rect 59564 1092 59626 1093
rect 59596 1062 59626 1092
rect 59872 1077 59902 1103
rect 59114 986 59200 1016
rect 59170 902 59200 986
rect 59248 983 59314 999
rect 59248 949 59264 983
rect 59298 949 59314 983
rect 59248 933 59314 949
rect 59266 902 59296 933
rect 58355 790 58409 806
rect 58620 821 58706 837
rect 58950 831 58980 862
rect 58283 768 58313 777
rect 57282 671 57312 702
rect 57378 676 57408 702
rect 57264 655 57330 671
rect 57264 621 57280 655
rect 57314 634 57330 655
rect 57314 621 57442 634
rect 58283 744 58319 768
rect 58289 729 58319 744
rect 58377 729 58407 790
rect 58620 787 58636 821
rect 58670 787 58706 821
rect 58620 771 58706 787
rect 58676 749 58706 771
rect 58932 815 58998 831
rect 58932 781 58948 815
rect 58982 781 58998 815
rect 58932 765 58998 781
rect 56788 593 56818 619
rect 57264 602 57442 621
rect 55488 540 55504 574
rect 55538 540 55554 574
rect 53618 502 53648 524
rect 55410 502 55440 528
rect 55488 524 55554 540
rect 57376 574 57442 602
rect 57984 601 58014 627
rect 58289 599 58319 625
rect 58377 599 58407 625
rect 60177 1075 60207 1101
rect 60265 1075 60295 1101
rect 60177 902 60207 917
rect 60171 878 60207 902
rect 59596 831 59626 862
rect 59872 845 59902 877
rect 59578 815 59644 831
rect 59578 781 59594 815
rect 59628 781 59644 815
rect 59578 765 59644 781
rect 59816 829 59902 845
rect 60171 843 60201 878
rect 60265 856 60295 917
rect 59816 795 59832 829
rect 59866 795 59902 829
rect 59816 779 59902 795
rect 59872 757 59902 779
rect 60125 827 60201 843
rect 60125 793 60135 827
rect 60169 793 60201 827
rect 60125 777 60201 793
rect 60243 840 60297 856
rect 60243 806 60253 840
rect 60287 806 60297 840
rect 60243 790 60297 806
rect 60171 768 60201 777
rect 59170 671 59200 702
rect 59266 676 59296 702
rect 59152 655 59218 671
rect 59152 621 59168 655
rect 59202 634 59218 655
rect 59202 621 59330 634
rect 60171 744 60207 768
rect 60177 729 60207 744
rect 60265 729 60295 790
rect 58676 593 58706 619
rect 59152 602 59330 621
rect 57376 540 57392 574
rect 57426 540 57442 574
rect 55506 502 55536 524
rect 57298 502 57328 528
rect 57376 524 57442 540
rect 59264 574 59330 602
rect 59872 601 59902 627
rect 60177 599 60207 625
rect 60265 599 60295 625
rect 59264 540 59280 574
rect 59314 540 59330 574
rect 57394 502 57424 524
rect 59186 502 59216 528
rect 59264 524 59330 540
rect 59282 502 59312 524
rect 670 350 700 372
rect 652 334 718 350
rect 766 346 796 372
rect 2558 350 2588 372
rect 652 300 668 334
rect 702 300 718 334
rect 652 284 718 300
rect 2540 334 2606 350
rect 2654 346 2684 372
rect 4446 350 4476 372
rect 2540 300 2556 334
rect 2590 300 2606 334
rect 2540 284 2606 300
rect 4428 334 4494 350
rect 4542 346 4572 372
rect 6334 350 6364 372
rect 4428 300 4444 334
rect 4478 300 4494 334
rect 4428 284 4494 300
rect 6316 334 6382 350
rect 6430 346 6460 372
rect 8222 350 8252 372
rect 6316 300 6332 334
rect 6366 300 6382 334
rect 6316 284 6382 300
rect 8204 334 8270 350
rect 8318 346 8348 372
rect 10110 350 10140 372
rect 8204 300 8220 334
rect 8254 300 8270 334
rect 8204 284 8270 300
rect 10092 334 10158 350
rect 10206 346 10236 372
rect 11998 350 12028 372
rect 10092 300 10108 334
rect 10142 300 10158 334
rect 10092 284 10158 300
rect 11980 334 12046 350
rect 12094 346 12124 372
rect 13886 350 13916 372
rect 11980 300 11996 334
rect 12030 300 12046 334
rect 11980 284 12046 300
rect 13868 334 13934 350
rect 13982 346 14012 372
rect 15768 350 15798 372
rect 13868 300 13884 334
rect 13918 300 13934 334
rect 13868 284 13934 300
rect 15750 334 15816 350
rect 15864 346 15894 372
rect 17656 350 17686 372
rect 15750 300 15766 334
rect 15800 300 15816 334
rect 15750 284 15816 300
rect 17638 334 17704 350
rect 17752 346 17782 372
rect 19544 350 19574 372
rect 17638 300 17654 334
rect 17688 300 17704 334
rect 17638 284 17704 300
rect 19526 334 19592 350
rect 19640 346 19670 372
rect 21432 350 21462 372
rect 19526 300 19542 334
rect 19576 300 19592 334
rect 19526 284 19592 300
rect 21414 334 21480 350
rect 21528 346 21558 372
rect 23320 350 23350 372
rect 21414 300 21430 334
rect 21464 300 21480 334
rect 21414 284 21480 300
rect 23302 334 23368 350
rect 23416 346 23446 372
rect 25208 350 25238 372
rect 23302 300 23318 334
rect 23352 300 23368 334
rect 23302 284 23368 300
rect 25190 334 25256 350
rect 25304 346 25334 372
rect 27096 350 27126 372
rect 25190 300 25206 334
rect 25240 300 25256 334
rect 25190 284 25256 300
rect 27078 334 27144 350
rect 27192 346 27222 372
rect 28984 350 29014 372
rect 27078 300 27094 334
rect 27128 300 27144 334
rect 27078 284 27144 300
rect 28966 334 29032 350
rect 29080 346 29110 372
rect 30872 350 30902 372
rect 28966 300 28982 334
rect 29016 300 29032 334
rect 28966 284 29032 300
rect 30854 334 30920 350
rect 30968 346 30998 372
rect 32760 350 32790 372
rect 30854 300 30870 334
rect 30904 300 30920 334
rect 30854 284 30920 300
rect 32742 334 32808 350
rect 32856 346 32886 372
rect 34648 350 34678 372
rect 32742 300 32758 334
rect 32792 300 32808 334
rect 32742 284 32808 300
rect 34630 334 34696 350
rect 34744 346 34774 372
rect 36536 350 36566 372
rect 34630 300 34646 334
rect 34680 300 34696 334
rect 34630 284 34696 300
rect 36518 334 36584 350
rect 36632 346 36662 372
rect 38424 350 38454 372
rect 36518 300 36534 334
rect 36568 300 36584 334
rect 36518 284 36584 300
rect 38406 334 38472 350
rect 38520 346 38550 372
rect 40312 350 40342 372
rect 38406 300 38422 334
rect 38456 300 38472 334
rect 38406 284 38472 300
rect 40294 334 40360 350
rect 40408 346 40438 372
rect 42200 350 42230 372
rect 40294 300 40310 334
rect 40344 300 40360 334
rect 40294 284 40360 300
rect 42182 334 42248 350
rect 42296 346 42326 372
rect 44088 350 44118 372
rect 42182 300 42198 334
rect 42232 300 42248 334
rect 42182 284 42248 300
rect 44070 334 44136 350
rect 44184 346 44214 372
rect 45970 350 46000 372
rect 44070 300 44086 334
rect 44120 300 44136 334
rect 44070 284 44136 300
rect 45952 334 46018 350
rect 46066 346 46096 372
rect 47858 350 47888 372
rect 45952 300 45968 334
rect 46002 300 46018 334
rect 45952 284 46018 300
rect 47840 334 47906 350
rect 47954 346 47984 372
rect 49746 350 49776 372
rect 47840 300 47856 334
rect 47890 300 47906 334
rect 47840 284 47906 300
rect 49728 334 49794 350
rect 49842 346 49872 372
rect 51634 350 51664 372
rect 49728 300 49744 334
rect 49778 300 49794 334
rect 49728 284 49794 300
rect 51616 334 51682 350
rect 51730 346 51760 372
rect 53522 350 53552 372
rect 51616 300 51632 334
rect 51666 300 51682 334
rect 51616 284 51682 300
rect 53504 334 53570 350
rect 53618 346 53648 372
rect 55410 350 55440 372
rect 53504 300 53520 334
rect 53554 300 53570 334
rect 53504 284 53570 300
rect 55392 334 55458 350
rect 55506 346 55536 372
rect 57298 350 57328 372
rect 55392 300 55408 334
rect 55442 300 55458 334
rect 55392 284 55458 300
rect 57280 334 57346 350
rect 57394 346 57424 372
rect 59186 350 59216 372
rect 57280 300 57296 334
rect 57330 300 57346 334
rect 57280 284 57346 300
rect 59168 334 59234 350
rect 59282 346 59312 372
rect 59168 300 59184 334
rect 59218 300 59234 334
rect 59168 284 59234 300
<< polycont >>
rect 764 7106 798 7140
rect 2652 7106 2686 7140
rect 4540 7106 4574 7140
rect 6428 7106 6462 7140
rect 8316 7106 8350 7140
rect 10204 7106 10238 7140
rect 12092 7106 12126 7140
rect 13980 7106 14014 7140
rect 15862 7106 15896 7140
rect 17750 7106 17784 7140
rect 19638 7106 19672 7140
rect 21526 7106 21560 7140
rect 23414 7106 23448 7140
rect 25302 7106 25336 7140
rect 27190 7106 27224 7140
rect 29078 7106 29112 7140
rect 30966 7106 31000 7140
rect 32854 7106 32888 7140
rect 34742 7106 34776 7140
rect 36630 7106 36664 7140
rect 38518 7106 38552 7140
rect 40406 7106 40440 7140
rect 42294 7106 42328 7140
rect 44182 7106 44216 7140
rect 46064 7106 46098 7140
rect 47952 7106 47986 7140
rect 49840 7106 49874 7140
rect 51728 7106 51762 7140
rect 53616 7106 53650 7140
rect 55504 7106 55538 7140
rect 57392 7106 57426 7140
rect 59280 7106 59314 7140
rect 668 6866 702 6900
rect 2556 6866 2590 6900
rect 780 6785 814 6819
rect -305 6600 -271 6634
rect -187 6613 -153 6647
rect 116 6611 150 6645
rect 354 6625 388 6659
rect 4444 6866 4478 6900
rect 1000 6625 1034 6659
rect 1312 6619 1346 6653
rect 2668 6785 2702 6819
rect 684 6457 718 6491
rect 354 6297 388 6331
rect 1583 6600 1617 6634
rect 1701 6613 1735 6647
rect 2004 6611 2038 6645
rect 2242 6625 2276 6659
rect 6332 6866 6366 6900
rect 2888 6625 2922 6659
rect 3200 6619 3234 6653
rect 4556 6785 4590 6819
rect 2572 6457 2606 6491
rect 1000 6297 1034 6331
rect 2242 6297 2276 6331
rect 3471 6600 3505 6634
rect 3589 6613 3623 6647
rect 3892 6611 3926 6645
rect 4130 6625 4164 6659
rect 8220 6866 8254 6900
rect 4776 6625 4810 6659
rect 5088 6619 5122 6653
rect 6444 6785 6478 6819
rect 4460 6457 4494 6491
rect 2888 6297 2922 6331
rect 4130 6297 4164 6331
rect 5359 6600 5393 6634
rect 5477 6613 5511 6647
rect 5780 6611 5814 6645
rect 6018 6625 6052 6659
rect 10108 6866 10142 6900
rect 6664 6625 6698 6659
rect 6976 6619 7010 6653
rect 8332 6785 8366 6819
rect 6348 6457 6382 6491
rect 4776 6297 4810 6331
rect 6018 6297 6052 6331
rect 7247 6600 7281 6634
rect 7365 6613 7399 6647
rect 7668 6611 7702 6645
rect 7906 6625 7940 6659
rect 11996 6866 12030 6900
rect 8552 6625 8586 6659
rect 8864 6619 8898 6653
rect 10220 6785 10254 6819
rect 8236 6457 8270 6491
rect 6664 6297 6698 6331
rect 7906 6297 7940 6331
rect 9135 6600 9169 6634
rect 9253 6613 9287 6647
rect 9556 6611 9590 6645
rect 9794 6625 9828 6659
rect 13884 6866 13918 6900
rect 10440 6625 10474 6659
rect 10752 6619 10786 6653
rect 12108 6785 12142 6819
rect 10124 6457 10158 6491
rect 8552 6297 8586 6331
rect 9794 6297 9828 6331
rect 11023 6600 11057 6634
rect 11141 6613 11175 6647
rect 11444 6611 11478 6645
rect 11682 6625 11716 6659
rect 15766 6866 15800 6900
rect 12328 6625 12362 6659
rect 12640 6619 12674 6653
rect 13996 6785 14030 6819
rect 12012 6457 12046 6491
rect 10440 6297 10474 6331
rect 11682 6297 11716 6331
rect 12911 6600 12945 6634
rect 13029 6613 13063 6647
rect 13332 6611 13366 6645
rect 13570 6625 13604 6659
rect 17654 6866 17688 6900
rect 14216 6625 14250 6659
rect 14528 6619 14562 6653
rect 15878 6785 15912 6819
rect 13900 6457 13934 6491
rect 12328 6297 12362 6331
rect 13570 6297 13604 6331
rect 14793 6600 14827 6634
rect 14911 6613 14945 6647
rect 15214 6611 15248 6645
rect 15452 6625 15486 6659
rect 19542 6866 19576 6900
rect 16098 6625 16132 6659
rect 16410 6619 16444 6653
rect 17766 6785 17800 6819
rect 15782 6457 15816 6491
rect 14216 6297 14250 6331
rect 15452 6297 15486 6331
rect 16681 6600 16715 6634
rect 16799 6613 16833 6647
rect 17102 6611 17136 6645
rect 17340 6625 17374 6659
rect 21430 6866 21464 6900
rect 17986 6625 18020 6659
rect 18298 6619 18332 6653
rect 19654 6785 19688 6819
rect 17670 6457 17704 6491
rect 16098 6297 16132 6331
rect 17340 6297 17374 6331
rect 18569 6600 18603 6634
rect 18687 6613 18721 6647
rect 18990 6611 19024 6645
rect 19228 6625 19262 6659
rect 23318 6866 23352 6900
rect 19874 6625 19908 6659
rect 20186 6619 20220 6653
rect 21542 6785 21576 6819
rect 19558 6457 19592 6491
rect 17986 6297 18020 6331
rect 19228 6297 19262 6331
rect 20457 6600 20491 6634
rect 20575 6613 20609 6647
rect 20878 6611 20912 6645
rect 21116 6625 21150 6659
rect 25206 6866 25240 6900
rect 21762 6625 21796 6659
rect 22074 6619 22108 6653
rect 23430 6785 23464 6819
rect 21446 6457 21480 6491
rect 19874 6297 19908 6331
rect 21116 6297 21150 6331
rect 22345 6600 22379 6634
rect 22463 6613 22497 6647
rect 22766 6611 22800 6645
rect 23004 6625 23038 6659
rect 27094 6866 27128 6900
rect 23650 6625 23684 6659
rect 23962 6619 23996 6653
rect 25318 6785 25352 6819
rect 23334 6457 23368 6491
rect 21762 6297 21796 6331
rect 23004 6297 23038 6331
rect 24233 6600 24267 6634
rect 24351 6613 24385 6647
rect 24654 6611 24688 6645
rect 24892 6625 24926 6659
rect 28982 6866 29016 6900
rect 25538 6625 25572 6659
rect 25850 6619 25884 6653
rect 27206 6785 27240 6819
rect 25222 6457 25256 6491
rect 23650 6297 23684 6331
rect 24892 6297 24926 6331
rect 26121 6600 26155 6634
rect 26239 6613 26273 6647
rect 26542 6611 26576 6645
rect 26780 6625 26814 6659
rect 30870 6866 30904 6900
rect 27426 6625 27460 6659
rect 27738 6619 27772 6653
rect 29094 6785 29128 6819
rect 27110 6457 27144 6491
rect 25538 6297 25572 6331
rect 26780 6297 26814 6331
rect 28009 6600 28043 6634
rect 28127 6613 28161 6647
rect 28430 6611 28464 6645
rect 28668 6625 28702 6659
rect 32758 6866 32792 6900
rect 29314 6625 29348 6659
rect 29626 6619 29660 6653
rect 30982 6785 31016 6819
rect 28998 6457 29032 6491
rect 27426 6297 27460 6331
rect 28668 6297 28702 6331
rect 29897 6600 29931 6634
rect 30015 6613 30049 6647
rect 30318 6611 30352 6645
rect 30556 6625 30590 6659
rect 34646 6866 34680 6900
rect 31202 6625 31236 6659
rect 31514 6619 31548 6653
rect 32870 6785 32904 6819
rect 30886 6457 30920 6491
rect 29314 6297 29348 6331
rect 30556 6297 30590 6331
rect 31785 6600 31819 6634
rect 31903 6613 31937 6647
rect 32206 6611 32240 6645
rect 32444 6625 32478 6659
rect 36534 6866 36568 6900
rect 33090 6625 33124 6659
rect 33402 6619 33436 6653
rect 34758 6785 34792 6819
rect 32774 6457 32808 6491
rect 31202 6297 31236 6331
rect 32444 6297 32478 6331
rect 33673 6600 33707 6634
rect 33791 6613 33825 6647
rect 34094 6611 34128 6645
rect 34332 6625 34366 6659
rect 38422 6866 38456 6900
rect 34978 6625 35012 6659
rect 35290 6619 35324 6653
rect 36646 6785 36680 6819
rect 34662 6457 34696 6491
rect 33090 6297 33124 6331
rect 34332 6297 34366 6331
rect 35561 6600 35595 6634
rect 35679 6613 35713 6647
rect 35982 6611 36016 6645
rect 36220 6625 36254 6659
rect 40310 6866 40344 6900
rect 36866 6625 36900 6659
rect 37178 6619 37212 6653
rect 38534 6785 38568 6819
rect 36550 6457 36584 6491
rect 34978 6297 35012 6331
rect 36220 6297 36254 6331
rect 37449 6600 37483 6634
rect 37567 6613 37601 6647
rect 37870 6611 37904 6645
rect 38108 6625 38142 6659
rect 42198 6866 42232 6900
rect 38754 6625 38788 6659
rect 39066 6619 39100 6653
rect 40422 6785 40456 6819
rect 38438 6457 38472 6491
rect 36866 6297 36900 6331
rect 38108 6297 38142 6331
rect 39337 6600 39371 6634
rect 39455 6613 39489 6647
rect 39758 6611 39792 6645
rect 39996 6625 40030 6659
rect 44086 6866 44120 6900
rect 40642 6625 40676 6659
rect 40954 6619 40988 6653
rect 42310 6785 42344 6819
rect 40326 6457 40360 6491
rect 38754 6297 38788 6331
rect 39996 6297 40030 6331
rect 41225 6600 41259 6634
rect 41343 6613 41377 6647
rect 41646 6611 41680 6645
rect 41884 6625 41918 6659
rect 45968 6866 46002 6900
rect 42530 6625 42564 6659
rect 42842 6619 42876 6653
rect 44198 6785 44232 6819
rect 42214 6457 42248 6491
rect 40642 6297 40676 6331
rect 41884 6297 41918 6331
rect 43113 6600 43147 6634
rect 43231 6613 43265 6647
rect 43534 6611 43568 6645
rect 43772 6625 43806 6659
rect 47856 6866 47890 6900
rect 44418 6625 44452 6659
rect 44730 6619 44764 6653
rect 46080 6785 46114 6819
rect 44102 6457 44136 6491
rect 42530 6297 42564 6331
rect 43772 6297 43806 6331
rect 44995 6600 45029 6634
rect 45113 6613 45147 6647
rect 45416 6611 45450 6645
rect 45654 6625 45688 6659
rect 49744 6866 49778 6900
rect 46300 6625 46334 6659
rect 46612 6619 46646 6653
rect 47968 6785 48002 6819
rect 45984 6457 46018 6491
rect 44418 6297 44452 6331
rect 45654 6297 45688 6331
rect 46883 6600 46917 6634
rect 47001 6613 47035 6647
rect 47304 6611 47338 6645
rect 47542 6625 47576 6659
rect 51632 6866 51666 6900
rect 48188 6625 48222 6659
rect 48500 6619 48534 6653
rect 49856 6785 49890 6819
rect 47872 6457 47906 6491
rect 46300 6297 46334 6331
rect 47542 6297 47576 6331
rect 48771 6600 48805 6634
rect 48889 6613 48923 6647
rect 49192 6611 49226 6645
rect 49430 6625 49464 6659
rect 53520 6866 53554 6900
rect 50076 6625 50110 6659
rect 50388 6619 50422 6653
rect 51744 6785 51778 6819
rect 49760 6457 49794 6491
rect 48188 6297 48222 6331
rect 49430 6297 49464 6331
rect 50659 6600 50693 6634
rect 50777 6613 50811 6647
rect 51080 6611 51114 6645
rect 51318 6625 51352 6659
rect 55408 6866 55442 6900
rect 51964 6625 51998 6659
rect 52276 6619 52310 6653
rect 53632 6785 53666 6819
rect 51648 6457 51682 6491
rect 50076 6297 50110 6331
rect 51318 6297 51352 6331
rect 52547 6600 52581 6634
rect 52665 6613 52699 6647
rect 52968 6611 53002 6645
rect 53206 6625 53240 6659
rect 57296 6866 57330 6900
rect 53852 6625 53886 6659
rect 54164 6619 54198 6653
rect 55520 6785 55554 6819
rect 53536 6457 53570 6491
rect 51964 6297 51998 6331
rect 53206 6297 53240 6331
rect 54435 6600 54469 6634
rect 54553 6613 54587 6647
rect 54856 6611 54890 6645
rect 55094 6625 55128 6659
rect 59184 6866 59218 6900
rect 55740 6625 55774 6659
rect 56052 6619 56086 6653
rect 57408 6785 57442 6819
rect 55424 6457 55458 6491
rect 53852 6297 53886 6331
rect 55094 6297 55128 6331
rect 56323 6600 56357 6634
rect 56441 6613 56475 6647
rect 56744 6611 56778 6645
rect 56982 6625 57016 6659
rect 57628 6625 57662 6659
rect 57940 6619 57974 6653
rect 59296 6785 59330 6819
rect 57312 6457 57346 6491
rect 55740 6297 55774 6331
rect 56982 6297 57016 6331
rect 58211 6600 58245 6634
rect 58329 6613 58363 6647
rect 58632 6611 58666 6645
rect 58870 6625 58904 6659
rect 59516 6625 59550 6659
rect 59828 6619 59862 6653
rect 59200 6457 59234 6491
rect 57628 6297 57662 6331
rect 58870 6297 58904 6331
rect 59516 6297 59550 6331
rect 762 6050 796 6084
rect 2650 6050 2684 6084
rect 4538 6050 4572 6084
rect 6426 6050 6460 6084
rect 8314 6050 8348 6084
rect 10202 6050 10236 6084
rect 12090 6050 12124 6084
rect 13978 6050 14012 6084
rect 15860 6050 15894 6084
rect 17748 6050 17782 6084
rect 19636 6050 19670 6084
rect 21524 6050 21558 6084
rect 23412 6050 23446 6084
rect 25300 6050 25334 6084
rect 27188 6050 27222 6084
rect 29076 6050 29110 6084
rect 30964 6050 30998 6084
rect 32852 6050 32886 6084
rect 34740 6050 34774 6084
rect 36628 6050 36662 6084
rect 38516 6050 38550 6084
rect 40404 6050 40438 6084
rect 42292 6050 42326 6084
rect 44180 6050 44214 6084
rect 46062 6050 46096 6084
rect 47950 6050 47984 6084
rect 49838 6050 49872 6084
rect 51726 6050 51760 6084
rect 53614 6050 53648 6084
rect 55502 6050 55536 6084
rect 57390 6050 57424 6084
rect 59278 6050 59312 6084
rect 666 5810 700 5844
rect 2554 5810 2588 5844
rect 4442 5810 4476 5844
rect 778 5729 812 5763
rect 195 5565 229 5599
rect 363 5565 397 5599
rect 6330 5810 6364 5844
rect 2666 5729 2700 5763
rect 1009 5565 1043 5599
rect 1177 5565 1211 5599
rect 2083 5565 2117 5599
rect 2251 5565 2285 5599
rect 682 5401 716 5435
rect 8218 5810 8252 5844
rect 4554 5729 4588 5763
rect 2897 5565 2931 5599
rect 3065 5565 3099 5599
rect 3971 5565 4005 5599
rect 4139 5565 4173 5599
rect 2570 5401 2604 5435
rect 10106 5810 10140 5844
rect 6442 5729 6476 5763
rect 4785 5565 4819 5599
rect 4953 5565 4987 5599
rect 5859 5565 5893 5599
rect 6027 5565 6061 5599
rect 4458 5401 4492 5435
rect 11994 5810 12028 5844
rect 8330 5729 8364 5763
rect 6673 5565 6707 5599
rect 6841 5565 6875 5599
rect 7747 5565 7781 5599
rect 7915 5565 7949 5599
rect 6346 5401 6380 5435
rect 13882 5810 13916 5844
rect 10218 5729 10252 5763
rect 8561 5565 8595 5599
rect 8729 5565 8763 5599
rect 9635 5565 9669 5599
rect 9803 5565 9837 5599
rect 8234 5401 8268 5435
rect 15764 5810 15798 5844
rect 12106 5729 12140 5763
rect 10449 5565 10483 5599
rect 10617 5565 10651 5599
rect 11523 5565 11557 5599
rect 11691 5565 11725 5599
rect 10122 5401 10156 5435
rect 17652 5810 17686 5844
rect 13994 5729 14028 5763
rect 12337 5565 12371 5599
rect 12505 5565 12539 5599
rect 13411 5565 13445 5599
rect 13579 5565 13613 5599
rect 12010 5401 12044 5435
rect 19540 5810 19574 5844
rect 15876 5729 15910 5763
rect 14225 5565 14259 5599
rect 14393 5565 14427 5599
rect 15293 5565 15327 5599
rect 15461 5565 15495 5599
rect 13898 5401 13932 5435
rect 21428 5810 21462 5844
rect 17764 5729 17798 5763
rect 16107 5565 16141 5599
rect 16275 5565 16309 5599
rect 17181 5565 17215 5599
rect 17349 5565 17383 5599
rect 15780 5401 15814 5435
rect 23316 5810 23350 5844
rect 19652 5729 19686 5763
rect 17995 5565 18029 5599
rect 18163 5565 18197 5599
rect 19069 5565 19103 5599
rect 19237 5565 19271 5599
rect 17668 5401 17702 5435
rect 25204 5810 25238 5844
rect 21540 5729 21574 5763
rect 19883 5565 19917 5599
rect 20051 5565 20085 5599
rect 20957 5565 20991 5599
rect 21125 5565 21159 5599
rect 19556 5401 19590 5435
rect 27092 5810 27126 5844
rect 23428 5729 23462 5763
rect 21771 5565 21805 5599
rect 21939 5565 21973 5599
rect 22845 5565 22879 5599
rect 23013 5565 23047 5599
rect 21444 5401 21478 5435
rect 28980 5810 29014 5844
rect 25316 5729 25350 5763
rect 23659 5565 23693 5599
rect 23827 5565 23861 5599
rect 24733 5565 24767 5599
rect 24901 5565 24935 5599
rect 23332 5401 23366 5435
rect 30868 5810 30902 5844
rect 27204 5729 27238 5763
rect 25547 5565 25581 5599
rect 25715 5565 25749 5599
rect 26621 5565 26655 5599
rect 26789 5565 26823 5599
rect 25220 5401 25254 5435
rect 32756 5810 32790 5844
rect 29092 5729 29126 5763
rect 27435 5565 27469 5599
rect 27603 5565 27637 5599
rect 28509 5565 28543 5599
rect 28677 5565 28711 5599
rect 27108 5401 27142 5435
rect 34644 5810 34678 5844
rect 30980 5729 31014 5763
rect 29323 5565 29357 5599
rect 29491 5565 29525 5599
rect 30397 5565 30431 5599
rect 30565 5565 30599 5599
rect 28996 5401 29030 5435
rect 36532 5810 36566 5844
rect 32868 5729 32902 5763
rect 31211 5565 31245 5599
rect 31379 5565 31413 5599
rect 32285 5565 32319 5599
rect 32453 5565 32487 5599
rect 30884 5401 30918 5435
rect 38420 5810 38454 5844
rect 34756 5729 34790 5763
rect 33099 5565 33133 5599
rect 33267 5565 33301 5599
rect 34173 5565 34207 5599
rect 34341 5565 34375 5599
rect 32772 5401 32806 5435
rect 40308 5810 40342 5844
rect 36644 5729 36678 5763
rect 34987 5565 35021 5599
rect 35155 5565 35189 5599
rect 36061 5565 36095 5599
rect 36229 5565 36263 5599
rect 34660 5401 34694 5435
rect 42196 5810 42230 5844
rect 38532 5729 38566 5763
rect 36875 5565 36909 5599
rect 37043 5565 37077 5599
rect 37949 5565 37983 5599
rect 38117 5565 38151 5599
rect 36548 5401 36582 5435
rect 44084 5810 44118 5844
rect 40420 5729 40454 5763
rect 38763 5565 38797 5599
rect 38931 5565 38965 5599
rect 39837 5565 39871 5599
rect 40005 5565 40039 5599
rect 38436 5401 38470 5435
rect 45966 5810 46000 5844
rect 42308 5729 42342 5763
rect 40651 5565 40685 5599
rect 40819 5565 40853 5599
rect 41725 5565 41759 5599
rect 41893 5565 41927 5599
rect 40324 5401 40358 5435
rect 47854 5810 47888 5844
rect 44196 5729 44230 5763
rect 42539 5565 42573 5599
rect 42707 5565 42741 5599
rect 43613 5565 43647 5599
rect 43781 5565 43815 5599
rect 42212 5401 42246 5435
rect 49742 5810 49776 5844
rect 46078 5729 46112 5763
rect 44427 5565 44461 5599
rect 44595 5565 44629 5599
rect 45495 5565 45529 5599
rect 45663 5565 45697 5599
rect 44100 5401 44134 5435
rect 51630 5810 51664 5844
rect 47966 5729 48000 5763
rect 46309 5565 46343 5599
rect 46477 5565 46511 5599
rect 47383 5565 47417 5599
rect 47551 5565 47585 5599
rect 45982 5401 46016 5435
rect 53518 5810 53552 5844
rect 49854 5729 49888 5763
rect 48197 5565 48231 5599
rect 48365 5565 48399 5599
rect 49271 5565 49305 5599
rect 49439 5565 49473 5599
rect 47870 5401 47904 5435
rect 55406 5810 55440 5844
rect 51742 5729 51776 5763
rect 50085 5565 50119 5599
rect 50253 5565 50287 5599
rect 51159 5565 51193 5599
rect 51327 5565 51361 5599
rect 49758 5401 49792 5435
rect 57294 5810 57328 5844
rect 53630 5729 53664 5763
rect 51973 5565 52007 5599
rect 52141 5565 52175 5599
rect 53047 5565 53081 5599
rect 53215 5565 53249 5599
rect 51646 5401 51680 5435
rect 59182 5810 59216 5844
rect 55518 5729 55552 5763
rect 53861 5565 53895 5599
rect 54029 5565 54063 5599
rect 54935 5565 54969 5599
rect 55103 5565 55137 5599
rect 53534 5401 53568 5435
rect 57406 5729 57440 5763
rect 55749 5565 55783 5599
rect 55917 5565 55951 5599
rect 56823 5565 56857 5599
rect 56991 5565 57025 5599
rect 55422 5401 55456 5435
rect 59294 5729 59328 5763
rect 57637 5565 57671 5599
rect 57805 5565 57839 5599
rect 58711 5565 58745 5599
rect 58879 5565 58913 5599
rect 57310 5401 57344 5435
rect 59525 5565 59559 5599
rect 59693 5565 59727 5599
rect 59198 5401 59232 5435
rect 6047 4863 6081 4897
rect 6214 4863 6248 4897
rect 6382 4863 6416 4897
rect 6549 4863 6583 4897
rect 6718 4863 6752 4897
rect 6886 4863 6920 4897
rect 7060 4863 7094 4897
rect 7929 4861 7963 4895
rect 8096 4861 8130 4895
rect 8264 4861 8298 4895
rect 8431 4861 8465 4895
rect 8600 4861 8634 4895
rect 8768 4861 8802 4895
rect 8942 4861 8976 4895
rect 21145 4863 21179 4897
rect 21312 4863 21346 4897
rect 21480 4863 21514 4897
rect 21647 4863 21681 4897
rect 21816 4863 21850 4897
rect 21984 4863 22018 4897
rect 22158 4863 22192 4897
rect 23027 4861 23061 4895
rect 23194 4861 23228 4895
rect 23362 4861 23396 4895
rect 23529 4861 23563 4895
rect 23698 4861 23732 4895
rect 23866 4861 23900 4895
rect 24040 4861 24074 4895
rect 36249 4863 36283 4897
rect 36416 4863 36450 4897
rect 36584 4863 36618 4897
rect 36751 4863 36785 4897
rect 36920 4863 36954 4897
rect 37088 4863 37122 4897
rect 37262 4863 37296 4897
rect 38131 4861 38165 4895
rect 38298 4861 38332 4895
rect 38466 4861 38500 4895
rect 38633 4861 38667 4895
rect 38802 4861 38836 4895
rect 38970 4861 39004 4895
rect 39144 4861 39178 4895
rect 51347 4863 51381 4897
rect 51514 4863 51548 4897
rect 51682 4863 51716 4897
rect 51849 4863 51883 4897
rect 52018 4863 52052 4897
rect 52186 4863 52220 4897
rect 52360 4863 52394 4897
rect 53229 4861 53263 4895
rect 53396 4861 53430 4895
rect 53564 4861 53598 4895
rect 53731 4861 53765 4895
rect 53900 4861 53934 4895
rect 54068 4861 54102 4895
rect 54242 4861 54276 4895
rect 30064 3786 30098 3820
rect 30156 3786 30190 3820
rect 30240 3786 30274 3820
rect 30324 3786 30358 3820
rect 30597 3786 30631 3820
rect 30771 3786 30805 3820
rect 30939 3786 30973 3820
rect 31108 3786 31142 3820
rect 31275 3786 31309 3820
rect 31443 3786 31477 3820
rect 31610 3786 31644 3820
rect 43423 3570 43457 3604
rect 43597 3570 43631 3604
rect 43765 3570 43799 3604
rect 43934 3570 43968 3604
rect 44101 3570 44135 3604
rect 44269 3570 44303 3604
rect 44436 3570 44470 3604
rect 45353 3570 45387 3604
rect 45527 3570 45561 3604
rect 45695 3570 45729 3604
rect 45864 3570 45898 3604
rect 46031 3570 46065 3604
rect 46199 3570 46233 3604
rect 46366 3570 46400 3604
rect 13281 3410 13315 3444
rect 13455 3410 13489 3444
rect 13623 3410 13657 3444
rect 13792 3410 13826 3444
rect 13959 3410 13993 3444
rect 14127 3410 14161 3444
rect 14294 3410 14328 3444
rect 15211 3410 15245 3444
rect 15385 3410 15419 3444
rect 15553 3410 15587 3444
rect 15722 3410 15756 3444
rect 15889 3410 15923 3444
rect 16057 3410 16091 3444
rect 16224 3410 16258 3444
rect 5706 2545 5740 2579
rect 5880 2545 5914 2579
rect 6048 2545 6082 2579
rect 6217 2545 6251 2579
rect 6384 2545 6418 2579
rect 6552 2545 6586 2579
rect 6719 2545 6753 2579
rect 7588 2543 7622 2577
rect 7762 2543 7796 2577
rect 7930 2543 7964 2577
rect 8099 2543 8133 2577
rect 8266 2543 8300 2577
rect 8434 2543 8468 2577
rect 8601 2543 8635 2577
rect 20804 2545 20838 2579
rect 20978 2545 21012 2579
rect 21146 2545 21180 2579
rect 21315 2545 21349 2579
rect 21482 2545 21516 2579
rect 21650 2545 21684 2579
rect 21817 2545 21851 2579
rect 22686 2543 22720 2577
rect 22860 2543 22894 2577
rect 23028 2543 23062 2577
rect 23197 2543 23231 2577
rect 23364 2543 23398 2577
rect 23532 2543 23566 2577
rect 23699 2543 23733 2577
rect 35908 2545 35942 2579
rect 36082 2545 36116 2579
rect 36250 2545 36284 2579
rect 36419 2545 36453 2579
rect 36586 2545 36620 2579
rect 36754 2545 36788 2579
rect 36921 2545 36955 2579
rect 37790 2543 37824 2577
rect 37964 2543 37998 2577
rect 38132 2543 38166 2577
rect 38301 2543 38335 2577
rect 38468 2543 38502 2577
rect 38636 2543 38670 2577
rect 38803 2543 38837 2577
rect 51006 2545 51040 2579
rect 51180 2545 51214 2579
rect 51348 2545 51382 2579
rect 51517 2545 51551 2579
rect 51684 2545 51718 2579
rect 51852 2545 51886 2579
rect 52019 2545 52053 2579
rect 52888 2543 52922 2577
rect 53062 2543 53096 2577
rect 53230 2543 53264 2577
rect 53399 2543 53433 2577
rect 53566 2543 53600 2577
rect 53734 2543 53768 2577
rect 53901 2543 53935 2577
rect 750 2005 784 2039
rect 255 1841 289 1875
rect 423 1841 457 1875
rect 2638 2005 2672 2039
rect 1069 1841 1103 1875
rect 1237 1841 1271 1875
rect 2143 1841 2177 1875
rect 2311 1841 2345 1875
rect 654 1677 688 1711
rect 4526 2005 4560 2039
rect 2957 1841 2991 1875
rect 3125 1841 3159 1875
rect 4031 1841 4065 1875
rect 4199 1841 4233 1875
rect 2542 1677 2576 1711
rect 6414 2005 6448 2039
rect 4845 1841 4879 1875
rect 5013 1841 5047 1875
rect 5919 1841 5953 1875
rect 6087 1841 6121 1875
rect 4430 1677 4464 1711
rect 766 1596 800 1630
rect 8302 2005 8336 2039
rect 6733 1841 6767 1875
rect 6901 1841 6935 1875
rect 7807 1841 7841 1875
rect 7975 1841 8009 1875
rect 6318 1677 6352 1711
rect 2654 1596 2688 1630
rect 10190 2005 10224 2039
rect 8621 1841 8655 1875
rect 8789 1841 8823 1875
rect 9695 1841 9729 1875
rect 9863 1841 9897 1875
rect 8206 1677 8240 1711
rect 4542 1596 4576 1630
rect 12078 2005 12112 2039
rect 10509 1841 10543 1875
rect 10677 1841 10711 1875
rect 11583 1841 11617 1875
rect 11751 1841 11785 1875
rect 10094 1677 10128 1711
rect 6430 1596 6464 1630
rect 13966 2005 14000 2039
rect 12397 1841 12431 1875
rect 12565 1841 12599 1875
rect 13471 1841 13505 1875
rect 13639 1841 13673 1875
rect 11982 1677 12016 1711
rect 8318 1596 8352 1630
rect 15848 2005 15882 2039
rect 14285 1841 14319 1875
rect 14453 1841 14487 1875
rect 15353 1841 15387 1875
rect 15521 1841 15555 1875
rect 13870 1677 13904 1711
rect 10206 1596 10240 1630
rect 17736 2005 17770 2039
rect 16167 1841 16201 1875
rect 16335 1841 16369 1875
rect 17241 1841 17275 1875
rect 17409 1841 17443 1875
rect 15752 1677 15786 1711
rect 12094 1596 12128 1630
rect 19624 2005 19658 2039
rect 18055 1841 18089 1875
rect 18223 1841 18257 1875
rect 19129 1841 19163 1875
rect 19297 1841 19331 1875
rect 17640 1677 17674 1711
rect 13982 1596 14016 1630
rect 21512 2005 21546 2039
rect 19943 1841 19977 1875
rect 20111 1841 20145 1875
rect 21017 1841 21051 1875
rect 21185 1841 21219 1875
rect 19528 1677 19562 1711
rect 15864 1596 15898 1630
rect 23400 2005 23434 2039
rect 21831 1841 21865 1875
rect 21999 1841 22033 1875
rect 22905 1841 22939 1875
rect 23073 1841 23107 1875
rect 21416 1677 21450 1711
rect 17752 1596 17786 1630
rect 25288 2005 25322 2039
rect 23719 1841 23753 1875
rect 23887 1841 23921 1875
rect 24793 1841 24827 1875
rect 24961 1841 24995 1875
rect 23304 1677 23338 1711
rect 19640 1596 19674 1630
rect 27176 2005 27210 2039
rect 25607 1841 25641 1875
rect 25775 1841 25809 1875
rect 26681 1841 26715 1875
rect 26849 1841 26883 1875
rect 25192 1677 25226 1711
rect 21528 1596 21562 1630
rect 29064 2005 29098 2039
rect 27495 1841 27529 1875
rect 27663 1841 27697 1875
rect 28569 1841 28603 1875
rect 28737 1841 28771 1875
rect 27080 1677 27114 1711
rect 23416 1596 23450 1630
rect 30952 2005 30986 2039
rect 29383 1841 29417 1875
rect 29551 1841 29585 1875
rect 30457 1841 30491 1875
rect 30625 1841 30659 1875
rect 28968 1677 29002 1711
rect 25304 1596 25338 1630
rect 32840 2005 32874 2039
rect 31271 1841 31305 1875
rect 31439 1841 31473 1875
rect 32345 1841 32379 1875
rect 32513 1841 32547 1875
rect 30856 1677 30890 1711
rect 27192 1596 27226 1630
rect 34728 2005 34762 2039
rect 33159 1841 33193 1875
rect 33327 1841 33361 1875
rect 34233 1841 34267 1875
rect 34401 1841 34435 1875
rect 32744 1677 32778 1711
rect 29080 1596 29114 1630
rect 36616 2005 36650 2039
rect 35047 1841 35081 1875
rect 35215 1841 35249 1875
rect 36121 1841 36155 1875
rect 36289 1841 36323 1875
rect 34632 1677 34666 1711
rect 30968 1596 31002 1630
rect 38504 2005 38538 2039
rect 36935 1841 36969 1875
rect 37103 1841 37137 1875
rect 38009 1841 38043 1875
rect 38177 1841 38211 1875
rect 36520 1677 36554 1711
rect 32856 1596 32890 1630
rect 40392 2005 40426 2039
rect 38823 1841 38857 1875
rect 38991 1841 39025 1875
rect 39897 1841 39931 1875
rect 40065 1841 40099 1875
rect 38408 1677 38442 1711
rect 34744 1596 34778 1630
rect 42280 2005 42314 2039
rect 40711 1841 40745 1875
rect 40879 1841 40913 1875
rect 41785 1841 41819 1875
rect 41953 1841 41987 1875
rect 40296 1677 40330 1711
rect 36632 1596 36666 1630
rect 44168 2005 44202 2039
rect 42599 1841 42633 1875
rect 42767 1841 42801 1875
rect 43673 1841 43707 1875
rect 43841 1841 43875 1875
rect 42184 1677 42218 1711
rect 38520 1596 38554 1630
rect 46050 2005 46084 2039
rect 44487 1841 44521 1875
rect 44655 1841 44689 1875
rect 45555 1841 45589 1875
rect 45723 1841 45757 1875
rect 44072 1677 44106 1711
rect 40408 1596 40442 1630
rect 47938 2005 47972 2039
rect 46369 1841 46403 1875
rect 46537 1841 46571 1875
rect 47443 1841 47477 1875
rect 47611 1841 47645 1875
rect 45954 1677 45988 1711
rect 42296 1596 42330 1630
rect 49826 2005 49860 2039
rect 48257 1841 48291 1875
rect 48425 1841 48459 1875
rect 49331 1841 49365 1875
rect 49499 1841 49533 1875
rect 47842 1677 47876 1711
rect 44184 1596 44218 1630
rect 51714 2005 51748 2039
rect 50145 1841 50179 1875
rect 50313 1841 50347 1875
rect 51219 1841 51253 1875
rect 51387 1841 51421 1875
rect 49730 1677 49764 1711
rect 46066 1596 46100 1630
rect 53602 2005 53636 2039
rect 52033 1841 52067 1875
rect 52201 1841 52235 1875
rect 53107 1841 53141 1875
rect 53275 1841 53309 1875
rect 51618 1677 51652 1711
rect 47954 1596 47988 1630
rect 55490 2005 55524 2039
rect 53921 1841 53955 1875
rect 54089 1841 54123 1875
rect 54995 1841 55029 1875
rect 55163 1841 55197 1875
rect 53506 1677 53540 1711
rect 49842 1596 49876 1630
rect 57378 2005 57412 2039
rect 55809 1841 55843 1875
rect 55977 1841 56011 1875
rect 56883 1841 56917 1875
rect 57051 1841 57085 1875
rect 55394 1677 55428 1711
rect 51730 1596 51764 1630
rect 59266 2005 59300 2039
rect 57697 1841 57731 1875
rect 57865 1841 57899 1875
rect 58771 1841 58805 1875
rect 58939 1841 58973 1875
rect 57282 1677 57316 1711
rect 53618 1596 53652 1630
rect 59585 1841 59619 1875
rect 59753 1841 59787 1875
rect 59170 1677 59204 1711
rect 55506 1596 55540 1630
rect 57394 1596 57428 1630
rect 59282 1596 59316 1630
rect 670 1356 704 1390
rect 2558 1356 2592 1390
rect 4446 1356 4480 1390
rect 6334 1356 6368 1390
rect 8222 1356 8256 1390
rect 10110 1356 10144 1390
rect 11998 1356 12032 1390
rect 13886 1356 13920 1390
rect 15768 1356 15802 1390
rect 17656 1356 17690 1390
rect 19544 1356 19578 1390
rect 21432 1356 21466 1390
rect 23320 1356 23354 1390
rect 25208 1356 25242 1390
rect 27096 1356 27130 1390
rect 28984 1356 29018 1390
rect 30872 1356 30906 1390
rect 32760 1356 32794 1390
rect 34648 1356 34682 1390
rect 36536 1356 36570 1390
rect 38424 1356 38458 1390
rect 40312 1356 40346 1390
rect 42200 1356 42234 1390
rect 44088 1356 44122 1390
rect 45970 1356 46004 1390
rect 47858 1356 47892 1390
rect 49746 1356 49780 1390
rect 51634 1356 51668 1390
rect 53522 1356 53556 1390
rect 55410 1356 55444 1390
rect 57298 1356 57332 1390
rect 59186 1356 59220 1390
rect 432 1109 466 1143
rect 1078 1109 1112 1143
rect 2320 1109 2354 1143
rect 748 949 782 983
rect 120 787 154 821
rect 432 781 466 815
rect 1078 781 1112 815
rect 1316 795 1350 829
rect 1619 793 1653 827
rect 1737 806 1771 840
rect 2966 1109 3000 1143
rect 4208 1109 4242 1143
rect 2636 949 2670 983
rect 652 621 686 655
rect 2008 787 2042 821
rect 2320 781 2354 815
rect 2966 781 3000 815
rect 3204 795 3238 829
rect 3507 793 3541 827
rect 3625 806 3659 840
rect 4854 1109 4888 1143
rect 6096 1109 6130 1143
rect 4524 949 4558 983
rect 2540 621 2574 655
rect 3896 787 3930 821
rect 4208 781 4242 815
rect 764 540 798 574
rect 4854 781 4888 815
rect 5092 795 5126 829
rect 5395 793 5429 827
rect 5513 806 5547 840
rect 6742 1109 6776 1143
rect 7984 1109 8018 1143
rect 6412 949 6446 983
rect 4428 621 4462 655
rect 5784 787 5818 821
rect 6096 781 6130 815
rect 2652 540 2686 574
rect 6742 781 6776 815
rect 6980 795 7014 829
rect 7283 793 7317 827
rect 7401 806 7435 840
rect 8630 1109 8664 1143
rect 9872 1109 9906 1143
rect 8300 949 8334 983
rect 6316 621 6350 655
rect 7672 787 7706 821
rect 7984 781 8018 815
rect 4540 540 4574 574
rect 8630 781 8664 815
rect 8868 795 8902 829
rect 9171 793 9205 827
rect 9289 806 9323 840
rect 10518 1109 10552 1143
rect 11760 1109 11794 1143
rect 10188 949 10222 983
rect 8204 621 8238 655
rect 9560 787 9594 821
rect 9872 781 9906 815
rect 6428 540 6462 574
rect 10518 781 10552 815
rect 10756 795 10790 829
rect 11059 793 11093 827
rect 11177 806 11211 840
rect 12406 1109 12440 1143
rect 13648 1109 13682 1143
rect 12076 949 12110 983
rect 10092 621 10126 655
rect 11448 787 11482 821
rect 11760 781 11794 815
rect 8316 540 8350 574
rect 12406 781 12440 815
rect 12644 795 12678 829
rect 12947 793 12981 827
rect 13065 806 13099 840
rect 14294 1109 14328 1143
rect 15530 1109 15564 1143
rect 13964 949 13998 983
rect 11980 621 12014 655
rect 13336 787 13370 821
rect 13648 781 13682 815
rect 10204 540 10238 574
rect 14294 781 14328 815
rect 14532 795 14566 829
rect 14835 793 14869 827
rect 14953 806 14987 840
rect 16176 1109 16210 1143
rect 17418 1109 17452 1143
rect 15846 949 15880 983
rect 13868 621 13902 655
rect 15218 787 15252 821
rect 15530 781 15564 815
rect 12092 540 12126 574
rect 16176 781 16210 815
rect 16414 795 16448 829
rect 16717 793 16751 827
rect 16835 806 16869 840
rect 18064 1109 18098 1143
rect 19306 1109 19340 1143
rect 17734 949 17768 983
rect 15750 621 15784 655
rect 17106 787 17140 821
rect 17418 781 17452 815
rect 13980 540 14014 574
rect 18064 781 18098 815
rect 18302 795 18336 829
rect 18605 793 18639 827
rect 18723 806 18757 840
rect 19952 1109 19986 1143
rect 21194 1109 21228 1143
rect 19622 949 19656 983
rect 17638 621 17672 655
rect 18994 787 19028 821
rect 19306 781 19340 815
rect 15862 540 15896 574
rect 19952 781 19986 815
rect 20190 795 20224 829
rect 20493 793 20527 827
rect 20611 806 20645 840
rect 21840 1109 21874 1143
rect 23082 1109 23116 1143
rect 21510 949 21544 983
rect 19526 621 19560 655
rect 20882 787 20916 821
rect 21194 781 21228 815
rect 17750 540 17784 574
rect 21840 781 21874 815
rect 22078 795 22112 829
rect 22381 793 22415 827
rect 22499 806 22533 840
rect 23728 1109 23762 1143
rect 24970 1109 25004 1143
rect 23398 949 23432 983
rect 21414 621 21448 655
rect 22770 787 22804 821
rect 23082 781 23116 815
rect 19638 540 19672 574
rect 23728 781 23762 815
rect 23966 795 24000 829
rect 24269 793 24303 827
rect 24387 806 24421 840
rect 25616 1109 25650 1143
rect 26858 1109 26892 1143
rect 25286 949 25320 983
rect 23302 621 23336 655
rect 24658 787 24692 821
rect 24970 781 25004 815
rect 21526 540 21560 574
rect 25616 781 25650 815
rect 25854 795 25888 829
rect 26157 793 26191 827
rect 26275 806 26309 840
rect 27504 1109 27538 1143
rect 28746 1109 28780 1143
rect 27174 949 27208 983
rect 25190 621 25224 655
rect 26546 787 26580 821
rect 26858 781 26892 815
rect 23414 540 23448 574
rect 27504 781 27538 815
rect 27742 795 27776 829
rect 28045 793 28079 827
rect 28163 806 28197 840
rect 29392 1109 29426 1143
rect 30634 1109 30668 1143
rect 29062 949 29096 983
rect 27078 621 27112 655
rect 28434 787 28468 821
rect 28746 781 28780 815
rect 25302 540 25336 574
rect 29392 781 29426 815
rect 29630 795 29664 829
rect 29933 793 29967 827
rect 30051 806 30085 840
rect 31280 1109 31314 1143
rect 32522 1109 32556 1143
rect 30950 949 30984 983
rect 28966 621 29000 655
rect 30322 787 30356 821
rect 30634 781 30668 815
rect 27190 540 27224 574
rect 31280 781 31314 815
rect 31518 795 31552 829
rect 31821 793 31855 827
rect 31939 806 31973 840
rect 33168 1109 33202 1143
rect 34410 1109 34444 1143
rect 32838 949 32872 983
rect 30854 621 30888 655
rect 32210 787 32244 821
rect 32522 781 32556 815
rect 29078 540 29112 574
rect 33168 781 33202 815
rect 33406 795 33440 829
rect 33709 793 33743 827
rect 33827 806 33861 840
rect 35056 1109 35090 1143
rect 36298 1109 36332 1143
rect 34726 949 34760 983
rect 32742 621 32776 655
rect 34098 787 34132 821
rect 34410 781 34444 815
rect 30966 540 31000 574
rect 35056 781 35090 815
rect 35294 795 35328 829
rect 35597 793 35631 827
rect 35715 806 35749 840
rect 36944 1109 36978 1143
rect 38186 1109 38220 1143
rect 36614 949 36648 983
rect 34630 621 34664 655
rect 35986 787 36020 821
rect 36298 781 36332 815
rect 32854 540 32888 574
rect 36944 781 36978 815
rect 37182 795 37216 829
rect 37485 793 37519 827
rect 37603 806 37637 840
rect 38832 1109 38866 1143
rect 40074 1109 40108 1143
rect 38502 949 38536 983
rect 36518 621 36552 655
rect 37874 787 37908 821
rect 38186 781 38220 815
rect 34742 540 34776 574
rect 38832 781 38866 815
rect 39070 795 39104 829
rect 39373 793 39407 827
rect 39491 806 39525 840
rect 40720 1109 40754 1143
rect 41962 1109 41996 1143
rect 40390 949 40424 983
rect 38406 621 38440 655
rect 39762 787 39796 821
rect 40074 781 40108 815
rect 36630 540 36664 574
rect 40720 781 40754 815
rect 40958 795 40992 829
rect 41261 793 41295 827
rect 41379 806 41413 840
rect 42608 1109 42642 1143
rect 43850 1109 43884 1143
rect 42278 949 42312 983
rect 40294 621 40328 655
rect 41650 787 41684 821
rect 41962 781 41996 815
rect 38518 540 38552 574
rect 42608 781 42642 815
rect 42846 795 42880 829
rect 43149 793 43183 827
rect 43267 806 43301 840
rect 44496 1109 44530 1143
rect 45732 1109 45766 1143
rect 44166 949 44200 983
rect 42182 621 42216 655
rect 43538 787 43572 821
rect 43850 781 43884 815
rect 40406 540 40440 574
rect 44496 781 44530 815
rect 44734 795 44768 829
rect 45037 793 45071 827
rect 45155 806 45189 840
rect 46378 1109 46412 1143
rect 47620 1109 47654 1143
rect 46048 949 46082 983
rect 44070 621 44104 655
rect 45420 787 45454 821
rect 45732 781 45766 815
rect 42294 540 42328 574
rect 46378 781 46412 815
rect 46616 795 46650 829
rect 46919 793 46953 827
rect 47037 806 47071 840
rect 48266 1109 48300 1143
rect 49508 1109 49542 1143
rect 47936 949 47970 983
rect 45952 621 45986 655
rect 47308 787 47342 821
rect 47620 781 47654 815
rect 44182 540 44216 574
rect 48266 781 48300 815
rect 48504 795 48538 829
rect 48807 793 48841 827
rect 48925 806 48959 840
rect 50154 1109 50188 1143
rect 51396 1109 51430 1143
rect 49824 949 49858 983
rect 47840 621 47874 655
rect 49196 787 49230 821
rect 49508 781 49542 815
rect 46064 540 46098 574
rect 50154 781 50188 815
rect 50392 795 50426 829
rect 50695 793 50729 827
rect 50813 806 50847 840
rect 52042 1109 52076 1143
rect 53284 1109 53318 1143
rect 51712 949 51746 983
rect 49728 621 49762 655
rect 51084 787 51118 821
rect 51396 781 51430 815
rect 47952 540 47986 574
rect 52042 781 52076 815
rect 52280 795 52314 829
rect 52583 793 52617 827
rect 52701 806 52735 840
rect 53930 1109 53964 1143
rect 55172 1109 55206 1143
rect 53600 949 53634 983
rect 51616 621 51650 655
rect 52972 787 53006 821
rect 53284 781 53318 815
rect 49840 540 49874 574
rect 53930 781 53964 815
rect 54168 795 54202 829
rect 54471 793 54505 827
rect 54589 806 54623 840
rect 55818 1109 55852 1143
rect 57060 1109 57094 1143
rect 55488 949 55522 983
rect 53504 621 53538 655
rect 54860 787 54894 821
rect 55172 781 55206 815
rect 51728 540 51762 574
rect 55818 781 55852 815
rect 56056 795 56090 829
rect 56359 793 56393 827
rect 56477 806 56511 840
rect 57706 1109 57740 1143
rect 58948 1109 58982 1143
rect 57376 949 57410 983
rect 55392 621 55426 655
rect 56748 787 56782 821
rect 57060 781 57094 815
rect 53616 540 53650 574
rect 57706 781 57740 815
rect 57944 795 57978 829
rect 58247 793 58281 827
rect 58365 806 58399 840
rect 59594 1109 59628 1143
rect 59264 949 59298 983
rect 57280 621 57314 655
rect 58636 787 58670 821
rect 58948 781 58982 815
rect 55504 540 55538 574
rect 59594 781 59628 815
rect 59832 795 59866 829
rect 60135 793 60169 827
rect 60253 806 60287 840
rect 59168 621 59202 655
rect 57392 540 57426 574
rect 59280 540 59314 574
rect 668 300 702 334
rect 2556 300 2590 334
rect 4444 300 4478 334
rect 6332 300 6366 334
rect 8220 300 8254 334
rect 10108 300 10142 334
rect 11996 300 12030 334
rect 13884 300 13918 334
rect 15766 300 15800 334
rect 17654 300 17688 334
rect 19542 300 19576 334
rect 21430 300 21464 334
rect 23318 300 23352 334
rect 25206 300 25240 334
rect 27094 300 27128 334
rect 28982 300 29016 334
rect 30870 300 30904 334
rect 32758 300 32792 334
rect 34646 300 34680 334
rect 36534 300 36568 334
rect 38422 300 38456 334
rect 40310 300 40344 334
rect 42198 300 42232 334
rect 44086 300 44120 334
rect 45968 300 46002 334
rect 47856 300 47890 334
rect 49744 300 49778 334
rect 51632 300 51666 334
rect 53520 300 53554 334
rect 55408 300 55442 334
rect 57296 300 57330 334
rect 59184 300 59218 334
<< locali >>
rect 624 7249 894 7268
rect 624 7244 844 7249
rect 624 7210 723 7244
rect 757 7215 844 7244
rect 878 7215 894 7249
rect 757 7210 894 7215
rect 624 7190 894 7210
rect 2512 7249 2782 7268
rect 2512 7244 2732 7249
rect 2512 7210 2611 7244
rect 2645 7215 2732 7244
rect 2766 7215 2782 7249
rect 2645 7210 2782 7215
rect 2512 7190 2782 7210
rect 4400 7249 4670 7268
rect 4400 7244 4620 7249
rect 4400 7210 4499 7244
rect 4533 7215 4620 7244
rect 4654 7215 4670 7249
rect 4533 7210 4670 7215
rect 4400 7190 4670 7210
rect 6288 7249 6558 7268
rect 6288 7244 6508 7249
rect 6288 7210 6387 7244
rect 6421 7215 6508 7244
rect 6542 7215 6558 7249
rect 6421 7210 6558 7215
rect 6288 7190 6558 7210
rect 8176 7249 8446 7268
rect 8176 7244 8396 7249
rect 8176 7210 8275 7244
rect 8309 7215 8396 7244
rect 8430 7215 8446 7249
rect 8309 7210 8446 7215
rect 8176 7190 8446 7210
rect 10064 7249 10334 7268
rect 10064 7244 10284 7249
rect 10064 7210 10163 7244
rect 10197 7215 10284 7244
rect 10318 7215 10334 7249
rect 10197 7210 10334 7215
rect 10064 7190 10334 7210
rect 11952 7249 12222 7268
rect 11952 7244 12172 7249
rect 11952 7210 12051 7244
rect 12085 7215 12172 7244
rect 12206 7215 12222 7249
rect 12085 7210 12222 7215
rect 11952 7190 12222 7210
rect 13840 7249 14110 7268
rect 13840 7244 14060 7249
rect 13840 7210 13939 7244
rect 13973 7215 14060 7244
rect 14094 7215 14110 7249
rect 13973 7210 14110 7215
rect 13840 7190 14110 7210
rect 15722 7249 15992 7268
rect 15722 7244 15942 7249
rect 15722 7210 15821 7244
rect 15855 7215 15942 7244
rect 15976 7215 15992 7249
rect 15855 7210 15992 7215
rect 15722 7190 15992 7210
rect 17610 7249 17880 7268
rect 17610 7244 17830 7249
rect 17610 7210 17709 7244
rect 17743 7215 17830 7244
rect 17864 7215 17880 7249
rect 17743 7210 17880 7215
rect 17610 7190 17880 7210
rect 19498 7249 19768 7268
rect 19498 7244 19718 7249
rect 19498 7210 19597 7244
rect 19631 7215 19718 7244
rect 19752 7215 19768 7249
rect 19631 7210 19768 7215
rect 19498 7190 19768 7210
rect 21386 7249 21656 7268
rect 21386 7244 21606 7249
rect 21386 7210 21485 7244
rect 21519 7215 21606 7244
rect 21640 7215 21656 7249
rect 21519 7210 21656 7215
rect 21386 7190 21656 7210
rect 23274 7249 23544 7268
rect 23274 7244 23494 7249
rect 23274 7210 23373 7244
rect 23407 7215 23494 7244
rect 23528 7215 23544 7249
rect 23407 7210 23544 7215
rect 23274 7190 23544 7210
rect 25162 7249 25432 7268
rect 25162 7244 25382 7249
rect 25162 7210 25261 7244
rect 25295 7215 25382 7244
rect 25416 7215 25432 7249
rect 25295 7210 25432 7215
rect 25162 7190 25432 7210
rect 27050 7249 27320 7268
rect 27050 7244 27270 7249
rect 27050 7210 27149 7244
rect 27183 7215 27270 7244
rect 27304 7215 27320 7249
rect 27183 7210 27320 7215
rect 27050 7190 27320 7210
rect 28938 7249 29208 7268
rect 28938 7244 29158 7249
rect 28938 7210 29037 7244
rect 29071 7215 29158 7244
rect 29192 7215 29208 7249
rect 29071 7210 29208 7215
rect 28938 7190 29208 7210
rect 30826 7249 31096 7268
rect 30826 7244 31046 7249
rect 30826 7210 30925 7244
rect 30959 7215 31046 7244
rect 31080 7215 31096 7249
rect 30959 7210 31096 7215
rect 30826 7190 31096 7210
rect 32714 7249 32984 7268
rect 32714 7244 32934 7249
rect 32714 7210 32813 7244
rect 32847 7215 32934 7244
rect 32968 7215 32984 7249
rect 32847 7210 32984 7215
rect 32714 7190 32984 7210
rect 34602 7249 34872 7268
rect 34602 7244 34822 7249
rect 34602 7210 34701 7244
rect 34735 7215 34822 7244
rect 34856 7215 34872 7249
rect 34735 7210 34872 7215
rect 34602 7190 34872 7210
rect 36490 7249 36760 7268
rect 36490 7244 36710 7249
rect 36490 7210 36589 7244
rect 36623 7215 36710 7244
rect 36744 7215 36760 7249
rect 36623 7210 36760 7215
rect 36490 7190 36760 7210
rect 38378 7249 38648 7268
rect 38378 7244 38598 7249
rect 38378 7210 38477 7244
rect 38511 7215 38598 7244
rect 38632 7215 38648 7249
rect 38511 7210 38648 7215
rect 38378 7190 38648 7210
rect 40266 7249 40536 7268
rect 40266 7244 40486 7249
rect 40266 7210 40365 7244
rect 40399 7215 40486 7244
rect 40520 7215 40536 7249
rect 40399 7210 40536 7215
rect 40266 7190 40536 7210
rect 42154 7249 42424 7268
rect 42154 7244 42374 7249
rect 42154 7210 42253 7244
rect 42287 7215 42374 7244
rect 42408 7215 42424 7249
rect 42287 7210 42424 7215
rect 42154 7190 42424 7210
rect 44042 7249 44312 7268
rect 44042 7244 44262 7249
rect 44042 7210 44141 7244
rect 44175 7215 44262 7244
rect 44296 7215 44312 7249
rect 44175 7210 44312 7215
rect 44042 7190 44312 7210
rect 45924 7249 46194 7268
rect 45924 7244 46144 7249
rect 45924 7210 46023 7244
rect 46057 7215 46144 7244
rect 46178 7215 46194 7249
rect 46057 7210 46194 7215
rect 45924 7190 46194 7210
rect 47812 7249 48082 7268
rect 47812 7244 48032 7249
rect 47812 7210 47911 7244
rect 47945 7215 48032 7244
rect 48066 7215 48082 7249
rect 47945 7210 48082 7215
rect 47812 7190 48082 7210
rect 49700 7249 49970 7268
rect 49700 7244 49920 7249
rect 49700 7210 49799 7244
rect 49833 7215 49920 7244
rect 49954 7215 49970 7249
rect 49833 7210 49970 7215
rect 49700 7190 49970 7210
rect 51588 7249 51858 7268
rect 51588 7244 51808 7249
rect 51588 7210 51687 7244
rect 51721 7215 51808 7244
rect 51842 7215 51858 7249
rect 51721 7210 51858 7215
rect 51588 7190 51858 7210
rect 53476 7249 53746 7268
rect 53476 7244 53696 7249
rect 53476 7210 53575 7244
rect 53609 7215 53696 7244
rect 53730 7215 53746 7249
rect 53609 7210 53746 7215
rect 53476 7190 53746 7210
rect 55364 7249 55634 7268
rect 55364 7244 55584 7249
rect 55364 7210 55463 7244
rect 55497 7215 55584 7244
rect 55618 7215 55634 7249
rect 55497 7210 55634 7215
rect 55364 7190 55634 7210
rect 57252 7249 57522 7268
rect 57252 7244 57472 7249
rect 57252 7210 57351 7244
rect 57385 7215 57472 7244
rect 57506 7215 57522 7249
rect 57385 7210 57522 7215
rect 57252 7190 57522 7210
rect 59140 7249 59410 7268
rect 59140 7244 59360 7249
rect 59140 7210 59239 7244
rect 59273 7215 59360 7244
rect 59394 7215 59410 7249
rect 59273 7210 59410 7215
rect 59140 7190 59410 7210
rect 748 7106 764 7140
rect 798 7106 814 7140
rect 2636 7106 2652 7140
rect 2686 7106 2702 7140
rect 4524 7106 4540 7140
rect 4574 7106 4590 7140
rect 6412 7106 6428 7140
rect 6462 7106 6478 7140
rect 8300 7106 8316 7140
rect 8350 7106 8366 7140
rect 10188 7106 10204 7140
rect 10238 7106 10254 7140
rect 12076 7106 12092 7140
rect 12126 7106 12142 7140
rect 13964 7106 13980 7140
rect 14014 7106 14030 7140
rect 15846 7106 15862 7140
rect 15896 7106 15912 7140
rect 17734 7106 17750 7140
rect 17784 7106 17800 7140
rect 19622 7106 19638 7140
rect 19672 7106 19688 7140
rect 21510 7106 21526 7140
rect 21560 7106 21576 7140
rect 23398 7106 23414 7140
rect 23448 7106 23464 7140
rect 25286 7106 25302 7140
rect 25336 7106 25352 7140
rect 27174 7106 27190 7140
rect 27224 7106 27240 7140
rect 29062 7106 29078 7140
rect 29112 7106 29128 7140
rect 30950 7106 30966 7140
rect 31000 7106 31016 7140
rect 32838 7106 32854 7140
rect 32888 7106 32904 7140
rect 34726 7106 34742 7140
rect 34776 7106 34792 7140
rect 36614 7106 36630 7140
rect 36664 7106 36680 7140
rect 38502 7106 38518 7140
rect 38552 7106 38568 7140
rect 40390 7106 40406 7140
rect 40440 7106 40456 7140
rect 42278 7106 42294 7140
rect 42328 7106 42344 7140
rect 44166 7106 44182 7140
rect 44216 7106 44232 7140
rect 46048 7106 46064 7140
rect 46098 7106 46114 7140
rect 47936 7106 47952 7140
rect 47986 7106 48002 7140
rect 49824 7106 49840 7140
rect 49874 7106 49890 7140
rect 51712 7106 51728 7140
rect 51762 7106 51778 7140
rect 53600 7106 53616 7140
rect 53650 7106 53666 7140
rect 55488 7106 55504 7140
rect 55538 7106 55554 7140
rect 57376 7106 57392 7140
rect 57426 7106 57442 7140
rect 59264 7106 59280 7140
rect 59314 7106 59330 7140
rect 620 7056 654 7072
rect 620 6986 654 7020
rect 620 6934 654 6950
rect 716 7056 750 7072
rect 812 7058 846 7072
rect 930 7058 1150 7080
rect 810 7056 1150 7058
rect 810 7022 812 7056
rect 846 7044 1150 7056
rect 846 7022 966 7044
rect 716 6986 750 7020
rect 811 7020 812 7022
rect 811 6986 846 7020
rect 1114 6996 1150 7044
rect 811 6985 812 6986
rect 716 6934 750 6950
rect 812 6934 846 6950
rect 1018 6960 1150 6996
rect 2508 7056 2542 7072
rect 2508 6986 2542 7020
rect -392 6845 -363 6879
rect -329 6845 -271 6879
rect -237 6845 -179 6879
rect -145 6845 -116 6879
rect -375 6773 -323 6811
rect -375 6739 -357 6773
rect -287 6803 -221 6845
rect -46 6843 -17 6877
rect 17 6843 75 6877
rect 109 6843 167 6877
rect 201 6843 230 6877
rect 390 6862 438 6874
rect 652 6866 668 6900
rect 702 6866 718 6900
rect 1018 6890 1068 6960
rect 2508 6934 2542 6950
rect 2604 7056 2638 7072
rect 2700 7058 2734 7072
rect 2818 7058 3038 7080
rect 2698 7056 3038 7058
rect 2698 7022 2700 7056
rect 2734 7044 3038 7056
rect 2734 7022 2854 7044
rect 2604 6986 2638 7020
rect 2699 7020 2700 7022
rect 2699 6986 2734 7020
rect 3002 6996 3038 7044
rect 2699 6985 2700 6986
rect 2604 6934 2638 6950
rect 2700 6934 2734 6950
rect 2906 6960 3038 6996
rect 4396 7056 4430 7072
rect 4396 6986 4430 7020
rect 1018 6876 1028 6890
rect -287 6769 -271 6803
rect -237 6769 -221 6803
rect -185 6790 -151 6811
rect -375 6710 -323 6739
rect -185 6735 -151 6756
rect -375 6638 -339 6710
rect -284 6701 -151 6735
rect 20 6797 86 6809
rect 20 6763 36 6797
rect 70 6763 86 6797
rect 20 6746 86 6763
rect -284 6650 -250 6701
rect 20 6695 36 6746
rect 70 6695 86 6746
rect 20 6683 86 6695
rect 120 6797 166 6843
rect 154 6763 166 6797
rect 120 6729 166 6763
rect 154 6695 166 6729
rect 390 6828 396 6862
rect 430 6828 438 6862
rect 1022 6856 1028 6876
rect 1062 6856 1068 6890
rect 1022 6846 1068 6856
rect 1150 6851 1179 6885
rect 1213 6851 1271 6885
rect 1305 6851 1363 6885
rect 1397 6851 1426 6885
rect 390 6740 438 6828
rect 764 6785 780 6819
rect 814 6818 830 6819
rect 814 6786 976 6818
rect 1216 6810 1282 6817
rect 1210 6805 1282 6810
rect 1210 6786 1232 6805
rect 814 6785 1232 6786
rect 764 6782 1232 6785
rect 940 6771 1232 6782
rect 1266 6771 1282 6805
rect 940 6750 1282 6771
rect 636 6740 670 6742
rect 390 6723 670 6740
rect 390 6706 636 6723
rect -380 6636 -339 6638
rect -380 6602 -378 6636
rect -344 6602 -339 6636
rect -380 6600 -339 6602
rect -375 6550 -339 6600
rect -305 6634 -250 6650
rect -271 6600 -250 6634
rect -305 6584 -250 6600
rect -205 6648 -137 6665
rect -205 6647 -185 6648
rect -205 6613 -187 6647
rect -151 6614 -137 6648
rect -153 6613 -137 6614
rect -205 6591 -137 6613
rect -284 6555 -250 6584
rect 20 6563 66 6683
rect 120 6679 166 6695
rect 338 6658 354 6659
rect 100 6611 116 6645
rect 150 6638 166 6645
rect 218 6638 354 6658
rect 150 6625 354 6638
rect 388 6625 404 6659
rect 150 6624 404 6625
rect 150 6611 258 6624
rect 338 6622 404 6624
rect 636 6655 670 6657
rect 100 6597 258 6611
rect 114 6596 258 6597
rect 636 6619 670 6621
rect 310 6563 344 6582
rect -375 6500 -321 6550
rect -284 6521 -149 6555
rect -375 6466 -357 6500
rect -323 6466 -321 6500
rect -185 6487 -149 6521
rect -375 6419 -321 6466
rect -375 6385 -357 6419
rect -323 6385 -321 6419
rect -375 6369 -321 6385
rect -287 6453 -271 6487
rect -237 6453 -221 6487
rect -287 6419 -221 6453
rect -287 6385 -271 6419
rect -237 6385 -221 6419
rect -287 6335 -221 6385
rect -151 6453 -149 6487
rect -185 6419 -149 6453
rect -151 6385 -149 6419
rect -185 6369 -149 6385
rect 20 6545 86 6563
rect 20 6511 36 6545
rect 70 6511 86 6545
rect 20 6477 86 6511
rect 20 6443 36 6477
rect 70 6443 86 6477
rect 20 6409 86 6443
rect 20 6375 36 6409
rect 70 6375 86 6409
rect 20 6367 86 6375
rect 120 6545 162 6561
rect 154 6511 162 6545
rect 120 6477 162 6511
rect 154 6443 162 6477
rect 120 6409 162 6443
rect 310 6495 344 6497
rect 310 6459 344 6461
rect 154 6375 162 6409
rect -392 6301 -363 6335
rect -329 6301 -271 6335
rect -237 6301 -179 6335
rect -145 6301 -116 6335
rect 120 6333 162 6375
rect 270 6393 310 6414
rect 398 6563 432 6582
rect 636 6534 670 6553
rect 732 6723 766 6742
rect 732 6655 766 6657
rect 732 6619 766 6621
rect 732 6534 766 6553
rect 828 6723 862 6742
rect 1216 6737 1282 6750
rect 1216 6703 1232 6737
rect 1266 6703 1282 6737
rect 1216 6691 1282 6703
rect 1316 6805 1362 6851
rect 1496 6845 1525 6879
rect 1559 6845 1617 6879
rect 1651 6845 1709 6879
rect 1743 6845 1772 6879
rect 1350 6771 1362 6805
rect 1316 6737 1362 6771
rect 1350 6703 1362 6737
rect 828 6655 862 6657
rect 984 6625 1000 6659
rect 1034 6625 1050 6659
rect 828 6619 862 6621
rect 828 6534 862 6553
rect 956 6563 990 6582
rect 398 6495 432 6497
rect 956 6495 990 6497
rect 398 6459 432 6461
rect 668 6457 684 6491
rect 718 6457 734 6491
rect 956 6459 990 6461
rect 344 6393 346 6414
rect 270 6374 346 6393
rect 432 6393 956 6418
rect 1044 6563 1078 6582
rect 1044 6495 1078 6497
rect 1044 6459 1078 6461
rect 990 6393 992 6418
rect 398 6385 992 6393
rect 398 6374 634 6385
rect -46 6299 -17 6333
rect 17 6299 75 6333
rect 109 6299 167 6333
rect 201 6299 230 6333
rect 270 6016 304 6374
rect 544 6351 634 6374
rect 668 6383 992 6385
rect 668 6351 753 6383
rect 544 6349 753 6351
rect 787 6374 992 6383
rect 1044 6374 1078 6393
rect 1216 6571 1262 6691
rect 1316 6687 1362 6703
rect 1513 6773 1565 6811
rect 1513 6739 1531 6773
rect 1601 6803 1667 6845
rect 1842 6843 1871 6877
rect 1905 6843 1963 6877
rect 1997 6843 2055 6877
rect 2089 6843 2118 6877
rect 2278 6862 2326 6874
rect 2540 6866 2556 6900
rect 2590 6866 2606 6900
rect 2906 6890 2956 6960
rect 4396 6934 4430 6950
rect 4492 7056 4526 7072
rect 4588 7058 4622 7072
rect 4706 7058 4926 7080
rect 4586 7056 4926 7058
rect 4586 7022 4588 7056
rect 4622 7044 4926 7056
rect 4622 7022 4742 7044
rect 4492 6986 4526 7020
rect 4587 7020 4588 7022
rect 4587 6986 4622 7020
rect 4890 6996 4926 7044
rect 4587 6985 4588 6986
rect 4492 6934 4526 6950
rect 4588 6934 4622 6950
rect 4794 6960 4926 6996
rect 6284 7056 6318 7072
rect 6284 6986 6318 7020
rect 2906 6876 2916 6890
rect 1601 6769 1617 6803
rect 1651 6769 1667 6803
rect 1703 6790 1737 6811
rect 1513 6710 1565 6739
rect 1703 6735 1737 6756
rect 1296 6619 1312 6653
rect 1346 6642 1362 6653
rect 1296 6608 1314 6619
rect 1348 6608 1362 6642
rect 1513 6638 1549 6710
rect 1604 6701 1737 6735
rect 1908 6797 1974 6809
rect 1908 6763 1924 6797
rect 1958 6763 1974 6797
rect 1908 6746 1974 6763
rect 1604 6650 1638 6701
rect 1908 6695 1924 6746
rect 1958 6695 1974 6746
rect 1908 6683 1974 6695
rect 2008 6797 2054 6843
rect 2042 6763 2054 6797
rect 2008 6729 2054 6763
rect 2042 6695 2054 6729
rect 2278 6828 2284 6862
rect 2318 6828 2326 6862
rect 2910 6856 2916 6876
rect 2950 6856 2956 6890
rect 2910 6846 2956 6856
rect 3038 6851 3067 6885
rect 3101 6851 3159 6885
rect 3193 6851 3251 6885
rect 3285 6851 3314 6885
rect 2278 6740 2326 6828
rect 2652 6785 2668 6819
rect 2702 6818 2718 6819
rect 2702 6786 2864 6818
rect 3104 6810 3170 6817
rect 3098 6805 3170 6810
rect 3098 6786 3120 6805
rect 2702 6785 3120 6786
rect 2652 6782 3120 6785
rect 2828 6771 3120 6782
rect 3154 6771 3170 6805
rect 2828 6750 3170 6771
rect 2524 6740 2558 6742
rect 2278 6723 2558 6740
rect 2278 6706 2524 6723
rect 1296 6605 1362 6608
rect 1508 6636 1549 6638
rect 1508 6602 1510 6636
rect 1544 6602 1549 6636
rect 1508 6600 1549 6602
rect 1216 6553 1282 6571
rect 1216 6519 1232 6553
rect 1266 6519 1282 6553
rect 1216 6485 1282 6519
rect 1216 6451 1232 6485
rect 1266 6451 1282 6485
rect 1216 6417 1282 6451
rect 1216 6383 1232 6417
rect 1266 6383 1282 6417
rect 1216 6375 1282 6383
rect 1316 6553 1358 6569
rect 1350 6519 1358 6553
rect 1316 6485 1358 6519
rect 1350 6451 1358 6485
rect 1316 6417 1358 6451
rect 1350 6383 1358 6417
rect 787 6349 826 6374
rect 338 6297 354 6331
rect 388 6297 404 6331
rect 544 6310 826 6349
rect 1316 6341 1358 6383
rect 1513 6550 1549 6600
rect 1583 6634 1638 6650
rect 1617 6600 1638 6634
rect 1583 6584 1638 6600
rect 1683 6648 1751 6665
rect 1683 6647 1703 6648
rect 1683 6613 1701 6647
rect 1737 6614 1751 6648
rect 1735 6613 1751 6614
rect 1683 6591 1751 6613
rect 1604 6555 1638 6584
rect 1908 6563 1954 6683
rect 2008 6679 2054 6695
rect 2226 6658 2242 6659
rect 1988 6611 2004 6645
rect 2038 6638 2054 6645
rect 2106 6638 2242 6658
rect 2038 6625 2242 6638
rect 2276 6625 2292 6659
rect 2038 6624 2292 6625
rect 2038 6611 2146 6624
rect 2226 6622 2292 6624
rect 2524 6655 2558 6657
rect 1988 6597 2146 6611
rect 2002 6596 2146 6597
rect 2524 6619 2558 6621
rect 2198 6563 2232 6582
rect 1513 6500 1567 6550
rect 1604 6521 1739 6555
rect 1513 6466 1531 6500
rect 1565 6466 1567 6500
rect 1703 6487 1739 6521
rect 1513 6419 1567 6466
rect 1513 6385 1531 6419
rect 1565 6385 1567 6419
rect 1513 6369 1567 6385
rect 1601 6453 1617 6487
rect 1651 6453 1667 6487
rect 1601 6419 1667 6453
rect 1601 6385 1617 6419
rect 1651 6385 1667 6419
rect 712 6308 826 6310
rect 984 6297 1000 6331
rect 1034 6297 1050 6331
rect 1150 6307 1179 6341
rect 1213 6307 1271 6341
rect 1305 6307 1363 6341
rect 1397 6307 1426 6341
rect 1601 6335 1667 6385
rect 1737 6453 1739 6487
rect 1703 6419 1739 6453
rect 1737 6385 1739 6419
rect 1703 6369 1739 6385
rect 1908 6545 1974 6563
rect 1908 6511 1924 6545
rect 1958 6511 1974 6545
rect 1908 6477 1974 6511
rect 1908 6443 1924 6477
rect 1958 6443 1974 6477
rect 1908 6409 1974 6443
rect 1908 6375 1924 6409
rect 1958 6375 1974 6409
rect 1908 6367 1974 6375
rect 2008 6545 2050 6561
rect 2042 6511 2050 6545
rect 2008 6477 2050 6511
rect 2042 6443 2050 6477
rect 2008 6409 2050 6443
rect 2198 6495 2232 6497
rect 2198 6459 2232 6461
rect 2042 6375 2050 6409
rect 1317 6300 1351 6307
rect 1496 6301 1525 6335
rect 1559 6301 1617 6335
rect 1651 6301 1709 6335
rect 1743 6301 1772 6335
rect 2008 6333 2050 6375
rect 2158 6393 2198 6414
rect 2286 6563 2320 6582
rect 2524 6534 2558 6553
rect 2620 6723 2654 6742
rect 2620 6655 2654 6657
rect 2620 6619 2654 6621
rect 2620 6534 2654 6553
rect 2716 6723 2750 6742
rect 3104 6737 3170 6750
rect 3104 6703 3120 6737
rect 3154 6703 3170 6737
rect 3104 6691 3170 6703
rect 3204 6805 3250 6851
rect 3384 6845 3413 6879
rect 3447 6845 3505 6879
rect 3539 6845 3597 6879
rect 3631 6845 3660 6879
rect 3238 6771 3250 6805
rect 3204 6737 3250 6771
rect 3238 6703 3250 6737
rect 2716 6655 2750 6657
rect 2872 6625 2888 6659
rect 2922 6625 2938 6659
rect 2716 6619 2750 6621
rect 2716 6534 2750 6553
rect 2844 6563 2878 6582
rect 2286 6495 2320 6497
rect 2844 6495 2878 6497
rect 2286 6459 2320 6461
rect 2556 6457 2572 6491
rect 2606 6457 2622 6491
rect 2844 6459 2878 6461
rect 2232 6393 2234 6414
rect 2158 6374 2234 6393
rect 2320 6393 2844 6418
rect 2932 6563 2966 6582
rect 2932 6495 2966 6497
rect 2932 6459 2966 6461
rect 2878 6393 2880 6418
rect 2286 6385 2880 6393
rect 2286 6374 2522 6385
rect 1842 6299 1871 6333
rect 1905 6299 1963 6333
rect 1997 6299 2055 6333
rect 2089 6299 2118 6333
rect 404 6212 450 6218
rect 404 6210 892 6212
rect 404 6176 412 6210
rect 446 6193 892 6210
rect 446 6188 842 6193
rect 446 6178 721 6188
rect 446 6176 450 6178
rect 404 6174 450 6176
rect 622 6154 721 6178
rect 755 6159 842 6188
rect 876 6168 892 6193
rect 876 6159 1017 6168
rect 755 6154 1017 6159
rect 622 6134 1017 6154
rect 746 6050 762 6084
rect 796 6050 932 6084
rect 270 6000 652 6016
rect 270 5976 618 6000
rect 618 5930 652 5964
rect 618 5878 652 5894
rect 714 6000 748 6016
rect 714 5930 748 5964
rect 714 5878 748 5894
rect 810 6000 844 6016
rect 810 5930 844 5964
rect 810 5878 844 5894
rect 158 5797 187 5831
rect 221 5797 279 5831
rect 313 5797 371 5831
rect 405 5797 434 5831
rect 650 5810 666 5844
rect 700 5810 716 5844
rect 177 5753 231 5797
rect 177 5719 197 5753
rect 177 5685 231 5719
rect 177 5651 197 5685
rect 177 5635 231 5651
rect 265 5753 331 5763
rect 265 5719 281 5753
rect 315 5719 331 5753
rect 265 5715 331 5719
rect 265 5681 279 5715
rect 313 5685 331 5715
rect 265 5651 281 5681
rect 315 5651 331 5685
rect 265 5635 331 5651
rect 365 5753 413 5797
rect 399 5719 413 5753
rect 762 5729 778 5763
rect 812 5729 828 5763
rect 365 5685 413 5719
rect 399 5651 413 5685
rect 365 5635 413 5651
rect 634 5667 668 5686
rect 175 5592 195 5599
rect 175 5558 193 5592
rect 229 5565 245 5599
rect 227 5558 245 5565
rect 175 5549 245 5558
rect 279 5515 313 5635
rect 634 5599 668 5601
rect 347 5565 363 5599
rect 397 5592 417 5599
rect 347 5558 367 5565
rect 401 5558 417 5592
rect 347 5549 417 5558
rect 634 5563 668 5565
rect 177 5499 243 5515
rect 177 5465 209 5499
rect 279 5499 415 5515
rect 279 5481 365 5499
rect 177 5431 243 5465
rect 177 5397 209 5431
rect 177 5363 243 5397
rect 177 5329 209 5363
rect 177 5287 243 5329
rect 349 5465 365 5481
rect 399 5465 415 5499
rect 634 5478 668 5497
rect 730 5667 764 5686
rect 730 5599 764 5601
rect 730 5563 764 5565
rect 730 5478 764 5497
rect 826 5667 860 5686
rect 826 5599 860 5601
rect 826 5563 860 5565
rect 826 5478 860 5497
rect 349 5431 415 5465
rect 349 5397 365 5431
rect 399 5397 415 5431
rect 666 5436 732 5438
rect 898 5436 932 6050
rect 983 5831 1017 6134
rect 1214 5831 1248 6042
rect 2158 6016 2192 6374
rect 2432 6351 2522 6374
rect 2556 6383 2880 6385
rect 2556 6351 2641 6383
rect 2432 6349 2641 6351
rect 2675 6374 2880 6383
rect 2932 6374 2966 6393
rect 3104 6571 3150 6691
rect 3204 6687 3250 6703
rect 3401 6773 3453 6811
rect 3401 6739 3419 6773
rect 3489 6803 3555 6845
rect 3730 6843 3759 6877
rect 3793 6843 3851 6877
rect 3885 6843 3943 6877
rect 3977 6843 4006 6877
rect 4166 6862 4214 6874
rect 4428 6866 4444 6900
rect 4478 6866 4494 6900
rect 4794 6890 4844 6960
rect 6284 6934 6318 6950
rect 6380 7056 6414 7072
rect 6476 7058 6510 7072
rect 6594 7058 6814 7080
rect 6474 7056 6814 7058
rect 6474 7022 6476 7056
rect 6510 7044 6814 7056
rect 6510 7022 6630 7044
rect 6380 6986 6414 7020
rect 6475 7020 6476 7022
rect 6475 6986 6510 7020
rect 6778 6996 6814 7044
rect 6475 6985 6476 6986
rect 6380 6934 6414 6950
rect 6476 6934 6510 6950
rect 6682 6960 6814 6996
rect 8172 7056 8206 7072
rect 8172 6986 8206 7020
rect 4794 6876 4804 6890
rect 3489 6769 3505 6803
rect 3539 6769 3555 6803
rect 3591 6790 3625 6811
rect 3401 6710 3453 6739
rect 3591 6735 3625 6756
rect 3184 6619 3200 6653
rect 3234 6642 3250 6653
rect 3184 6608 3202 6619
rect 3236 6608 3250 6642
rect 3401 6638 3437 6710
rect 3492 6701 3625 6735
rect 3796 6797 3862 6809
rect 3796 6763 3812 6797
rect 3846 6763 3862 6797
rect 3796 6746 3862 6763
rect 3492 6650 3526 6701
rect 3796 6695 3812 6746
rect 3846 6695 3862 6746
rect 3796 6683 3862 6695
rect 3896 6797 3942 6843
rect 3930 6763 3942 6797
rect 3896 6729 3942 6763
rect 3930 6695 3942 6729
rect 4166 6828 4172 6862
rect 4206 6828 4214 6862
rect 4798 6856 4804 6876
rect 4838 6856 4844 6890
rect 4798 6846 4844 6856
rect 4926 6851 4955 6885
rect 4989 6851 5047 6885
rect 5081 6851 5139 6885
rect 5173 6851 5202 6885
rect 4166 6740 4214 6828
rect 4540 6785 4556 6819
rect 4590 6818 4606 6819
rect 4590 6786 4752 6818
rect 4992 6810 5058 6817
rect 4986 6805 5058 6810
rect 4986 6786 5008 6805
rect 4590 6785 5008 6786
rect 4540 6782 5008 6785
rect 4716 6771 5008 6782
rect 5042 6771 5058 6805
rect 4716 6750 5058 6771
rect 4412 6740 4446 6742
rect 4166 6723 4446 6740
rect 4166 6706 4412 6723
rect 3184 6605 3250 6608
rect 3396 6636 3437 6638
rect 3396 6602 3398 6636
rect 3432 6602 3437 6636
rect 3396 6600 3437 6602
rect 3104 6553 3170 6571
rect 3104 6519 3120 6553
rect 3154 6519 3170 6553
rect 3104 6485 3170 6519
rect 3104 6451 3120 6485
rect 3154 6451 3170 6485
rect 3104 6417 3170 6451
rect 3104 6383 3120 6417
rect 3154 6383 3170 6417
rect 3104 6375 3170 6383
rect 3204 6553 3246 6569
rect 3238 6519 3246 6553
rect 3204 6485 3246 6519
rect 3238 6451 3246 6485
rect 3204 6417 3246 6451
rect 3238 6383 3246 6417
rect 2675 6349 2714 6374
rect 2226 6297 2242 6331
rect 2276 6297 2292 6331
rect 2432 6310 2714 6349
rect 3204 6341 3246 6383
rect 3401 6550 3437 6600
rect 3471 6634 3526 6650
rect 3505 6600 3526 6634
rect 3471 6584 3526 6600
rect 3571 6648 3639 6665
rect 3571 6647 3591 6648
rect 3571 6613 3589 6647
rect 3625 6614 3639 6648
rect 3623 6613 3639 6614
rect 3571 6591 3639 6613
rect 3492 6555 3526 6584
rect 3796 6563 3842 6683
rect 3896 6679 3942 6695
rect 4114 6658 4130 6659
rect 3876 6611 3892 6645
rect 3926 6638 3942 6645
rect 3994 6638 4130 6658
rect 3926 6625 4130 6638
rect 4164 6625 4180 6659
rect 3926 6624 4180 6625
rect 3926 6611 4034 6624
rect 4114 6622 4180 6624
rect 4412 6655 4446 6657
rect 3876 6597 4034 6611
rect 3890 6596 4034 6597
rect 4412 6619 4446 6621
rect 4086 6563 4120 6582
rect 3401 6500 3455 6550
rect 3492 6521 3627 6555
rect 3401 6466 3419 6500
rect 3453 6466 3455 6500
rect 3591 6487 3627 6521
rect 3401 6419 3455 6466
rect 3401 6385 3419 6419
rect 3453 6385 3455 6419
rect 3401 6369 3455 6385
rect 3489 6453 3505 6487
rect 3539 6453 3555 6487
rect 3489 6419 3555 6453
rect 3489 6385 3505 6419
rect 3539 6385 3555 6419
rect 2600 6308 2714 6310
rect 2872 6297 2888 6331
rect 2922 6297 2938 6331
rect 3038 6307 3067 6341
rect 3101 6307 3159 6341
rect 3193 6307 3251 6341
rect 3285 6307 3314 6341
rect 3489 6335 3555 6385
rect 3625 6453 3627 6487
rect 3591 6419 3627 6453
rect 3625 6385 3627 6419
rect 3591 6369 3627 6385
rect 3796 6545 3862 6563
rect 3796 6511 3812 6545
rect 3846 6511 3862 6545
rect 3796 6477 3862 6511
rect 3796 6443 3812 6477
rect 3846 6443 3862 6477
rect 3796 6409 3862 6443
rect 3796 6375 3812 6409
rect 3846 6375 3862 6409
rect 3796 6367 3862 6375
rect 3896 6545 3938 6561
rect 3930 6511 3938 6545
rect 3896 6477 3938 6511
rect 3930 6443 3938 6477
rect 3896 6409 3938 6443
rect 4086 6495 4120 6497
rect 4086 6459 4120 6461
rect 3930 6375 3938 6409
rect 3205 6300 3239 6307
rect 3384 6301 3413 6335
rect 3447 6301 3505 6335
rect 3539 6301 3597 6335
rect 3631 6301 3660 6335
rect 3896 6333 3938 6375
rect 4046 6393 4086 6414
rect 4174 6563 4208 6582
rect 4412 6534 4446 6553
rect 4508 6723 4542 6742
rect 4508 6655 4542 6657
rect 4508 6619 4542 6621
rect 4508 6534 4542 6553
rect 4604 6723 4638 6742
rect 4992 6737 5058 6750
rect 4992 6703 5008 6737
rect 5042 6703 5058 6737
rect 4992 6691 5058 6703
rect 5092 6805 5138 6851
rect 5272 6845 5301 6879
rect 5335 6845 5393 6879
rect 5427 6845 5485 6879
rect 5519 6845 5548 6879
rect 5126 6771 5138 6805
rect 5092 6737 5138 6771
rect 5126 6703 5138 6737
rect 4604 6655 4638 6657
rect 4760 6625 4776 6659
rect 4810 6625 4826 6659
rect 4604 6619 4638 6621
rect 4604 6534 4638 6553
rect 4732 6563 4766 6582
rect 4174 6495 4208 6497
rect 4732 6495 4766 6497
rect 4174 6459 4208 6461
rect 4444 6457 4460 6491
rect 4494 6457 4510 6491
rect 4732 6459 4766 6461
rect 4120 6393 4122 6414
rect 4046 6374 4122 6393
rect 4208 6393 4732 6418
rect 4820 6563 4854 6582
rect 4820 6495 4854 6497
rect 4820 6459 4854 6461
rect 4766 6393 4768 6418
rect 4174 6385 4768 6393
rect 4174 6374 4410 6385
rect 3730 6299 3759 6333
rect 3793 6299 3851 6333
rect 3885 6299 3943 6333
rect 3977 6299 4006 6333
rect 2292 6212 2338 6218
rect 2292 6210 2780 6212
rect 2292 6176 2300 6210
rect 2334 6193 2780 6210
rect 2334 6188 2730 6193
rect 2334 6178 2609 6188
rect 2334 6176 2338 6178
rect 2292 6174 2338 6176
rect 2510 6154 2609 6178
rect 2643 6159 2730 6188
rect 2764 6168 2780 6193
rect 2764 6159 2905 6168
rect 2643 6154 2905 6159
rect 2510 6134 2905 6154
rect 2634 6050 2650 6084
rect 2684 6050 2820 6084
rect 2158 6000 2540 6016
rect 2158 5976 2506 6000
rect 2506 5930 2540 5964
rect 2506 5878 2540 5894
rect 2602 6000 2636 6016
rect 2602 5930 2636 5964
rect 2602 5878 2636 5894
rect 2698 6000 2732 6016
rect 2698 5930 2732 5964
rect 2698 5878 2732 5894
rect 972 5797 1001 5831
rect 1035 5797 1093 5831
rect 1127 5797 1185 5831
rect 1219 5797 1248 5831
rect 2046 5797 2075 5831
rect 2109 5797 2167 5831
rect 2201 5797 2259 5831
rect 2293 5797 2322 5831
rect 2538 5810 2554 5844
rect 2588 5810 2604 5844
rect 991 5753 1045 5797
rect 991 5719 1011 5753
rect 991 5685 1045 5719
rect 991 5651 1011 5685
rect 991 5635 1045 5651
rect 1079 5753 1145 5763
rect 1079 5719 1095 5753
rect 1129 5719 1145 5753
rect 1079 5710 1145 5719
rect 1079 5685 1097 5710
rect 1079 5651 1095 5685
rect 1131 5676 1145 5710
rect 1129 5651 1145 5676
rect 1079 5635 1145 5651
rect 1179 5753 1227 5797
rect 1213 5719 1227 5753
rect 1179 5685 1227 5719
rect 1213 5651 1227 5685
rect 1179 5635 1227 5651
rect 2065 5753 2119 5797
rect 2065 5719 2085 5753
rect 2065 5685 2119 5719
rect 2065 5651 2085 5685
rect 2065 5635 2119 5651
rect 2153 5753 2219 5763
rect 2153 5719 2169 5753
rect 2203 5719 2219 5753
rect 2153 5715 2219 5719
rect 2153 5681 2167 5715
rect 2201 5685 2219 5715
rect 2153 5651 2169 5681
rect 2203 5651 2219 5685
rect 2153 5635 2219 5651
rect 2253 5753 2301 5797
rect 2287 5719 2301 5753
rect 2650 5729 2666 5763
rect 2700 5729 2716 5763
rect 2253 5685 2301 5719
rect 2287 5651 2301 5685
rect 2253 5635 2301 5651
rect 2522 5667 2556 5686
rect 989 5594 1009 5599
rect 989 5560 1006 5594
rect 1043 5565 1059 5599
rect 1040 5560 1059 5565
rect 989 5549 1059 5560
rect 1093 5515 1127 5635
rect 1161 5565 1177 5599
rect 1211 5590 1231 5599
rect 1161 5556 1179 5565
rect 1213 5556 1231 5590
rect 1161 5549 1231 5556
rect 2063 5592 2083 5599
rect 2063 5558 2081 5592
rect 2117 5565 2133 5599
rect 2115 5558 2133 5565
rect 2063 5549 2133 5558
rect 2167 5515 2201 5635
rect 2522 5599 2556 5601
rect 2235 5565 2251 5599
rect 2285 5592 2305 5599
rect 2235 5558 2255 5565
rect 2289 5558 2305 5592
rect 2235 5549 2305 5558
rect 2522 5563 2556 5565
rect 666 5435 932 5436
rect 666 5401 682 5435
rect 716 5401 932 5435
rect 666 5400 932 5401
rect 991 5499 1057 5515
rect 991 5465 1023 5499
rect 1093 5499 1229 5515
rect 1093 5481 1179 5499
rect 991 5431 1057 5465
rect 349 5363 415 5397
rect 349 5329 365 5363
rect 399 5329 415 5363
rect 991 5397 1023 5431
rect 991 5363 1057 5397
rect 349 5324 415 5329
rect 542 5329 824 5362
rect 542 5295 632 5329
rect 666 5327 824 5329
rect 666 5295 751 5327
rect 542 5293 751 5295
rect 785 5293 824 5327
rect 542 5287 824 5293
rect 991 5329 1023 5363
rect 991 5287 1057 5329
rect 1163 5465 1179 5481
rect 1213 5465 1229 5499
rect 1163 5431 1229 5465
rect 1163 5397 1179 5431
rect 1213 5397 1229 5431
rect 1163 5363 1229 5397
rect 1163 5329 1179 5363
rect 1213 5329 1229 5363
rect 1163 5324 1229 5329
rect 2065 5499 2131 5515
rect 2065 5465 2097 5499
rect 2167 5499 2303 5515
rect 2167 5481 2253 5499
rect 2065 5431 2131 5465
rect 2065 5397 2097 5431
rect 2065 5363 2131 5397
rect 2065 5329 2097 5363
rect 2065 5287 2131 5329
rect 2237 5465 2253 5481
rect 2287 5465 2303 5499
rect 2522 5478 2556 5497
rect 2618 5667 2652 5686
rect 2618 5599 2652 5601
rect 2618 5563 2652 5565
rect 2618 5478 2652 5497
rect 2714 5667 2748 5686
rect 2714 5599 2748 5601
rect 2714 5563 2748 5565
rect 2714 5478 2748 5497
rect 2237 5431 2303 5465
rect 2237 5397 2253 5431
rect 2287 5397 2303 5431
rect 2554 5436 2620 5438
rect 2786 5436 2820 6050
rect 2871 5831 2905 6134
rect 3102 5831 3136 6042
rect 4046 6016 4080 6374
rect 4320 6351 4410 6374
rect 4444 6383 4768 6385
rect 4444 6351 4529 6383
rect 4320 6349 4529 6351
rect 4563 6374 4768 6383
rect 4820 6374 4854 6393
rect 4992 6571 5038 6691
rect 5092 6687 5138 6703
rect 5289 6773 5341 6811
rect 5289 6739 5307 6773
rect 5377 6803 5443 6845
rect 5618 6843 5647 6877
rect 5681 6843 5739 6877
rect 5773 6843 5831 6877
rect 5865 6843 5894 6877
rect 6054 6862 6102 6874
rect 6316 6866 6332 6900
rect 6366 6866 6382 6900
rect 6682 6890 6732 6960
rect 8172 6934 8206 6950
rect 8268 7056 8302 7072
rect 8364 7058 8398 7072
rect 8482 7058 8702 7080
rect 8362 7056 8702 7058
rect 8362 7022 8364 7056
rect 8398 7044 8702 7056
rect 8398 7022 8518 7044
rect 8268 6986 8302 7020
rect 8363 7020 8364 7022
rect 8363 6986 8398 7020
rect 8666 6996 8702 7044
rect 8363 6985 8364 6986
rect 8268 6934 8302 6950
rect 8364 6934 8398 6950
rect 8570 6960 8702 6996
rect 10060 7056 10094 7072
rect 10060 6986 10094 7020
rect 6682 6876 6692 6890
rect 5377 6769 5393 6803
rect 5427 6769 5443 6803
rect 5479 6790 5513 6811
rect 5289 6710 5341 6739
rect 5479 6735 5513 6756
rect 5072 6619 5088 6653
rect 5122 6642 5138 6653
rect 5072 6608 5090 6619
rect 5124 6608 5138 6642
rect 5289 6638 5325 6710
rect 5380 6701 5513 6735
rect 5684 6797 5750 6809
rect 5684 6763 5700 6797
rect 5734 6763 5750 6797
rect 5684 6746 5750 6763
rect 5380 6650 5414 6701
rect 5684 6695 5700 6746
rect 5734 6695 5750 6746
rect 5684 6683 5750 6695
rect 5784 6797 5830 6843
rect 5818 6763 5830 6797
rect 5784 6729 5830 6763
rect 5818 6695 5830 6729
rect 6054 6828 6060 6862
rect 6094 6828 6102 6862
rect 6686 6856 6692 6876
rect 6726 6856 6732 6890
rect 6686 6846 6732 6856
rect 6814 6851 6843 6885
rect 6877 6851 6935 6885
rect 6969 6851 7027 6885
rect 7061 6851 7090 6885
rect 6054 6740 6102 6828
rect 6428 6785 6444 6819
rect 6478 6818 6494 6819
rect 6478 6786 6640 6818
rect 6880 6810 6946 6817
rect 6874 6805 6946 6810
rect 6874 6786 6896 6805
rect 6478 6785 6896 6786
rect 6428 6782 6896 6785
rect 6604 6771 6896 6782
rect 6930 6771 6946 6805
rect 6604 6750 6946 6771
rect 6300 6740 6334 6742
rect 6054 6723 6334 6740
rect 6054 6706 6300 6723
rect 5072 6605 5138 6608
rect 5284 6636 5325 6638
rect 5284 6602 5286 6636
rect 5320 6602 5325 6636
rect 5284 6600 5325 6602
rect 4992 6553 5058 6571
rect 4992 6519 5008 6553
rect 5042 6519 5058 6553
rect 4992 6485 5058 6519
rect 4992 6451 5008 6485
rect 5042 6451 5058 6485
rect 4992 6417 5058 6451
rect 4992 6383 5008 6417
rect 5042 6383 5058 6417
rect 4992 6375 5058 6383
rect 5092 6553 5134 6569
rect 5126 6519 5134 6553
rect 5092 6485 5134 6519
rect 5126 6451 5134 6485
rect 5092 6417 5134 6451
rect 5126 6383 5134 6417
rect 4563 6349 4602 6374
rect 4114 6297 4130 6331
rect 4164 6297 4180 6331
rect 4320 6310 4602 6349
rect 5092 6341 5134 6383
rect 5289 6550 5325 6600
rect 5359 6634 5414 6650
rect 5393 6600 5414 6634
rect 5359 6584 5414 6600
rect 5459 6648 5527 6665
rect 5459 6647 5479 6648
rect 5459 6613 5477 6647
rect 5513 6614 5527 6648
rect 5511 6613 5527 6614
rect 5459 6591 5527 6613
rect 5380 6555 5414 6584
rect 5684 6563 5730 6683
rect 5784 6679 5830 6695
rect 6002 6658 6018 6659
rect 5764 6611 5780 6645
rect 5814 6638 5830 6645
rect 5882 6638 6018 6658
rect 5814 6625 6018 6638
rect 6052 6625 6068 6659
rect 5814 6624 6068 6625
rect 5814 6611 5922 6624
rect 6002 6622 6068 6624
rect 6300 6655 6334 6657
rect 5764 6597 5922 6611
rect 5778 6596 5922 6597
rect 6300 6619 6334 6621
rect 5974 6563 6008 6582
rect 5289 6500 5343 6550
rect 5380 6521 5515 6555
rect 5289 6466 5307 6500
rect 5341 6466 5343 6500
rect 5479 6487 5515 6521
rect 5289 6419 5343 6466
rect 5289 6385 5307 6419
rect 5341 6385 5343 6419
rect 5289 6369 5343 6385
rect 5377 6453 5393 6487
rect 5427 6453 5443 6487
rect 5377 6419 5443 6453
rect 5377 6385 5393 6419
rect 5427 6385 5443 6419
rect 4488 6308 4602 6310
rect 4760 6297 4776 6331
rect 4810 6297 4826 6331
rect 4926 6307 4955 6341
rect 4989 6307 5047 6341
rect 5081 6307 5139 6341
rect 5173 6307 5202 6341
rect 5377 6335 5443 6385
rect 5513 6453 5515 6487
rect 5479 6419 5515 6453
rect 5513 6385 5515 6419
rect 5479 6369 5515 6385
rect 5684 6545 5750 6563
rect 5684 6511 5700 6545
rect 5734 6511 5750 6545
rect 5684 6477 5750 6511
rect 5684 6443 5700 6477
rect 5734 6443 5750 6477
rect 5684 6409 5750 6443
rect 5684 6375 5700 6409
rect 5734 6375 5750 6409
rect 5684 6367 5750 6375
rect 5784 6545 5826 6561
rect 5818 6511 5826 6545
rect 5784 6477 5826 6511
rect 5818 6443 5826 6477
rect 5784 6409 5826 6443
rect 5974 6495 6008 6497
rect 5974 6459 6008 6461
rect 5818 6375 5826 6409
rect 5093 6300 5127 6307
rect 5272 6301 5301 6335
rect 5335 6301 5393 6335
rect 5427 6301 5485 6335
rect 5519 6301 5548 6335
rect 5784 6333 5826 6375
rect 5934 6393 5974 6414
rect 6062 6563 6096 6582
rect 6300 6534 6334 6553
rect 6396 6723 6430 6742
rect 6396 6655 6430 6657
rect 6396 6619 6430 6621
rect 6396 6534 6430 6553
rect 6492 6723 6526 6742
rect 6880 6737 6946 6750
rect 6880 6703 6896 6737
rect 6930 6703 6946 6737
rect 6880 6691 6946 6703
rect 6980 6805 7026 6851
rect 7160 6845 7189 6879
rect 7223 6845 7281 6879
rect 7315 6845 7373 6879
rect 7407 6845 7436 6879
rect 7014 6771 7026 6805
rect 6980 6737 7026 6771
rect 7014 6703 7026 6737
rect 6492 6655 6526 6657
rect 6648 6625 6664 6659
rect 6698 6625 6714 6659
rect 6492 6619 6526 6621
rect 6492 6534 6526 6553
rect 6620 6563 6654 6582
rect 6062 6495 6096 6497
rect 6620 6495 6654 6497
rect 6062 6459 6096 6461
rect 6332 6457 6348 6491
rect 6382 6457 6398 6491
rect 6620 6459 6654 6461
rect 6008 6393 6010 6414
rect 5934 6374 6010 6393
rect 6096 6393 6620 6418
rect 6708 6563 6742 6582
rect 6708 6495 6742 6497
rect 6708 6459 6742 6461
rect 6654 6393 6656 6418
rect 6062 6385 6656 6393
rect 6062 6374 6298 6385
rect 5618 6299 5647 6333
rect 5681 6299 5739 6333
rect 5773 6299 5831 6333
rect 5865 6299 5894 6333
rect 4180 6212 4226 6218
rect 4180 6210 4668 6212
rect 4180 6176 4188 6210
rect 4222 6193 4668 6210
rect 4222 6188 4618 6193
rect 4222 6178 4497 6188
rect 4222 6176 4226 6178
rect 4180 6174 4226 6176
rect 4398 6154 4497 6178
rect 4531 6159 4618 6188
rect 4652 6168 4668 6193
rect 4652 6159 4793 6168
rect 4531 6154 4793 6159
rect 4398 6134 4793 6154
rect 4522 6050 4538 6084
rect 4572 6050 4708 6084
rect 4046 6000 4428 6016
rect 4046 5976 4394 6000
rect 4394 5930 4428 5964
rect 4394 5878 4428 5894
rect 4490 6000 4524 6016
rect 4490 5930 4524 5964
rect 4490 5878 4524 5894
rect 4586 6000 4620 6016
rect 4586 5930 4620 5964
rect 4586 5878 4620 5894
rect 2860 5797 2889 5831
rect 2923 5797 2981 5831
rect 3015 5797 3073 5831
rect 3107 5797 3136 5831
rect 3934 5797 3963 5831
rect 3997 5797 4055 5831
rect 4089 5797 4147 5831
rect 4181 5797 4210 5831
rect 4426 5810 4442 5844
rect 4476 5810 4492 5844
rect 2879 5753 2933 5797
rect 2879 5719 2899 5753
rect 2879 5685 2933 5719
rect 2879 5651 2899 5685
rect 2879 5635 2933 5651
rect 2967 5753 3033 5763
rect 2967 5719 2983 5753
rect 3017 5719 3033 5753
rect 2967 5710 3033 5719
rect 2967 5685 2985 5710
rect 2967 5651 2983 5685
rect 3019 5676 3033 5710
rect 3017 5651 3033 5676
rect 2967 5635 3033 5651
rect 3067 5753 3115 5797
rect 3101 5719 3115 5753
rect 3067 5685 3115 5719
rect 3101 5651 3115 5685
rect 3067 5635 3115 5651
rect 3953 5753 4007 5797
rect 3953 5719 3973 5753
rect 3953 5685 4007 5719
rect 3953 5651 3973 5685
rect 3953 5635 4007 5651
rect 4041 5753 4107 5763
rect 4041 5719 4057 5753
rect 4091 5719 4107 5753
rect 4041 5715 4107 5719
rect 4041 5681 4055 5715
rect 4089 5685 4107 5715
rect 4041 5651 4057 5681
rect 4091 5651 4107 5685
rect 4041 5635 4107 5651
rect 4141 5753 4189 5797
rect 4175 5719 4189 5753
rect 4538 5729 4554 5763
rect 4588 5729 4604 5763
rect 4141 5685 4189 5719
rect 4175 5651 4189 5685
rect 4141 5635 4189 5651
rect 4410 5667 4444 5686
rect 2877 5594 2897 5599
rect 2877 5560 2894 5594
rect 2931 5565 2947 5599
rect 2928 5560 2947 5565
rect 2877 5549 2947 5560
rect 2981 5515 3015 5635
rect 3049 5565 3065 5599
rect 3099 5590 3119 5599
rect 3049 5556 3067 5565
rect 3101 5556 3119 5590
rect 3049 5549 3119 5556
rect 3951 5592 3971 5599
rect 3951 5558 3969 5592
rect 4005 5565 4021 5599
rect 4003 5558 4021 5565
rect 3951 5549 4021 5558
rect 4055 5515 4089 5635
rect 4410 5599 4444 5601
rect 4123 5565 4139 5599
rect 4173 5592 4193 5599
rect 4123 5558 4143 5565
rect 4177 5558 4193 5592
rect 4123 5549 4193 5558
rect 4410 5563 4444 5565
rect 2554 5435 2820 5436
rect 2554 5401 2570 5435
rect 2604 5401 2820 5435
rect 2554 5400 2820 5401
rect 2879 5499 2945 5515
rect 2879 5465 2911 5499
rect 2981 5499 3117 5515
rect 2981 5481 3067 5499
rect 2879 5431 2945 5465
rect 2237 5363 2303 5397
rect 2237 5329 2253 5363
rect 2287 5329 2303 5363
rect 2879 5397 2911 5431
rect 2879 5363 2945 5397
rect 2237 5324 2303 5329
rect 2430 5329 2712 5362
rect 2430 5295 2520 5329
rect 2554 5327 2712 5329
rect 2554 5295 2639 5327
rect 2430 5293 2639 5295
rect 2673 5293 2712 5327
rect 2430 5287 2712 5293
rect 2879 5329 2911 5363
rect 2879 5287 2945 5329
rect 3051 5465 3067 5481
rect 3101 5465 3117 5499
rect 3051 5431 3117 5465
rect 3051 5397 3067 5431
rect 3101 5397 3117 5431
rect 3051 5363 3117 5397
rect 3051 5329 3067 5363
rect 3101 5329 3117 5363
rect 3051 5324 3117 5329
rect 3953 5499 4019 5515
rect 3953 5465 3985 5499
rect 4055 5499 4191 5515
rect 4055 5481 4141 5499
rect 3953 5431 4019 5465
rect 3953 5397 3985 5431
rect 3953 5363 4019 5397
rect 3953 5329 3985 5363
rect 3953 5287 4019 5329
rect 4125 5465 4141 5481
rect 4175 5465 4191 5499
rect 4410 5478 4444 5497
rect 4506 5667 4540 5686
rect 4506 5599 4540 5601
rect 4506 5563 4540 5565
rect 4506 5478 4540 5497
rect 4602 5667 4636 5686
rect 4602 5599 4636 5601
rect 4602 5563 4636 5565
rect 4602 5478 4636 5497
rect 4125 5431 4191 5465
rect 4125 5397 4141 5431
rect 4175 5397 4191 5431
rect 4442 5436 4508 5438
rect 4674 5436 4708 6050
rect 4759 5831 4793 6134
rect 4990 5831 5024 6042
rect 5934 6016 5968 6374
rect 6208 6351 6298 6374
rect 6332 6383 6656 6385
rect 6332 6351 6417 6383
rect 6208 6349 6417 6351
rect 6451 6374 6656 6383
rect 6708 6374 6742 6393
rect 6880 6571 6926 6691
rect 6980 6687 7026 6703
rect 7177 6773 7229 6811
rect 7177 6739 7195 6773
rect 7265 6803 7331 6845
rect 7506 6843 7535 6877
rect 7569 6843 7627 6877
rect 7661 6843 7719 6877
rect 7753 6843 7782 6877
rect 7942 6862 7990 6874
rect 8204 6866 8220 6900
rect 8254 6866 8270 6900
rect 8570 6890 8620 6960
rect 10060 6934 10094 6950
rect 10156 7056 10190 7072
rect 10252 7058 10286 7072
rect 10370 7058 10590 7080
rect 10250 7056 10590 7058
rect 10250 7022 10252 7056
rect 10286 7044 10590 7056
rect 10286 7022 10406 7044
rect 10156 6986 10190 7020
rect 10251 7020 10252 7022
rect 10251 6986 10286 7020
rect 10554 6996 10590 7044
rect 10251 6985 10252 6986
rect 10156 6934 10190 6950
rect 10252 6934 10286 6950
rect 10458 6960 10590 6996
rect 11948 7056 11982 7072
rect 11948 6986 11982 7020
rect 8570 6876 8580 6890
rect 7265 6769 7281 6803
rect 7315 6769 7331 6803
rect 7367 6790 7401 6811
rect 7177 6710 7229 6739
rect 7367 6735 7401 6756
rect 6960 6619 6976 6653
rect 7010 6642 7026 6653
rect 6960 6608 6978 6619
rect 7012 6608 7026 6642
rect 7177 6638 7213 6710
rect 7268 6701 7401 6735
rect 7572 6797 7638 6809
rect 7572 6763 7588 6797
rect 7622 6763 7638 6797
rect 7572 6746 7638 6763
rect 7268 6650 7302 6701
rect 7572 6695 7588 6746
rect 7622 6695 7638 6746
rect 7572 6683 7638 6695
rect 7672 6797 7718 6843
rect 7706 6763 7718 6797
rect 7672 6729 7718 6763
rect 7706 6695 7718 6729
rect 7942 6828 7948 6862
rect 7982 6828 7990 6862
rect 8574 6856 8580 6876
rect 8614 6856 8620 6890
rect 8574 6846 8620 6856
rect 8702 6851 8731 6885
rect 8765 6851 8823 6885
rect 8857 6851 8915 6885
rect 8949 6851 8978 6885
rect 7942 6740 7990 6828
rect 8316 6785 8332 6819
rect 8366 6818 8382 6819
rect 8366 6786 8528 6818
rect 8768 6810 8834 6817
rect 8762 6805 8834 6810
rect 8762 6786 8784 6805
rect 8366 6785 8784 6786
rect 8316 6782 8784 6785
rect 8492 6771 8784 6782
rect 8818 6771 8834 6805
rect 8492 6750 8834 6771
rect 8188 6740 8222 6742
rect 7942 6723 8222 6740
rect 7942 6706 8188 6723
rect 6960 6605 7026 6608
rect 7172 6636 7213 6638
rect 7172 6602 7174 6636
rect 7208 6602 7213 6636
rect 7172 6600 7213 6602
rect 6880 6553 6946 6571
rect 6880 6519 6896 6553
rect 6930 6519 6946 6553
rect 6880 6485 6946 6519
rect 6880 6451 6896 6485
rect 6930 6451 6946 6485
rect 6880 6417 6946 6451
rect 6880 6383 6896 6417
rect 6930 6383 6946 6417
rect 6880 6375 6946 6383
rect 6980 6553 7022 6569
rect 7014 6519 7022 6553
rect 6980 6485 7022 6519
rect 7014 6451 7022 6485
rect 6980 6417 7022 6451
rect 7014 6383 7022 6417
rect 6451 6349 6490 6374
rect 6002 6297 6018 6331
rect 6052 6297 6068 6331
rect 6208 6310 6490 6349
rect 6980 6341 7022 6383
rect 7177 6550 7213 6600
rect 7247 6634 7302 6650
rect 7281 6600 7302 6634
rect 7247 6584 7302 6600
rect 7347 6648 7415 6665
rect 7347 6647 7367 6648
rect 7347 6613 7365 6647
rect 7401 6614 7415 6648
rect 7399 6613 7415 6614
rect 7347 6591 7415 6613
rect 7268 6555 7302 6584
rect 7572 6563 7618 6683
rect 7672 6679 7718 6695
rect 7890 6658 7906 6659
rect 7652 6611 7668 6645
rect 7702 6638 7718 6645
rect 7770 6638 7906 6658
rect 7702 6625 7906 6638
rect 7940 6625 7956 6659
rect 7702 6624 7956 6625
rect 7702 6611 7810 6624
rect 7890 6622 7956 6624
rect 8188 6655 8222 6657
rect 7652 6597 7810 6611
rect 7666 6596 7810 6597
rect 8188 6619 8222 6621
rect 7862 6563 7896 6582
rect 7177 6500 7231 6550
rect 7268 6521 7403 6555
rect 7177 6466 7195 6500
rect 7229 6466 7231 6500
rect 7367 6487 7403 6521
rect 7177 6419 7231 6466
rect 7177 6385 7195 6419
rect 7229 6385 7231 6419
rect 7177 6369 7231 6385
rect 7265 6453 7281 6487
rect 7315 6453 7331 6487
rect 7265 6419 7331 6453
rect 7265 6385 7281 6419
rect 7315 6385 7331 6419
rect 6376 6308 6490 6310
rect 6648 6297 6664 6331
rect 6698 6297 6714 6331
rect 6814 6307 6843 6341
rect 6877 6307 6935 6341
rect 6969 6307 7027 6341
rect 7061 6307 7090 6341
rect 7265 6335 7331 6385
rect 7401 6453 7403 6487
rect 7367 6419 7403 6453
rect 7401 6385 7403 6419
rect 7367 6369 7403 6385
rect 7572 6545 7638 6563
rect 7572 6511 7588 6545
rect 7622 6511 7638 6545
rect 7572 6477 7638 6511
rect 7572 6443 7588 6477
rect 7622 6443 7638 6477
rect 7572 6409 7638 6443
rect 7572 6375 7588 6409
rect 7622 6375 7638 6409
rect 7572 6367 7638 6375
rect 7672 6545 7714 6561
rect 7706 6511 7714 6545
rect 7672 6477 7714 6511
rect 7706 6443 7714 6477
rect 7672 6409 7714 6443
rect 7862 6495 7896 6497
rect 7862 6459 7896 6461
rect 7706 6375 7714 6409
rect 6981 6300 7015 6307
rect 7160 6301 7189 6335
rect 7223 6301 7281 6335
rect 7315 6301 7373 6335
rect 7407 6301 7436 6335
rect 7672 6333 7714 6375
rect 7822 6393 7862 6414
rect 7950 6563 7984 6582
rect 8188 6534 8222 6553
rect 8284 6723 8318 6742
rect 8284 6655 8318 6657
rect 8284 6619 8318 6621
rect 8284 6534 8318 6553
rect 8380 6723 8414 6742
rect 8768 6737 8834 6750
rect 8768 6703 8784 6737
rect 8818 6703 8834 6737
rect 8768 6691 8834 6703
rect 8868 6805 8914 6851
rect 9048 6845 9077 6879
rect 9111 6845 9169 6879
rect 9203 6845 9261 6879
rect 9295 6845 9324 6879
rect 8902 6771 8914 6805
rect 8868 6737 8914 6771
rect 8902 6703 8914 6737
rect 8380 6655 8414 6657
rect 8536 6625 8552 6659
rect 8586 6625 8602 6659
rect 8380 6619 8414 6621
rect 8380 6534 8414 6553
rect 8508 6563 8542 6582
rect 7950 6495 7984 6497
rect 8508 6495 8542 6497
rect 7950 6459 7984 6461
rect 8220 6457 8236 6491
rect 8270 6457 8286 6491
rect 8508 6459 8542 6461
rect 7896 6393 7898 6414
rect 7822 6374 7898 6393
rect 7984 6393 8508 6418
rect 8596 6563 8630 6582
rect 8596 6495 8630 6497
rect 8596 6459 8630 6461
rect 8542 6393 8544 6418
rect 7950 6385 8544 6393
rect 7950 6374 8186 6385
rect 7506 6299 7535 6333
rect 7569 6299 7627 6333
rect 7661 6299 7719 6333
rect 7753 6299 7782 6333
rect 6068 6212 6114 6218
rect 6068 6210 6556 6212
rect 6068 6176 6076 6210
rect 6110 6193 6556 6210
rect 6110 6188 6506 6193
rect 6110 6178 6385 6188
rect 6110 6176 6114 6178
rect 6068 6174 6114 6176
rect 6286 6154 6385 6178
rect 6419 6159 6506 6188
rect 6540 6168 6556 6193
rect 6540 6159 6681 6168
rect 6419 6154 6681 6159
rect 6286 6134 6681 6154
rect 6410 6050 6426 6084
rect 6460 6050 6596 6084
rect 5934 6000 6316 6016
rect 5934 5976 6282 6000
rect 6282 5930 6316 5964
rect 6282 5878 6316 5894
rect 6378 6000 6412 6016
rect 6378 5930 6412 5964
rect 6378 5878 6412 5894
rect 6474 6000 6508 6016
rect 6474 5930 6508 5964
rect 6474 5878 6508 5894
rect 4748 5797 4777 5831
rect 4811 5797 4869 5831
rect 4903 5797 4961 5831
rect 4995 5797 5024 5831
rect 5822 5797 5851 5831
rect 5885 5797 5943 5831
rect 5977 5797 6035 5831
rect 6069 5797 6098 5831
rect 6314 5810 6330 5844
rect 6364 5810 6380 5844
rect 4767 5753 4821 5797
rect 4767 5719 4787 5753
rect 4767 5685 4821 5719
rect 4767 5651 4787 5685
rect 4767 5635 4821 5651
rect 4855 5753 4921 5763
rect 4855 5719 4871 5753
rect 4905 5719 4921 5753
rect 4855 5710 4921 5719
rect 4855 5685 4873 5710
rect 4855 5651 4871 5685
rect 4907 5676 4921 5710
rect 4905 5651 4921 5676
rect 4855 5635 4921 5651
rect 4955 5753 5003 5797
rect 4989 5719 5003 5753
rect 4955 5685 5003 5719
rect 4989 5651 5003 5685
rect 4955 5635 5003 5651
rect 5841 5753 5895 5797
rect 5841 5719 5861 5753
rect 5841 5685 5895 5719
rect 5841 5651 5861 5685
rect 5841 5635 5895 5651
rect 5929 5753 5995 5763
rect 5929 5719 5945 5753
rect 5979 5719 5995 5753
rect 5929 5715 5995 5719
rect 5929 5681 5943 5715
rect 5977 5685 5995 5715
rect 5929 5651 5945 5681
rect 5979 5651 5995 5685
rect 5929 5635 5995 5651
rect 6029 5753 6077 5797
rect 6063 5719 6077 5753
rect 6426 5729 6442 5763
rect 6476 5729 6492 5763
rect 6029 5685 6077 5719
rect 6063 5651 6077 5685
rect 6029 5635 6077 5651
rect 6298 5667 6332 5686
rect 4765 5594 4785 5599
rect 4765 5560 4782 5594
rect 4819 5565 4835 5599
rect 4816 5560 4835 5565
rect 4765 5549 4835 5560
rect 4869 5515 4903 5635
rect 4937 5565 4953 5599
rect 4987 5590 5007 5599
rect 4937 5556 4955 5565
rect 4989 5556 5007 5590
rect 4937 5549 5007 5556
rect 5839 5592 5859 5599
rect 5839 5558 5857 5592
rect 5893 5565 5909 5599
rect 5891 5558 5909 5565
rect 5839 5549 5909 5558
rect 5943 5515 5977 5635
rect 6298 5599 6332 5601
rect 6011 5565 6027 5599
rect 6061 5592 6081 5599
rect 6011 5558 6031 5565
rect 6065 5558 6081 5592
rect 6011 5549 6081 5558
rect 6298 5563 6332 5565
rect 4442 5435 4708 5436
rect 4442 5401 4458 5435
rect 4492 5401 4708 5435
rect 4442 5400 4708 5401
rect 4767 5499 4833 5515
rect 4767 5465 4799 5499
rect 4869 5499 5005 5515
rect 4869 5481 4955 5499
rect 4767 5431 4833 5465
rect 4125 5363 4191 5397
rect 4125 5329 4141 5363
rect 4175 5329 4191 5363
rect 4767 5397 4799 5431
rect 4767 5363 4833 5397
rect 4125 5324 4191 5329
rect 4318 5329 4600 5362
rect 4318 5295 4408 5329
rect 4442 5327 4600 5329
rect 4442 5295 4527 5327
rect 4318 5293 4527 5295
rect 4561 5293 4600 5327
rect 4318 5287 4600 5293
rect 4767 5329 4799 5363
rect 4767 5287 4833 5329
rect 4939 5465 4955 5481
rect 4989 5465 5005 5499
rect 4939 5431 5005 5465
rect 4939 5397 4955 5431
rect 4989 5397 5005 5431
rect 4939 5363 5005 5397
rect 4939 5329 4955 5363
rect 4989 5329 5005 5363
rect 4939 5324 5005 5329
rect 5841 5499 5907 5515
rect 5841 5465 5873 5499
rect 5943 5499 6079 5515
rect 5943 5481 6029 5499
rect 5841 5431 5907 5465
rect 5841 5397 5873 5431
rect 5841 5363 5907 5397
rect 5841 5329 5873 5363
rect 5841 5287 5907 5329
rect 6013 5465 6029 5481
rect 6063 5465 6079 5499
rect 6298 5478 6332 5497
rect 6394 5667 6428 5686
rect 6394 5599 6428 5601
rect 6394 5563 6428 5565
rect 6394 5478 6428 5497
rect 6490 5667 6524 5686
rect 6490 5599 6524 5601
rect 6490 5563 6524 5565
rect 6490 5478 6524 5497
rect 6013 5431 6079 5465
rect 6013 5397 6029 5431
rect 6063 5397 6079 5431
rect 6330 5436 6396 5438
rect 6562 5436 6596 6050
rect 6647 5831 6681 6134
rect 6878 5831 6912 6042
rect 7822 6016 7856 6374
rect 8096 6351 8186 6374
rect 8220 6383 8544 6385
rect 8220 6351 8305 6383
rect 8096 6349 8305 6351
rect 8339 6374 8544 6383
rect 8596 6374 8630 6393
rect 8768 6571 8814 6691
rect 8868 6687 8914 6703
rect 9065 6773 9117 6811
rect 9065 6739 9083 6773
rect 9153 6803 9219 6845
rect 9394 6843 9423 6877
rect 9457 6843 9515 6877
rect 9549 6843 9607 6877
rect 9641 6843 9670 6877
rect 9830 6862 9878 6874
rect 10092 6866 10108 6900
rect 10142 6866 10158 6900
rect 10458 6890 10508 6960
rect 11948 6934 11982 6950
rect 12044 7056 12078 7072
rect 12140 7058 12174 7072
rect 12258 7058 12478 7080
rect 12138 7056 12478 7058
rect 12138 7022 12140 7056
rect 12174 7044 12478 7056
rect 12174 7022 12294 7044
rect 12044 6986 12078 7020
rect 12139 7020 12140 7022
rect 12139 6986 12174 7020
rect 12442 6996 12478 7044
rect 12139 6985 12140 6986
rect 12044 6934 12078 6950
rect 12140 6934 12174 6950
rect 12346 6960 12478 6996
rect 13836 7056 13870 7072
rect 13836 6986 13870 7020
rect 10458 6876 10468 6890
rect 9153 6769 9169 6803
rect 9203 6769 9219 6803
rect 9255 6790 9289 6811
rect 9065 6710 9117 6739
rect 9255 6735 9289 6756
rect 8848 6619 8864 6653
rect 8898 6642 8914 6653
rect 8848 6608 8866 6619
rect 8900 6608 8914 6642
rect 9065 6638 9101 6710
rect 9156 6701 9289 6735
rect 9460 6797 9526 6809
rect 9460 6763 9476 6797
rect 9510 6763 9526 6797
rect 9460 6746 9526 6763
rect 9156 6650 9190 6701
rect 9460 6695 9476 6746
rect 9510 6695 9526 6746
rect 9460 6683 9526 6695
rect 9560 6797 9606 6843
rect 9594 6763 9606 6797
rect 9560 6729 9606 6763
rect 9594 6695 9606 6729
rect 9830 6828 9836 6862
rect 9870 6828 9878 6862
rect 10462 6856 10468 6876
rect 10502 6856 10508 6890
rect 10462 6846 10508 6856
rect 10590 6851 10619 6885
rect 10653 6851 10711 6885
rect 10745 6851 10803 6885
rect 10837 6851 10866 6885
rect 9830 6740 9878 6828
rect 10204 6785 10220 6819
rect 10254 6818 10270 6819
rect 10254 6786 10416 6818
rect 10656 6810 10722 6817
rect 10650 6805 10722 6810
rect 10650 6786 10672 6805
rect 10254 6785 10672 6786
rect 10204 6782 10672 6785
rect 10380 6771 10672 6782
rect 10706 6771 10722 6805
rect 10380 6750 10722 6771
rect 10076 6740 10110 6742
rect 9830 6723 10110 6740
rect 9830 6706 10076 6723
rect 8848 6605 8914 6608
rect 9060 6636 9101 6638
rect 9060 6602 9062 6636
rect 9096 6602 9101 6636
rect 9060 6600 9101 6602
rect 8768 6553 8834 6571
rect 8768 6519 8784 6553
rect 8818 6519 8834 6553
rect 8768 6485 8834 6519
rect 8768 6451 8784 6485
rect 8818 6451 8834 6485
rect 8768 6417 8834 6451
rect 8768 6383 8784 6417
rect 8818 6383 8834 6417
rect 8768 6375 8834 6383
rect 8868 6553 8910 6569
rect 8902 6519 8910 6553
rect 8868 6485 8910 6519
rect 8902 6451 8910 6485
rect 8868 6417 8910 6451
rect 8902 6383 8910 6417
rect 8339 6349 8378 6374
rect 7890 6297 7906 6331
rect 7940 6297 7956 6331
rect 8096 6310 8378 6349
rect 8868 6341 8910 6383
rect 9065 6550 9101 6600
rect 9135 6634 9190 6650
rect 9169 6600 9190 6634
rect 9135 6584 9190 6600
rect 9235 6648 9303 6665
rect 9235 6647 9255 6648
rect 9235 6613 9253 6647
rect 9289 6614 9303 6648
rect 9287 6613 9303 6614
rect 9235 6591 9303 6613
rect 9156 6555 9190 6584
rect 9460 6563 9506 6683
rect 9560 6679 9606 6695
rect 9778 6658 9794 6659
rect 9540 6611 9556 6645
rect 9590 6638 9606 6645
rect 9658 6638 9794 6658
rect 9590 6625 9794 6638
rect 9828 6625 9844 6659
rect 9590 6624 9844 6625
rect 9590 6611 9698 6624
rect 9778 6622 9844 6624
rect 10076 6655 10110 6657
rect 9540 6597 9698 6611
rect 9554 6596 9698 6597
rect 10076 6619 10110 6621
rect 9750 6563 9784 6582
rect 9065 6500 9119 6550
rect 9156 6521 9291 6555
rect 9065 6466 9083 6500
rect 9117 6466 9119 6500
rect 9255 6487 9291 6521
rect 9065 6419 9119 6466
rect 9065 6385 9083 6419
rect 9117 6385 9119 6419
rect 9065 6369 9119 6385
rect 9153 6453 9169 6487
rect 9203 6453 9219 6487
rect 9153 6419 9219 6453
rect 9153 6385 9169 6419
rect 9203 6385 9219 6419
rect 8264 6308 8378 6310
rect 8536 6297 8552 6331
rect 8586 6297 8602 6331
rect 8702 6307 8731 6341
rect 8765 6307 8823 6341
rect 8857 6307 8915 6341
rect 8949 6307 8978 6341
rect 9153 6335 9219 6385
rect 9289 6453 9291 6487
rect 9255 6419 9291 6453
rect 9289 6385 9291 6419
rect 9255 6369 9291 6385
rect 9460 6545 9526 6563
rect 9460 6511 9476 6545
rect 9510 6511 9526 6545
rect 9460 6477 9526 6511
rect 9460 6443 9476 6477
rect 9510 6443 9526 6477
rect 9460 6409 9526 6443
rect 9460 6375 9476 6409
rect 9510 6375 9526 6409
rect 9460 6367 9526 6375
rect 9560 6545 9602 6561
rect 9594 6511 9602 6545
rect 9560 6477 9602 6511
rect 9594 6443 9602 6477
rect 9560 6409 9602 6443
rect 9750 6495 9784 6497
rect 9750 6459 9784 6461
rect 9594 6375 9602 6409
rect 8869 6300 8903 6307
rect 9048 6301 9077 6335
rect 9111 6301 9169 6335
rect 9203 6301 9261 6335
rect 9295 6301 9324 6335
rect 9560 6333 9602 6375
rect 9710 6393 9750 6414
rect 9838 6563 9872 6582
rect 10076 6534 10110 6553
rect 10172 6723 10206 6742
rect 10172 6655 10206 6657
rect 10172 6619 10206 6621
rect 10172 6534 10206 6553
rect 10268 6723 10302 6742
rect 10656 6737 10722 6750
rect 10656 6703 10672 6737
rect 10706 6703 10722 6737
rect 10656 6691 10722 6703
rect 10756 6805 10802 6851
rect 10936 6845 10965 6879
rect 10999 6845 11057 6879
rect 11091 6845 11149 6879
rect 11183 6845 11212 6879
rect 10790 6771 10802 6805
rect 10756 6737 10802 6771
rect 10790 6703 10802 6737
rect 10268 6655 10302 6657
rect 10424 6625 10440 6659
rect 10474 6625 10490 6659
rect 10268 6619 10302 6621
rect 10268 6534 10302 6553
rect 10396 6563 10430 6582
rect 9838 6495 9872 6497
rect 10396 6495 10430 6497
rect 9838 6459 9872 6461
rect 10108 6457 10124 6491
rect 10158 6457 10174 6491
rect 10396 6459 10430 6461
rect 9784 6393 9786 6414
rect 9710 6374 9786 6393
rect 9872 6393 10396 6418
rect 10484 6563 10518 6582
rect 10484 6495 10518 6497
rect 10484 6459 10518 6461
rect 10430 6393 10432 6418
rect 9838 6385 10432 6393
rect 9838 6374 10074 6385
rect 9394 6299 9423 6333
rect 9457 6299 9515 6333
rect 9549 6299 9607 6333
rect 9641 6299 9670 6333
rect 7956 6212 8002 6218
rect 7956 6210 8444 6212
rect 7956 6176 7964 6210
rect 7998 6193 8444 6210
rect 7998 6188 8394 6193
rect 7998 6178 8273 6188
rect 7998 6176 8002 6178
rect 7956 6174 8002 6176
rect 8174 6154 8273 6178
rect 8307 6159 8394 6188
rect 8428 6168 8444 6193
rect 8428 6159 8569 6168
rect 8307 6154 8569 6159
rect 8174 6134 8569 6154
rect 8298 6050 8314 6084
rect 8348 6050 8484 6084
rect 7822 6000 8204 6016
rect 7822 5976 8170 6000
rect 8170 5930 8204 5964
rect 8170 5878 8204 5894
rect 8266 6000 8300 6016
rect 8266 5930 8300 5964
rect 8266 5878 8300 5894
rect 8362 6000 8396 6016
rect 8362 5930 8396 5964
rect 8362 5878 8396 5894
rect 6636 5797 6665 5831
rect 6699 5797 6757 5831
rect 6791 5797 6849 5831
rect 6883 5797 6912 5831
rect 7710 5797 7739 5831
rect 7773 5797 7831 5831
rect 7865 5797 7923 5831
rect 7957 5797 7986 5831
rect 8202 5810 8218 5844
rect 8252 5810 8268 5844
rect 6655 5753 6709 5797
rect 6655 5719 6675 5753
rect 6655 5685 6709 5719
rect 6655 5651 6675 5685
rect 6655 5635 6709 5651
rect 6743 5753 6809 5763
rect 6743 5719 6759 5753
rect 6793 5719 6809 5753
rect 6743 5710 6809 5719
rect 6743 5685 6761 5710
rect 6743 5651 6759 5685
rect 6795 5676 6809 5710
rect 6793 5651 6809 5676
rect 6743 5635 6809 5651
rect 6843 5753 6891 5797
rect 6877 5719 6891 5753
rect 6843 5685 6891 5719
rect 6877 5651 6891 5685
rect 6843 5635 6891 5651
rect 7729 5753 7783 5797
rect 7729 5719 7749 5753
rect 7729 5685 7783 5719
rect 7729 5651 7749 5685
rect 7729 5635 7783 5651
rect 7817 5753 7883 5763
rect 7817 5719 7833 5753
rect 7867 5719 7883 5753
rect 7817 5715 7883 5719
rect 7817 5681 7831 5715
rect 7865 5685 7883 5715
rect 7817 5651 7833 5681
rect 7867 5651 7883 5685
rect 7817 5635 7883 5651
rect 7917 5753 7965 5797
rect 7951 5719 7965 5753
rect 8314 5729 8330 5763
rect 8364 5729 8380 5763
rect 7917 5685 7965 5719
rect 7951 5651 7965 5685
rect 7917 5635 7965 5651
rect 8186 5667 8220 5686
rect 6653 5594 6673 5599
rect 6653 5560 6670 5594
rect 6707 5565 6723 5599
rect 6704 5560 6723 5565
rect 6653 5549 6723 5560
rect 6757 5515 6791 5635
rect 6825 5565 6841 5599
rect 6875 5590 6895 5599
rect 6825 5556 6843 5565
rect 6877 5556 6895 5590
rect 6825 5549 6895 5556
rect 7727 5592 7747 5599
rect 7727 5558 7745 5592
rect 7781 5565 7797 5599
rect 7779 5558 7797 5565
rect 7727 5549 7797 5558
rect 7831 5515 7865 5635
rect 8186 5599 8220 5601
rect 7899 5565 7915 5599
rect 7949 5592 7969 5599
rect 7899 5558 7919 5565
rect 7953 5558 7969 5592
rect 7899 5549 7969 5558
rect 8186 5563 8220 5565
rect 6330 5435 6596 5436
rect 6330 5401 6346 5435
rect 6380 5401 6596 5435
rect 6330 5400 6596 5401
rect 6655 5499 6721 5515
rect 6655 5465 6687 5499
rect 6757 5499 6893 5515
rect 6757 5481 6843 5499
rect 6655 5431 6721 5465
rect 6013 5363 6079 5397
rect 6013 5329 6029 5363
rect 6063 5329 6079 5363
rect 6655 5397 6687 5431
rect 6655 5363 6721 5397
rect 6013 5324 6079 5329
rect 6206 5329 6488 5362
rect 6206 5295 6296 5329
rect 6330 5327 6488 5329
rect 6330 5295 6415 5327
rect 6206 5293 6415 5295
rect 6449 5293 6488 5327
rect 6206 5287 6488 5293
rect 6655 5329 6687 5363
rect 6655 5287 6721 5329
rect 6827 5465 6843 5481
rect 6877 5465 6893 5499
rect 6827 5431 6893 5465
rect 6827 5397 6843 5431
rect 6877 5397 6893 5431
rect 6827 5363 6893 5397
rect 6827 5329 6843 5363
rect 6877 5329 6893 5363
rect 6827 5324 6893 5329
rect 7729 5499 7795 5515
rect 7729 5465 7761 5499
rect 7831 5499 7967 5515
rect 7831 5481 7917 5499
rect 7729 5431 7795 5465
rect 7729 5397 7761 5431
rect 7729 5363 7795 5397
rect 7729 5329 7761 5363
rect 7729 5287 7795 5329
rect 7901 5465 7917 5481
rect 7951 5465 7967 5499
rect 8186 5478 8220 5497
rect 8282 5667 8316 5686
rect 8282 5599 8316 5601
rect 8282 5563 8316 5565
rect 8282 5478 8316 5497
rect 8378 5667 8412 5686
rect 8378 5599 8412 5601
rect 8378 5563 8412 5565
rect 8378 5478 8412 5497
rect 7901 5431 7967 5465
rect 7901 5397 7917 5431
rect 7951 5397 7967 5431
rect 8218 5436 8284 5438
rect 8450 5436 8484 6050
rect 8535 5831 8569 6134
rect 8766 5831 8800 6042
rect 9710 6016 9744 6374
rect 9984 6351 10074 6374
rect 10108 6383 10432 6385
rect 10108 6351 10193 6383
rect 9984 6349 10193 6351
rect 10227 6374 10432 6383
rect 10484 6374 10518 6393
rect 10656 6571 10702 6691
rect 10756 6687 10802 6703
rect 10953 6773 11005 6811
rect 10953 6739 10971 6773
rect 11041 6803 11107 6845
rect 11282 6843 11311 6877
rect 11345 6843 11403 6877
rect 11437 6843 11495 6877
rect 11529 6843 11558 6877
rect 11718 6862 11766 6874
rect 11980 6866 11996 6900
rect 12030 6866 12046 6900
rect 12346 6890 12396 6960
rect 13836 6934 13870 6950
rect 13932 7056 13966 7072
rect 14028 7058 14062 7072
rect 14146 7058 14366 7080
rect 14026 7056 14366 7058
rect 14026 7022 14028 7056
rect 14062 7044 14366 7056
rect 14062 7022 14182 7044
rect 13932 6986 13966 7020
rect 14027 7020 14028 7022
rect 14027 6986 14062 7020
rect 14330 6996 14366 7044
rect 14027 6985 14028 6986
rect 13932 6934 13966 6950
rect 14028 6934 14062 6950
rect 14234 6960 14366 6996
rect 15718 7056 15752 7072
rect 15718 6986 15752 7020
rect 12346 6876 12356 6890
rect 11041 6769 11057 6803
rect 11091 6769 11107 6803
rect 11143 6790 11177 6811
rect 10953 6710 11005 6739
rect 11143 6735 11177 6756
rect 10736 6619 10752 6653
rect 10786 6642 10802 6653
rect 10736 6608 10754 6619
rect 10788 6608 10802 6642
rect 10953 6638 10989 6710
rect 11044 6701 11177 6735
rect 11348 6797 11414 6809
rect 11348 6763 11364 6797
rect 11398 6763 11414 6797
rect 11348 6746 11414 6763
rect 11044 6650 11078 6701
rect 11348 6695 11364 6746
rect 11398 6695 11414 6746
rect 11348 6683 11414 6695
rect 11448 6797 11494 6843
rect 11482 6763 11494 6797
rect 11448 6729 11494 6763
rect 11482 6695 11494 6729
rect 11718 6828 11724 6862
rect 11758 6828 11766 6862
rect 12350 6856 12356 6876
rect 12390 6856 12396 6890
rect 12350 6846 12396 6856
rect 12478 6851 12507 6885
rect 12541 6851 12599 6885
rect 12633 6851 12691 6885
rect 12725 6851 12754 6885
rect 11718 6740 11766 6828
rect 12092 6785 12108 6819
rect 12142 6818 12158 6819
rect 12142 6786 12304 6818
rect 12544 6810 12610 6817
rect 12538 6805 12610 6810
rect 12538 6786 12560 6805
rect 12142 6785 12560 6786
rect 12092 6782 12560 6785
rect 12268 6771 12560 6782
rect 12594 6771 12610 6805
rect 12268 6750 12610 6771
rect 11964 6740 11998 6742
rect 11718 6723 11998 6740
rect 11718 6706 11964 6723
rect 10736 6605 10802 6608
rect 10948 6636 10989 6638
rect 10948 6602 10950 6636
rect 10984 6602 10989 6636
rect 10948 6600 10989 6602
rect 10656 6553 10722 6571
rect 10656 6519 10672 6553
rect 10706 6519 10722 6553
rect 10656 6485 10722 6519
rect 10656 6451 10672 6485
rect 10706 6451 10722 6485
rect 10656 6417 10722 6451
rect 10656 6383 10672 6417
rect 10706 6383 10722 6417
rect 10656 6375 10722 6383
rect 10756 6553 10798 6569
rect 10790 6519 10798 6553
rect 10756 6485 10798 6519
rect 10790 6451 10798 6485
rect 10756 6417 10798 6451
rect 10790 6383 10798 6417
rect 10227 6349 10266 6374
rect 9778 6297 9794 6331
rect 9828 6297 9844 6331
rect 9984 6310 10266 6349
rect 10756 6341 10798 6383
rect 10953 6550 10989 6600
rect 11023 6634 11078 6650
rect 11057 6600 11078 6634
rect 11023 6584 11078 6600
rect 11123 6648 11191 6665
rect 11123 6647 11143 6648
rect 11123 6613 11141 6647
rect 11177 6614 11191 6648
rect 11175 6613 11191 6614
rect 11123 6591 11191 6613
rect 11044 6555 11078 6584
rect 11348 6563 11394 6683
rect 11448 6679 11494 6695
rect 11666 6658 11682 6659
rect 11428 6611 11444 6645
rect 11478 6638 11494 6645
rect 11546 6638 11682 6658
rect 11478 6625 11682 6638
rect 11716 6625 11732 6659
rect 11478 6624 11732 6625
rect 11478 6611 11586 6624
rect 11666 6622 11732 6624
rect 11964 6655 11998 6657
rect 11428 6597 11586 6611
rect 11442 6596 11586 6597
rect 11964 6619 11998 6621
rect 11638 6563 11672 6582
rect 10953 6500 11007 6550
rect 11044 6521 11179 6555
rect 10953 6466 10971 6500
rect 11005 6466 11007 6500
rect 11143 6487 11179 6521
rect 10953 6419 11007 6466
rect 10953 6385 10971 6419
rect 11005 6385 11007 6419
rect 10953 6369 11007 6385
rect 11041 6453 11057 6487
rect 11091 6453 11107 6487
rect 11041 6419 11107 6453
rect 11041 6385 11057 6419
rect 11091 6385 11107 6419
rect 10152 6308 10266 6310
rect 10424 6297 10440 6331
rect 10474 6297 10490 6331
rect 10590 6307 10619 6341
rect 10653 6307 10711 6341
rect 10745 6307 10803 6341
rect 10837 6307 10866 6341
rect 11041 6335 11107 6385
rect 11177 6453 11179 6487
rect 11143 6419 11179 6453
rect 11177 6385 11179 6419
rect 11143 6369 11179 6385
rect 11348 6545 11414 6563
rect 11348 6511 11364 6545
rect 11398 6511 11414 6545
rect 11348 6477 11414 6511
rect 11348 6443 11364 6477
rect 11398 6443 11414 6477
rect 11348 6409 11414 6443
rect 11348 6375 11364 6409
rect 11398 6375 11414 6409
rect 11348 6367 11414 6375
rect 11448 6545 11490 6561
rect 11482 6511 11490 6545
rect 11448 6477 11490 6511
rect 11482 6443 11490 6477
rect 11448 6409 11490 6443
rect 11638 6495 11672 6497
rect 11638 6459 11672 6461
rect 11482 6375 11490 6409
rect 10757 6300 10791 6307
rect 10936 6301 10965 6335
rect 10999 6301 11057 6335
rect 11091 6301 11149 6335
rect 11183 6301 11212 6335
rect 11448 6333 11490 6375
rect 11598 6393 11638 6414
rect 11726 6563 11760 6582
rect 11964 6534 11998 6553
rect 12060 6723 12094 6742
rect 12060 6655 12094 6657
rect 12060 6619 12094 6621
rect 12060 6534 12094 6553
rect 12156 6723 12190 6742
rect 12544 6737 12610 6750
rect 12544 6703 12560 6737
rect 12594 6703 12610 6737
rect 12544 6691 12610 6703
rect 12644 6805 12690 6851
rect 12824 6845 12853 6879
rect 12887 6845 12945 6879
rect 12979 6845 13037 6879
rect 13071 6845 13100 6879
rect 12678 6771 12690 6805
rect 12644 6737 12690 6771
rect 12678 6703 12690 6737
rect 12156 6655 12190 6657
rect 12312 6625 12328 6659
rect 12362 6625 12378 6659
rect 12156 6619 12190 6621
rect 12156 6534 12190 6553
rect 12284 6563 12318 6582
rect 11726 6495 11760 6497
rect 12284 6495 12318 6497
rect 11726 6459 11760 6461
rect 11996 6457 12012 6491
rect 12046 6457 12062 6491
rect 12284 6459 12318 6461
rect 11672 6393 11674 6414
rect 11598 6374 11674 6393
rect 11760 6393 12284 6418
rect 12372 6563 12406 6582
rect 12372 6495 12406 6497
rect 12372 6459 12406 6461
rect 12318 6393 12320 6418
rect 11726 6385 12320 6393
rect 11726 6374 11962 6385
rect 11282 6299 11311 6333
rect 11345 6299 11403 6333
rect 11437 6299 11495 6333
rect 11529 6299 11558 6333
rect 9844 6212 9890 6218
rect 9844 6210 10332 6212
rect 9844 6176 9852 6210
rect 9886 6193 10332 6210
rect 9886 6188 10282 6193
rect 9886 6178 10161 6188
rect 9886 6176 9890 6178
rect 9844 6174 9890 6176
rect 10062 6154 10161 6178
rect 10195 6159 10282 6188
rect 10316 6168 10332 6193
rect 10316 6159 10457 6168
rect 10195 6154 10457 6159
rect 10062 6134 10457 6154
rect 10186 6050 10202 6084
rect 10236 6050 10372 6084
rect 9710 6000 10092 6016
rect 9710 5976 10058 6000
rect 10058 5930 10092 5964
rect 10058 5878 10092 5894
rect 10154 6000 10188 6016
rect 10154 5930 10188 5964
rect 10154 5878 10188 5894
rect 10250 6000 10284 6016
rect 10250 5930 10284 5964
rect 10250 5878 10284 5894
rect 8524 5797 8553 5831
rect 8587 5797 8645 5831
rect 8679 5797 8737 5831
rect 8771 5797 8800 5831
rect 9598 5797 9627 5831
rect 9661 5797 9719 5831
rect 9753 5797 9811 5831
rect 9845 5797 9874 5831
rect 10090 5810 10106 5844
rect 10140 5810 10156 5844
rect 8543 5753 8597 5797
rect 8543 5719 8563 5753
rect 8543 5685 8597 5719
rect 8543 5651 8563 5685
rect 8543 5635 8597 5651
rect 8631 5753 8697 5763
rect 8631 5719 8647 5753
rect 8681 5719 8697 5753
rect 8631 5710 8697 5719
rect 8631 5685 8649 5710
rect 8631 5651 8647 5685
rect 8683 5676 8697 5710
rect 8681 5651 8697 5676
rect 8631 5635 8697 5651
rect 8731 5753 8779 5797
rect 8765 5719 8779 5753
rect 8731 5685 8779 5719
rect 8765 5651 8779 5685
rect 8731 5635 8779 5651
rect 9617 5753 9671 5797
rect 9617 5719 9637 5753
rect 9617 5685 9671 5719
rect 9617 5651 9637 5685
rect 9617 5635 9671 5651
rect 9705 5753 9771 5763
rect 9705 5719 9721 5753
rect 9755 5719 9771 5753
rect 9705 5715 9771 5719
rect 9705 5681 9719 5715
rect 9753 5685 9771 5715
rect 9705 5651 9721 5681
rect 9755 5651 9771 5685
rect 9705 5635 9771 5651
rect 9805 5753 9853 5797
rect 9839 5719 9853 5753
rect 10202 5729 10218 5763
rect 10252 5729 10268 5763
rect 9805 5685 9853 5719
rect 9839 5651 9853 5685
rect 9805 5635 9853 5651
rect 10074 5667 10108 5686
rect 8541 5594 8561 5599
rect 8541 5560 8558 5594
rect 8595 5565 8611 5599
rect 8592 5560 8611 5565
rect 8541 5549 8611 5560
rect 8645 5515 8679 5635
rect 8713 5565 8729 5599
rect 8763 5590 8783 5599
rect 8713 5556 8731 5565
rect 8765 5556 8783 5590
rect 8713 5549 8783 5556
rect 9615 5592 9635 5599
rect 9615 5558 9633 5592
rect 9669 5565 9685 5599
rect 9667 5558 9685 5565
rect 9615 5549 9685 5558
rect 9719 5515 9753 5635
rect 10074 5599 10108 5601
rect 9787 5565 9803 5599
rect 9837 5592 9857 5599
rect 9787 5558 9807 5565
rect 9841 5558 9857 5592
rect 9787 5549 9857 5558
rect 10074 5563 10108 5565
rect 8218 5435 8484 5436
rect 8218 5401 8234 5435
rect 8268 5401 8484 5435
rect 8218 5400 8484 5401
rect 8543 5499 8609 5515
rect 8543 5465 8575 5499
rect 8645 5499 8781 5515
rect 8645 5481 8731 5499
rect 8543 5431 8609 5465
rect 7901 5363 7967 5397
rect 7901 5329 7917 5363
rect 7951 5329 7967 5363
rect 8543 5397 8575 5431
rect 8543 5363 8609 5397
rect 7901 5324 7967 5329
rect 8094 5329 8376 5362
rect 8094 5295 8184 5329
rect 8218 5327 8376 5329
rect 8218 5295 8303 5327
rect 8094 5293 8303 5295
rect 8337 5293 8376 5327
rect 8094 5287 8376 5293
rect 8543 5329 8575 5363
rect 8543 5287 8609 5329
rect 8715 5465 8731 5481
rect 8765 5465 8781 5499
rect 8715 5431 8781 5465
rect 8715 5397 8731 5431
rect 8765 5397 8781 5431
rect 8715 5363 8781 5397
rect 8715 5329 8731 5363
rect 8765 5329 8781 5363
rect 8715 5324 8781 5329
rect 9617 5499 9683 5515
rect 9617 5465 9649 5499
rect 9719 5499 9855 5515
rect 9719 5481 9805 5499
rect 9617 5431 9683 5465
rect 9617 5397 9649 5431
rect 9617 5363 9683 5397
rect 9617 5329 9649 5363
rect 9617 5287 9683 5329
rect 9789 5465 9805 5481
rect 9839 5465 9855 5499
rect 10074 5478 10108 5497
rect 10170 5667 10204 5686
rect 10170 5599 10204 5601
rect 10170 5563 10204 5565
rect 10170 5478 10204 5497
rect 10266 5667 10300 5686
rect 10266 5599 10300 5601
rect 10266 5563 10300 5565
rect 10266 5478 10300 5497
rect 9789 5431 9855 5465
rect 9789 5397 9805 5431
rect 9839 5397 9855 5431
rect 10106 5436 10172 5438
rect 10338 5436 10372 6050
rect 10423 5831 10457 6134
rect 10654 5831 10688 6042
rect 11598 6016 11632 6374
rect 11872 6351 11962 6374
rect 11996 6383 12320 6385
rect 11996 6351 12081 6383
rect 11872 6349 12081 6351
rect 12115 6374 12320 6383
rect 12372 6374 12406 6393
rect 12544 6571 12590 6691
rect 12644 6687 12690 6703
rect 12841 6773 12893 6811
rect 12841 6739 12859 6773
rect 12929 6803 12995 6845
rect 13170 6843 13199 6877
rect 13233 6843 13291 6877
rect 13325 6843 13383 6877
rect 13417 6843 13446 6877
rect 13606 6862 13654 6874
rect 13868 6866 13884 6900
rect 13918 6866 13934 6900
rect 14234 6890 14284 6960
rect 15718 6934 15752 6950
rect 15814 7056 15848 7072
rect 15910 7058 15944 7072
rect 16028 7058 16248 7080
rect 15908 7056 16248 7058
rect 15908 7022 15910 7056
rect 15944 7044 16248 7056
rect 15944 7022 16064 7044
rect 15814 6986 15848 7020
rect 15909 7020 15910 7022
rect 15909 6986 15944 7020
rect 16212 6996 16248 7044
rect 15909 6985 15910 6986
rect 15814 6934 15848 6950
rect 15910 6934 15944 6950
rect 16116 6960 16248 6996
rect 17606 7056 17640 7072
rect 17606 6986 17640 7020
rect 14234 6876 14244 6890
rect 12929 6769 12945 6803
rect 12979 6769 12995 6803
rect 13031 6790 13065 6811
rect 12841 6710 12893 6739
rect 13031 6735 13065 6756
rect 12624 6619 12640 6653
rect 12674 6642 12690 6653
rect 12624 6608 12642 6619
rect 12676 6608 12690 6642
rect 12841 6638 12877 6710
rect 12932 6701 13065 6735
rect 13236 6797 13302 6809
rect 13236 6763 13252 6797
rect 13286 6763 13302 6797
rect 13236 6746 13302 6763
rect 12932 6650 12966 6701
rect 13236 6695 13252 6746
rect 13286 6695 13302 6746
rect 13236 6683 13302 6695
rect 13336 6797 13382 6843
rect 13370 6763 13382 6797
rect 13336 6729 13382 6763
rect 13370 6695 13382 6729
rect 13606 6828 13612 6862
rect 13646 6828 13654 6862
rect 14238 6856 14244 6876
rect 14278 6856 14284 6890
rect 14238 6846 14284 6856
rect 14366 6851 14395 6885
rect 14429 6851 14487 6885
rect 14521 6851 14579 6885
rect 14613 6851 14642 6885
rect 13606 6740 13654 6828
rect 13980 6785 13996 6819
rect 14030 6818 14046 6819
rect 14030 6786 14192 6818
rect 14432 6810 14498 6817
rect 14426 6805 14498 6810
rect 14426 6786 14448 6805
rect 14030 6785 14448 6786
rect 13980 6782 14448 6785
rect 14156 6771 14448 6782
rect 14482 6771 14498 6805
rect 14156 6750 14498 6771
rect 13852 6740 13886 6742
rect 13606 6723 13886 6740
rect 13606 6706 13852 6723
rect 12624 6605 12690 6608
rect 12836 6636 12877 6638
rect 12836 6602 12838 6636
rect 12872 6602 12877 6636
rect 12836 6600 12877 6602
rect 12544 6553 12610 6571
rect 12544 6519 12560 6553
rect 12594 6519 12610 6553
rect 12544 6485 12610 6519
rect 12544 6451 12560 6485
rect 12594 6451 12610 6485
rect 12544 6417 12610 6451
rect 12544 6383 12560 6417
rect 12594 6383 12610 6417
rect 12544 6375 12610 6383
rect 12644 6553 12686 6569
rect 12678 6519 12686 6553
rect 12644 6485 12686 6519
rect 12678 6451 12686 6485
rect 12644 6417 12686 6451
rect 12678 6383 12686 6417
rect 12115 6349 12154 6374
rect 11666 6297 11682 6331
rect 11716 6297 11732 6331
rect 11872 6310 12154 6349
rect 12644 6341 12686 6383
rect 12841 6550 12877 6600
rect 12911 6634 12966 6650
rect 12945 6600 12966 6634
rect 12911 6584 12966 6600
rect 13011 6648 13079 6665
rect 13011 6647 13031 6648
rect 13011 6613 13029 6647
rect 13065 6614 13079 6648
rect 13063 6613 13079 6614
rect 13011 6591 13079 6613
rect 12932 6555 12966 6584
rect 13236 6563 13282 6683
rect 13336 6679 13382 6695
rect 13554 6658 13570 6659
rect 13316 6611 13332 6645
rect 13366 6638 13382 6645
rect 13434 6638 13570 6658
rect 13366 6625 13570 6638
rect 13604 6625 13620 6659
rect 13366 6624 13620 6625
rect 13366 6611 13474 6624
rect 13554 6622 13620 6624
rect 13852 6655 13886 6657
rect 13316 6597 13474 6611
rect 13330 6596 13474 6597
rect 13852 6619 13886 6621
rect 13526 6563 13560 6582
rect 12841 6500 12895 6550
rect 12932 6521 13067 6555
rect 12841 6466 12859 6500
rect 12893 6466 12895 6500
rect 13031 6487 13067 6521
rect 12841 6419 12895 6466
rect 12841 6385 12859 6419
rect 12893 6385 12895 6419
rect 12841 6369 12895 6385
rect 12929 6453 12945 6487
rect 12979 6453 12995 6487
rect 12929 6419 12995 6453
rect 12929 6385 12945 6419
rect 12979 6385 12995 6419
rect 12040 6308 12154 6310
rect 12312 6297 12328 6331
rect 12362 6297 12378 6331
rect 12478 6307 12507 6341
rect 12541 6307 12599 6341
rect 12633 6307 12691 6341
rect 12725 6307 12754 6341
rect 12929 6335 12995 6385
rect 13065 6453 13067 6487
rect 13031 6419 13067 6453
rect 13065 6385 13067 6419
rect 13031 6369 13067 6385
rect 13236 6545 13302 6563
rect 13236 6511 13252 6545
rect 13286 6511 13302 6545
rect 13236 6477 13302 6511
rect 13236 6443 13252 6477
rect 13286 6443 13302 6477
rect 13236 6409 13302 6443
rect 13236 6375 13252 6409
rect 13286 6375 13302 6409
rect 13236 6367 13302 6375
rect 13336 6545 13378 6561
rect 13370 6511 13378 6545
rect 13336 6477 13378 6511
rect 13370 6443 13378 6477
rect 13336 6409 13378 6443
rect 13526 6495 13560 6497
rect 13526 6459 13560 6461
rect 13370 6375 13378 6409
rect 12645 6300 12679 6307
rect 12824 6301 12853 6335
rect 12887 6301 12945 6335
rect 12979 6301 13037 6335
rect 13071 6301 13100 6335
rect 13336 6333 13378 6375
rect 13486 6393 13526 6414
rect 13614 6563 13648 6582
rect 13852 6534 13886 6553
rect 13948 6723 13982 6742
rect 13948 6655 13982 6657
rect 13948 6619 13982 6621
rect 13948 6534 13982 6553
rect 14044 6723 14078 6742
rect 14432 6737 14498 6750
rect 14432 6703 14448 6737
rect 14482 6703 14498 6737
rect 14432 6691 14498 6703
rect 14532 6805 14578 6851
rect 14706 6845 14735 6879
rect 14769 6845 14827 6879
rect 14861 6845 14919 6879
rect 14953 6845 14982 6879
rect 14566 6771 14578 6805
rect 14532 6737 14578 6771
rect 14566 6703 14578 6737
rect 14044 6655 14078 6657
rect 14200 6625 14216 6659
rect 14250 6625 14266 6659
rect 14044 6619 14078 6621
rect 14044 6534 14078 6553
rect 14172 6563 14206 6582
rect 13614 6495 13648 6497
rect 14172 6495 14206 6497
rect 13614 6459 13648 6461
rect 13884 6457 13900 6491
rect 13934 6457 13950 6491
rect 14172 6459 14206 6461
rect 13560 6393 13562 6414
rect 13486 6374 13562 6393
rect 13648 6393 14172 6418
rect 14260 6563 14294 6582
rect 14260 6495 14294 6497
rect 14260 6459 14294 6461
rect 14206 6393 14208 6418
rect 13614 6385 14208 6393
rect 13614 6374 13850 6385
rect 13170 6299 13199 6333
rect 13233 6299 13291 6333
rect 13325 6299 13383 6333
rect 13417 6299 13446 6333
rect 11732 6212 11778 6218
rect 11732 6210 12220 6212
rect 11732 6176 11740 6210
rect 11774 6193 12220 6210
rect 11774 6188 12170 6193
rect 11774 6178 12049 6188
rect 11774 6176 11778 6178
rect 11732 6174 11778 6176
rect 11950 6154 12049 6178
rect 12083 6159 12170 6188
rect 12204 6168 12220 6193
rect 12204 6159 12345 6168
rect 12083 6154 12345 6159
rect 11950 6134 12345 6154
rect 12074 6050 12090 6084
rect 12124 6050 12260 6084
rect 11598 6000 11980 6016
rect 11598 5976 11946 6000
rect 11946 5930 11980 5964
rect 11946 5878 11980 5894
rect 12042 6000 12076 6016
rect 12042 5930 12076 5964
rect 12042 5878 12076 5894
rect 12138 6000 12172 6016
rect 12138 5930 12172 5964
rect 12138 5878 12172 5894
rect 10412 5797 10441 5831
rect 10475 5797 10533 5831
rect 10567 5797 10625 5831
rect 10659 5797 10688 5831
rect 11486 5797 11515 5831
rect 11549 5797 11607 5831
rect 11641 5797 11699 5831
rect 11733 5797 11762 5831
rect 11978 5810 11994 5844
rect 12028 5810 12044 5844
rect 10431 5753 10485 5797
rect 10431 5719 10451 5753
rect 10431 5685 10485 5719
rect 10431 5651 10451 5685
rect 10431 5635 10485 5651
rect 10519 5753 10585 5763
rect 10519 5719 10535 5753
rect 10569 5719 10585 5753
rect 10519 5710 10585 5719
rect 10519 5685 10537 5710
rect 10519 5651 10535 5685
rect 10571 5676 10585 5710
rect 10569 5651 10585 5676
rect 10519 5635 10585 5651
rect 10619 5753 10667 5797
rect 10653 5719 10667 5753
rect 10619 5685 10667 5719
rect 10653 5651 10667 5685
rect 10619 5635 10667 5651
rect 11505 5753 11559 5797
rect 11505 5719 11525 5753
rect 11505 5685 11559 5719
rect 11505 5651 11525 5685
rect 11505 5635 11559 5651
rect 11593 5753 11659 5763
rect 11593 5719 11609 5753
rect 11643 5719 11659 5753
rect 11593 5715 11659 5719
rect 11593 5681 11607 5715
rect 11641 5685 11659 5715
rect 11593 5651 11609 5681
rect 11643 5651 11659 5685
rect 11593 5635 11659 5651
rect 11693 5753 11741 5797
rect 11727 5719 11741 5753
rect 12090 5729 12106 5763
rect 12140 5729 12156 5763
rect 11693 5685 11741 5719
rect 11727 5651 11741 5685
rect 11693 5635 11741 5651
rect 11962 5667 11996 5686
rect 10429 5594 10449 5599
rect 10429 5560 10446 5594
rect 10483 5565 10499 5599
rect 10480 5560 10499 5565
rect 10429 5549 10499 5560
rect 10533 5515 10567 5635
rect 10601 5565 10617 5599
rect 10651 5590 10671 5599
rect 10601 5556 10619 5565
rect 10653 5556 10671 5590
rect 10601 5549 10671 5556
rect 11503 5592 11523 5599
rect 11503 5558 11521 5592
rect 11557 5565 11573 5599
rect 11555 5558 11573 5565
rect 11503 5549 11573 5558
rect 11607 5515 11641 5635
rect 11962 5599 11996 5601
rect 11675 5565 11691 5599
rect 11725 5592 11745 5599
rect 11675 5558 11695 5565
rect 11729 5558 11745 5592
rect 11675 5549 11745 5558
rect 11962 5563 11996 5565
rect 10106 5435 10372 5436
rect 10106 5401 10122 5435
rect 10156 5401 10372 5435
rect 10106 5400 10372 5401
rect 10431 5499 10497 5515
rect 10431 5465 10463 5499
rect 10533 5499 10669 5515
rect 10533 5481 10619 5499
rect 10431 5431 10497 5465
rect 9789 5363 9855 5397
rect 9789 5329 9805 5363
rect 9839 5329 9855 5363
rect 10431 5397 10463 5431
rect 10431 5363 10497 5397
rect 9789 5324 9855 5329
rect 9982 5329 10264 5362
rect 9982 5295 10072 5329
rect 10106 5327 10264 5329
rect 10106 5295 10191 5327
rect 9982 5293 10191 5295
rect 10225 5293 10264 5327
rect 9982 5287 10264 5293
rect 10431 5329 10463 5363
rect 10431 5287 10497 5329
rect 10603 5465 10619 5481
rect 10653 5465 10669 5499
rect 10603 5431 10669 5465
rect 10603 5397 10619 5431
rect 10653 5397 10669 5431
rect 10603 5363 10669 5397
rect 10603 5329 10619 5363
rect 10653 5329 10669 5363
rect 10603 5324 10669 5329
rect 11505 5499 11571 5515
rect 11505 5465 11537 5499
rect 11607 5499 11743 5515
rect 11607 5481 11693 5499
rect 11505 5431 11571 5465
rect 11505 5397 11537 5431
rect 11505 5363 11571 5397
rect 11505 5329 11537 5363
rect 11505 5287 11571 5329
rect 11677 5465 11693 5481
rect 11727 5465 11743 5499
rect 11962 5478 11996 5497
rect 12058 5667 12092 5686
rect 12058 5599 12092 5601
rect 12058 5563 12092 5565
rect 12058 5478 12092 5497
rect 12154 5667 12188 5686
rect 12154 5599 12188 5601
rect 12154 5563 12188 5565
rect 12154 5478 12188 5497
rect 11677 5431 11743 5465
rect 11677 5397 11693 5431
rect 11727 5397 11743 5431
rect 11994 5436 12060 5438
rect 12226 5436 12260 6050
rect 12311 5831 12345 6134
rect 12542 5831 12576 6042
rect 13486 6016 13520 6374
rect 13760 6351 13850 6374
rect 13884 6383 14208 6385
rect 13884 6351 13969 6383
rect 13760 6349 13969 6351
rect 14003 6374 14208 6383
rect 14260 6374 14294 6393
rect 14432 6571 14478 6691
rect 14532 6687 14578 6703
rect 14723 6773 14775 6811
rect 14723 6739 14741 6773
rect 14811 6803 14877 6845
rect 15052 6843 15081 6877
rect 15115 6843 15173 6877
rect 15207 6843 15265 6877
rect 15299 6843 15328 6877
rect 15488 6862 15536 6874
rect 15750 6866 15766 6900
rect 15800 6866 15816 6900
rect 16116 6890 16166 6960
rect 17606 6934 17640 6950
rect 17702 7056 17736 7072
rect 17798 7058 17832 7072
rect 17916 7058 18136 7080
rect 17796 7056 18136 7058
rect 17796 7022 17798 7056
rect 17832 7044 18136 7056
rect 17832 7022 17952 7044
rect 17702 6986 17736 7020
rect 17797 7020 17798 7022
rect 17797 6986 17832 7020
rect 18100 6996 18136 7044
rect 17797 6985 17798 6986
rect 17702 6934 17736 6950
rect 17798 6934 17832 6950
rect 18004 6960 18136 6996
rect 19494 7056 19528 7072
rect 19494 6986 19528 7020
rect 16116 6876 16126 6890
rect 14811 6769 14827 6803
rect 14861 6769 14877 6803
rect 14913 6790 14947 6811
rect 14723 6710 14775 6739
rect 14913 6735 14947 6756
rect 14512 6619 14528 6653
rect 14562 6642 14578 6653
rect 14512 6608 14530 6619
rect 14564 6608 14578 6642
rect 14723 6638 14759 6710
rect 14814 6701 14947 6735
rect 15118 6797 15184 6809
rect 15118 6763 15134 6797
rect 15168 6763 15184 6797
rect 15118 6746 15184 6763
rect 14814 6650 14848 6701
rect 15118 6695 15134 6746
rect 15168 6695 15184 6746
rect 15118 6683 15184 6695
rect 15218 6797 15264 6843
rect 15252 6763 15264 6797
rect 15218 6729 15264 6763
rect 15252 6695 15264 6729
rect 15488 6828 15494 6862
rect 15528 6828 15536 6862
rect 16120 6856 16126 6876
rect 16160 6856 16166 6890
rect 16120 6846 16166 6856
rect 16248 6851 16277 6885
rect 16311 6851 16369 6885
rect 16403 6851 16461 6885
rect 16495 6851 16524 6885
rect 15488 6740 15536 6828
rect 15862 6785 15878 6819
rect 15912 6818 15928 6819
rect 15912 6786 16074 6818
rect 16314 6810 16380 6817
rect 16308 6805 16380 6810
rect 16308 6786 16330 6805
rect 15912 6785 16330 6786
rect 15862 6782 16330 6785
rect 16038 6771 16330 6782
rect 16364 6771 16380 6805
rect 16038 6750 16380 6771
rect 15734 6740 15768 6742
rect 15488 6723 15768 6740
rect 15488 6706 15734 6723
rect 14512 6605 14578 6608
rect 14718 6636 14759 6638
rect 14718 6602 14720 6636
rect 14754 6602 14759 6636
rect 14718 6600 14759 6602
rect 14432 6553 14498 6571
rect 14432 6519 14448 6553
rect 14482 6519 14498 6553
rect 14432 6485 14498 6519
rect 14432 6451 14448 6485
rect 14482 6451 14498 6485
rect 14432 6417 14498 6451
rect 14432 6383 14448 6417
rect 14482 6383 14498 6417
rect 14432 6375 14498 6383
rect 14532 6553 14574 6569
rect 14566 6519 14574 6553
rect 14532 6485 14574 6519
rect 14566 6451 14574 6485
rect 14532 6417 14574 6451
rect 14566 6383 14574 6417
rect 14003 6349 14042 6374
rect 13554 6297 13570 6331
rect 13604 6297 13620 6331
rect 13760 6310 14042 6349
rect 14532 6341 14574 6383
rect 14723 6550 14759 6600
rect 14793 6634 14848 6650
rect 14827 6600 14848 6634
rect 14793 6584 14848 6600
rect 14893 6648 14961 6665
rect 14893 6647 14913 6648
rect 14893 6613 14911 6647
rect 14947 6614 14961 6648
rect 14945 6613 14961 6614
rect 14893 6591 14961 6613
rect 14814 6555 14848 6584
rect 15118 6563 15164 6683
rect 15218 6679 15264 6695
rect 15436 6658 15452 6659
rect 15198 6611 15214 6645
rect 15248 6638 15264 6645
rect 15316 6638 15452 6658
rect 15248 6625 15452 6638
rect 15486 6625 15502 6659
rect 15248 6624 15502 6625
rect 15248 6611 15356 6624
rect 15436 6622 15502 6624
rect 15734 6655 15768 6657
rect 15198 6597 15356 6611
rect 15212 6596 15356 6597
rect 15734 6619 15768 6621
rect 15408 6563 15442 6582
rect 14723 6500 14777 6550
rect 14814 6521 14949 6555
rect 14723 6466 14741 6500
rect 14775 6466 14777 6500
rect 14913 6487 14949 6521
rect 14723 6419 14777 6466
rect 14723 6385 14741 6419
rect 14775 6385 14777 6419
rect 14723 6369 14777 6385
rect 14811 6453 14827 6487
rect 14861 6453 14877 6487
rect 14811 6419 14877 6453
rect 14811 6385 14827 6419
rect 14861 6385 14877 6419
rect 13928 6308 14042 6310
rect 14200 6297 14216 6331
rect 14250 6297 14266 6331
rect 14366 6307 14395 6341
rect 14429 6307 14487 6341
rect 14521 6307 14579 6341
rect 14613 6307 14642 6341
rect 14811 6335 14877 6385
rect 14947 6453 14949 6487
rect 14913 6419 14949 6453
rect 14947 6385 14949 6419
rect 14913 6369 14949 6385
rect 15118 6545 15184 6563
rect 15118 6511 15134 6545
rect 15168 6511 15184 6545
rect 15118 6477 15184 6511
rect 15118 6443 15134 6477
rect 15168 6443 15184 6477
rect 15118 6409 15184 6443
rect 15118 6375 15134 6409
rect 15168 6375 15184 6409
rect 15118 6367 15184 6375
rect 15218 6545 15260 6561
rect 15252 6511 15260 6545
rect 15218 6477 15260 6511
rect 15252 6443 15260 6477
rect 15218 6409 15260 6443
rect 15408 6495 15442 6497
rect 15408 6459 15442 6461
rect 15252 6375 15260 6409
rect 14533 6300 14567 6307
rect 14706 6301 14735 6335
rect 14769 6301 14827 6335
rect 14861 6301 14919 6335
rect 14953 6301 14982 6335
rect 15218 6333 15260 6375
rect 15368 6393 15408 6414
rect 15496 6563 15530 6582
rect 15734 6534 15768 6553
rect 15830 6723 15864 6742
rect 15830 6655 15864 6657
rect 15830 6619 15864 6621
rect 15830 6534 15864 6553
rect 15926 6723 15960 6742
rect 16314 6737 16380 6750
rect 16314 6703 16330 6737
rect 16364 6703 16380 6737
rect 16314 6691 16380 6703
rect 16414 6805 16460 6851
rect 16594 6845 16623 6879
rect 16657 6845 16715 6879
rect 16749 6845 16807 6879
rect 16841 6845 16870 6879
rect 16448 6771 16460 6805
rect 16414 6737 16460 6771
rect 16448 6703 16460 6737
rect 15926 6655 15960 6657
rect 16082 6625 16098 6659
rect 16132 6625 16148 6659
rect 15926 6619 15960 6621
rect 15926 6534 15960 6553
rect 16054 6563 16088 6582
rect 15496 6495 15530 6497
rect 16054 6495 16088 6497
rect 15496 6459 15530 6461
rect 15766 6457 15782 6491
rect 15816 6457 15832 6491
rect 16054 6459 16088 6461
rect 15442 6393 15444 6414
rect 15368 6374 15444 6393
rect 15530 6393 16054 6418
rect 16142 6563 16176 6582
rect 16142 6495 16176 6497
rect 16142 6459 16176 6461
rect 16088 6393 16090 6418
rect 15496 6385 16090 6393
rect 15496 6374 15732 6385
rect 15052 6299 15081 6333
rect 15115 6299 15173 6333
rect 15207 6299 15265 6333
rect 15299 6299 15328 6333
rect 13620 6212 13666 6218
rect 13620 6210 14108 6212
rect 13620 6176 13628 6210
rect 13662 6193 14108 6210
rect 13662 6188 14058 6193
rect 13662 6178 13937 6188
rect 13662 6176 13666 6178
rect 13620 6174 13666 6176
rect 13838 6154 13937 6178
rect 13971 6159 14058 6188
rect 14092 6168 14108 6193
rect 14092 6159 14233 6168
rect 13971 6154 14233 6159
rect 13838 6134 14233 6154
rect 13962 6050 13978 6084
rect 14012 6050 14148 6084
rect 13486 6000 13868 6016
rect 13486 5976 13834 6000
rect 13834 5930 13868 5964
rect 13834 5878 13868 5894
rect 13930 6000 13964 6016
rect 13930 5930 13964 5964
rect 13930 5878 13964 5894
rect 14026 6000 14060 6016
rect 14026 5930 14060 5964
rect 14026 5878 14060 5894
rect 12300 5797 12329 5831
rect 12363 5797 12421 5831
rect 12455 5797 12513 5831
rect 12547 5797 12576 5831
rect 13374 5797 13403 5831
rect 13437 5797 13495 5831
rect 13529 5797 13587 5831
rect 13621 5797 13650 5831
rect 13866 5810 13882 5844
rect 13916 5810 13932 5844
rect 12319 5753 12373 5797
rect 12319 5719 12339 5753
rect 12319 5685 12373 5719
rect 12319 5651 12339 5685
rect 12319 5635 12373 5651
rect 12407 5753 12473 5763
rect 12407 5719 12423 5753
rect 12457 5719 12473 5753
rect 12407 5710 12473 5719
rect 12407 5685 12425 5710
rect 12407 5651 12423 5685
rect 12459 5676 12473 5710
rect 12457 5651 12473 5676
rect 12407 5635 12473 5651
rect 12507 5753 12555 5797
rect 12541 5719 12555 5753
rect 12507 5685 12555 5719
rect 12541 5651 12555 5685
rect 12507 5635 12555 5651
rect 13393 5753 13447 5797
rect 13393 5719 13413 5753
rect 13393 5685 13447 5719
rect 13393 5651 13413 5685
rect 13393 5635 13447 5651
rect 13481 5753 13547 5763
rect 13481 5719 13497 5753
rect 13531 5719 13547 5753
rect 13481 5715 13547 5719
rect 13481 5681 13495 5715
rect 13529 5685 13547 5715
rect 13481 5651 13497 5681
rect 13531 5651 13547 5685
rect 13481 5635 13547 5651
rect 13581 5753 13629 5797
rect 13615 5719 13629 5753
rect 13978 5729 13994 5763
rect 14028 5729 14044 5763
rect 13581 5685 13629 5719
rect 13615 5651 13629 5685
rect 13581 5635 13629 5651
rect 13850 5667 13884 5686
rect 12317 5594 12337 5599
rect 12317 5560 12334 5594
rect 12371 5565 12387 5599
rect 12368 5560 12387 5565
rect 12317 5549 12387 5560
rect 12421 5515 12455 5635
rect 12489 5565 12505 5599
rect 12539 5590 12559 5599
rect 12489 5556 12507 5565
rect 12541 5556 12559 5590
rect 12489 5549 12559 5556
rect 13391 5592 13411 5599
rect 13391 5558 13409 5592
rect 13445 5565 13461 5599
rect 13443 5558 13461 5565
rect 13391 5549 13461 5558
rect 13495 5515 13529 5635
rect 13850 5599 13884 5601
rect 13563 5565 13579 5599
rect 13613 5592 13633 5599
rect 13563 5558 13583 5565
rect 13617 5558 13633 5592
rect 13563 5549 13633 5558
rect 13850 5563 13884 5565
rect 11994 5435 12260 5436
rect 11994 5401 12010 5435
rect 12044 5401 12260 5435
rect 11994 5400 12260 5401
rect 12319 5499 12385 5515
rect 12319 5465 12351 5499
rect 12421 5499 12557 5515
rect 12421 5481 12507 5499
rect 12319 5431 12385 5465
rect 11677 5363 11743 5397
rect 11677 5329 11693 5363
rect 11727 5329 11743 5363
rect 12319 5397 12351 5431
rect 12319 5363 12385 5397
rect 11677 5324 11743 5329
rect 11870 5329 12152 5362
rect 11870 5295 11960 5329
rect 11994 5327 12152 5329
rect 11994 5295 12079 5327
rect 11870 5293 12079 5295
rect 12113 5293 12152 5327
rect 11870 5287 12152 5293
rect 12319 5329 12351 5363
rect 12319 5287 12385 5329
rect 12491 5465 12507 5481
rect 12541 5465 12557 5499
rect 12491 5431 12557 5465
rect 12491 5397 12507 5431
rect 12541 5397 12557 5431
rect 12491 5363 12557 5397
rect 12491 5329 12507 5363
rect 12541 5329 12557 5363
rect 12491 5324 12557 5329
rect 13393 5499 13459 5515
rect 13393 5465 13425 5499
rect 13495 5499 13631 5515
rect 13495 5481 13581 5499
rect 13393 5431 13459 5465
rect 13393 5397 13425 5431
rect 13393 5363 13459 5397
rect 13393 5329 13425 5363
rect 13393 5287 13459 5329
rect 13565 5465 13581 5481
rect 13615 5465 13631 5499
rect 13850 5478 13884 5497
rect 13946 5667 13980 5686
rect 13946 5599 13980 5601
rect 13946 5563 13980 5565
rect 13946 5478 13980 5497
rect 14042 5667 14076 5686
rect 14042 5599 14076 5601
rect 14042 5563 14076 5565
rect 14042 5478 14076 5497
rect 13565 5431 13631 5465
rect 13565 5397 13581 5431
rect 13615 5397 13631 5431
rect 13882 5436 13948 5438
rect 14114 5436 14148 6050
rect 14199 5831 14233 6134
rect 14430 5831 14464 6042
rect 15368 6016 15402 6374
rect 15642 6351 15732 6374
rect 15766 6383 16090 6385
rect 15766 6351 15851 6383
rect 15642 6349 15851 6351
rect 15885 6374 16090 6383
rect 16142 6374 16176 6393
rect 16314 6571 16360 6691
rect 16414 6687 16460 6703
rect 16611 6773 16663 6811
rect 16611 6739 16629 6773
rect 16699 6803 16765 6845
rect 16940 6843 16969 6877
rect 17003 6843 17061 6877
rect 17095 6843 17153 6877
rect 17187 6843 17216 6877
rect 17376 6862 17424 6874
rect 17638 6866 17654 6900
rect 17688 6866 17704 6900
rect 18004 6890 18054 6960
rect 19494 6934 19528 6950
rect 19590 7056 19624 7072
rect 19686 7058 19720 7072
rect 19804 7058 20024 7080
rect 19684 7056 20024 7058
rect 19684 7022 19686 7056
rect 19720 7044 20024 7056
rect 19720 7022 19840 7044
rect 19590 6986 19624 7020
rect 19685 7020 19686 7022
rect 19685 6986 19720 7020
rect 19988 6996 20024 7044
rect 19685 6985 19686 6986
rect 19590 6934 19624 6950
rect 19686 6934 19720 6950
rect 19892 6960 20024 6996
rect 21382 7056 21416 7072
rect 21382 6986 21416 7020
rect 18004 6876 18014 6890
rect 16699 6769 16715 6803
rect 16749 6769 16765 6803
rect 16801 6790 16835 6811
rect 16611 6710 16663 6739
rect 16801 6735 16835 6756
rect 16394 6619 16410 6653
rect 16444 6642 16460 6653
rect 16394 6608 16412 6619
rect 16446 6608 16460 6642
rect 16611 6638 16647 6710
rect 16702 6701 16835 6735
rect 17006 6797 17072 6809
rect 17006 6763 17022 6797
rect 17056 6763 17072 6797
rect 17006 6746 17072 6763
rect 16702 6650 16736 6701
rect 17006 6695 17022 6746
rect 17056 6695 17072 6746
rect 17006 6683 17072 6695
rect 17106 6797 17152 6843
rect 17140 6763 17152 6797
rect 17106 6729 17152 6763
rect 17140 6695 17152 6729
rect 17376 6828 17382 6862
rect 17416 6828 17424 6862
rect 18008 6856 18014 6876
rect 18048 6856 18054 6890
rect 18008 6846 18054 6856
rect 18136 6851 18165 6885
rect 18199 6851 18257 6885
rect 18291 6851 18349 6885
rect 18383 6851 18412 6885
rect 17376 6740 17424 6828
rect 17750 6785 17766 6819
rect 17800 6818 17816 6819
rect 17800 6786 17962 6818
rect 18202 6810 18268 6817
rect 18196 6805 18268 6810
rect 18196 6786 18218 6805
rect 17800 6785 18218 6786
rect 17750 6782 18218 6785
rect 17926 6771 18218 6782
rect 18252 6771 18268 6805
rect 17926 6750 18268 6771
rect 17622 6740 17656 6742
rect 17376 6723 17656 6740
rect 17376 6706 17622 6723
rect 16394 6605 16460 6608
rect 16606 6636 16647 6638
rect 16606 6602 16608 6636
rect 16642 6602 16647 6636
rect 16606 6600 16647 6602
rect 16314 6553 16380 6571
rect 16314 6519 16330 6553
rect 16364 6519 16380 6553
rect 16314 6485 16380 6519
rect 16314 6451 16330 6485
rect 16364 6451 16380 6485
rect 16314 6417 16380 6451
rect 16314 6383 16330 6417
rect 16364 6383 16380 6417
rect 16314 6375 16380 6383
rect 16414 6553 16456 6569
rect 16448 6519 16456 6553
rect 16414 6485 16456 6519
rect 16448 6451 16456 6485
rect 16414 6417 16456 6451
rect 16448 6383 16456 6417
rect 15885 6349 15924 6374
rect 15436 6297 15452 6331
rect 15486 6297 15502 6331
rect 15642 6310 15924 6349
rect 16414 6341 16456 6383
rect 16611 6550 16647 6600
rect 16681 6634 16736 6650
rect 16715 6600 16736 6634
rect 16681 6584 16736 6600
rect 16781 6648 16849 6665
rect 16781 6647 16801 6648
rect 16781 6613 16799 6647
rect 16835 6614 16849 6648
rect 16833 6613 16849 6614
rect 16781 6591 16849 6613
rect 16702 6555 16736 6584
rect 17006 6563 17052 6683
rect 17106 6679 17152 6695
rect 17324 6658 17340 6659
rect 17086 6611 17102 6645
rect 17136 6638 17152 6645
rect 17204 6638 17340 6658
rect 17136 6625 17340 6638
rect 17374 6625 17390 6659
rect 17136 6624 17390 6625
rect 17136 6611 17244 6624
rect 17324 6622 17390 6624
rect 17622 6655 17656 6657
rect 17086 6597 17244 6611
rect 17100 6596 17244 6597
rect 17622 6619 17656 6621
rect 17296 6563 17330 6582
rect 16611 6500 16665 6550
rect 16702 6521 16837 6555
rect 16611 6466 16629 6500
rect 16663 6466 16665 6500
rect 16801 6487 16837 6521
rect 16611 6419 16665 6466
rect 16611 6385 16629 6419
rect 16663 6385 16665 6419
rect 16611 6369 16665 6385
rect 16699 6453 16715 6487
rect 16749 6453 16765 6487
rect 16699 6419 16765 6453
rect 16699 6385 16715 6419
rect 16749 6385 16765 6419
rect 15810 6308 15924 6310
rect 16082 6297 16098 6331
rect 16132 6297 16148 6331
rect 16248 6307 16277 6341
rect 16311 6307 16369 6341
rect 16403 6307 16461 6341
rect 16495 6307 16524 6341
rect 16699 6335 16765 6385
rect 16835 6453 16837 6487
rect 16801 6419 16837 6453
rect 16835 6385 16837 6419
rect 16801 6369 16837 6385
rect 17006 6545 17072 6563
rect 17006 6511 17022 6545
rect 17056 6511 17072 6545
rect 17006 6477 17072 6511
rect 17006 6443 17022 6477
rect 17056 6443 17072 6477
rect 17006 6409 17072 6443
rect 17006 6375 17022 6409
rect 17056 6375 17072 6409
rect 17006 6367 17072 6375
rect 17106 6545 17148 6561
rect 17140 6511 17148 6545
rect 17106 6477 17148 6511
rect 17140 6443 17148 6477
rect 17106 6409 17148 6443
rect 17296 6495 17330 6497
rect 17296 6459 17330 6461
rect 17140 6375 17148 6409
rect 16415 6300 16449 6307
rect 16594 6301 16623 6335
rect 16657 6301 16715 6335
rect 16749 6301 16807 6335
rect 16841 6301 16870 6335
rect 17106 6333 17148 6375
rect 17256 6393 17296 6414
rect 17384 6563 17418 6582
rect 17622 6534 17656 6553
rect 17718 6723 17752 6742
rect 17718 6655 17752 6657
rect 17718 6619 17752 6621
rect 17718 6534 17752 6553
rect 17814 6723 17848 6742
rect 18202 6737 18268 6750
rect 18202 6703 18218 6737
rect 18252 6703 18268 6737
rect 18202 6691 18268 6703
rect 18302 6805 18348 6851
rect 18482 6845 18511 6879
rect 18545 6845 18603 6879
rect 18637 6845 18695 6879
rect 18729 6845 18758 6879
rect 18336 6771 18348 6805
rect 18302 6737 18348 6771
rect 18336 6703 18348 6737
rect 17814 6655 17848 6657
rect 17970 6625 17986 6659
rect 18020 6625 18036 6659
rect 17814 6619 17848 6621
rect 17814 6534 17848 6553
rect 17942 6563 17976 6582
rect 17384 6495 17418 6497
rect 17942 6495 17976 6497
rect 17384 6459 17418 6461
rect 17654 6457 17670 6491
rect 17704 6457 17720 6491
rect 17942 6459 17976 6461
rect 17330 6393 17332 6414
rect 17256 6374 17332 6393
rect 17418 6393 17942 6418
rect 18030 6563 18064 6582
rect 18030 6495 18064 6497
rect 18030 6459 18064 6461
rect 17976 6393 17978 6418
rect 17384 6385 17978 6393
rect 17384 6374 17620 6385
rect 16940 6299 16969 6333
rect 17003 6299 17061 6333
rect 17095 6299 17153 6333
rect 17187 6299 17216 6333
rect 15502 6212 15548 6218
rect 15502 6210 15990 6212
rect 15502 6176 15510 6210
rect 15544 6193 15990 6210
rect 15544 6188 15940 6193
rect 15544 6178 15819 6188
rect 15544 6176 15548 6178
rect 15502 6174 15548 6176
rect 15720 6154 15819 6178
rect 15853 6159 15940 6188
rect 15974 6168 15990 6193
rect 15974 6159 16115 6168
rect 15853 6154 16115 6159
rect 15720 6134 16115 6154
rect 15844 6050 15860 6084
rect 15894 6050 16030 6084
rect 15368 6000 15750 6016
rect 15368 5976 15716 6000
rect 15716 5930 15750 5964
rect 15716 5878 15750 5894
rect 15812 6000 15846 6016
rect 15812 5930 15846 5964
rect 15812 5878 15846 5894
rect 15908 6000 15942 6016
rect 15908 5930 15942 5964
rect 15908 5878 15942 5894
rect 14188 5797 14217 5831
rect 14251 5797 14309 5831
rect 14343 5797 14401 5831
rect 14435 5797 14464 5831
rect 15256 5797 15285 5831
rect 15319 5797 15377 5831
rect 15411 5797 15469 5831
rect 15503 5797 15532 5831
rect 15748 5810 15764 5844
rect 15798 5810 15814 5844
rect 14207 5753 14261 5797
rect 14207 5719 14227 5753
rect 14207 5685 14261 5719
rect 14207 5651 14227 5685
rect 14207 5635 14261 5651
rect 14295 5753 14361 5763
rect 14295 5719 14311 5753
rect 14345 5719 14361 5753
rect 14295 5710 14361 5719
rect 14295 5685 14313 5710
rect 14295 5651 14311 5685
rect 14347 5676 14361 5710
rect 14345 5651 14361 5676
rect 14295 5635 14361 5651
rect 14395 5753 14443 5797
rect 14429 5719 14443 5753
rect 14395 5685 14443 5719
rect 14429 5651 14443 5685
rect 14395 5635 14443 5651
rect 15275 5753 15329 5797
rect 15275 5719 15295 5753
rect 15275 5685 15329 5719
rect 15275 5651 15295 5685
rect 15275 5635 15329 5651
rect 15363 5753 15429 5763
rect 15363 5719 15379 5753
rect 15413 5719 15429 5753
rect 15363 5715 15429 5719
rect 15363 5681 15377 5715
rect 15411 5685 15429 5715
rect 15363 5651 15379 5681
rect 15413 5651 15429 5685
rect 15363 5635 15429 5651
rect 15463 5753 15511 5797
rect 15497 5719 15511 5753
rect 15860 5729 15876 5763
rect 15910 5729 15926 5763
rect 15463 5685 15511 5719
rect 15497 5651 15511 5685
rect 15463 5635 15511 5651
rect 15732 5667 15766 5686
rect 14205 5594 14225 5599
rect 14205 5560 14222 5594
rect 14259 5565 14275 5599
rect 14256 5560 14275 5565
rect 14205 5549 14275 5560
rect 14309 5515 14343 5635
rect 14377 5565 14393 5599
rect 14427 5590 14447 5599
rect 14377 5556 14395 5565
rect 14429 5556 14447 5590
rect 14377 5549 14447 5556
rect 15273 5592 15293 5599
rect 15273 5558 15291 5592
rect 15327 5565 15343 5599
rect 15325 5558 15343 5565
rect 15273 5549 15343 5558
rect 15377 5515 15411 5635
rect 15732 5599 15766 5601
rect 15445 5565 15461 5599
rect 15495 5592 15515 5599
rect 15445 5558 15465 5565
rect 15499 5558 15515 5592
rect 15445 5549 15515 5558
rect 15732 5563 15766 5565
rect 13882 5435 14148 5436
rect 13882 5401 13898 5435
rect 13932 5401 14148 5435
rect 13882 5400 14148 5401
rect 14207 5499 14273 5515
rect 14207 5465 14239 5499
rect 14309 5499 14445 5515
rect 14309 5481 14395 5499
rect 14207 5431 14273 5465
rect 13565 5363 13631 5397
rect 13565 5329 13581 5363
rect 13615 5329 13631 5363
rect 14207 5397 14239 5431
rect 14207 5363 14273 5397
rect 13565 5324 13631 5329
rect 13758 5329 14040 5362
rect 13758 5295 13848 5329
rect 13882 5327 14040 5329
rect 13882 5295 13967 5327
rect 13758 5293 13967 5295
rect 14001 5293 14040 5327
rect 13758 5287 14040 5293
rect 14207 5329 14239 5363
rect 14207 5287 14273 5329
rect 14379 5465 14395 5481
rect 14429 5465 14445 5499
rect 14379 5431 14445 5465
rect 14379 5397 14395 5431
rect 14429 5397 14445 5431
rect 14379 5363 14445 5397
rect 14379 5329 14395 5363
rect 14429 5329 14445 5363
rect 14379 5324 14445 5329
rect 15275 5499 15341 5515
rect 15275 5465 15307 5499
rect 15377 5499 15513 5515
rect 15377 5481 15463 5499
rect 15275 5431 15341 5465
rect 15275 5397 15307 5431
rect 15275 5363 15341 5397
rect 15275 5329 15307 5363
rect 15275 5287 15341 5329
rect 15447 5465 15463 5481
rect 15497 5465 15513 5499
rect 15732 5478 15766 5497
rect 15828 5667 15862 5686
rect 15828 5599 15862 5601
rect 15828 5563 15862 5565
rect 15828 5478 15862 5497
rect 15924 5667 15958 5686
rect 15924 5599 15958 5601
rect 15924 5563 15958 5565
rect 15924 5478 15958 5497
rect 15447 5431 15513 5465
rect 15447 5397 15463 5431
rect 15497 5397 15513 5431
rect 15764 5436 15830 5438
rect 15996 5436 16030 6050
rect 16081 5831 16115 6134
rect 16312 5831 16346 6042
rect 17256 6016 17290 6374
rect 17530 6351 17620 6374
rect 17654 6383 17978 6385
rect 17654 6351 17739 6383
rect 17530 6349 17739 6351
rect 17773 6374 17978 6383
rect 18030 6374 18064 6393
rect 18202 6571 18248 6691
rect 18302 6687 18348 6703
rect 18499 6773 18551 6811
rect 18499 6739 18517 6773
rect 18587 6803 18653 6845
rect 18828 6843 18857 6877
rect 18891 6843 18949 6877
rect 18983 6843 19041 6877
rect 19075 6843 19104 6877
rect 19264 6862 19312 6874
rect 19526 6866 19542 6900
rect 19576 6866 19592 6900
rect 19892 6890 19942 6960
rect 21382 6934 21416 6950
rect 21478 7056 21512 7072
rect 21574 7058 21608 7072
rect 21692 7058 21912 7080
rect 21572 7056 21912 7058
rect 21572 7022 21574 7056
rect 21608 7044 21912 7056
rect 21608 7022 21728 7044
rect 21478 6986 21512 7020
rect 21573 7020 21574 7022
rect 21573 6986 21608 7020
rect 21876 6996 21912 7044
rect 21573 6985 21574 6986
rect 21478 6934 21512 6950
rect 21574 6934 21608 6950
rect 21780 6960 21912 6996
rect 23270 7056 23304 7072
rect 23270 6986 23304 7020
rect 19892 6876 19902 6890
rect 18587 6769 18603 6803
rect 18637 6769 18653 6803
rect 18689 6790 18723 6811
rect 18499 6710 18551 6739
rect 18689 6735 18723 6756
rect 18282 6619 18298 6653
rect 18332 6642 18348 6653
rect 18282 6608 18300 6619
rect 18334 6608 18348 6642
rect 18499 6638 18535 6710
rect 18590 6701 18723 6735
rect 18894 6797 18960 6809
rect 18894 6763 18910 6797
rect 18944 6763 18960 6797
rect 18894 6746 18960 6763
rect 18590 6650 18624 6701
rect 18894 6695 18910 6746
rect 18944 6695 18960 6746
rect 18894 6683 18960 6695
rect 18994 6797 19040 6843
rect 19028 6763 19040 6797
rect 18994 6729 19040 6763
rect 19028 6695 19040 6729
rect 19264 6828 19270 6862
rect 19304 6828 19312 6862
rect 19896 6856 19902 6876
rect 19936 6856 19942 6890
rect 19896 6846 19942 6856
rect 20024 6851 20053 6885
rect 20087 6851 20145 6885
rect 20179 6851 20237 6885
rect 20271 6851 20300 6885
rect 19264 6740 19312 6828
rect 19638 6785 19654 6819
rect 19688 6818 19704 6819
rect 19688 6786 19850 6818
rect 20090 6810 20156 6817
rect 20084 6805 20156 6810
rect 20084 6786 20106 6805
rect 19688 6785 20106 6786
rect 19638 6782 20106 6785
rect 19814 6771 20106 6782
rect 20140 6771 20156 6805
rect 19814 6750 20156 6771
rect 19510 6740 19544 6742
rect 19264 6723 19544 6740
rect 19264 6706 19510 6723
rect 18282 6605 18348 6608
rect 18494 6636 18535 6638
rect 18494 6602 18496 6636
rect 18530 6602 18535 6636
rect 18494 6600 18535 6602
rect 18202 6553 18268 6571
rect 18202 6519 18218 6553
rect 18252 6519 18268 6553
rect 18202 6485 18268 6519
rect 18202 6451 18218 6485
rect 18252 6451 18268 6485
rect 18202 6417 18268 6451
rect 18202 6383 18218 6417
rect 18252 6383 18268 6417
rect 18202 6375 18268 6383
rect 18302 6553 18344 6569
rect 18336 6519 18344 6553
rect 18302 6485 18344 6519
rect 18336 6451 18344 6485
rect 18302 6417 18344 6451
rect 18336 6383 18344 6417
rect 17773 6349 17812 6374
rect 17324 6297 17340 6331
rect 17374 6297 17390 6331
rect 17530 6310 17812 6349
rect 18302 6341 18344 6383
rect 18499 6550 18535 6600
rect 18569 6634 18624 6650
rect 18603 6600 18624 6634
rect 18569 6584 18624 6600
rect 18669 6648 18737 6665
rect 18669 6647 18689 6648
rect 18669 6613 18687 6647
rect 18723 6614 18737 6648
rect 18721 6613 18737 6614
rect 18669 6591 18737 6613
rect 18590 6555 18624 6584
rect 18894 6563 18940 6683
rect 18994 6679 19040 6695
rect 19212 6658 19228 6659
rect 18974 6611 18990 6645
rect 19024 6638 19040 6645
rect 19092 6638 19228 6658
rect 19024 6625 19228 6638
rect 19262 6625 19278 6659
rect 19024 6624 19278 6625
rect 19024 6611 19132 6624
rect 19212 6622 19278 6624
rect 19510 6655 19544 6657
rect 18974 6597 19132 6611
rect 18988 6596 19132 6597
rect 19510 6619 19544 6621
rect 19184 6563 19218 6582
rect 18499 6500 18553 6550
rect 18590 6521 18725 6555
rect 18499 6466 18517 6500
rect 18551 6466 18553 6500
rect 18689 6487 18725 6521
rect 18499 6419 18553 6466
rect 18499 6385 18517 6419
rect 18551 6385 18553 6419
rect 18499 6369 18553 6385
rect 18587 6453 18603 6487
rect 18637 6453 18653 6487
rect 18587 6419 18653 6453
rect 18587 6385 18603 6419
rect 18637 6385 18653 6419
rect 17698 6308 17812 6310
rect 17970 6297 17986 6331
rect 18020 6297 18036 6331
rect 18136 6307 18165 6341
rect 18199 6307 18257 6341
rect 18291 6307 18349 6341
rect 18383 6307 18412 6341
rect 18587 6335 18653 6385
rect 18723 6453 18725 6487
rect 18689 6419 18725 6453
rect 18723 6385 18725 6419
rect 18689 6369 18725 6385
rect 18894 6545 18960 6563
rect 18894 6511 18910 6545
rect 18944 6511 18960 6545
rect 18894 6477 18960 6511
rect 18894 6443 18910 6477
rect 18944 6443 18960 6477
rect 18894 6409 18960 6443
rect 18894 6375 18910 6409
rect 18944 6375 18960 6409
rect 18894 6367 18960 6375
rect 18994 6545 19036 6561
rect 19028 6511 19036 6545
rect 18994 6477 19036 6511
rect 19028 6443 19036 6477
rect 18994 6409 19036 6443
rect 19184 6495 19218 6497
rect 19184 6459 19218 6461
rect 19028 6375 19036 6409
rect 18303 6300 18337 6307
rect 18482 6301 18511 6335
rect 18545 6301 18603 6335
rect 18637 6301 18695 6335
rect 18729 6301 18758 6335
rect 18994 6333 19036 6375
rect 19144 6393 19184 6414
rect 19272 6563 19306 6582
rect 19510 6534 19544 6553
rect 19606 6723 19640 6742
rect 19606 6655 19640 6657
rect 19606 6619 19640 6621
rect 19606 6534 19640 6553
rect 19702 6723 19736 6742
rect 20090 6737 20156 6750
rect 20090 6703 20106 6737
rect 20140 6703 20156 6737
rect 20090 6691 20156 6703
rect 20190 6805 20236 6851
rect 20370 6845 20399 6879
rect 20433 6845 20491 6879
rect 20525 6845 20583 6879
rect 20617 6845 20646 6879
rect 20224 6771 20236 6805
rect 20190 6737 20236 6771
rect 20224 6703 20236 6737
rect 19702 6655 19736 6657
rect 19858 6625 19874 6659
rect 19908 6625 19924 6659
rect 19702 6619 19736 6621
rect 19702 6534 19736 6553
rect 19830 6563 19864 6582
rect 19272 6495 19306 6497
rect 19830 6495 19864 6497
rect 19272 6459 19306 6461
rect 19542 6457 19558 6491
rect 19592 6457 19608 6491
rect 19830 6459 19864 6461
rect 19218 6393 19220 6414
rect 19144 6374 19220 6393
rect 19306 6393 19830 6418
rect 19918 6563 19952 6582
rect 19918 6495 19952 6497
rect 19918 6459 19952 6461
rect 19864 6393 19866 6418
rect 19272 6385 19866 6393
rect 19272 6374 19508 6385
rect 18828 6299 18857 6333
rect 18891 6299 18949 6333
rect 18983 6299 19041 6333
rect 19075 6299 19104 6333
rect 17390 6212 17436 6218
rect 17390 6210 17878 6212
rect 17390 6176 17398 6210
rect 17432 6193 17878 6210
rect 17432 6188 17828 6193
rect 17432 6178 17707 6188
rect 17432 6176 17436 6178
rect 17390 6174 17436 6176
rect 17608 6154 17707 6178
rect 17741 6159 17828 6188
rect 17862 6168 17878 6193
rect 17862 6159 18003 6168
rect 17741 6154 18003 6159
rect 17608 6134 18003 6154
rect 17732 6050 17748 6084
rect 17782 6050 17918 6084
rect 17256 6000 17638 6016
rect 17256 5976 17604 6000
rect 17604 5930 17638 5964
rect 17604 5878 17638 5894
rect 17700 6000 17734 6016
rect 17700 5930 17734 5964
rect 17700 5878 17734 5894
rect 17796 6000 17830 6016
rect 17796 5930 17830 5964
rect 17796 5878 17830 5894
rect 16070 5797 16099 5831
rect 16133 5797 16191 5831
rect 16225 5797 16283 5831
rect 16317 5797 16346 5831
rect 17144 5797 17173 5831
rect 17207 5797 17265 5831
rect 17299 5797 17357 5831
rect 17391 5797 17420 5831
rect 17636 5810 17652 5844
rect 17686 5810 17702 5844
rect 16089 5753 16143 5797
rect 16089 5719 16109 5753
rect 16089 5685 16143 5719
rect 16089 5651 16109 5685
rect 16089 5635 16143 5651
rect 16177 5753 16243 5763
rect 16177 5719 16193 5753
rect 16227 5719 16243 5753
rect 16177 5710 16243 5719
rect 16177 5685 16195 5710
rect 16177 5651 16193 5685
rect 16229 5676 16243 5710
rect 16227 5651 16243 5676
rect 16177 5635 16243 5651
rect 16277 5753 16325 5797
rect 16311 5719 16325 5753
rect 16277 5685 16325 5719
rect 16311 5651 16325 5685
rect 16277 5635 16325 5651
rect 17163 5753 17217 5797
rect 17163 5719 17183 5753
rect 17163 5685 17217 5719
rect 17163 5651 17183 5685
rect 17163 5635 17217 5651
rect 17251 5753 17317 5763
rect 17251 5719 17267 5753
rect 17301 5719 17317 5753
rect 17251 5715 17317 5719
rect 17251 5681 17265 5715
rect 17299 5685 17317 5715
rect 17251 5651 17267 5681
rect 17301 5651 17317 5685
rect 17251 5635 17317 5651
rect 17351 5753 17399 5797
rect 17385 5719 17399 5753
rect 17748 5729 17764 5763
rect 17798 5729 17814 5763
rect 17351 5685 17399 5719
rect 17385 5651 17399 5685
rect 17351 5635 17399 5651
rect 17620 5667 17654 5686
rect 16087 5594 16107 5599
rect 16087 5560 16104 5594
rect 16141 5565 16157 5599
rect 16138 5560 16157 5565
rect 16087 5549 16157 5560
rect 16191 5515 16225 5635
rect 16259 5565 16275 5599
rect 16309 5590 16329 5599
rect 16259 5556 16277 5565
rect 16311 5556 16329 5590
rect 16259 5549 16329 5556
rect 17161 5592 17181 5599
rect 17161 5558 17179 5592
rect 17215 5565 17231 5599
rect 17213 5558 17231 5565
rect 17161 5549 17231 5558
rect 17265 5515 17299 5635
rect 17620 5599 17654 5601
rect 17333 5565 17349 5599
rect 17383 5592 17403 5599
rect 17333 5558 17353 5565
rect 17387 5558 17403 5592
rect 17333 5549 17403 5558
rect 17620 5563 17654 5565
rect 15764 5435 16030 5436
rect 15764 5401 15780 5435
rect 15814 5401 16030 5435
rect 15764 5400 16030 5401
rect 16089 5499 16155 5515
rect 16089 5465 16121 5499
rect 16191 5499 16327 5515
rect 16191 5481 16277 5499
rect 16089 5431 16155 5465
rect 15447 5363 15513 5397
rect 15447 5329 15463 5363
rect 15497 5329 15513 5363
rect 16089 5397 16121 5431
rect 16089 5363 16155 5397
rect 15447 5324 15513 5329
rect 15640 5329 15922 5362
rect 15640 5295 15730 5329
rect 15764 5327 15922 5329
rect 15764 5295 15849 5327
rect 15640 5293 15849 5295
rect 15883 5293 15922 5327
rect 15640 5287 15922 5293
rect 16089 5329 16121 5363
rect 16089 5287 16155 5329
rect 16261 5465 16277 5481
rect 16311 5465 16327 5499
rect 16261 5431 16327 5465
rect 16261 5397 16277 5431
rect 16311 5397 16327 5431
rect 16261 5363 16327 5397
rect 16261 5329 16277 5363
rect 16311 5329 16327 5363
rect 16261 5324 16327 5329
rect 17163 5499 17229 5515
rect 17163 5465 17195 5499
rect 17265 5499 17401 5515
rect 17265 5481 17351 5499
rect 17163 5431 17229 5465
rect 17163 5397 17195 5431
rect 17163 5363 17229 5397
rect 17163 5329 17195 5363
rect 17163 5287 17229 5329
rect 17335 5465 17351 5481
rect 17385 5465 17401 5499
rect 17620 5478 17654 5497
rect 17716 5667 17750 5686
rect 17716 5599 17750 5601
rect 17716 5563 17750 5565
rect 17716 5478 17750 5497
rect 17812 5667 17846 5686
rect 17812 5599 17846 5601
rect 17812 5563 17846 5565
rect 17812 5478 17846 5497
rect 17335 5431 17401 5465
rect 17335 5397 17351 5431
rect 17385 5397 17401 5431
rect 17652 5436 17718 5438
rect 17884 5436 17918 6050
rect 17969 5831 18003 6134
rect 18200 5831 18234 6042
rect 19144 6016 19178 6374
rect 19418 6351 19508 6374
rect 19542 6383 19866 6385
rect 19542 6351 19627 6383
rect 19418 6349 19627 6351
rect 19661 6374 19866 6383
rect 19918 6374 19952 6393
rect 20090 6571 20136 6691
rect 20190 6687 20236 6703
rect 20387 6773 20439 6811
rect 20387 6739 20405 6773
rect 20475 6803 20541 6845
rect 20716 6843 20745 6877
rect 20779 6843 20837 6877
rect 20871 6843 20929 6877
rect 20963 6843 20992 6877
rect 21152 6862 21200 6874
rect 21414 6866 21430 6900
rect 21464 6866 21480 6900
rect 21780 6890 21830 6960
rect 23270 6934 23304 6950
rect 23366 7056 23400 7072
rect 23462 7058 23496 7072
rect 23580 7058 23800 7080
rect 23460 7056 23800 7058
rect 23460 7022 23462 7056
rect 23496 7044 23800 7056
rect 23496 7022 23616 7044
rect 23366 6986 23400 7020
rect 23461 7020 23462 7022
rect 23461 6986 23496 7020
rect 23764 6996 23800 7044
rect 23461 6985 23462 6986
rect 23366 6934 23400 6950
rect 23462 6934 23496 6950
rect 23668 6960 23800 6996
rect 25158 7056 25192 7072
rect 25158 6986 25192 7020
rect 21780 6876 21790 6890
rect 20475 6769 20491 6803
rect 20525 6769 20541 6803
rect 20577 6790 20611 6811
rect 20387 6710 20439 6739
rect 20577 6735 20611 6756
rect 20170 6619 20186 6653
rect 20220 6642 20236 6653
rect 20170 6608 20188 6619
rect 20222 6608 20236 6642
rect 20387 6638 20423 6710
rect 20478 6701 20611 6735
rect 20782 6797 20848 6809
rect 20782 6763 20798 6797
rect 20832 6763 20848 6797
rect 20782 6746 20848 6763
rect 20478 6650 20512 6701
rect 20782 6695 20798 6746
rect 20832 6695 20848 6746
rect 20782 6683 20848 6695
rect 20882 6797 20928 6843
rect 20916 6763 20928 6797
rect 20882 6729 20928 6763
rect 20916 6695 20928 6729
rect 21152 6828 21158 6862
rect 21192 6828 21200 6862
rect 21784 6856 21790 6876
rect 21824 6856 21830 6890
rect 21784 6846 21830 6856
rect 21912 6851 21941 6885
rect 21975 6851 22033 6885
rect 22067 6851 22125 6885
rect 22159 6851 22188 6885
rect 21152 6740 21200 6828
rect 21526 6785 21542 6819
rect 21576 6818 21592 6819
rect 21576 6786 21738 6818
rect 21978 6810 22044 6817
rect 21972 6805 22044 6810
rect 21972 6786 21994 6805
rect 21576 6785 21994 6786
rect 21526 6782 21994 6785
rect 21702 6771 21994 6782
rect 22028 6771 22044 6805
rect 21702 6750 22044 6771
rect 21398 6740 21432 6742
rect 21152 6723 21432 6740
rect 21152 6706 21398 6723
rect 20170 6605 20236 6608
rect 20382 6636 20423 6638
rect 20382 6602 20384 6636
rect 20418 6602 20423 6636
rect 20382 6600 20423 6602
rect 20090 6553 20156 6571
rect 20090 6519 20106 6553
rect 20140 6519 20156 6553
rect 20090 6485 20156 6519
rect 20090 6451 20106 6485
rect 20140 6451 20156 6485
rect 20090 6417 20156 6451
rect 20090 6383 20106 6417
rect 20140 6383 20156 6417
rect 20090 6375 20156 6383
rect 20190 6553 20232 6569
rect 20224 6519 20232 6553
rect 20190 6485 20232 6519
rect 20224 6451 20232 6485
rect 20190 6417 20232 6451
rect 20224 6383 20232 6417
rect 19661 6349 19700 6374
rect 19212 6297 19228 6331
rect 19262 6297 19278 6331
rect 19418 6310 19700 6349
rect 20190 6341 20232 6383
rect 20387 6550 20423 6600
rect 20457 6634 20512 6650
rect 20491 6600 20512 6634
rect 20457 6584 20512 6600
rect 20557 6648 20625 6665
rect 20557 6647 20577 6648
rect 20557 6613 20575 6647
rect 20611 6614 20625 6648
rect 20609 6613 20625 6614
rect 20557 6591 20625 6613
rect 20478 6555 20512 6584
rect 20782 6563 20828 6683
rect 20882 6679 20928 6695
rect 21100 6658 21116 6659
rect 20862 6611 20878 6645
rect 20912 6638 20928 6645
rect 20980 6638 21116 6658
rect 20912 6625 21116 6638
rect 21150 6625 21166 6659
rect 20912 6624 21166 6625
rect 20912 6611 21020 6624
rect 21100 6622 21166 6624
rect 21398 6655 21432 6657
rect 20862 6597 21020 6611
rect 20876 6596 21020 6597
rect 21398 6619 21432 6621
rect 21072 6563 21106 6582
rect 20387 6500 20441 6550
rect 20478 6521 20613 6555
rect 20387 6466 20405 6500
rect 20439 6466 20441 6500
rect 20577 6487 20613 6521
rect 20387 6419 20441 6466
rect 20387 6385 20405 6419
rect 20439 6385 20441 6419
rect 20387 6369 20441 6385
rect 20475 6453 20491 6487
rect 20525 6453 20541 6487
rect 20475 6419 20541 6453
rect 20475 6385 20491 6419
rect 20525 6385 20541 6419
rect 19586 6308 19700 6310
rect 19858 6297 19874 6331
rect 19908 6297 19924 6331
rect 20024 6307 20053 6341
rect 20087 6307 20145 6341
rect 20179 6307 20237 6341
rect 20271 6307 20300 6341
rect 20475 6335 20541 6385
rect 20611 6453 20613 6487
rect 20577 6419 20613 6453
rect 20611 6385 20613 6419
rect 20577 6369 20613 6385
rect 20782 6545 20848 6563
rect 20782 6511 20798 6545
rect 20832 6511 20848 6545
rect 20782 6477 20848 6511
rect 20782 6443 20798 6477
rect 20832 6443 20848 6477
rect 20782 6409 20848 6443
rect 20782 6375 20798 6409
rect 20832 6375 20848 6409
rect 20782 6367 20848 6375
rect 20882 6545 20924 6561
rect 20916 6511 20924 6545
rect 20882 6477 20924 6511
rect 20916 6443 20924 6477
rect 20882 6409 20924 6443
rect 21072 6495 21106 6497
rect 21072 6459 21106 6461
rect 20916 6375 20924 6409
rect 20191 6300 20225 6307
rect 20370 6301 20399 6335
rect 20433 6301 20491 6335
rect 20525 6301 20583 6335
rect 20617 6301 20646 6335
rect 20882 6333 20924 6375
rect 21032 6393 21072 6414
rect 21160 6563 21194 6582
rect 21398 6534 21432 6553
rect 21494 6723 21528 6742
rect 21494 6655 21528 6657
rect 21494 6619 21528 6621
rect 21494 6534 21528 6553
rect 21590 6723 21624 6742
rect 21978 6737 22044 6750
rect 21978 6703 21994 6737
rect 22028 6703 22044 6737
rect 21978 6691 22044 6703
rect 22078 6805 22124 6851
rect 22258 6845 22287 6879
rect 22321 6845 22379 6879
rect 22413 6845 22471 6879
rect 22505 6845 22534 6879
rect 22112 6771 22124 6805
rect 22078 6737 22124 6771
rect 22112 6703 22124 6737
rect 21590 6655 21624 6657
rect 21746 6625 21762 6659
rect 21796 6625 21812 6659
rect 21590 6619 21624 6621
rect 21590 6534 21624 6553
rect 21718 6563 21752 6582
rect 21160 6495 21194 6497
rect 21718 6495 21752 6497
rect 21160 6459 21194 6461
rect 21430 6457 21446 6491
rect 21480 6457 21496 6491
rect 21718 6459 21752 6461
rect 21106 6393 21108 6414
rect 21032 6374 21108 6393
rect 21194 6393 21718 6418
rect 21806 6563 21840 6582
rect 21806 6495 21840 6497
rect 21806 6459 21840 6461
rect 21752 6393 21754 6418
rect 21160 6385 21754 6393
rect 21160 6374 21396 6385
rect 20716 6299 20745 6333
rect 20779 6299 20837 6333
rect 20871 6299 20929 6333
rect 20963 6299 20992 6333
rect 19278 6212 19324 6218
rect 19278 6210 19766 6212
rect 19278 6176 19286 6210
rect 19320 6193 19766 6210
rect 19320 6188 19716 6193
rect 19320 6178 19595 6188
rect 19320 6176 19324 6178
rect 19278 6174 19324 6176
rect 19496 6154 19595 6178
rect 19629 6159 19716 6188
rect 19750 6168 19766 6193
rect 19750 6159 19891 6168
rect 19629 6154 19891 6159
rect 19496 6134 19891 6154
rect 19620 6050 19636 6084
rect 19670 6050 19806 6084
rect 19144 6000 19526 6016
rect 19144 5976 19492 6000
rect 19492 5930 19526 5964
rect 19492 5878 19526 5894
rect 19588 6000 19622 6016
rect 19588 5930 19622 5964
rect 19588 5878 19622 5894
rect 19684 6000 19718 6016
rect 19684 5930 19718 5964
rect 19684 5878 19718 5894
rect 17958 5797 17987 5831
rect 18021 5797 18079 5831
rect 18113 5797 18171 5831
rect 18205 5797 18234 5831
rect 19032 5797 19061 5831
rect 19095 5797 19153 5831
rect 19187 5797 19245 5831
rect 19279 5797 19308 5831
rect 19524 5810 19540 5844
rect 19574 5810 19590 5844
rect 17977 5753 18031 5797
rect 17977 5719 17997 5753
rect 17977 5685 18031 5719
rect 17977 5651 17997 5685
rect 17977 5635 18031 5651
rect 18065 5753 18131 5763
rect 18065 5719 18081 5753
rect 18115 5719 18131 5753
rect 18065 5710 18131 5719
rect 18065 5685 18083 5710
rect 18065 5651 18081 5685
rect 18117 5676 18131 5710
rect 18115 5651 18131 5676
rect 18065 5635 18131 5651
rect 18165 5753 18213 5797
rect 18199 5719 18213 5753
rect 18165 5685 18213 5719
rect 18199 5651 18213 5685
rect 18165 5635 18213 5651
rect 19051 5753 19105 5797
rect 19051 5719 19071 5753
rect 19051 5685 19105 5719
rect 19051 5651 19071 5685
rect 19051 5635 19105 5651
rect 19139 5753 19205 5763
rect 19139 5719 19155 5753
rect 19189 5719 19205 5753
rect 19139 5715 19205 5719
rect 19139 5681 19153 5715
rect 19187 5685 19205 5715
rect 19139 5651 19155 5681
rect 19189 5651 19205 5685
rect 19139 5635 19205 5651
rect 19239 5753 19287 5797
rect 19273 5719 19287 5753
rect 19636 5729 19652 5763
rect 19686 5729 19702 5763
rect 19239 5685 19287 5719
rect 19273 5651 19287 5685
rect 19239 5635 19287 5651
rect 19508 5667 19542 5686
rect 17975 5594 17995 5599
rect 17975 5560 17992 5594
rect 18029 5565 18045 5599
rect 18026 5560 18045 5565
rect 17975 5549 18045 5560
rect 18079 5515 18113 5635
rect 18147 5565 18163 5599
rect 18197 5590 18217 5599
rect 18147 5556 18165 5565
rect 18199 5556 18217 5590
rect 18147 5549 18217 5556
rect 19049 5592 19069 5599
rect 19049 5558 19067 5592
rect 19103 5565 19119 5599
rect 19101 5558 19119 5565
rect 19049 5549 19119 5558
rect 19153 5515 19187 5635
rect 19508 5599 19542 5601
rect 19221 5565 19237 5599
rect 19271 5592 19291 5599
rect 19221 5558 19241 5565
rect 19275 5558 19291 5592
rect 19221 5549 19291 5558
rect 19508 5563 19542 5565
rect 17652 5435 17918 5436
rect 17652 5401 17668 5435
rect 17702 5401 17918 5435
rect 17652 5400 17918 5401
rect 17977 5499 18043 5515
rect 17977 5465 18009 5499
rect 18079 5499 18215 5515
rect 18079 5481 18165 5499
rect 17977 5431 18043 5465
rect 17335 5363 17401 5397
rect 17335 5329 17351 5363
rect 17385 5329 17401 5363
rect 17977 5397 18009 5431
rect 17977 5363 18043 5397
rect 17335 5324 17401 5329
rect 17528 5329 17810 5362
rect 17528 5295 17618 5329
rect 17652 5327 17810 5329
rect 17652 5295 17737 5327
rect 17528 5293 17737 5295
rect 17771 5293 17810 5327
rect 17528 5287 17810 5293
rect 17977 5329 18009 5363
rect 17977 5287 18043 5329
rect 18149 5465 18165 5481
rect 18199 5465 18215 5499
rect 18149 5431 18215 5465
rect 18149 5397 18165 5431
rect 18199 5397 18215 5431
rect 18149 5363 18215 5397
rect 18149 5329 18165 5363
rect 18199 5329 18215 5363
rect 18149 5324 18215 5329
rect 19051 5499 19117 5515
rect 19051 5465 19083 5499
rect 19153 5499 19289 5515
rect 19153 5481 19239 5499
rect 19051 5431 19117 5465
rect 19051 5397 19083 5431
rect 19051 5363 19117 5397
rect 19051 5329 19083 5363
rect 19051 5287 19117 5329
rect 19223 5465 19239 5481
rect 19273 5465 19289 5499
rect 19508 5478 19542 5497
rect 19604 5667 19638 5686
rect 19604 5599 19638 5601
rect 19604 5563 19638 5565
rect 19604 5478 19638 5497
rect 19700 5667 19734 5686
rect 19700 5599 19734 5601
rect 19700 5563 19734 5565
rect 19700 5478 19734 5497
rect 19223 5431 19289 5465
rect 19223 5397 19239 5431
rect 19273 5397 19289 5431
rect 19540 5436 19606 5438
rect 19772 5436 19806 6050
rect 19857 5831 19891 6134
rect 20088 5831 20122 6042
rect 21032 6016 21066 6374
rect 21306 6351 21396 6374
rect 21430 6383 21754 6385
rect 21430 6351 21515 6383
rect 21306 6349 21515 6351
rect 21549 6374 21754 6383
rect 21806 6374 21840 6393
rect 21978 6571 22024 6691
rect 22078 6687 22124 6703
rect 22275 6773 22327 6811
rect 22275 6739 22293 6773
rect 22363 6803 22429 6845
rect 22604 6843 22633 6877
rect 22667 6843 22725 6877
rect 22759 6843 22817 6877
rect 22851 6843 22880 6877
rect 23040 6862 23088 6874
rect 23302 6866 23318 6900
rect 23352 6866 23368 6900
rect 23668 6890 23718 6960
rect 25158 6934 25192 6950
rect 25254 7056 25288 7072
rect 25350 7058 25384 7072
rect 25468 7058 25688 7080
rect 25348 7056 25688 7058
rect 25348 7022 25350 7056
rect 25384 7044 25688 7056
rect 25384 7022 25504 7044
rect 25254 6986 25288 7020
rect 25349 7020 25350 7022
rect 25349 6986 25384 7020
rect 25652 6996 25688 7044
rect 25349 6985 25350 6986
rect 25254 6934 25288 6950
rect 25350 6934 25384 6950
rect 25556 6960 25688 6996
rect 27046 7056 27080 7072
rect 27046 6986 27080 7020
rect 23668 6876 23678 6890
rect 22363 6769 22379 6803
rect 22413 6769 22429 6803
rect 22465 6790 22499 6811
rect 22275 6710 22327 6739
rect 22465 6735 22499 6756
rect 22058 6619 22074 6653
rect 22108 6642 22124 6653
rect 22058 6608 22076 6619
rect 22110 6608 22124 6642
rect 22275 6638 22311 6710
rect 22366 6701 22499 6735
rect 22670 6797 22736 6809
rect 22670 6763 22686 6797
rect 22720 6763 22736 6797
rect 22670 6746 22736 6763
rect 22366 6650 22400 6701
rect 22670 6695 22686 6746
rect 22720 6695 22736 6746
rect 22670 6683 22736 6695
rect 22770 6797 22816 6843
rect 22804 6763 22816 6797
rect 22770 6729 22816 6763
rect 22804 6695 22816 6729
rect 23040 6828 23046 6862
rect 23080 6828 23088 6862
rect 23672 6856 23678 6876
rect 23712 6856 23718 6890
rect 23672 6846 23718 6856
rect 23800 6851 23829 6885
rect 23863 6851 23921 6885
rect 23955 6851 24013 6885
rect 24047 6851 24076 6885
rect 23040 6740 23088 6828
rect 23414 6785 23430 6819
rect 23464 6818 23480 6819
rect 23464 6786 23626 6818
rect 23866 6810 23932 6817
rect 23860 6805 23932 6810
rect 23860 6786 23882 6805
rect 23464 6785 23882 6786
rect 23414 6782 23882 6785
rect 23590 6771 23882 6782
rect 23916 6771 23932 6805
rect 23590 6750 23932 6771
rect 23286 6740 23320 6742
rect 23040 6723 23320 6740
rect 23040 6706 23286 6723
rect 22058 6605 22124 6608
rect 22270 6636 22311 6638
rect 22270 6602 22272 6636
rect 22306 6602 22311 6636
rect 22270 6600 22311 6602
rect 21978 6553 22044 6571
rect 21978 6519 21994 6553
rect 22028 6519 22044 6553
rect 21978 6485 22044 6519
rect 21978 6451 21994 6485
rect 22028 6451 22044 6485
rect 21978 6417 22044 6451
rect 21978 6383 21994 6417
rect 22028 6383 22044 6417
rect 21978 6375 22044 6383
rect 22078 6553 22120 6569
rect 22112 6519 22120 6553
rect 22078 6485 22120 6519
rect 22112 6451 22120 6485
rect 22078 6417 22120 6451
rect 22112 6383 22120 6417
rect 21549 6349 21588 6374
rect 21100 6297 21116 6331
rect 21150 6297 21166 6331
rect 21306 6310 21588 6349
rect 22078 6341 22120 6383
rect 22275 6550 22311 6600
rect 22345 6634 22400 6650
rect 22379 6600 22400 6634
rect 22345 6584 22400 6600
rect 22445 6648 22513 6665
rect 22445 6647 22465 6648
rect 22445 6613 22463 6647
rect 22499 6614 22513 6648
rect 22497 6613 22513 6614
rect 22445 6591 22513 6613
rect 22366 6555 22400 6584
rect 22670 6563 22716 6683
rect 22770 6679 22816 6695
rect 22988 6658 23004 6659
rect 22750 6611 22766 6645
rect 22800 6638 22816 6645
rect 22868 6638 23004 6658
rect 22800 6625 23004 6638
rect 23038 6625 23054 6659
rect 22800 6624 23054 6625
rect 22800 6611 22908 6624
rect 22988 6622 23054 6624
rect 23286 6655 23320 6657
rect 22750 6597 22908 6611
rect 22764 6596 22908 6597
rect 23286 6619 23320 6621
rect 22960 6563 22994 6582
rect 22275 6500 22329 6550
rect 22366 6521 22501 6555
rect 22275 6466 22293 6500
rect 22327 6466 22329 6500
rect 22465 6487 22501 6521
rect 22275 6419 22329 6466
rect 22275 6385 22293 6419
rect 22327 6385 22329 6419
rect 22275 6369 22329 6385
rect 22363 6453 22379 6487
rect 22413 6453 22429 6487
rect 22363 6419 22429 6453
rect 22363 6385 22379 6419
rect 22413 6385 22429 6419
rect 21474 6308 21588 6310
rect 21746 6297 21762 6331
rect 21796 6297 21812 6331
rect 21912 6307 21941 6341
rect 21975 6307 22033 6341
rect 22067 6307 22125 6341
rect 22159 6307 22188 6341
rect 22363 6335 22429 6385
rect 22499 6453 22501 6487
rect 22465 6419 22501 6453
rect 22499 6385 22501 6419
rect 22465 6369 22501 6385
rect 22670 6545 22736 6563
rect 22670 6511 22686 6545
rect 22720 6511 22736 6545
rect 22670 6477 22736 6511
rect 22670 6443 22686 6477
rect 22720 6443 22736 6477
rect 22670 6409 22736 6443
rect 22670 6375 22686 6409
rect 22720 6375 22736 6409
rect 22670 6367 22736 6375
rect 22770 6545 22812 6561
rect 22804 6511 22812 6545
rect 22770 6477 22812 6511
rect 22804 6443 22812 6477
rect 22770 6409 22812 6443
rect 22960 6495 22994 6497
rect 22960 6459 22994 6461
rect 22804 6375 22812 6409
rect 22079 6300 22113 6307
rect 22258 6301 22287 6335
rect 22321 6301 22379 6335
rect 22413 6301 22471 6335
rect 22505 6301 22534 6335
rect 22770 6333 22812 6375
rect 22920 6393 22960 6414
rect 23048 6563 23082 6582
rect 23286 6534 23320 6553
rect 23382 6723 23416 6742
rect 23382 6655 23416 6657
rect 23382 6619 23416 6621
rect 23382 6534 23416 6553
rect 23478 6723 23512 6742
rect 23866 6737 23932 6750
rect 23866 6703 23882 6737
rect 23916 6703 23932 6737
rect 23866 6691 23932 6703
rect 23966 6805 24012 6851
rect 24146 6845 24175 6879
rect 24209 6845 24267 6879
rect 24301 6845 24359 6879
rect 24393 6845 24422 6879
rect 24000 6771 24012 6805
rect 23966 6737 24012 6771
rect 24000 6703 24012 6737
rect 23478 6655 23512 6657
rect 23634 6625 23650 6659
rect 23684 6625 23700 6659
rect 23478 6619 23512 6621
rect 23478 6534 23512 6553
rect 23606 6563 23640 6582
rect 23048 6495 23082 6497
rect 23606 6495 23640 6497
rect 23048 6459 23082 6461
rect 23318 6457 23334 6491
rect 23368 6457 23384 6491
rect 23606 6459 23640 6461
rect 22994 6393 22996 6414
rect 22920 6374 22996 6393
rect 23082 6393 23606 6418
rect 23694 6563 23728 6582
rect 23694 6495 23728 6497
rect 23694 6459 23728 6461
rect 23640 6393 23642 6418
rect 23048 6385 23642 6393
rect 23048 6374 23284 6385
rect 22604 6299 22633 6333
rect 22667 6299 22725 6333
rect 22759 6299 22817 6333
rect 22851 6299 22880 6333
rect 21166 6212 21212 6218
rect 21166 6210 21654 6212
rect 21166 6176 21174 6210
rect 21208 6193 21654 6210
rect 21208 6188 21604 6193
rect 21208 6178 21483 6188
rect 21208 6176 21212 6178
rect 21166 6174 21212 6176
rect 21384 6154 21483 6178
rect 21517 6159 21604 6188
rect 21638 6168 21654 6193
rect 21638 6159 21779 6168
rect 21517 6154 21779 6159
rect 21384 6134 21779 6154
rect 21508 6050 21524 6084
rect 21558 6050 21694 6084
rect 21032 6000 21414 6016
rect 21032 5976 21380 6000
rect 21380 5930 21414 5964
rect 21380 5878 21414 5894
rect 21476 6000 21510 6016
rect 21476 5930 21510 5964
rect 21476 5878 21510 5894
rect 21572 6000 21606 6016
rect 21572 5930 21606 5964
rect 21572 5878 21606 5894
rect 19846 5797 19875 5831
rect 19909 5797 19967 5831
rect 20001 5797 20059 5831
rect 20093 5797 20122 5831
rect 20920 5797 20949 5831
rect 20983 5797 21041 5831
rect 21075 5797 21133 5831
rect 21167 5797 21196 5831
rect 21412 5810 21428 5844
rect 21462 5810 21478 5844
rect 19865 5753 19919 5797
rect 19865 5719 19885 5753
rect 19865 5685 19919 5719
rect 19865 5651 19885 5685
rect 19865 5635 19919 5651
rect 19953 5753 20019 5763
rect 19953 5719 19969 5753
rect 20003 5719 20019 5753
rect 19953 5710 20019 5719
rect 19953 5685 19971 5710
rect 19953 5651 19969 5685
rect 20005 5676 20019 5710
rect 20003 5651 20019 5676
rect 19953 5635 20019 5651
rect 20053 5753 20101 5797
rect 20087 5719 20101 5753
rect 20053 5685 20101 5719
rect 20087 5651 20101 5685
rect 20053 5635 20101 5651
rect 20939 5753 20993 5797
rect 20939 5719 20959 5753
rect 20939 5685 20993 5719
rect 20939 5651 20959 5685
rect 20939 5635 20993 5651
rect 21027 5753 21093 5763
rect 21027 5719 21043 5753
rect 21077 5719 21093 5753
rect 21027 5715 21093 5719
rect 21027 5681 21041 5715
rect 21075 5685 21093 5715
rect 21027 5651 21043 5681
rect 21077 5651 21093 5685
rect 21027 5635 21093 5651
rect 21127 5753 21175 5797
rect 21161 5719 21175 5753
rect 21524 5729 21540 5763
rect 21574 5729 21590 5763
rect 21127 5685 21175 5719
rect 21161 5651 21175 5685
rect 21127 5635 21175 5651
rect 21396 5667 21430 5686
rect 19863 5594 19883 5599
rect 19863 5560 19880 5594
rect 19917 5565 19933 5599
rect 19914 5560 19933 5565
rect 19863 5549 19933 5560
rect 19967 5515 20001 5635
rect 20035 5565 20051 5599
rect 20085 5590 20105 5599
rect 20035 5556 20053 5565
rect 20087 5556 20105 5590
rect 20035 5549 20105 5556
rect 20937 5592 20957 5599
rect 20937 5558 20955 5592
rect 20991 5565 21007 5599
rect 20989 5558 21007 5565
rect 20937 5549 21007 5558
rect 21041 5515 21075 5635
rect 21396 5599 21430 5601
rect 21109 5565 21125 5599
rect 21159 5592 21179 5599
rect 21109 5558 21129 5565
rect 21163 5558 21179 5592
rect 21109 5549 21179 5558
rect 21396 5563 21430 5565
rect 19540 5435 19806 5436
rect 19540 5401 19556 5435
rect 19590 5401 19806 5435
rect 19540 5400 19806 5401
rect 19865 5499 19931 5515
rect 19865 5465 19897 5499
rect 19967 5499 20103 5515
rect 19967 5481 20053 5499
rect 19865 5431 19931 5465
rect 19223 5363 19289 5397
rect 19223 5329 19239 5363
rect 19273 5329 19289 5363
rect 19865 5397 19897 5431
rect 19865 5363 19931 5397
rect 19223 5324 19289 5329
rect 19416 5329 19698 5362
rect 19416 5295 19506 5329
rect 19540 5327 19698 5329
rect 19540 5295 19625 5327
rect 19416 5293 19625 5295
rect 19659 5293 19698 5327
rect 19416 5287 19698 5293
rect 19865 5329 19897 5363
rect 19865 5287 19931 5329
rect 20037 5465 20053 5481
rect 20087 5465 20103 5499
rect 20037 5431 20103 5465
rect 20037 5397 20053 5431
rect 20087 5397 20103 5431
rect 20037 5363 20103 5397
rect 20037 5329 20053 5363
rect 20087 5329 20103 5363
rect 20037 5324 20103 5329
rect 20939 5499 21005 5515
rect 20939 5465 20971 5499
rect 21041 5499 21177 5515
rect 21041 5481 21127 5499
rect 20939 5431 21005 5465
rect 20939 5397 20971 5431
rect 20939 5363 21005 5397
rect 20939 5329 20971 5363
rect 20939 5287 21005 5329
rect 21111 5465 21127 5481
rect 21161 5465 21177 5499
rect 21396 5478 21430 5497
rect 21492 5667 21526 5686
rect 21492 5599 21526 5601
rect 21492 5563 21526 5565
rect 21492 5478 21526 5497
rect 21588 5667 21622 5686
rect 21588 5599 21622 5601
rect 21588 5563 21622 5565
rect 21588 5478 21622 5497
rect 21111 5431 21177 5465
rect 21111 5397 21127 5431
rect 21161 5397 21177 5431
rect 21428 5436 21494 5438
rect 21660 5436 21694 6050
rect 21745 5831 21779 6134
rect 21976 5831 22010 6042
rect 22920 6016 22954 6374
rect 23194 6351 23284 6374
rect 23318 6383 23642 6385
rect 23318 6351 23403 6383
rect 23194 6349 23403 6351
rect 23437 6374 23642 6383
rect 23694 6374 23728 6393
rect 23866 6571 23912 6691
rect 23966 6687 24012 6703
rect 24163 6773 24215 6811
rect 24163 6739 24181 6773
rect 24251 6803 24317 6845
rect 24492 6843 24521 6877
rect 24555 6843 24613 6877
rect 24647 6843 24705 6877
rect 24739 6843 24768 6877
rect 24928 6862 24976 6874
rect 25190 6866 25206 6900
rect 25240 6866 25256 6900
rect 25556 6890 25606 6960
rect 27046 6934 27080 6950
rect 27142 7056 27176 7072
rect 27238 7058 27272 7072
rect 27356 7058 27576 7080
rect 27236 7056 27576 7058
rect 27236 7022 27238 7056
rect 27272 7044 27576 7056
rect 27272 7022 27392 7044
rect 27142 6986 27176 7020
rect 27237 7020 27238 7022
rect 27237 6986 27272 7020
rect 27540 6996 27576 7044
rect 27237 6985 27238 6986
rect 27142 6934 27176 6950
rect 27238 6934 27272 6950
rect 27444 6960 27576 6996
rect 28934 7056 28968 7072
rect 28934 6986 28968 7020
rect 25556 6876 25566 6890
rect 24251 6769 24267 6803
rect 24301 6769 24317 6803
rect 24353 6790 24387 6811
rect 24163 6710 24215 6739
rect 24353 6735 24387 6756
rect 23946 6619 23962 6653
rect 23996 6642 24012 6653
rect 23946 6608 23964 6619
rect 23998 6608 24012 6642
rect 24163 6638 24199 6710
rect 24254 6701 24387 6735
rect 24558 6797 24624 6809
rect 24558 6763 24574 6797
rect 24608 6763 24624 6797
rect 24558 6746 24624 6763
rect 24254 6650 24288 6701
rect 24558 6695 24574 6746
rect 24608 6695 24624 6746
rect 24558 6683 24624 6695
rect 24658 6797 24704 6843
rect 24692 6763 24704 6797
rect 24658 6729 24704 6763
rect 24692 6695 24704 6729
rect 24928 6828 24934 6862
rect 24968 6828 24976 6862
rect 25560 6856 25566 6876
rect 25600 6856 25606 6890
rect 25560 6846 25606 6856
rect 25688 6851 25717 6885
rect 25751 6851 25809 6885
rect 25843 6851 25901 6885
rect 25935 6851 25964 6885
rect 24928 6740 24976 6828
rect 25302 6785 25318 6819
rect 25352 6818 25368 6819
rect 25352 6786 25514 6818
rect 25754 6810 25820 6817
rect 25748 6805 25820 6810
rect 25748 6786 25770 6805
rect 25352 6785 25770 6786
rect 25302 6782 25770 6785
rect 25478 6771 25770 6782
rect 25804 6771 25820 6805
rect 25478 6750 25820 6771
rect 25174 6740 25208 6742
rect 24928 6723 25208 6740
rect 24928 6706 25174 6723
rect 23946 6605 24012 6608
rect 24158 6636 24199 6638
rect 24158 6602 24160 6636
rect 24194 6602 24199 6636
rect 24158 6600 24199 6602
rect 23866 6553 23932 6571
rect 23866 6519 23882 6553
rect 23916 6519 23932 6553
rect 23866 6485 23932 6519
rect 23866 6451 23882 6485
rect 23916 6451 23932 6485
rect 23866 6417 23932 6451
rect 23866 6383 23882 6417
rect 23916 6383 23932 6417
rect 23866 6375 23932 6383
rect 23966 6553 24008 6569
rect 24000 6519 24008 6553
rect 23966 6485 24008 6519
rect 24000 6451 24008 6485
rect 23966 6417 24008 6451
rect 24000 6383 24008 6417
rect 23437 6349 23476 6374
rect 22988 6297 23004 6331
rect 23038 6297 23054 6331
rect 23194 6310 23476 6349
rect 23966 6341 24008 6383
rect 24163 6550 24199 6600
rect 24233 6634 24288 6650
rect 24267 6600 24288 6634
rect 24233 6584 24288 6600
rect 24333 6648 24401 6665
rect 24333 6647 24353 6648
rect 24333 6613 24351 6647
rect 24387 6614 24401 6648
rect 24385 6613 24401 6614
rect 24333 6591 24401 6613
rect 24254 6555 24288 6584
rect 24558 6563 24604 6683
rect 24658 6679 24704 6695
rect 24876 6658 24892 6659
rect 24638 6611 24654 6645
rect 24688 6638 24704 6645
rect 24756 6638 24892 6658
rect 24688 6625 24892 6638
rect 24926 6625 24942 6659
rect 24688 6624 24942 6625
rect 24688 6611 24796 6624
rect 24876 6622 24942 6624
rect 25174 6655 25208 6657
rect 24638 6597 24796 6611
rect 24652 6596 24796 6597
rect 25174 6619 25208 6621
rect 24848 6563 24882 6582
rect 24163 6500 24217 6550
rect 24254 6521 24389 6555
rect 24163 6466 24181 6500
rect 24215 6466 24217 6500
rect 24353 6487 24389 6521
rect 24163 6419 24217 6466
rect 24163 6385 24181 6419
rect 24215 6385 24217 6419
rect 24163 6369 24217 6385
rect 24251 6453 24267 6487
rect 24301 6453 24317 6487
rect 24251 6419 24317 6453
rect 24251 6385 24267 6419
rect 24301 6385 24317 6419
rect 23362 6308 23476 6310
rect 23634 6297 23650 6331
rect 23684 6297 23700 6331
rect 23800 6307 23829 6341
rect 23863 6307 23921 6341
rect 23955 6307 24013 6341
rect 24047 6307 24076 6341
rect 24251 6335 24317 6385
rect 24387 6453 24389 6487
rect 24353 6419 24389 6453
rect 24387 6385 24389 6419
rect 24353 6369 24389 6385
rect 24558 6545 24624 6563
rect 24558 6511 24574 6545
rect 24608 6511 24624 6545
rect 24558 6477 24624 6511
rect 24558 6443 24574 6477
rect 24608 6443 24624 6477
rect 24558 6409 24624 6443
rect 24558 6375 24574 6409
rect 24608 6375 24624 6409
rect 24558 6367 24624 6375
rect 24658 6545 24700 6561
rect 24692 6511 24700 6545
rect 24658 6477 24700 6511
rect 24692 6443 24700 6477
rect 24658 6409 24700 6443
rect 24848 6495 24882 6497
rect 24848 6459 24882 6461
rect 24692 6375 24700 6409
rect 23967 6300 24001 6307
rect 24146 6301 24175 6335
rect 24209 6301 24267 6335
rect 24301 6301 24359 6335
rect 24393 6301 24422 6335
rect 24658 6333 24700 6375
rect 24808 6393 24848 6414
rect 24936 6563 24970 6582
rect 25174 6534 25208 6553
rect 25270 6723 25304 6742
rect 25270 6655 25304 6657
rect 25270 6619 25304 6621
rect 25270 6534 25304 6553
rect 25366 6723 25400 6742
rect 25754 6737 25820 6750
rect 25754 6703 25770 6737
rect 25804 6703 25820 6737
rect 25754 6691 25820 6703
rect 25854 6805 25900 6851
rect 26034 6845 26063 6879
rect 26097 6845 26155 6879
rect 26189 6845 26247 6879
rect 26281 6845 26310 6879
rect 25888 6771 25900 6805
rect 25854 6737 25900 6771
rect 25888 6703 25900 6737
rect 25366 6655 25400 6657
rect 25522 6625 25538 6659
rect 25572 6625 25588 6659
rect 25366 6619 25400 6621
rect 25366 6534 25400 6553
rect 25494 6563 25528 6582
rect 24936 6495 24970 6497
rect 25494 6495 25528 6497
rect 24936 6459 24970 6461
rect 25206 6457 25222 6491
rect 25256 6457 25272 6491
rect 25494 6459 25528 6461
rect 24882 6393 24884 6414
rect 24808 6374 24884 6393
rect 24970 6393 25494 6418
rect 25582 6563 25616 6582
rect 25582 6495 25616 6497
rect 25582 6459 25616 6461
rect 25528 6393 25530 6418
rect 24936 6385 25530 6393
rect 24936 6374 25172 6385
rect 24492 6299 24521 6333
rect 24555 6299 24613 6333
rect 24647 6299 24705 6333
rect 24739 6299 24768 6333
rect 23054 6212 23100 6218
rect 23054 6210 23542 6212
rect 23054 6176 23062 6210
rect 23096 6193 23542 6210
rect 23096 6188 23492 6193
rect 23096 6178 23371 6188
rect 23096 6176 23100 6178
rect 23054 6174 23100 6176
rect 23272 6154 23371 6178
rect 23405 6159 23492 6188
rect 23526 6168 23542 6193
rect 23526 6159 23667 6168
rect 23405 6154 23667 6159
rect 23272 6134 23667 6154
rect 23396 6050 23412 6084
rect 23446 6050 23582 6084
rect 22920 6000 23302 6016
rect 22920 5976 23268 6000
rect 23268 5930 23302 5964
rect 23268 5878 23302 5894
rect 23364 6000 23398 6016
rect 23364 5930 23398 5964
rect 23364 5878 23398 5894
rect 23460 6000 23494 6016
rect 23460 5930 23494 5964
rect 23460 5878 23494 5894
rect 21734 5797 21763 5831
rect 21797 5797 21855 5831
rect 21889 5797 21947 5831
rect 21981 5797 22010 5831
rect 22808 5797 22837 5831
rect 22871 5797 22929 5831
rect 22963 5797 23021 5831
rect 23055 5797 23084 5831
rect 23300 5810 23316 5844
rect 23350 5810 23366 5844
rect 21753 5753 21807 5797
rect 21753 5719 21773 5753
rect 21753 5685 21807 5719
rect 21753 5651 21773 5685
rect 21753 5635 21807 5651
rect 21841 5753 21907 5763
rect 21841 5719 21857 5753
rect 21891 5719 21907 5753
rect 21841 5710 21907 5719
rect 21841 5685 21859 5710
rect 21841 5651 21857 5685
rect 21893 5676 21907 5710
rect 21891 5651 21907 5676
rect 21841 5635 21907 5651
rect 21941 5753 21989 5797
rect 21975 5719 21989 5753
rect 21941 5685 21989 5719
rect 21975 5651 21989 5685
rect 21941 5635 21989 5651
rect 22827 5753 22881 5797
rect 22827 5719 22847 5753
rect 22827 5685 22881 5719
rect 22827 5651 22847 5685
rect 22827 5635 22881 5651
rect 22915 5753 22981 5763
rect 22915 5719 22931 5753
rect 22965 5719 22981 5753
rect 22915 5715 22981 5719
rect 22915 5681 22929 5715
rect 22963 5685 22981 5715
rect 22915 5651 22931 5681
rect 22965 5651 22981 5685
rect 22915 5635 22981 5651
rect 23015 5753 23063 5797
rect 23049 5719 23063 5753
rect 23412 5729 23428 5763
rect 23462 5729 23478 5763
rect 23015 5685 23063 5719
rect 23049 5651 23063 5685
rect 23015 5635 23063 5651
rect 23284 5667 23318 5686
rect 21751 5594 21771 5599
rect 21751 5560 21768 5594
rect 21805 5565 21821 5599
rect 21802 5560 21821 5565
rect 21751 5549 21821 5560
rect 21855 5515 21889 5635
rect 21923 5565 21939 5599
rect 21973 5590 21993 5599
rect 21923 5556 21941 5565
rect 21975 5556 21993 5590
rect 21923 5549 21993 5556
rect 22825 5592 22845 5599
rect 22825 5558 22843 5592
rect 22879 5565 22895 5599
rect 22877 5558 22895 5565
rect 22825 5549 22895 5558
rect 22929 5515 22963 5635
rect 23284 5599 23318 5601
rect 22997 5565 23013 5599
rect 23047 5592 23067 5599
rect 22997 5558 23017 5565
rect 23051 5558 23067 5592
rect 22997 5549 23067 5558
rect 23284 5563 23318 5565
rect 21428 5435 21694 5436
rect 21428 5401 21444 5435
rect 21478 5401 21694 5435
rect 21428 5400 21694 5401
rect 21753 5499 21819 5515
rect 21753 5465 21785 5499
rect 21855 5499 21991 5515
rect 21855 5481 21941 5499
rect 21753 5431 21819 5465
rect 21111 5363 21177 5397
rect 21111 5329 21127 5363
rect 21161 5329 21177 5363
rect 21753 5397 21785 5431
rect 21753 5363 21819 5397
rect 21111 5324 21177 5329
rect 21304 5329 21586 5362
rect 21304 5295 21394 5329
rect 21428 5327 21586 5329
rect 21428 5295 21513 5327
rect 21304 5293 21513 5295
rect 21547 5293 21586 5327
rect 21304 5287 21586 5293
rect 21753 5329 21785 5363
rect 21753 5287 21819 5329
rect 21925 5465 21941 5481
rect 21975 5465 21991 5499
rect 21925 5431 21991 5465
rect 21925 5397 21941 5431
rect 21975 5397 21991 5431
rect 21925 5363 21991 5397
rect 21925 5329 21941 5363
rect 21975 5329 21991 5363
rect 21925 5324 21991 5329
rect 22827 5499 22893 5515
rect 22827 5465 22859 5499
rect 22929 5499 23065 5515
rect 22929 5481 23015 5499
rect 22827 5431 22893 5465
rect 22827 5397 22859 5431
rect 22827 5363 22893 5397
rect 22827 5329 22859 5363
rect 22827 5287 22893 5329
rect 22999 5465 23015 5481
rect 23049 5465 23065 5499
rect 23284 5478 23318 5497
rect 23380 5667 23414 5686
rect 23380 5599 23414 5601
rect 23380 5563 23414 5565
rect 23380 5478 23414 5497
rect 23476 5667 23510 5686
rect 23476 5599 23510 5601
rect 23476 5563 23510 5565
rect 23476 5478 23510 5497
rect 22999 5431 23065 5465
rect 22999 5397 23015 5431
rect 23049 5397 23065 5431
rect 23316 5436 23382 5438
rect 23548 5436 23582 6050
rect 23633 5831 23667 6134
rect 23864 5831 23898 6042
rect 24808 6016 24842 6374
rect 25082 6351 25172 6374
rect 25206 6383 25530 6385
rect 25206 6351 25291 6383
rect 25082 6349 25291 6351
rect 25325 6374 25530 6383
rect 25582 6374 25616 6393
rect 25754 6571 25800 6691
rect 25854 6687 25900 6703
rect 26051 6773 26103 6811
rect 26051 6739 26069 6773
rect 26139 6803 26205 6845
rect 26380 6843 26409 6877
rect 26443 6843 26501 6877
rect 26535 6843 26593 6877
rect 26627 6843 26656 6877
rect 26816 6862 26864 6874
rect 27078 6866 27094 6900
rect 27128 6866 27144 6900
rect 27444 6890 27494 6960
rect 28934 6934 28968 6950
rect 29030 7056 29064 7072
rect 29126 7058 29160 7072
rect 29244 7058 29464 7080
rect 29124 7056 29464 7058
rect 29124 7022 29126 7056
rect 29160 7044 29464 7056
rect 29160 7022 29280 7044
rect 29030 6986 29064 7020
rect 29125 7020 29126 7022
rect 29125 6986 29160 7020
rect 29428 6996 29464 7044
rect 29125 6985 29126 6986
rect 29030 6934 29064 6950
rect 29126 6934 29160 6950
rect 29332 6960 29464 6996
rect 30822 7056 30856 7072
rect 30822 6986 30856 7020
rect 27444 6876 27454 6890
rect 26139 6769 26155 6803
rect 26189 6769 26205 6803
rect 26241 6790 26275 6811
rect 26051 6710 26103 6739
rect 26241 6735 26275 6756
rect 25834 6619 25850 6653
rect 25884 6642 25900 6653
rect 25834 6608 25852 6619
rect 25886 6608 25900 6642
rect 26051 6638 26087 6710
rect 26142 6701 26275 6735
rect 26446 6797 26512 6809
rect 26446 6763 26462 6797
rect 26496 6763 26512 6797
rect 26446 6746 26512 6763
rect 26142 6650 26176 6701
rect 26446 6695 26462 6746
rect 26496 6695 26512 6746
rect 26446 6683 26512 6695
rect 26546 6797 26592 6843
rect 26580 6763 26592 6797
rect 26546 6729 26592 6763
rect 26580 6695 26592 6729
rect 26816 6828 26822 6862
rect 26856 6828 26864 6862
rect 27448 6856 27454 6876
rect 27488 6856 27494 6890
rect 27448 6846 27494 6856
rect 27576 6851 27605 6885
rect 27639 6851 27697 6885
rect 27731 6851 27789 6885
rect 27823 6851 27852 6885
rect 26816 6740 26864 6828
rect 27190 6785 27206 6819
rect 27240 6818 27256 6819
rect 27240 6786 27402 6818
rect 27642 6810 27708 6817
rect 27636 6805 27708 6810
rect 27636 6786 27658 6805
rect 27240 6785 27658 6786
rect 27190 6782 27658 6785
rect 27366 6771 27658 6782
rect 27692 6771 27708 6805
rect 27366 6750 27708 6771
rect 27062 6740 27096 6742
rect 26816 6723 27096 6740
rect 26816 6706 27062 6723
rect 25834 6605 25900 6608
rect 26046 6636 26087 6638
rect 26046 6602 26048 6636
rect 26082 6602 26087 6636
rect 26046 6600 26087 6602
rect 25754 6553 25820 6571
rect 25754 6519 25770 6553
rect 25804 6519 25820 6553
rect 25754 6485 25820 6519
rect 25754 6451 25770 6485
rect 25804 6451 25820 6485
rect 25754 6417 25820 6451
rect 25754 6383 25770 6417
rect 25804 6383 25820 6417
rect 25754 6375 25820 6383
rect 25854 6553 25896 6569
rect 25888 6519 25896 6553
rect 25854 6485 25896 6519
rect 25888 6451 25896 6485
rect 25854 6417 25896 6451
rect 25888 6383 25896 6417
rect 25325 6349 25364 6374
rect 24876 6297 24892 6331
rect 24926 6297 24942 6331
rect 25082 6310 25364 6349
rect 25854 6341 25896 6383
rect 26051 6550 26087 6600
rect 26121 6634 26176 6650
rect 26155 6600 26176 6634
rect 26121 6584 26176 6600
rect 26221 6648 26289 6665
rect 26221 6647 26241 6648
rect 26221 6613 26239 6647
rect 26275 6614 26289 6648
rect 26273 6613 26289 6614
rect 26221 6591 26289 6613
rect 26142 6555 26176 6584
rect 26446 6563 26492 6683
rect 26546 6679 26592 6695
rect 26764 6658 26780 6659
rect 26526 6611 26542 6645
rect 26576 6638 26592 6645
rect 26644 6638 26780 6658
rect 26576 6625 26780 6638
rect 26814 6625 26830 6659
rect 26576 6624 26830 6625
rect 26576 6611 26684 6624
rect 26764 6622 26830 6624
rect 27062 6655 27096 6657
rect 26526 6597 26684 6611
rect 26540 6596 26684 6597
rect 27062 6619 27096 6621
rect 26736 6563 26770 6582
rect 26051 6500 26105 6550
rect 26142 6521 26277 6555
rect 26051 6466 26069 6500
rect 26103 6466 26105 6500
rect 26241 6487 26277 6521
rect 26051 6419 26105 6466
rect 26051 6385 26069 6419
rect 26103 6385 26105 6419
rect 26051 6369 26105 6385
rect 26139 6453 26155 6487
rect 26189 6453 26205 6487
rect 26139 6419 26205 6453
rect 26139 6385 26155 6419
rect 26189 6385 26205 6419
rect 25250 6308 25364 6310
rect 25522 6297 25538 6331
rect 25572 6297 25588 6331
rect 25688 6307 25717 6341
rect 25751 6307 25809 6341
rect 25843 6307 25901 6341
rect 25935 6307 25964 6341
rect 26139 6335 26205 6385
rect 26275 6453 26277 6487
rect 26241 6419 26277 6453
rect 26275 6385 26277 6419
rect 26241 6369 26277 6385
rect 26446 6545 26512 6563
rect 26446 6511 26462 6545
rect 26496 6511 26512 6545
rect 26446 6477 26512 6511
rect 26446 6443 26462 6477
rect 26496 6443 26512 6477
rect 26446 6409 26512 6443
rect 26446 6375 26462 6409
rect 26496 6375 26512 6409
rect 26446 6367 26512 6375
rect 26546 6545 26588 6561
rect 26580 6511 26588 6545
rect 26546 6477 26588 6511
rect 26580 6443 26588 6477
rect 26546 6409 26588 6443
rect 26736 6495 26770 6497
rect 26736 6459 26770 6461
rect 26580 6375 26588 6409
rect 25855 6300 25889 6307
rect 26034 6301 26063 6335
rect 26097 6301 26155 6335
rect 26189 6301 26247 6335
rect 26281 6301 26310 6335
rect 26546 6333 26588 6375
rect 26696 6393 26736 6414
rect 26824 6563 26858 6582
rect 27062 6534 27096 6553
rect 27158 6723 27192 6742
rect 27158 6655 27192 6657
rect 27158 6619 27192 6621
rect 27158 6534 27192 6553
rect 27254 6723 27288 6742
rect 27642 6737 27708 6750
rect 27642 6703 27658 6737
rect 27692 6703 27708 6737
rect 27642 6691 27708 6703
rect 27742 6805 27788 6851
rect 27922 6845 27951 6879
rect 27985 6845 28043 6879
rect 28077 6845 28135 6879
rect 28169 6845 28198 6879
rect 27776 6771 27788 6805
rect 27742 6737 27788 6771
rect 27776 6703 27788 6737
rect 27254 6655 27288 6657
rect 27410 6625 27426 6659
rect 27460 6625 27476 6659
rect 27254 6619 27288 6621
rect 27254 6534 27288 6553
rect 27382 6563 27416 6582
rect 26824 6495 26858 6497
rect 27382 6495 27416 6497
rect 26824 6459 26858 6461
rect 27094 6457 27110 6491
rect 27144 6457 27160 6491
rect 27382 6459 27416 6461
rect 26770 6393 26772 6414
rect 26696 6374 26772 6393
rect 26858 6393 27382 6418
rect 27470 6563 27504 6582
rect 27470 6495 27504 6497
rect 27470 6459 27504 6461
rect 27416 6393 27418 6418
rect 26824 6385 27418 6393
rect 26824 6374 27060 6385
rect 26380 6299 26409 6333
rect 26443 6299 26501 6333
rect 26535 6299 26593 6333
rect 26627 6299 26656 6333
rect 24942 6212 24988 6218
rect 24942 6210 25430 6212
rect 24942 6176 24950 6210
rect 24984 6193 25430 6210
rect 24984 6188 25380 6193
rect 24984 6178 25259 6188
rect 24984 6176 24988 6178
rect 24942 6174 24988 6176
rect 25160 6154 25259 6178
rect 25293 6159 25380 6188
rect 25414 6168 25430 6193
rect 25414 6159 25555 6168
rect 25293 6154 25555 6159
rect 25160 6134 25555 6154
rect 25284 6050 25300 6084
rect 25334 6050 25470 6084
rect 24808 6000 25190 6016
rect 24808 5976 25156 6000
rect 25156 5930 25190 5964
rect 25156 5878 25190 5894
rect 25252 6000 25286 6016
rect 25252 5930 25286 5964
rect 25252 5878 25286 5894
rect 25348 6000 25382 6016
rect 25348 5930 25382 5964
rect 25348 5878 25382 5894
rect 23622 5797 23651 5831
rect 23685 5797 23743 5831
rect 23777 5797 23835 5831
rect 23869 5797 23898 5831
rect 24696 5797 24725 5831
rect 24759 5797 24817 5831
rect 24851 5797 24909 5831
rect 24943 5797 24972 5831
rect 25188 5810 25204 5844
rect 25238 5810 25254 5844
rect 23641 5753 23695 5797
rect 23641 5719 23661 5753
rect 23641 5685 23695 5719
rect 23641 5651 23661 5685
rect 23641 5635 23695 5651
rect 23729 5753 23795 5763
rect 23729 5719 23745 5753
rect 23779 5719 23795 5753
rect 23729 5710 23795 5719
rect 23729 5685 23747 5710
rect 23729 5651 23745 5685
rect 23781 5676 23795 5710
rect 23779 5651 23795 5676
rect 23729 5635 23795 5651
rect 23829 5753 23877 5797
rect 23863 5719 23877 5753
rect 23829 5685 23877 5719
rect 23863 5651 23877 5685
rect 23829 5635 23877 5651
rect 24715 5753 24769 5797
rect 24715 5719 24735 5753
rect 24715 5685 24769 5719
rect 24715 5651 24735 5685
rect 24715 5635 24769 5651
rect 24803 5753 24869 5763
rect 24803 5719 24819 5753
rect 24853 5719 24869 5753
rect 24803 5715 24869 5719
rect 24803 5681 24817 5715
rect 24851 5685 24869 5715
rect 24803 5651 24819 5681
rect 24853 5651 24869 5685
rect 24803 5635 24869 5651
rect 24903 5753 24951 5797
rect 24937 5719 24951 5753
rect 25300 5729 25316 5763
rect 25350 5729 25366 5763
rect 24903 5685 24951 5719
rect 24937 5651 24951 5685
rect 24903 5635 24951 5651
rect 25172 5667 25206 5686
rect 23639 5594 23659 5599
rect 23639 5560 23656 5594
rect 23693 5565 23709 5599
rect 23690 5560 23709 5565
rect 23639 5549 23709 5560
rect 23743 5515 23777 5635
rect 23811 5565 23827 5599
rect 23861 5590 23881 5599
rect 23811 5556 23829 5565
rect 23863 5556 23881 5590
rect 23811 5549 23881 5556
rect 24713 5592 24733 5599
rect 24713 5558 24731 5592
rect 24767 5565 24783 5599
rect 24765 5558 24783 5565
rect 24713 5549 24783 5558
rect 24817 5515 24851 5635
rect 25172 5599 25206 5601
rect 24885 5565 24901 5599
rect 24935 5592 24955 5599
rect 24885 5558 24905 5565
rect 24939 5558 24955 5592
rect 24885 5549 24955 5558
rect 25172 5563 25206 5565
rect 23316 5435 23582 5436
rect 23316 5401 23332 5435
rect 23366 5401 23582 5435
rect 23316 5400 23582 5401
rect 23641 5499 23707 5515
rect 23641 5465 23673 5499
rect 23743 5499 23879 5515
rect 23743 5481 23829 5499
rect 23641 5431 23707 5465
rect 22999 5363 23065 5397
rect 22999 5329 23015 5363
rect 23049 5329 23065 5363
rect 23641 5397 23673 5431
rect 23641 5363 23707 5397
rect 22999 5324 23065 5329
rect 23192 5329 23474 5362
rect 23192 5295 23282 5329
rect 23316 5327 23474 5329
rect 23316 5295 23401 5327
rect 23192 5293 23401 5295
rect 23435 5293 23474 5327
rect 23192 5287 23474 5293
rect 23641 5329 23673 5363
rect 23641 5287 23707 5329
rect 23813 5465 23829 5481
rect 23863 5465 23879 5499
rect 23813 5431 23879 5465
rect 23813 5397 23829 5431
rect 23863 5397 23879 5431
rect 23813 5363 23879 5397
rect 23813 5329 23829 5363
rect 23863 5329 23879 5363
rect 23813 5324 23879 5329
rect 24715 5499 24781 5515
rect 24715 5465 24747 5499
rect 24817 5499 24953 5515
rect 24817 5481 24903 5499
rect 24715 5431 24781 5465
rect 24715 5397 24747 5431
rect 24715 5363 24781 5397
rect 24715 5329 24747 5363
rect 24715 5287 24781 5329
rect 24887 5465 24903 5481
rect 24937 5465 24953 5499
rect 25172 5478 25206 5497
rect 25268 5667 25302 5686
rect 25268 5599 25302 5601
rect 25268 5563 25302 5565
rect 25268 5478 25302 5497
rect 25364 5667 25398 5686
rect 25364 5599 25398 5601
rect 25364 5563 25398 5565
rect 25364 5478 25398 5497
rect 24887 5431 24953 5465
rect 24887 5397 24903 5431
rect 24937 5397 24953 5431
rect 25204 5436 25270 5438
rect 25436 5436 25470 6050
rect 25521 5831 25555 6134
rect 25752 5831 25786 6042
rect 26696 6016 26730 6374
rect 26970 6351 27060 6374
rect 27094 6383 27418 6385
rect 27094 6351 27179 6383
rect 26970 6349 27179 6351
rect 27213 6374 27418 6383
rect 27470 6374 27504 6393
rect 27642 6571 27688 6691
rect 27742 6687 27788 6703
rect 27939 6773 27991 6811
rect 27939 6739 27957 6773
rect 28027 6803 28093 6845
rect 28268 6843 28297 6877
rect 28331 6843 28389 6877
rect 28423 6843 28481 6877
rect 28515 6843 28544 6877
rect 28704 6862 28752 6874
rect 28966 6866 28982 6900
rect 29016 6866 29032 6900
rect 29332 6890 29382 6960
rect 30822 6934 30856 6950
rect 30918 7056 30952 7072
rect 31014 7058 31048 7072
rect 31132 7058 31352 7080
rect 31012 7056 31352 7058
rect 31012 7022 31014 7056
rect 31048 7044 31352 7056
rect 31048 7022 31168 7044
rect 30918 6986 30952 7020
rect 31013 7020 31014 7022
rect 31013 6986 31048 7020
rect 31316 6996 31352 7044
rect 31013 6985 31014 6986
rect 30918 6934 30952 6950
rect 31014 6934 31048 6950
rect 31220 6960 31352 6996
rect 32710 7056 32744 7072
rect 32710 6986 32744 7020
rect 29332 6876 29342 6890
rect 28027 6769 28043 6803
rect 28077 6769 28093 6803
rect 28129 6790 28163 6811
rect 27939 6710 27991 6739
rect 28129 6735 28163 6756
rect 27722 6619 27738 6653
rect 27772 6642 27788 6653
rect 27722 6608 27740 6619
rect 27774 6608 27788 6642
rect 27939 6638 27975 6710
rect 28030 6701 28163 6735
rect 28334 6797 28400 6809
rect 28334 6763 28350 6797
rect 28384 6763 28400 6797
rect 28334 6746 28400 6763
rect 28030 6650 28064 6701
rect 28334 6695 28350 6746
rect 28384 6695 28400 6746
rect 28334 6683 28400 6695
rect 28434 6797 28480 6843
rect 28468 6763 28480 6797
rect 28434 6729 28480 6763
rect 28468 6695 28480 6729
rect 28704 6828 28710 6862
rect 28744 6828 28752 6862
rect 29336 6856 29342 6876
rect 29376 6856 29382 6890
rect 29336 6846 29382 6856
rect 29464 6851 29493 6885
rect 29527 6851 29585 6885
rect 29619 6851 29677 6885
rect 29711 6851 29740 6885
rect 28704 6740 28752 6828
rect 29078 6785 29094 6819
rect 29128 6818 29144 6819
rect 29128 6786 29290 6818
rect 29530 6810 29596 6817
rect 29524 6805 29596 6810
rect 29524 6786 29546 6805
rect 29128 6785 29546 6786
rect 29078 6782 29546 6785
rect 29254 6771 29546 6782
rect 29580 6771 29596 6805
rect 29254 6750 29596 6771
rect 28950 6740 28984 6742
rect 28704 6723 28984 6740
rect 28704 6706 28950 6723
rect 27722 6605 27788 6608
rect 27934 6636 27975 6638
rect 27934 6602 27936 6636
rect 27970 6602 27975 6636
rect 27934 6600 27975 6602
rect 27642 6553 27708 6571
rect 27642 6519 27658 6553
rect 27692 6519 27708 6553
rect 27642 6485 27708 6519
rect 27642 6451 27658 6485
rect 27692 6451 27708 6485
rect 27642 6417 27708 6451
rect 27642 6383 27658 6417
rect 27692 6383 27708 6417
rect 27642 6375 27708 6383
rect 27742 6553 27784 6569
rect 27776 6519 27784 6553
rect 27742 6485 27784 6519
rect 27776 6451 27784 6485
rect 27742 6417 27784 6451
rect 27776 6383 27784 6417
rect 27213 6349 27252 6374
rect 26764 6297 26780 6331
rect 26814 6297 26830 6331
rect 26970 6310 27252 6349
rect 27742 6341 27784 6383
rect 27939 6550 27975 6600
rect 28009 6634 28064 6650
rect 28043 6600 28064 6634
rect 28009 6584 28064 6600
rect 28109 6648 28177 6665
rect 28109 6647 28129 6648
rect 28109 6613 28127 6647
rect 28163 6614 28177 6648
rect 28161 6613 28177 6614
rect 28109 6591 28177 6613
rect 28030 6555 28064 6584
rect 28334 6563 28380 6683
rect 28434 6679 28480 6695
rect 28652 6658 28668 6659
rect 28414 6611 28430 6645
rect 28464 6638 28480 6645
rect 28532 6638 28668 6658
rect 28464 6625 28668 6638
rect 28702 6625 28718 6659
rect 28464 6624 28718 6625
rect 28464 6611 28572 6624
rect 28652 6622 28718 6624
rect 28950 6655 28984 6657
rect 28414 6597 28572 6611
rect 28428 6596 28572 6597
rect 28950 6619 28984 6621
rect 28624 6563 28658 6582
rect 27939 6500 27993 6550
rect 28030 6521 28165 6555
rect 27939 6466 27957 6500
rect 27991 6466 27993 6500
rect 28129 6487 28165 6521
rect 27939 6419 27993 6466
rect 27939 6385 27957 6419
rect 27991 6385 27993 6419
rect 27939 6369 27993 6385
rect 28027 6453 28043 6487
rect 28077 6453 28093 6487
rect 28027 6419 28093 6453
rect 28027 6385 28043 6419
rect 28077 6385 28093 6419
rect 27138 6308 27252 6310
rect 27410 6297 27426 6331
rect 27460 6297 27476 6331
rect 27576 6307 27605 6341
rect 27639 6307 27697 6341
rect 27731 6307 27789 6341
rect 27823 6307 27852 6341
rect 28027 6335 28093 6385
rect 28163 6453 28165 6487
rect 28129 6419 28165 6453
rect 28163 6385 28165 6419
rect 28129 6369 28165 6385
rect 28334 6545 28400 6563
rect 28334 6511 28350 6545
rect 28384 6511 28400 6545
rect 28334 6477 28400 6511
rect 28334 6443 28350 6477
rect 28384 6443 28400 6477
rect 28334 6409 28400 6443
rect 28334 6375 28350 6409
rect 28384 6375 28400 6409
rect 28334 6367 28400 6375
rect 28434 6545 28476 6561
rect 28468 6511 28476 6545
rect 28434 6477 28476 6511
rect 28468 6443 28476 6477
rect 28434 6409 28476 6443
rect 28624 6495 28658 6497
rect 28624 6459 28658 6461
rect 28468 6375 28476 6409
rect 27743 6300 27777 6307
rect 27922 6301 27951 6335
rect 27985 6301 28043 6335
rect 28077 6301 28135 6335
rect 28169 6301 28198 6335
rect 28434 6333 28476 6375
rect 28584 6393 28624 6414
rect 28712 6563 28746 6582
rect 28950 6534 28984 6553
rect 29046 6723 29080 6742
rect 29046 6655 29080 6657
rect 29046 6619 29080 6621
rect 29046 6534 29080 6553
rect 29142 6723 29176 6742
rect 29530 6737 29596 6750
rect 29530 6703 29546 6737
rect 29580 6703 29596 6737
rect 29530 6691 29596 6703
rect 29630 6805 29676 6851
rect 29810 6845 29839 6879
rect 29873 6845 29931 6879
rect 29965 6845 30023 6879
rect 30057 6845 30086 6879
rect 29664 6771 29676 6805
rect 29630 6737 29676 6771
rect 29664 6703 29676 6737
rect 29142 6655 29176 6657
rect 29298 6625 29314 6659
rect 29348 6625 29364 6659
rect 29142 6619 29176 6621
rect 29142 6534 29176 6553
rect 29270 6563 29304 6582
rect 28712 6495 28746 6497
rect 29270 6495 29304 6497
rect 28712 6459 28746 6461
rect 28982 6457 28998 6491
rect 29032 6457 29048 6491
rect 29270 6459 29304 6461
rect 28658 6393 28660 6414
rect 28584 6374 28660 6393
rect 28746 6393 29270 6418
rect 29358 6563 29392 6582
rect 29358 6495 29392 6497
rect 29358 6459 29392 6461
rect 29304 6393 29306 6418
rect 28712 6385 29306 6393
rect 28712 6374 28948 6385
rect 28268 6299 28297 6333
rect 28331 6299 28389 6333
rect 28423 6299 28481 6333
rect 28515 6299 28544 6333
rect 26830 6212 26876 6218
rect 26830 6210 27318 6212
rect 26830 6176 26838 6210
rect 26872 6193 27318 6210
rect 26872 6188 27268 6193
rect 26872 6178 27147 6188
rect 26872 6176 26876 6178
rect 26830 6174 26876 6176
rect 27048 6154 27147 6178
rect 27181 6159 27268 6188
rect 27302 6168 27318 6193
rect 27302 6159 27443 6168
rect 27181 6154 27443 6159
rect 27048 6134 27443 6154
rect 27172 6050 27188 6084
rect 27222 6050 27358 6084
rect 26696 6000 27078 6016
rect 26696 5976 27044 6000
rect 27044 5930 27078 5964
rect 27044 5878 27078 5894
rect 27140 6000 27174 6016
rect 27140 5930 27174 5964
rect 27140 5878 27174 5894
rect 27236 6000 27270 6016
rect 27236 5930 27270 5964
rect 27236 5878 27270 5894
rect 25510 5797 25539 5831
rect 25573 5797 25631 5831
rect 25665 5797 25723 5831
rect 25757 5797 25786 5831
rect 26584 5797 26613 5831
rect 26647 5797 26705 5831
rect 26739 5797 26797 5831
rect 26831 5797 26860 5831
rect 27076 5810 27092 5844
rect 27126 5810 27142 5844
rect 25529 5753 25583 5797
rect 25529 5719 25549 5753
rect 25529 5685 25583 5719
rect 25529 5651 25549 5685
rect 25529 5635 25583 5651
rect 25617 5753 25683 5763
rect 25617 5719 25633 5753
rect 25667 5719 25683 5753
rect 25617 5710 25683 5719
rect 25617 5685 25635 5710
rect 25617 5651 25633 5685
rect 25669 5676 25683 5710
rect 25667 5651 25683 5676
rect 25617 5635 25683 5651
rect 25717 5753 25765 5797
rect 25751 5719 25765 5753
rect 25717 5685 25765 5719
rect 25751 5651 25765 5685
rect 25717 5635 25765 5651
rect 26603 5753 26657 5797
rect 26603 5719 26623 5753
rect 26603 5685 26657 5719
rect 26603 5651 26623 5685
rect 26603 5635 26657 5651
rect 26691 5753 26757 5763
rect 26691 5719 26707 5753
rect 26741 5719 26757 5753
rect 26691 5715 26757 5719
rect 26691 5681 26705 5715
rect 26739 5685 26757 5715
rect 26691 5651 26707 5681
rect 26741 5651 26757 5685
rect 26691 5635 26757 5651
rect 26791 5753 26839 5797
rect 26825 5719 26839 5753
rect 27188 5729 27204 5763
rect 27238 5729 27254 5763
rect 26791 5685 26839 5719
rect 26825 5651 26839 5685
rect 26791 5635 26839 5651
rect 27060 5667 27094 5686
rect 25527 5594 25547 5599
rect 25527 5560 25544 5594
rect 25581 5565 25597 5599
rect 25578 5560 25597 5565
rect 25527 5549 25597 5560
rect 25631 5515 25665 5635
rect 25699 5565 25715 5599
rect 25749 5590 25769 5599
rect 25699 5556 25717 5565
rect 25751 5556 25769 5590
rect 25699 5549 25769 5556
rect 26601 5592 26621 5599
rect 26601 5558 26619 5592
rect 26655 5565 26671 5599
rect 26653 5558 26671 5565
rect 26601 5549 26671 5558
rect 26705 5515 26739 5635
rect 27060 5599 27094 5601
rect 26773 5565 26789 5599
rect 26823 5592 26843 5599
rect 26773 5558 26793 5565
rect 26827 5558 26843 5592
rect 26773 5549 26843 5558
rect 27060 5563 27094 5565
rect 25204 5435 25470 5436
rect 25204 5401 25220 5435
rect 25254 5401 25470 5435
rect 25204 5400 25470 5401
rect 25529 5499 25595 5515
rect 25529 5465 25561 5499
rect 25631 5499 25767 5515
rect 25631 5481 25717 5499
rect 25529 5431 25595 5465
rect 24887 5363 24953 5397
rect 24887 5329 24903 5363
rect 24937 5329 24953 5363
rect 25529 5397 25561 5431
rect 25529 5363 25595 5397
rect 24887 5324 24953 5329
rect 25080 5329 25362 5362
rect 25080 5295 25170 5329
rect 25204 5327 25362 5329
rect 25204 5295 25289 5327
rect 25080 5293 25289 5295
rect 25323 5293 25362 5327
rect 25080 5287 25362 5293
rect 25529 5329 25561 5363
rect 25529 5287 25595 5329
rect 25701 5465 25717 5481
rect 25751 5465 25767 5499
rect 25701 5431 25767 5465
rect 25701 5397 25717 5431
rect 25751 5397 25767 5431
rect 25701 5363 25767 5397
rect 25701 5329 25717 5363
rect 25751 5329 25767 5363
rect 25701 5324 25767 5329
rect 26603 5499 26669 5515
rect 26603 5465 26635 5499
rect 26705 5499 26841 5515
rect 26705 5481 26791 5499
rect 26603 5431 26669 5465
rect 26603 5397 26635 5431
rect 26603 5363 26669 5397
rect 26603 5329 26635 5363
rect 26603 5287 26669 5329
rect 26775 5465 26791 5481
rect 26825 5465 26841 5499
rect 27060 5478 27094 5497
rect 27156 5667 27190 5686
rect 27156 5599 27190 5601
rect 27156 5563 27190 5565
rect 27156 5478 27190 5497
rect 27252 5667 27286 5686
rect 27252 5599 27286 5601
rect 27252 5563 27286 5565
rect 27252 5478 27286 5497
rect 26775 5431 26841 5465
rect 26775 5397 26791 5431
rect 26825 5397 26841 5431
rect 27092 5436 27158 5438
rect 27324 5436 27358 6050
rect 27409 5831 27443 6134
rect 27640 5831 27674 6042
rect 28584 6016 28618 6374
rect 28858 6351 28948 6374
rect 28982 6383 29306 6385
rect 28982 6351 29067 6383
rect 28858 6349 29067 6351
rect 29101 6374 29306 6383
rect 29358 6374 29392 6393
rect 29530 6571 29576 6691
rect 29630 6687 29676 6703
rect 29827 6773 29879 6811
rect 29827 6739 29845 6773
rect 29915 6803 29981 6845
rect 30156 6843 30185 6877
rect 30219 6843 30277 6877
rect 30311 6843 30369 6877
rect 30403 6843 30432 6877
rect 30592 6862 30640 6874
rect 30854 6866 30870 6900
rect 30904 6866 30920 6900
rect 31220 6890 31270 6960
rect 32710 6934 32744 6950
rect 32806 7056 32840 7072
rect 32902 7058 32936 7072
rect 33020 7058 33240 7080
rect 32900 7056 33240 7058
rect 32900 7022 32902 7056
rect 32936 7044 33240 7056
rect 32936 7022 33056 7044
rect 32806 6986 32840 7020
rect 32901 7020 32902 7022
rect 32901 6986 32936 7020
rect 33204 6996 33240 7044
rect 32901 6985 32902 6986
rect 32806 6934 32840 6950
rect 32902 6934 32936 6950
rect 33108 6960 33240 6996
rect 34598 7056 34632 7072
rect 34598 6986 34632 7020
rect 31220 6876 31230 6890
rect 29915 6769 29931 6803
rect 29965 6769 29981 6803
rect 30017 6790 30051 6811
rect 29827 6710 29879 6739
rect 30017 6735 30051 6756
rect 29610 6619 29626 6653
rect 29660 6642 29676 6653
rect 29610 6608 29628 6619
rect 29662 6608 29676 6642
rect 29827 6638 29863 6710
rect 29918 6701 30051 6735
rect 30222 6797 30288 6809
rect 30222 6763 30238 6797
rect 30272 6763 30288 6797
rect 30222 6746 30288 6763
rect 29918 6650 29952 6701
rect 30222 6695 30238 6746
rect 30272 6695 30288 6746
rect 30222 6683 30288 6695
rect 30322 6797 30368 6843
rect 30356 6763 30368 6797
rect 30322 6729 30368 6763
rect 30356 6695 30368 6729
rect 30592 6828 30598 6862
rect 30632 6828 30640 6862
rect 31224 6856 31230 6876
rect 31264 6856 31270 6890
rect 31224 6846 31270 6856
rect 31352 6851 31381 6885
rect 31415 6851 31473 6885
rect 31507 6851 31565 6885
rect 31599 6851 31628 6885
rect 30592 6740 30640 6828
rect 30966 6785 30982 6819
rect 31016 6818 31032 6819
rect 31016 6786 31178 6818
rect 31418 6810 31484 6817
rect 31412 6805 31484 6810
rect 31412 6786 31434 6805
rect 31016 6785 31434 6786
rect 30966 6782 31434 6785
rect 31142 6771 31434 6782
rect 31468 6771 31484 6805
rect 31142 6750 31484 6771
rect 30838 6740 30872 6742
rect 30592 6723 30872 6740
rect 30592 6706 30838 6723
rect 29610 6605 29676 6608
rect 29822 6636 29863 6638
rect 29822 6602 29824 6636
rect 29858 6602 29863 6636
rect 29822 6600 29863 6602
rect 29530 6553 29596 6571
rect 29530 6519 29546 6553
rect 29580 6519 29596 6553
rect 29530 6485 29596 6519
rect 29530 6451 29546 6485
rect 29580 6451 29596 6485
rect 29530 6417 29596 6451
rect 29530 6383 29546 6417
rect 29580 6383 29596 6417
rect 29530 6375 29596 6383
rect 29630 6553 29672 6569
rect 29664 6519 29672 6553
rect 29630 6485 29672 6519
rect 29664 6451 29672 6485
rect 29630 6417 29672 6451
rect 29664 6383 29672 6417
rect 29101 6349 29140 6374
rect 28652 6297 28668 6331
rect 28702 6297 28718 6331
rect 28858 6310 29140 6349
rect 29630 6341 29672 6383
rect 29827 6550 29863 6600
rect 29897 6634 29952 6650
rect 29931 6600 29952 6634
rect 29897 6584 29952 6600
rect 29997 6648 30065 6665
rect 29997 6647 30017 6648
rect 29997 6613 30015 6647
rect 30051 6614 30065 6648
rect 30049 6613 30065 6614
rect 29997 6591 30065 6613
rect 29918 6555 29952 6584
rect 30222 6563 30268 6683
rect 30322 6679 30368 6695
rect 30540 6658 30556 6659
rect 30302 6611 30318 6645
rect 30352 6638 30368 6645
rect 30420 6638 30556 6658
rect 30352 6625 30556 6638
rect 30590 6625 30606 6659
rect 30352 6624 30606 6625
rect 30352 6611 30460 6624
rect 30540 6622 30606 6624
rect 30838 6655 30872 6657
rect 30302 6597 30460 6611
rect 30316 6596 30460 6597
rect 30838 6619 30872 6621
rect 30512 6563 30546 6582
rect 29827 6500 29881 6550
rect 29918 6521 30053 6555
rect 29827 6466 29845 6500
rect 29879 6466 29881 6500
rect 30017 6487 30053 6521
rect 29827 6419 29881 6466
rect 29827 6385 29845 6419
rect 29879 6385 29881 6419
rect 29827 6369 29881 6385
rect 29915 6453 29931 6487
rect 29965 6453 29981 6487
rect 29915 6419 29981 6453
rect 29915 6385 29931 6419
rect 29965 6385 29981 6419
rect 29026 6308 29140 6310
rect 29298 6297 29314 6331
rect 29348 6297 29364 6331
rect 29464 6307 29493 6341
rect 29527 6307 29585 6341
rect 29619 6307 29677 6341
rect 29711 6307 29740 6341
rect 29915 6335 29981 6385
rect 30051 6453 30053 6487
rect 30017 6419 30053 6453
rect 30051 6385 30053 6419
rect 30017 6369 30053 6385
rect 30222 6545 30288 6563
rect 30222 6511 30238 6545
rect 30272 6511 30288 6545
rect 30222 6477 30288 6511
rect 30222 6443 30238 6477
rect 30272 6443 30288 6477
rect 30222 6409 30288 6443
rect 30222 6375 30238 6409
rect 30272 6375 30288 6409
rect 30222 6367 30288 6375
rect 30322 6545 30364 6561
rect 30356 6511 30364 6545
rect 30322 6477 30364 6511
rect 30356 6443 30364 6477
rect 30322 6409 30364 6443
rect 30512 6495 30546 6497
rect 30512 6459 30546 6461
rect 30356 6375 30364 6409
rect 29631 6300 29665 6307
rect 29810 6301 29839 6335
rect 29873 6301 29931 6335
rect 29965 6301 30023 6335
rect 30057 6301 30086 6335
rect 30322 6333 30364 6375
rect 30472 6393 30512 6414
rect 30600 6563 30634 6582
rect 30838 6534 30872 6553
rect 30934 6723 30968 6742
rect 30934 6655 30968 6657
rect 30934 6619 30968 6621
rect 30934 6534 30968 6553
rect 31030 6723 31064 6742
rect 31418 6737 31484 6750
rect 31418 6703 31434 6737
rect 31468 6703 31484 6737
rect 31418 6691 31484 6703
rect 31518 6805 31564 6851
rect 31698 6845 31727 6879
rect 31761 6845 31819 6879
rect 31853 6845 31911 6879
rect 31945 6845 31974 6879
rect 31552 6771 31564 6805
rect 31518 6737 31564 6771
rect 31552 6703 31564 6737
rect 31030 6655 31064 6657
rect 31186 6625 31202 6659
rect 31236 6625 31252 6659
rect 31030 6619 31064 6621
rect 31030 6534 31064 6553
rect 31158 6563 31192 6582
rect 30600 6495 30634 6497
rect 31158 6495 31192 6497
rect 30600 6459 30634 6461
rect 30870 6457 30886 6491
rect 30920 6457 30936 6491
rect 31158 6459 31192 6461
rect 30546 6393 30548 6414
rect 30472 6374 30548 6393
rect 30634 6393 31158 6418
rect 31246 6563 31280 6582
rect 31246 6495 31280 6497
rect 31246 6459 31280 6461
rect 31192 6393 31194 6418
rect 30600 6385 31194 6393
rect 30600 6374 30836 6385
rect 30156 6299 30185 6333
rect 30219 6299 30277 6333
rect 30311 6299 30369 6333
rect 30403 6299 30432 6333
rect 28718 6212 28764 6218
rect 28718 6210 29206 6212
rect 28718 6176 28726 6210
rect 28760 6193 29206 6210
rect 28760 6188 29156 6193
rect 28760 6178 29035 6188
rect 28760 6176 28764 6178
rect 28718 6174 28764 6176
rect 28936 6154 29035 6178
rect 29069 6159 29156 6188
rect 29190 6168 29206 6193
rect 29190 6159 29331 6168
rect 29069 6154 29331 6159
rect 28936 6134 29331 6154
rect 29060 6050 29076 6084
rect 29110 6050 29246 6084
rect 28584 6000 28966 6016
rect 28584 5976 28932 6000
rect 28932 5930 28966 5964
rect 28932 5878 28966 5894
rect 29028 6000 29062 6016
rect 29028 5930 29062 5964
rect 29028 5878 29062 5894
rect 29124 6000 29158 6016
rect 29124 5930 29158 5964
rect 29124 5878 29158 5894
rect 27398 5797 27427 5831
rect 27461 5797 27519 5831
rect 27553 5797 27611 5831
rect 27645 5797 27674 5831
rect 28472 5797 28501 5831
rect 28535 5797 28593 5831
rect 28627 5797 28685 5831
rect 28719 5797 28748 5831
rect 28964 5810 28980 5844
rect 29014 5810 29030 5844
rect 27417 5753 27471 5797
rect 27417 5719 27437 5753
rect 27417 5685 27471 5719
rect 27417 5651 27437 5685
rect 27417 5635 27471 5651
rect 27505 5753 27571 5763
rect 27505 5719 27521 5753
rect 27555 5719 27571 5753
rect 27505 5710 27571 5719
rect 27505 5685 27523 5710
rect 27505 5651 27521 5685
rect 27557 5676 27571 5710
rect 27555 5651 27571 5676
rect 27505 5635 27571 5651
rect 27605 5753 27653 5797
rect 27639 5719 27653 5753
rect 27605 5685 27653 5719
rect 27639 5651 27653 5685
rect 27605 5635 27653 5651
rect 28491 5753 28545 5797
rect 28491 5719 28511 5753
rect 28491 5685 28545 5719
rect 28491 5651 28511 5685
rect 28491 5635 28545 5651
rect 28579 5753 28645 5763
rect 28579 5719 28595 5753
rect 28629 5719 28645 5753
rect 28579 5715 28645 5719
rect 28579 5681 28593 5715
rect 28627 5685 28645 5715
rect 28579 5651 28595 5681
rect 28629 5651 28645 5685
rect 28579 5635 28645 5651
rect 28679 5753 28727 5797
rect 28713 5719 28727 5753
rect 29076 5729 29092 5763
rect 29126 5729 29142 5763
rect 28679 5685 28727 5719
rect 28713 5651 28727 5685
rect 28679 5635 28727 5651
rect 28948 5667 28982 5686
rect 27415 5594 27435 5599
rect 27415 5560 27432 5594
rect 27469 5565 27485 5599
rect 27466 5560 27485 5565
rect 27415 5549 27485 5560
rect 27519 5515 27553 5635
rect 27587 5565 27603 5599
rect 27637 5590 27657 5599
rect 27587 5556 27605 5565
rect 27639 5556 27657 5590
rect 27587 5549 27657 5556
rect 28489 5592 28509 5599
rect 28489 5558 28507 5592
rect 28543 5565 28559 5599
rect 28541 5558 28559 5565
rect 28489 5549 28559 5558
rect 28593 5515 28627 5635
rect 28948 5599 28982 5601
rect 28661 5565 28677 5599
rect 28711 5592 28731 5599
rect 28661 5558 28681 5565
rect 28715 5558 28731 5592
rect 28661 5549 28731 5558
rect 28948 5563 28982 5565
rect 27092 5435 27358 5436
rect 27092 5401 27108 5435
rect 27142 5401 27358 5435
rect 27092 5400 27358 5401
rect 27417 5499 27483 5515
rect 27417 5465 27449 5499
rect 27519 5499 27655 5515
rect 27519 5481 27605 5499
rect 27417 5431 27483 5465
rect 26775 5363 26841 5397
rect 26775 5329 26791 5363
rect 26825 5329 26841 5363
rect 27417 5397 27449 5431
rect 27417 5363 27483 5397
rect 26775 5324 26841 5329
rect 26968 5329 27250 5362
rect 26968 5295 27058 5329
rect 27092 5327 27250 5329
rect 27092 5295 27177 5327
rect 26968 5293 27177 5295
rect 27211 5293 27250 5327
rect 26968 5287 27250 5293
rect 27417 5329 27449 5363
rect 27417 5287 27483 5329
rect 27589 5465 27605 5481
rect 27639 5465 27655 5499
rect 27589 5431 27655 5465
rect 27589 5397 27605 5431
rect 27639 5397 27655 5431
rect 27589 5363 27655 5397
rect 27589 5329 27605 5363
rect 27639 5329 27655 5363
rect 27589 5324 27655 5329
rect 28491 5499 28557 5515
rect 28491 5465 28523 5499
rect 28593 5499 28729 5515
rect 28593 5481 28679 5499
rect 28491 5431 28557 5465
rect 28491 5397 28523 5431
rect 28491 5363 28557 5397
rect 28491 5329 28523 5363
rect 28491 5287 28557 5329
rect 28663 5465 28679 5481
rect 28713 5465 28729 5499
rect 28948 5478 28982 5497
rect 29044 5667 29078 5686
rect 29044 5599 29078 5601
rect 29044 5563 29078 5565
rect 29044 5478 29078 5497
rect 29140 5667 29174 5686
rect 29140 5599 29174 5601
rect 29140 5563 29174 5565
rect 29140 5478 29174 5497
rect 28663 5431 28729 5465
rect 28663 5397 28679 5431
rect 28713 5397 28729 5431
rect 28980 5436 29046 5438
rect 29212 5436 29246 6050
rect 29297 5831 29331 6134
rect 29528 5831 29562 6042
rect 30472 6016 30506 6374
rect 30746 6351 30836 6374
rect 30870 6383 31194 6385
rect 30870 6351 30955 6383
rect 30746 6349 30955 6351
rect 30989 6374 31194 6383
rect 31246 6374 31280 6393
rect 31418 6571 31464 6691
rect 31518 6687 31564 6703
rect 31715 6773 31767 6811
rect 31715 6739 31733 6773
rect 31803 6803 31869 6845
rect 32044 6843 32073 6877
rect 32107 6843 32165 6877
rect 32199 6843 32257 6877
rect 32291 6843 32320 6877
rect 32480 6862 32528 6874
rect 32742 6866 32758 6900
rect 32792 6866 32808 6900
rect 33108 6890 33158 6960
rect 34598 6934 34632 6950
rect 34694 7056 34728 7072
rect 34790 7058 34824 7072
rect 34908 7058 35128 7080
rect 34788 7056 35128 7058
rect 34788 7022 34790 7056
rect 34824 7044 35128 7056
rect 34824 7022 34944 7044
rect 34694 6986 34728 7020
rect 34789 7020 34790 7022
rect 34789 6986 34824 7020
rect 35092 6996 35128 7044
rect 34789 6985 34790 6986
rect 34694 6934 34728 6950
rect 34790 6934 34824 6950
rect 34996 6960 35128 6996
rect 36486 7056 36520 7072
rect 36486 6986 36520 7020
rect 33108 6876 33118 6890
rect 31803 6769 31819 6803
rect 31853 6769 31869 6803
rect 31905 6790 31939 6811
rect 31715 6710 31767 6739
rect 31905 6735 31939 6756
rect 31498 6619 31514 6653
rect 31548 6642 31564 6653
rect 31498 6608 31516 6619
rect 31550 6608 31564 6642
rect 31715 6638 31751 6710
rect 31806 6701 31939 6735
rect 32110 6797 32176 6809
rect 32110 6763 32126 6797
rect 32160 6763 32176 6797
rect 32110 6746 32176 6763
rect 31806 6650 31840 6701
rect 32110 6695 32126 6746
rect 32160 6695 32176 6746
rect 32110 6683 32176 6695
rect 32210 6797 32256 6843
rect 32244 6763 32256 6797
rect 32210 6729 32256 6763
rect 32244 6695 32256 6729
rect 32480 6828 32486 6862
rect 32520 6828 32528 6862
rect 33112 6856 33118 6876
rect 33152 6856 33158 6890
rect 33112 6846 33158 6856
rect 33240 6851 33269 6885
rect 33303 6851 33361 6885
rect 33395 6851 33453 6885
rect 33487 6851 33516 6885
rect 32480 6740 32528 6828
rect 32854 6785 32870 6819
rect 32904 6818 32920 6819
rect 32904 6786 33066 6818
rect 33306 6810 33372 6817
rect 33300 6805 33372 6810
rect 33300 6786 33322 6805
rect 32904 6785 33322 6786
rect 32854 6782 33322 6785
rect 33030 6771 33322 6782
rect 33356 6771 33372 6805
rect 33030 6750 33372 6771
rect 32726 6740 32760 6742
rect 32480 6723 32760 6740
rect 32480 6706 32726 6723
rect 31498 6605 31564 6608
rect 31710 6636 31751 6638
rect 31710 6602 31712 6636
rect 31746 6602 31751 6636
rect 31710 6600 31751 6602
rect 31418 6553 31484 6571
rect 31418 6519 31434 6553
rect 31468 6519 31484 6553
rect 31418 6485 31484 6519
rect 31418 6451 31434 6485
rect 31468 6451 31484 6485
rect 31418 6417 31484 6451
rect 31418 6383 31434 6417
rect 31468 6383 31484 6417
rect 31418 6375 31484 6383
rect 31518 6553 31560 6569
rect 31552 6519 31560 6553
rect 31518 6485 31560 6519
rect 31552 6451 31560 6485
rect 31518 6417 31560 6451
rect 31552 6383 31560 6417
rect 30989 6349 31028 6374
rect 30540 6297 30556 6331
rect 30590 6297 30606 6331
rect 30746 6310 31028 6349
rect 31518 6341 31560 6383
rect 31715 6550 31751 6600
rect 31785 6634 31840 6650
rect 31819 6600 31840 6634
rect 31785 6584 31840 6600
rect 31885 6648 31953 6665
rect 31885 6647 31905 6648
rect 31885 6613 31903 6647
rect 31939 6614 31953 6648
rect 31937 6613 31953 6614
rect 31885 6591 31953 6613
rect 31806 6555 31840 6584
rect 32110 6563 32156 6683
rect 32210 6679 32256 6695
rect 32428 6658 32444 6659
rect 32190 6611 32206 6645
rect 32240 6638 32256 6645
rect 32308 6638 32444 6658
rect 32240 6625 32444 6638
rect 32478 6625 32494 6659
rect 32240 6624 32494 6625
rect 32240 6611 32348 6624
rect 32428 6622 32494 6624
rect 32726 6655 32760 6657
rect 32190 6597 32348 6611
rect 32204 6596 32348 6597
rect 32726 6619 32760 6621
rect 32400 6563 32434 6582
rect 31715 6500 31769 6550
rect 31806 6521 31941 6555
rect 31715 6466 31733 6500
rect 31767 6466 31769 6500
rect 31905 6487 31941 6521
rect 31715 6419 31769 6466
rect 31715 6385 31733 6419
rect 31767 6385 31769 6419
rect 31715 6369 31769 6385
rect 31803 6453 31819 6487
rect 31853 6453 31869 6487
rect 31803 6419 31869 6453
rect 31803 6385 31819 6419
rect 31853 6385 31869 6419
rect 30914 6308 31028 6310
rect 31186 6297 31202 6331
rect 31236 6297 31252 6331
rect 31352 6307 31381 6341
rect 31415 6307 31473 6341
rect 31507 6307 31565 6341
rect 31599 6307 31628 6341
rect 31803 6335 31869 6385
rect 31939 6453 31941 6487
rect 31905 6419 31941 6453
rect 31939 6385 31941 6419
rect 31905 6369 31941 6385
rect 32110 6545 32176 6563
rect 32110 6511 32126 6545
rect 32160 6511 32176 6545
rect 32110 6477 32176 6511
rect 32110 6443 32126 6477
rect 32160 6443 32176 6477
rect 32110 6409 32176 6443
rect 32110 6375 32126 6409
rect 32160 6375 32176 6409
rect 32110 6367 32176 6375
rect 32210 6545 32252 6561
rect 32244 6511 32252 6545
rect 32210 6477 32252 6511
rect 32244 6443 32252 6477
rect 32210 6409 32252 6443
rect 32400 6495 32434 6497
rect 32400 6459 32434 6461
rect 32244 6375 32252 6409
rect 31519 6300 31553 6307
rect 31698 6301 31727 6335
rect 31761 6301 31819 6335
rect 31853 6301 31911 6335
rect 31945 6301 31974 6335
rect 32210 6333 32252 6375
rect 32360 6393 32400 6414
rect 32488 6563 32522 6582
rect 32726 6534 32760 6553
rect 32822 6723 32856 6742
rect 32822 6655 32856 6657
rect 32822 6619 32856 6621
rect 32822 6534 32856 6553
rect 32918 6723 32952 6742
rect 33306 6737 33372 6750
rect 33306 6703 33322 6737
rect 33356 6703 33372 6737
rect 33306 6691 33372 6703
rect 33406 6805 33452 6851
rect 33586 6845 33615 6879
rect 33649 6845 33707 6879
rect 33741 6845 33799 6879
rect 33833 6845 33862 6879
rect 33440 6771 33452 6805
rect 33406 6737 33452 6771
rect 33440 6703 33452 6737
rect 32918 6655 32952 6657
rect 33074 6625 33090 6659
rect 33124 6625 33140 6659
rect 32918 6619 32952 6621
rect 32918 6534 32952 6553
rect 33046 6563 33080 6582
rect 32488 6495 32522 6497
rect 33046 6495 33080 6497
rect 32488 6459 32522 6461
rect 32758 6457 32774 6491
rect 32808 6457 32824 6491
rect 33046 6459 33080 6461
rect 32434 6393 32436 6414
rect 32360 6374 32436 6393
rect 32522 6393 33046 6418
rect 33134 6563 33168 6582
rect 33134 6495 33168 6497
rect 33134 6459 33168 6461
rect 33080 6393 33082 6418
rect 32488 6385 33082 6393
rect 32488 6374 32724 6385
rect 32044 6299 32073 6333
rect 32107 6299 32165 6333
rect 32199 6299 32257 6333
rect 32291 6299 32320 6333
rect 30606 6212 30652 6218
rect 30606 6210 31094 6212
rect 30606 6176 30614 6210
rect 30648 6193 31094 6210
rect 30648 6188 31044 6193
rect 30648 6178 30923 6188
rect 30648 6176 30652 6178
rect 30606 6174 30652 6176
rect 30824 6154 30923 6178
rect 30957 6159 31044 6188
rect 31078 6168 31094 6193
rect 31078 6159 31219 6168
rect 30957 6154 31219 6159
rect 30824 6134 31219 6154
rect 30948 6050 30964 6084
rect 30998 6050 31134 6084
rect 30472 6000 30854 6016
rect 30472 5976 30820 6000
rect 30820 5930 30854 5964
rect 30820 5878 30854 5894
rect 30916 6000 30950 6016
rect 30916 5930 30950 5964
rect 30916 5878 30950 5894
rect 31012 6000 31046 6016
rect 31012 5930 31046 5964
rect 31012 5878 31046 5894
rect 29286 5797 29315 5831
rect 29349 5797 29407 5831
rect 29441 5797 29499 5831
rect 29533 5797 29562 5831
rect 30360 5797 30389 5831
rect 30423 5797 30481 5831
rect 30515 5797 30573 5831
rect 30607 5797 30636 5831
rect 30852 5810 30868 5844
rect 30902 5810 30918 5844
rect 29305 5753 29359 5797
rect 29305 5719 29325 5753
rect 29305 5685 29359 5719
rect 29305 5651 29325 5685
rect 29305 5635 29359 5651
rect 29393 5753 29459 5763
rect 29393 5719 29409 5753
rect 29443 5719 29459 5753
rect 29393 5710 29459 5719
rect 29393 5685 29411 5710
rect 29393 5651 29409 5685
rect 29445 5676 29459 5710
rect 29443 5651 29459 5676
rect 29393 5635 29459 5651
rect 29493 5753 29541 5797
rect 29527 5719 29541 5753
rect 29493 5685 29541 5719
rect 29527 5651 29541 5685
rect 29493 5635 29541 5651
rect 30379 5753 30433 5797
rect 30379 5719 30399 5753
rect 30379 5685 30433 5719
rect 30379 5651 30399 5685
rect 30379 5635 30433 5651
rect 30467 5753 30533 5763
rect 30467 5719 30483 5753
rect 30517 5719 30533 5753
rect 30467 5715 30533 5719
rect 30467 5681 30481 5715
rect 30515 5685 30533 5715
rect 30467 5651 30483 5681
rect 30517 5651 30533 5685
rect 30467 5635 30533 5651
rect 30567 5753 30615 5797
rect 30601 5719 30615 5753
rect 30964 5729 30980 5763
rect 31014 5729 31030 5763
rect 30567 5685 30615 5719
rect 30601 5651 30615 5685
rect 30567 5635 30615 5651
rect 30836 5667 30870 5686
rect 29303 5594 29323 5599
rect 29303 5560 29320 5594
rect 29357 5565 29373 5599
rect 29354 5560 29373 5565
rect 29303 5549 29373 5560
rect 29407 5515 29441 5635
rect 29475 5565 29491 5599
rect 29525 5590 29545 5599
rect 29475 5556 29493 5565
rect 29527 5556 29545 5590
rect 29475 5549 29545 5556
rect 30377 5592 30397 5599
rect 30377 5558 30395 5592
rect 30431 5565 30447 5599
rect 30429 5558 30447 5565
rect 30377 5549 30447 5558
rect 30481 5515 30515 5635
rect 30836 5599 30870 5601
rect 30549 5565 30565 5599
rect 30599 5592 30619 5599
rect 30549 5558 30569 5565
rect 30603 5558 30619 5592
rect 30549 5549 30619 5558
rect 30836 5563 30870 5565
rect 28980 5435 29246 5436
rect 28980 5401 28996 5435
rect 29030 5401 29246 5435
rect 28980 5400 29246 5401
rect 29305 5499 29371 5515
rect 29305 5465 29337 5499
rect 29407 5499 29543 5515
rect 29407 5481 29493 5499
rect 29305 5431 29371 5465
rect 28663 5363 28729 5397
rect 28663 5329 28679 5363
rect 28713 5329 28729 5363
rect 29305 5397 29337 5431
rect 29305 5363 29371 5397
rect 28663 5324 28729 5329
rect 28856 5329 29138 5362
rect 28856 5295 28946 5329
rect 28980 5327 29138 5329
rect 28980 5295 29065 5327
rect 28856 5293 29065 5295
rect 29099 5293 29138 5327
rect 28856 5287 29138 5293
rect 29305 5329 29337 5363
rect 29305 5287 29371 5329
rect 29477 5465 29493 5481
rect 29527 5465 29543 5499
rect 29477 5431 29543 5465
rect 29477 5397 29493 5431
rect 29527 5397 29543 5431
rect 29477 5363 29543 5397
rect 29477 5329 29493 5363
rect 29527 5329 29543 5363
rect 29477 5324 29543 5329
rect 30379 5499 30445 5515
rect 30379 5465 30411 5499
rect 30481 5499 30617 5515
rect 30481 5481 30567 5499
rect 30379 5431 30445 5465
rect 30379 5397 30411 5431
rect 30379 5363 30445 5397
rect 30379 5329 30411 5363
rect 30379 5287 30445 5329
rect 30551 5465 30567 5481
rect 30601 5465 30617 5499
rect 30836 5478 30870 5497
rect 30932 5667 30966 5686
rect 30932 5599 30966 5601
rect 30932 5563 30966 5565
rect 30932 5478 30966 5497
rect 31028 5667 31062 5686
rect 31028 5599 31062 5601
rect 31028 5563 31062 5565
rect 31028 5478 31062 5497
rect 30551 5431 30617 5465
rect 30551 5397 30567 5431
rect 30601 5397 30617 5431
rect 30868 5436 30934 5438
rect 31100 5436 31134 6050
rect 31185 5831 31219 6134
rect 31416 5831 31450 6042
rect 32360 6016 32394 6374
rect 32634 6351 32724 6374
rect 32758 6383 33082 6385
rect 32758 6351 32843 6383
rect 32634 6349 32843 6351
rect 32877 6374 33082 6383
rect 33134 6374 33168 6393
rect 33306 6571 33352 6691
rect 33406 6687 33452 6703
rect 33603 6773 33655 6811
rect 33603 6739 33621 6773
rect 33691 6803 33757 6845
rect 33932 6843 33961 6877
rect 33995 6843 34053 6877
rect 34087 6843 34145 6877
rect 34179 6843 34208 6877
rect 34368 6862 34416 6874
rect 34630 6866 34646 6900
rect 34680 6866 34696 6900
rect 34996 6890 35046 6960
rect 36486 6934 36520 6950
rect 36582 7056 36616 7072
rect 36678 7058 36712 7072
rect 36796 7058 37016 7080
rect 36676 7056 37016 7058
rect 36676 7022 36678 7056
rect 36712 7044 37016 7056
rect 36712 7022 36832 7044
rect 36582 6986 36616 7020
rect 36677 7020 36678 7022
rect 36677 6986 36712 7020
rect 36980 6996 37016 7044
rect 36677 6985 36678 6986
rect 36582 6934 36616 6950
rect 36678 6934 36712 6950
rect 36884 6960 37016 6996
rect 38374 7056 38408 7072
rect 38374 6986 38408 7020
rect 34996 6876 35006 6890
rect 33691 6769 33707 6803
rect 33741 6769 33757 6803
rect 33793 6790 33827 6811
rect 33603 6710 33655 6739
rect 33793 6735 33827 6756
rect 33386 6619 33402 6653
rect 33436 6642 33452 6653
rect 33386 6608 33404 6619
rect 33438 6608 33452 6642
rect 33603 6638 33639 6710
rect 33694 6701 33827 6735
rect 33998 6797 34064 6809
rect 33998 6763 34014 6797
rect 34048 6763 34064 6797
rect 33998 6746 34064 6763
rect 33694 6650 33728 6701
rect 33998 6695 34014 6746
rect 34048 6695 34064 6746
rect 33998 6683 34064 6695
rect 34098 6797 34144 6843
rect 34132 6763 34144 6797
rect 34098 6729 34144 6763
rect 34132 6695 34144 6729
rect 34368 6828 34374 6862
rect 34408 6828 34416 6862
rect 35000 6856 35006 6876
rect 35040 6856 35046 6890
rect 35000 6846 35046 6856
rect 35128 6851 35157 6885
rect 35191 6851 35249 6885
rect 35283 6851 35341 6885
rect 35375 6851 35404 6885
rect 34368 6740 34416 6828
rect 34742 6785 34758 6819
rect 34792 6818 34808 6819
rect 34792 6786 34954 6818
rect 35194 6810 35260 6817
rect 35188 6805 35260 6810
rect 35188 6786 35210 6805
rect 34792 6785 35210 6786
rect 34742 6782 35210 6785
rect 34918 6771 35210 6782
rect 35244 6771 35260 6805
rect 34918 6750 35260 6771
rect 34614 6740 34648 6742
rect 34368 6723 34648 6740
rect 34368 6706 34614 6723
rect 33386 6605 33452 6608
rect 33598 6636 33639 6638
rect 33598 6602 33600 6636
rect 33634 6602 33639 6636
rect 33598 6600 33639 6602
rect 33306 6553 33372 6571
rect 33306 6519 33322 6553
rect 33356 6519 33372 6553
rect 33306 6485 33372 6519
rect 33306 6451 33322 6485
rect 33356 6451 33372 6485
rect 33306 6417 33372 6451
rect 33306 6383 33322 6417
rect 33356 6383 33372 6417
rect 33306 6375 33372 6383
rect 33406 6553 33448 6569
rect 33440 6519 33448 6553
rect 33406 6485 33448 6519
rect 33440 6451 33448 6485
rect 33406 6417 33448 6451
rect 33440 6383 33448 6417
rect 32877 6349 32916 6374
rect 32428 6297 32444 6331
rect 32478 6297 32494 6331
rect 32634 6310 32916 6349
rect 33406 6341 33448 6383
rect 33603 6550 33639 6600
rect 33673 6634 33728 6650
rect 33707 6600 33728 6634
rect 33673 6584 33728 6600
rect 33773 6648 33841 6665
rect 33773 6647 33793 6648
rect 33773 6613 33791 6647
rect 33827 6614 33841 6648
rect 33825 6613 33841 6614
rect 33773 6591 33841 6613
rect 33694 6555 33728 6584
rect 33998 6563 34044 6683
rect 34098 6679 34144 6695
rect 34316 6658 34332 6659
rect 34078 6611 34094 6645
rect 34128 6638 34144 6645
rect 34196 6638 34332 6658
rect 34128 6625 34332 6638
rect 34366 6625 34382 6659
rect 34128 6624 34382 6625
rect 34128 6611 34236 6624
rect 34316 6622 34382 6624
rect 34614 6655 34648 6657
rect 34078 6597 34236 6611
rect 34092 6596 34236 6597
rect 34614 6619 34648 6621
rect 34288 6563 34322 6582
rect 33603 6500 33657 6550
rect 33694 6521 33829 6555
rect 33603 6466 33621 6500
rect 33655 6466 33657 6500
rect 33793 6487 33829 6521
rect 33603 6419 33657 6466
rect 33603 6385 33621 6419
rect 33655 6385 33657 6419
rect 33603 6369 33657 6385
rect 33691 6453 33707 6487
rect 33741 6453 33757 6487
rect 33691 6419 33757 6453
rect 33691 6385 33707 6419
rect 33741 6385 33757 6419
rect 32802 6308 32916 6310
rect 33074 6297 33090 6331
rect 33124 6297 33140 6331
rect 33240 6307 33269 6341
rect 33303 6307 33361 6341
rect 33395 6307 33453 6341
rect 33487 6307 33516 6341
rect 33691 6335 33757 6385
rect 33827 6453 33829 6487
rect 33793 6419 33829 6453
rect 33827 6385 33829 6419
rect 33793 6369 33829 6385
rect 33998 6545 34064 6563
rect 33998 6511 34014 6545
rect 34048 6511 34064 6545
rect 33998 6477 34064 6511
rect 33998 6443 34014 6477
rect 34048 6443 34064 6477
rect 33998 6409 34064 6443
rect 33998 6375 34014 6409
rect 34048 6375 34064 6409
rect 33998 6367 34064 6375
rect 34098 6545 34140 6561
rect 34132 6511 34140 6545
rect 34098 6477 34140 6511
rect 34132 6443 34140 6477
rect 34098 6409 34140 6443
rect 34288 6495 34322 6497
rect 34288 6459 34322 6461
rect 34132 6375 34140 6409
rect 33407 6300 33441 6307
rect 33586 6301 33615 6335
rect 33649 6301 33707 6335
rect 33741 6301 33799 6335
rect 33833 6301 33862 6335
rect 34098 6333 34140 6375
rect 34248 6393 34288 6414
rect 34376 6563 34410 6582
rect 34614 6534 34648 6553
rect 34710 6723 34744 6742
rect 34710 6655 34744 6657
rect 34710 6619 34744 6621
rect 34710 6534 34744 6553
rect 34806 6723 34840 6742
rect 35194 6737 35260 6750
rect 35194 6703 35210 6737
rect 35244 6703 35260 6737
rect 35194 6691 35260 6703
rect 35294 6805 35340 6851
rect 35474 6845 35503 6879
rect 35537 6845 35595 6879
rect 35629 6845 35687 6879
rect 35721 6845 35750 6879
rect 35328 6771 35340 6805
rect 35294 6737 35340 6771
rect 35328 6703 35340 6737
rect 34806 6655 34840 6657
rect 34962 6625 34978 6659
rect 35012 6625 35028 6659
rect 34806 6619 34840 6621
rect 34806 6534 34840 6553
rect 34934 6563 34968 6582
rect 34376 6495 34410 6497
rect 34934 6495 34968 6497
rect 34376 6459 34410 6461
rect 34646 6457 34662 6491
rect 34696 6457 34712 6491
rect 34934 6459 34968 6461
rect 34322 6393 34324 6414
rect 34248 6374 34324 6393
rect 34410 6393 34934 6418
rect 35022 6563 35056 6582
rect 35022 6495 35056 6497
rect 35022 6459 35056 6461
rect 34968 6393 34970 6418
rect 34376 6385 34970 6393
rect 34376 6374 34612 6385
rect 33932 6299 33961 6333
rect 33995 6299 34053 6333
rect 34087 6299 34145 6333
rect 34179 6299 34208 6333
rect 32494 6212 32540 6218
rect 32494 6210 32982 6212
rect 32494 6176 32502 6210
rect 32536 6193 32982 6210
rect 32536 6188 32932 6193
rect 32536 6178 32811 6188
rect 32536 6176 32540 6178
rect 32494 6174 32540 6176
rect 32712 6154 32811 6178
rect 32845 6159 32932 6188
rect 32966 6168 32982 6193
rect 32966 6159 33107 6168
rect 32845 6154 33107 6159
rect 32712 6134 33107 6154
rect 32836 6050 32852 6084
rect 32886 6050 33022 6084
rect 32360 6000 32742 6016
rect 32360 5976 32708 6000
rect 32708 5930 32742 5964
rect 32708 5878 32742 5894
rect 32804 6000 32838 6016
rect 32804 5930 32838 5964
rect 32804 5878 32838 5894
rect 32900 6000 32934 6016
rect 32900 5930 32934 5964
rect 32900 5878 32934 5894
rect 31174 5797 31203 5831
rect 31237 5797 31295 5831
rect 31329 5797 31387 5831
rect 31421 5797 31450 5831
rect 32248 5797 32277 5831
rect 32311 5797 32369 5831
rect 32403 5797 32461 5831
rect 32495 5797 32524 5831
rect 32740 5810 32756 5844
rect 32790 5810 32806 5844
rect 31193 5753 31247 5797
rect 31193 5719 31213 5753
rect 31193 5685 31247 5719
rect 31193 5651 31213 5685
rect 31193 5635 31247 5651
rect 31281 5753 31347 5763
rect 31281 5719 31297 5753
rect 31331 5719 31347 5753
rect 31281 5710 31347 5719
rect 31281 5685 31299 5710
rect 31281 5651 31297 5685
rect 31333 5676 31347 5710
rect 31331 5651 31347 5676
rect 31281 5635 31347 5651
rect 31381 5753 31429 5797
rect 31415 5719 31429 5753
rect 31381 5685 31429 5719
rect 31415 5651 31429 5685
rect 31381 5635 31429 5651
rect 32267 5753 32321 5797
rect 32267 5719 32287 5753
rect 32267 5685 32321 5719
rect 32267 5651 32287 5685
rect 32267 5635 32321 5651
rect 32355 5753 32421 5763
rect 32355 5719 32371 5753
rect 32405 5719 32421 5753
rect 32355 5715 32421 5719
rect 32355 5681 32369 5715
rect 32403 5685 32421 5715
rect 32355 5651 32371 5681
rect 32405 5651 32421 5685
rect 32355 5635 32421 5651
rect 32455 5753 32503 5797
rect 32489 5719 32503 5753
rect 32852 5729 32868 5763
rect 32902 5729 32918 5763
rect 32455 5685 32503 5719
rect 32489 5651 32503 5685
rect 32455 5635 32503 5651
rect 32724 5667 32758 5686
rect 31191 5594 31211 5599
rect 31191 5560 31208 5594
rect 31245 5565 31261 5599
rect 31242 5560 31261 5565
rect 31191 5549 31261 5560
rect 31295 5515 31329 5635
rect 31363 5565 31379 5599
rect 31413 5590 31433 5599
rect 31363 5556 31381 5565
rect 31415 5556 31433 5590
rect 31363 5549 31433 5556
rect 32265 5592 32285 5599
rect 32265 5558 32283 5592
rect 32319 5565 32335 5599
rect 32317 5558 32335 5565
rect 32265 5549 32335 5558
rect 32369 5515 32403 5635
rect 32724 5599 32758 5601
rect 32437 5565 32453 5599
rect 32487 5592 32507 5599
rect 32437 5558 32457 5565
rect 32491 5558 32507 5592
rect 32437 5549 32507 5558
rect 32724 5563 32758 5565
rect 30868 5435 31134 5436
rect 30868 5401 30884 5435
rect 30918 5401 31134 5435
rect 30868 5400 31134 5401
rect 31193 5499 31259 5515
rect 31193 5465 31225 5499
rect 31295 5499 31431 5515
rect 31295 5481 31381 5499
rect 31193 5431 31259 5465
rect 30551 5363 30617 5397
rect 30551 5329 30567 5363
rect 30601 5329 30617 5363
rect 31193 5397 31225 5431
rect 31193 5363 31259 5397
rect 30551 5324 30617 5329
rect 30744 5329 31026 5362
rect 30744 5295 30834 5329
rect 30868 5327 31026 5329
rect 30868 5295 30953 5327
rect 30744 5293 30953 5295
rect 30987 5293 31026 5327
rect 30744 5287 31026 5293
rect 31193 5329 31225 5363
rect 31193 5287 31259 5329
rect 31365 5465 31381 5481
rect 31415 5465 31431 5499
rect 31365 5431 31431 5465
rect 31365 5397 31381 5431
rect 31415 5397 31431 5431
rect 31365 5363 31431 5397
rect 31365 5329 31381 5363
rect 31415 5329 31431 5363
rect 31365 5324 31431 5329
rect 32267 5499 32333 5515
rect 32267 5465 32299 5499
rect 32369 5499 32505 5515
rect 32369 5481 32455 5499
rect 32267 5431 32333 5465
rect 32267 5397 32299 5431
rect 32267 5363 32333 5397
rect 32267 5329 32299 5363
rect 32267 5287 32333 5329
rect 32439 5465 32455 5481
rect 32489 5465 32505 5499
rect 32724 5478 32758 5497
rect 32820 5667 32854 5686
rect 32820 5599 32854 5601
rect 32820 5563 32854 5565
rect 32820 5478 32854 5497
rect 32916 5667 32950 5686
rect 32916 5599 32950 5601
rect 32916 5563 32950 5565
rect 32916 5478 32950 5497
rect 32439 5431 32505 5465
rect 32439 5397 32455 5431
rect 32489 5397 32505 5431
rect 32756 5436 32822 5438
rect 32988 5436 33022 6050
rect 33073 5831 33107 6134
rect 33304 5831 33338 6042
rect 34248 6016 34282 6374
rect 34522 6351 34612 6374
rect 34646 6383 34970 6385
rect 34646 6351 34731 6383
rect 34522 6349 34731 6351
rect 34765 6374 34970 6383
rect 35022 6374 35056 6393
rect 35194 6571 35240 6691
rect 35294 6687 35340 6703
rect 35491 6773 35543 6811
rect 35491 6739 35509 6773
rect 35579 6803 35645 6845
rect 35820 6843 35849 6877
rect 35883 6843 35941 6877
rect 35975 6843 36033 6877
rect 36067 6843 36096 6877
rect 36256 6862 36304 6874
rect 36518 6866 36534 6900
rect 36568 6866 36584 6900
rect 36884 6890 36934 6960
rect 38374 6934 38408 6950
rect 38470 7056 38504 7072
rect 38566 7058 38600 7072
rect 38684 7058 38904 7080
rect 38564 7056 38904 7058
rect 38564 7022 38566 7056
rect 38600 7044 38904 7056
rect 38600 7022 38720 7044
rect 38470 6986 38504 7020
rect 38565 7020 38566 7022
rect 38565 6986 38600 7020
rect 38868 6996 38904 7044
rect 38565 6985 38566 6986
rect 38470 6934 38504 6950
rect 38566 6934 38600 6950
rect 38772 6960 38904 6996
rect 40262 7056 40296 7072
rect 40262 6986 40296 7020
rect 36884 6876 36894 6890
rect 35579 6769 35595 6803
rect 35629 6769 35645 6803
rect 35681 6790 35715 6811
rect 35491 6710 35543 6739
rect 35681 6735 35715 6756
rect 35274 6619 35290 6653
rect 35324 6642 35340 6653
rect 35274 6608 35292 6619
rect 35326 6608 35340 6642
rect 35491 6638 35527 6710
rect 35582 6701 35715 6735
rect 35886 6797 35952 6809
rect 35886 6763 35902 6797
rect 35936 6763 35952 6797
rect 35886 6746 35952 6763
rect 35582 6650 35616 6701
rect 35886 6695 35902 6746
rect 35936 6695 35952 6746
rect 35886 6683 35952 6695
rect 35986 6797 36032 6843
rect 36020 6763 36032 6797
rect 35986 6729 36032 6763
rect 36020 6695 36032 6729
rect 36256 6828 36262 6862
rect 36296 6828 36304 6862
rect 36888 6856 36894 6876
rect 36928 6856 36934 6890
rect 36888 6846 36934 6856
rect 37016 6851 37045 6885
rect 37079 6851 37137 6885
rect 37171 6851 37229 6885
rect 37263 6851 37292 6885
rect 36256 6740 36304 6828
rect 36630 6785 36646 6819
rect 36680 6818 36696 6819
rect 36680 6786 36842 6818
rect 37082 6810 37148 6817
rect 37076 6805 37148 6810
rect 37076 6786 37098 6805
rect 36680 6785 37098 6786
rect 36630 6782 37098 6785
rect 36806 6771 37098 6782
rect 37132 6771 37148 6805
rect 36806 6750 37148 6771
rect 36502 6740 36536 6742
rect 36256 6723 36536 6740
rect 36256 6706 36502 6723
rect 35274 6605 35340 6608
rect 35486 6636 35527 6638
rect 35486 6602 35488 6636
rect 35522 6602 35527 6636
rect 35486 6600 35527 6602
rect 35194 6553 35260 6571
rect 35194 6519 35210 6553
rect 35244 6519 35260 6553
rect 35194 6485 35260 6519
rect 35194 6451 35210 6485
rect 35244 6451 35260 6485
rect 35194 6417 35260 6451
rect 35194 6383 35210 6417
rect 35244 6383 35260 6417
rect 35194 6375 35260 6383
rect 35294 6553 35336 6569
rect 35328 6519 35336 6553
rect 35294 6485 35336 6519
rect 35328 6451 35336 6485
rect 35294 6417 35336 6451
rect 35328 6383 35336 6417
rect 34765 6349 34804 6374
rect 34316 6297 34332 6331
rect 34366 6297 34382 6331
rect 34522 6310 34804 6349
rect 35294 6341 35336 6383
rect 35491 6550 35527 6600
rect 35561 6634 35616 6650
rect 35595 6600 35616 6634
rect 35561 6584 35616 6600
rect 35661 6648 35729 6665
rect 35661 6647 35681 6648
rect 35661 6613 35679 6647
rect 35715 6614 35729 6648
rect 35713 6613 35729 6614
rect 35661 6591 35729 6613
rect 35582 6555 35616 6584
rect 35886 6563 35932 6683
rect 35986 6679 36032 6695
rect 36204 6658 36220 6659
rect 35966 6611 35982 6645
rect 36016 6638 36032 6645
rect 36084 6638 36220 6658
rect 36016 6625 36220 6638
rect 36254 6625 36270 6659
rect 36016 6624 36270 6625
rect 36016 6611 36124 6624
rect 36204 6622 36270 6624
rect 36502 6655 36536 6657
rect 35966 6597 36124 6611
rect 35980 6596 36124 6597
rect 36502 6619 36536 6621
rect 36176 6563 36210 6582
rect 35491 6500 35545 6550
rect 35582 6521 35717 6555
rect 35491 6466 35509 6500
rect 35543 6466 35545 6500
rect 35681 6487 35717 6521
rect 35491 6419 35545 6466
rect 35491 6385 35509 6419
rect 35543 6385 35545 6419
rect 35491 6369 35545 6385
rect 35579 6453 35595 6487
rect 35629 6453 35645 6487
rect 35579 6419 35645 6453
rect 35579 6385 35595 6419
rect 35629 6385 35645 6419
rect 34690 6308 34804 6310
rect 34962 6297 34978 6331
rect 35012 6297 35028 6331
rect 35128 6307 35157 6341
rect 35191 6307 35249 6341
rect 35283 6307 35341 6341
rect 35375 6307 35404 6341
rect 35579 6335 35645 6385
rect 35715 6453 35717 6487
rect 35681 6419 35717 6453
rect 35715 6385 35717 6419
rect 35681 6369 35717 6385
rect 35886 6545 35952 6563
rect 35886 6511 35902 6545
rect 35936 6511 35952 6545
rect 35886 6477 35952 6511
rect 35886 6443 35902 6477
rect 35936 6443 35952 6477
rect 35886 6409 35952 6443
rect 35886 6375 35902 6409
rect 35936 6375 35952 6409
rect 35886 6367 35952 6375
rect 35986 6545 36028 6561
rect 36020 6511 36028 6545
rect 35986 6477 36028 6511
rect 36020 6443 36028 6477
rect 35986 6409 36028 6443
rect 36176 6495 36210 6497
rect 36176 6459 36210 6461
rect 36020 6375 36028 6409
rect 35295 6300 35329 6307
rect 35474 6301 35503 6335
rect 35537 6301 35595 6335
rect 35629 6301 35687 6335
rect 35721 6301 35750 6335
rect 35986 6333 36028 6375
rect 36136 6393 36176 6414
rect 36264 6563 36298 6582
rect 36502 6534 36536 6553
rect 36598 6723 36632 6742
rect 36598 6655 36632 6657
rect 36598 6619 36632 6621
rect 36598 6534 36632 6553
rect 36694 6723 36728 6742
rect 37082 6737 37148 6750
rect 37082 6703 37098 6737
rect 37132 6703 37148 6737
rect 37082 6691 37148 6703
rect 37182 6805 37228 6851
rect 37362 6845 37391 6879
rect 37425 6845 37483 6879
rect 37517 6845 37575 6879
rect 37609 6845 37638 6879
rect 37216 6771 37228 6805
rect 37182 6737 37228 6771
rect 37216 6703 37228 6737
rect 36694 6655 36728 6657
rect 36850 6625 36866 6659
rect 36900 6625 36916 6659
rect 36694 6619 36728 6621
rect 36694 6534 36728 6553
rect 36822 6563 36856 6582
rect 36264 6495 36298 6497
rect 36822 6495 36856 6497
rect 36264 6459 36298 6461
rect 36534 6457 36550 6491
rect 36584 6457 36600 6491
rect 36822 6459 36856 6461
rect 36210 6393 36212 6414
rect 36136 6374 36212 6393
rect 36298 6393 36822 6418
rect 36910 6563 36944 6582
rect 36910 6495 36944 6497
rect 36910 6459 36944 6461
rect 36856 6393 36858 6418
rect 36264 6385 36858 6393
rect 36264 6374 36500 6385
rect 35820 6299 35849 6333
rect 35883 6299 35941 6333
rect 35975 6299 36033 6333
rect 36067 6299 36096 6333
rect 34382 6212 34428 6218
rect 34382 6210 34870 6212
rect 34382 6176 34390 6210
rect 34424 6193 34870 6210
rect 34424 6188 34820 6193
rect 34424 6178 34699 6188
rect 34424 6176 34428 6178
rect 34382 6174 34428 6176
rect 34600 6154 34699 6178
rect 34733 6159 34820 6188
rect 34854 6168 34870 6193
rect 34854 6159 34995 6168
rect 34733 6154 34995 6159
rect 34600 6134 34995 6154
rect 34724 6050 34740 6084
rect 34774 6050 34910 6084
rect 34248 6000 34630 6016
rect 34248 5976 34596 6000
rect 34596 5930 34630 5964
rect 34596 5878 34630 5894
rect 34692 6000 34726 6016
rect 34692 5930 34726 5964
rect 34692 5878 34726 5894
rect 34788 6000 34822 6016
rect 34788 5930 34822 5964
rect 34788 5878 34822 5894
rect 33062 5797 33091 5831
rect 33125 5797 33183 5831
rect 33217 5797 33275 5831
rect 33309 5797 33338 5831
rect 34136 5797 34165 5831
rect 34199 5797 34257 5831
rect 34291 5797 34349 5831
rect 34383 5797 34412 5831
rect 34628 5810 34644 5844
rect 34678 5810 34694 5844
rect 33081 5753 33135 5797
rect 33081 5719 33101 5753
rect 33081 5685 33135 5719
rect 33081 5651 33101 5685
rect 33081 5635 33135 5651
rect 33169 5753 33235 5763
rect 33169 5719 33185 5753
rect 33219 5719 33235 5753
rect 33169 5710 33235 5719
rect 33169 5685 33187 5710
rect 33169 5651 33185 5685
rect 33221 5676 33235 5710
rect 33219 5651 33235 5676
rect 33169 5635 33235 5651
rect 33269 5753 33317 5797
rect 33303 5719 33317 5753
rect 33269 5685 33317 5719
rect 33303 5651 33317 5685
rect 33269 5635 33317 5651
rect 34155 5753 34209 5797
rect 34155 5719 34175 5753
rect 34155 5685 34209 5719
rect 34155 5651 34175 5685
rect 34155 5635 34209 5651
rect 34243 5753 34309 5763
rect 34243 5719 34259 5753
rect 34293 5719 34309 5753
rect 34243 5715 34309 5719
rect 34243 5681 34257 5715
rect 34291 5685 34309 5715
rect 34243 5651 34259 5681
rect 34293 5651 34309 5685
rect 34243 5635 34309 5651
rect 34343 5753 34391 5797
rect 34377 5719 34391 5753
rect 34740 5729 34756 5763
rect 34790 5729 34806 5763
rect 34343 5685 34391 5719
rect 34377 5651 34391 5685
rect 34343 5635 34391 5651
rect 34612 5667 34646 5686
rect 33079 5594 33099 5599
rect 33079 5560 33096 5594
rect 33133 5565 33149 5599
rect 33130 5560 33149 5565
rect 33079 5549 33149 5560
rect 33183 5515 33217 5635
rect 33251 5565 33267 5599
rect 33301 5590 33321 5599
rect 33251 5556 33269 5565
rect 33303 5556 33321 5590
rect 33251 5549 33321 5556
rect 34153 5592 34173 5599
rect 34153 5558 34171 5592
rect 34207 5565 34223 5599
rect 34205 5558 34223 5565
rect 34153 5549 34223 5558
rect 34257 5515 34291 5635
rect 34612 5599 34646 5601
rect 34325 5565 34341 5599
rect 34375 5592 34395 5599
rect 34325 5558 34345 5565
rect 34379 5558 34395 5592
rect 34325 5549 34395 5558
rect 34612 5563 34646 5565
rect 32756 5435 33022 5436
rect 32756 5401 32772 5435
rect 32806 5401 33022 5435
rect 32756 5400 33022 5401
rect 33081 5499 33147 5515
rect 33081 5465 33113 5499
rect 33183 5499 33319 5515
rect 33183 5481 33269 5499
rect 33081 5431 33147 5465
rect 32439 5363 32505 5397
rect 32439 5329 32455 5363
rect 32489 5329 32505 5363
rect 33081 5397 33113 5431
rect 33081 5363 33147 5397
rect 32439 5324 32505 5329
rect 32632 5329 32914 5362
rect 32632 5295 32722 5329
rect 32756 5327 32914 5329
rect 32756 5295 32841 5327
rect 32632 5293 32841 5295
rect 32875 5293 32914 5327
rect 32632 5287 32914 5293
rect 33081 5329 33113 5363
rect 33081 5287 33147 5329
rect 33253 5465 33269 5481
rect 33303 5465 33319 5499
rect 33253 5431 33319 5465
rect 33253 5397 33269 5431
rect 33303 5397 33319 5431
rect 33253 5363 33319 5397
rect 33253 5329 33269 5363
rect 33303 5329 33319 5363
rect 33253 5324 33319 5329
rect 34155 5499 34221 5515
rect 34155 5465 34187 5499
rect 34257 5499 34393 5515
rect 34257 5481 34343 5499
rect 34155 5431 34221 5465
rect 34155 5397 34187 5431
rect 34155 5363 34221 5397
rect 34155 5329 34187 5363
rect 34155 5287 34221 5329
rect 34327 5465 34343 5481
rect 34377 5465 34393 5499
rect 34612 5478 34646 5497
rect 34708 5667 34742 5686
rect 34708 5599 34742 5601
rect 34708 5563 34742 5565
rect 34708 5478 34742 5497
rect 34804 5667 34838 5686
rect 34804 5599 34838 5601
rect 34804 5563 34838 5565
rect 34804 5478 34838 5497
rect 34327 5431 34393 5465
rect 34327 5397 34343 5431
rect 34377 5397 34393 5431
rect 34644 5436 34710 5438
rect 34876 5436 34910 6050
rect 34961 5831 34995 6134
rect 35192 5831 35226 6042
rect 36136 6016 36170 6374
rect 36410 6351 36500 6374
rect 36534 6383 36858 6385
rect 36534 6351 36619 6383
rect 36410 6349 36619 6351
rect 36653 6374 36858 6383
rect 36910 6374 36944 6393
rect 37082 6571 37128 6691
rect 37182 6687 37228 6703
rect 37379 6773 37431 6811
rect 37379 6739 37397 6773
rect 37467 6803 37533 6845
rect 37708 6843 37737 6877
rect 37771 6843 37829 6877
rect 37863 6843 37921 6877
rect 37955 6843 37984 6877
rect 38144 6862 38192 6874
rect 38406 6866 38422 6900
rect 38456 6866 38472 6900
rect 38772 6890 38822 6960
rect 40262 6934 40296 6950
rect 40358 7056 40392 7072
rect 40454 7058 40488 7072
rect 40572 7058 40792 7080
rect 40452 7056 40792 7058
rect 40452 7022 40454 7056
rect 40488 7044 40792 7056
rect 40488 7022 40608 7044
rect 40358 6986 40392 7020
rect 40453 7020 40454 7022
rect 40453 6986 40488 7020
rect 40756 6996 40792 7044
rect 40453 6985 40454 6986
rect 40358 6934 40392 6950
rect 40454 6934 40488 6950
rect 40660 6960 40792 6996
rect 42150 7056 42184 7072
rect 42150 6986 42184 7020
rect 38772 6876 38782 6890
rect 37467 6769 37483 6803
rect 37517 6769 37533 6803
rect 37569 6790 37603 6811
rect 37379 6710 37431 6739
rect 37569 6735 37603 6756
rect 37162 6619 37178 6653
rect 37212 6642 37228 6653
rect 37162 6608 37180 6619
rect 37214 6608 37228 6642
rect 37379 6638 37415 6710
rect 37470 6701 37603 6735
rect 37774 6797 37840 6809
rect 37774 6763 37790 6797
rect 37824 6763 37840 6797
rect 37774 6746 37840 6763
rect 37470 6650 37504 6701
rect 37774 6695 37790 6746
rect 37824 6695 37840 6746
rect 37774 6683 37840 6695
rect 37874 6797 37920 6843
rect 37908 6763 37920 6797
rect 37874 6729 37920 6763
rect 37908 6695 37920 6729
rect 38144 6828 38150 6862
rect 38184 6828 38192 6862
rect 38776 6856 38782 6876
rect 38816 6856 38822 6890
rect 38776 6846 38822 6856
rect 38904 6851 38933 6885
rect 38967 6851 39025 6885
rect 39059 6851 39117 6885
rect 39151 6851 39180 6885
rect 38144 6740 38192 6828
rect 38518 6785 38534 6819
rect 38568 6818 38584 6819
rect 38568 6786 38730 6818
rect 38970 6810 39036 6817
rect 38964 6805 39036 6810
rect 38964 6786 38986 6805
rect 38568 6785 38986 6786
rect 38518 6782 38986 6785
rect 38694 6771 38986 6782
rect 39020 6771 39036 6805
rect 38694 6750 39036 6771
rect 38390 6740 38424 6742
rect 38144 6723 38424 6740
rect 38144 6706 38390 6723
rect 37162 6605 37228 6608
rect 37374 6636 37415 6638
rect 37374 6602 37376 6636
rect 37410 6602 37415 6636
rect 37374 6600 37415 6602
rect 37082 6553 37148 6571
rect 37082 6519 37098 6553
rect 37132 6519 37148 6553
rect 37082 6485 37148 6519
rect 37082 6451 37098 6485
rect 37132 6451 37148 6485
rect 37082 6417 37148 6451
rect 37082 6383 37098 6417
rect 37132 6383 37148 6417
rect 37082 6375 37148 6383
rect 37182 6553 37224 6569
rect 37216 6519 37224 6553
rect 37182 6485 37224 6519
rect 37216 6451 37224 6485
rect 37182 6417 37224 6451
rect 37216 6383 37224 6417
rect 36653 6349 36692 6374
rect 36204 6297 36220 6331
rect 36254 6297 36270 6331
rect 36410 6310 36692 6349
rect 37182 6341 37224 6383
rect 37379 6550 37415 6600
rect 37449 6634 37504 6650
rect 37483 6600 37504 6634
rect 37449 6584 37504 6600
rect 37549 6648 37617 6665
rect 37549 6647 37569 6648
rect 37549 6613 37567 6647
rect 37603 6614 37617 6648
rect 37601 6613 37617 6614
rect 37549 6591 37617 6613
rect 37470 6555 37504 6584
rect 37774 6563 37820 6683
rect 37874 6679 37920 6695
rect 38092 6658 38108 6659
rect 37854 6611 37870 6645
rect 37904 6638 37920 6645
rect 37972 6638 38108 6658
rect 37904 6625 38108 6638
rect 38142 6625 38158 6659
rect 37904 6624 38158 6625
rect 37904 6611 38012 6624
rect 38092 6622 38158 6624
rect 38390 6655 38424 6657
rect 37854 6597 38012 6611
rect 37868 6596 38012 6597
rect 38390 6619 38424 6621
rect 38064 6563 38098 6582
rect 37379 6500 37433 6550
rect 37470 6521 37605 6555
rect 37379 6466 37397 6500
rect 37431 6466 37433 6500
rect 37569 6487 37605 6521
rect 37379 6419 37433 6466
rect 37379 6385 37397 6419
rect 37431 6385 37433 6419
rect 37379 6369 37433 6385
rect 37467 6453 37483 6487
rect 37517 6453 37533 6487
rect 37467 6419 37533 6453
rect 37467 6385 37483 6419
rect 37517 6385 37533 6419
rect 36578 6308 36692 6310
rect 36850 6297 36866 6331
rect 36900 6297 36916 6331
rect 37016 6307 37045 6341
rect 37079 6307 37137 6341
rect 37171 6307 37229 6341
rect 37263 6307 37292 6341
rect 37467 6335 37533 6385
rect 37603 6453 37605 6487
rect 37569 6419 37605 6453
rect 37603 6385 37605 6419
rect 37569 6369 37605 6385
rect 37774 6545 37840 6563
rect 37774 6511 37790 6545
rect 37824 6511 37840 6545
rect 37774 6477 37840 6511
rect 37774 6443 37790 6477
rect 37824 6443 37840 6477
rect 37774 6409 37840 6443
rect 37774 6375 37790 6409
rect 37824 6375 37840 6409
rect 37774 6367 37840 6375
rect 37874 6545 37916 6561
rect 37908 6511 37916 6545
rect 37874 6477 37916 6511
rect 37908 6443 37916 6477
rect 37874 6409 37916 6443
rect 38064 6495 38098 6497
rect 38064 6459 38098 6461
rect 37908 6375 37916 6409
rect 37183 6300 37217 6307
rect 37362 6301 37391 6335
rect 37425 6301 37483 6335
rect 37517 6301 37575 6335
rect 37609 6301 37638 6335
rect 37874 6333 37916 6375
rect 38024 6393 38064 6414
rect 38152 6563 38186 6582
rect 38390 6534 38424 6553
rect 38486 6723 38520 6742
rect 38486 6655 38520 6657
rect 38486 6619 38520 6621
rect 38486 6534 38520 6553
rect 38582 6723 38616 6742
rect 38970 6737 39036 6750
rect 38970 6703 38986 6737
rect 39020 6703 39036 6737
rect 38970 6691 39036 6703
rect 39070 6805 39116 6851
rect 39250 6845 39279 6879
rect 39313 6845 39371 6879
rect 39405 6845 39463 6879
rect 39497 6845 39526 6879
rect 39104 6771 39116 6805
rect 39070 6737 39116 6771
rect 39104 6703 39116 6737
rect 38582 6655 38616 6657
rect 38738 6625 38754 6659
rect 38788 6625 38804 6659
rect 38582 6619 38616 6621
rect 38582 6534 38616 6553
rect 38710 6563 38744 6582
rect 38152 6495 38186 6497
rect 38710 6495 38744 6497
rect 38152 6459 38186 6461
rect 38422 6457 38438 6491
rect 38472 6457 38488 6491
rect 38710 6459 38744 6461
rect 38098 6393 38100 6414
rect 38024 6374 38100 6393
rect 38186 6393 38710 6418
rect 38798 6563 38832 6582
rect 38798 6495 38832 6497
rect 38798 6459 38832 6461
rect 38744 6393 38746 6418
rect 38152 6385 38746 6393
rect 38152 6374 38388 6385
rect 37708 6299 37737 6333
rect 37771 6299 37829 6333
rect 37863 6299 37921 6333
rect 37955 6299 37984 6333
rect 36270 6212 36316 6218
rect 36270 6210 36758 6212
rect 36270 6176 36278 6210
rect 36312 6193 36758 6210
rect 36312 6188 36708 6193
rect 36312 6178 36587 6188
rect 36312 6176 36316 6178
rect 36270 6174 36316 6176
rect 36488 6154 36587 6178
rect 36621 6159 36708 6188
rect 36742 6168 36758 6193
rect 36742 6159 36883 6168
rect 36621 6154 36883 6159
rect 36488 6134 36883 6154
rect 36612 6050 36628 6084
rect 36662 6050 36798 6084
rect 36136 6000 36518 6016
rect 36136 5976 36484 6000
rect 36484 5930 36518 5964
rect 36484 5878 36518 5894
rect 36580 6000 36614 6016
rect 36580 5930 36614 5964
rect 36580 5878 36614 5894
rect 36676 6000 36710 6016
rect 36676 5930 36710 5964
rect 36676 5878 36710 5894
rect 34950 5797 34979 5831
rect 35013 5797 35071 5831
rect 35105 5797 35163 5831
rect 35197 5797 35226 5831
rect 36024 5797 36053 5831
rect 36087 5797 36145 5831
rect 36179 5797 36237 5831
rect 36271 5797 36300 5831
rect 36516 5810 36532 5844
rect 36566 5810 36582 5844
rect 34969 5753 35023 5797
rect 34969 5719 34989 5753
rect 34969 5685 35023 5719
rect 34969 5651 34989 5685
rect 34969 5635 35023 5651
rect 35057 5753 35123 5763
rect 35057 5719 35073 5753
rect 35107 5719 35123 5753
rect 35057 5710 35123 5719
rect 35057 5685 35075 5710
rect 35057 5651 35073 5685
rect 35109 5676 35123 5710
rect 35107 5651 35123 5676
rect 35057 5635 35123 5651
rect 35157 5753 35205 5797
rect 35191 5719 35205 5753
rect 35157 5685 35205 5719
rect 35191 5651 35205 5685
rect 35157 5635 35205 5651
rect 36043 5753 36097 5797
rect 36043 5719 36063 5753
rect 36043 5685 36097 5719
rect 36043 5651 36063 5685
rect 36043 5635 36097 5651
rect 36131 5753 36197 5763
rect 36131 5719 36147 5753
rect 36181 5719 36197 5753
rect 36131 5715 36197 5719
rect 36131 5681 36145 5715
rect 36179 5685 36197 5715
rect 36131 5651 36147 5681
rect 36181 5651 36197 5685
rect 36131 5635 36197 5651
rect 36231 5753 36279 5797
rect 36265 5719 36279 5753
rect 36628 5729 36644 5763
rect 36678 5729 36694 5763
rect 36231 5685 36279 5719
rect 36265 5651 36279 5685
rect 36231 5635 36279 5651
rect 36500 5667 36534 5686
rect 34967 5594 34987 5599
rect 34967 5560 34984 5594
rect 35021 5565 35037 5599
rect 35018 5560 35037 5565
rect 34967 5549 35037 5560
rect 35071 5515 35105 5635
rect 35139 5565 35155 5599
rect 35189 5590 35209 5599
rect 35139 5556 35157 5565
rect 35191 5556 35209 5590
rect 35139 5549 35209 5556
rect 36041 5592 36061 5599
rect 36041 5558 36059 5592
rect 36095 5565 36111 5599
rect 36093 5558 36111 5565
rect 36041 5549 36111 5558
rect 36145 5515 36179 5635
rect 36500 5599 36534 5601
rect 36213 5565 36229 5599
rect 36263 5592 36283 5599
rect 36213 5558 36233 5565
rect 36267 5558 36283 5592
rect 36213 5549 36283 5558
rect 36500 5563 36534 5565
rect 34644 5435 34910 5436
rect 34644 5401 34660 5435
rect 34694 5401 34910 5435
rect 34644 5400 34910 5401
rect 34969 5499 35035 5515
rect 34969 5465 35001 5499
rect 35071 5499 35207 5515
rect 35071 5481 35157 5499
rect 34969 5431 35035 5465
rect 34327 5363 34393 5397
rect 34327 5329 34343 5363
rect 34377 5329 34393 5363
rect 34969 5397 35001 5431
rect 34969 5363 35035 5397
rect 34327 5324 34393 5329
rect 34520 5329 34802 5362
rect 34520 5295 34610 5329
rect 34644 5327 34802 5329
rect 34644 5295 34729 5327
rect 34520 5293 34729 5295
rect 34763 5293 34802 5327
rect 34520 5287 34802 5293
rect 34969 5329 35001 5363
rect 34969 5287 35035 5329
rect 35141 5465 35157 5481
rect 35191 5465 35207 5499
rect 35141 5431 35207 5465
rect 35141 5397 35157 5431
rect 35191 5397 35207 5431
rect 35141 5363 35207 5397
rect 35141 5329 35157 5363
rect 35191 5329 35207 5363
rect 35141 5324 35207 5329
rect 36043 5499 36109 5515
rect 36043 5465 36075 5499
rect 36145 5499 36281 5515
rect 36145 5481 36231 5499
rect 36043 5431 36109 5465
rect 36043 5397 36075 5431
rect 36043 5363 36109 5397
rect 36043 5329 36075 5363
rect 36043 5287 36109 5329
rect 36215 5465 36231 5481
rect 36265 5465 36281 5499
rect 36500 5478 36534 5497
rect 36596 5667 36630 5686
rect 36596 5599 36630 5601
rect 36596 5563 36630 5565
rect 36596 5478 36630 5497
rect 36692 5667 36726 5686
rect 36692 5599 36726 5601
rect 36692 5563 36726 5565
rect 36692 5478 36726 5497
rect 36215 5431 36281 5465
rect 36215 5397 36231 5431
rect 36265 5397 36281 5431
rect 36532 5436 36598 5438
rect 36764 5436 36798 6050
rect 36849 5831 36883 6134
rect 37080 5831 37114 6042
rect 38024 6016 38058 6374
rect 38298 6351 38388 6374
rect 38422 6383 38746 6385
rect 38422 6351 38507 6383
rect 38298 6349 38507 6351
rect 38541 6374 38746 6383
rect 38798 6374 38832 6393
rect 38970 6571 39016 6691
rect 39070 6687 39116 6703
rect 39267 6773 39319 6811
rect 39267 6739 39285 6773
rect 39355 6803 39421 6845
rect 39596 6843 39625 6877
rect 39659 6843 39717 6877
rect 39751 6843 39809 6877
rect 39843 6843 39872 6877
rect 40032 6862 40080 6874
rect 40294 6866 40310 6900
rect 40344 6866 40360 6900
rect 40660 6890 40710 6960
rect 42150 6934 42184 6950
rect 42246 7056 42280 7072
rect 42342 7058 42376 7072
rect 42460 7058 42680 7080
rect 42340 7056 42680 7058
rect 42340 7022 42342 7056
rect 42376 7044 42680 7056
rect 42376 7022 42496 7044
rect 42246 6986 42280 7020
rect 42341 7020 42342 7022
rect 42341 6986 42376 7020
rect 42644 6996 42680 7044
rect 42341 6985 42342 6986
rect 42246 6934 42280 6950
rect 42342 6934 42376 6950
rect 42548 6960 42680 6996
rect 44038 7056 44072 7072
rect 44038 6986 44072 7020
rect 40660 6876 40670 6890
rect 39355 6769 39371 6803
rect 39405 6769 39421 6803
rect 39457 6790 39491 6811
rect 39267 6710 39319 6739
rect 39457 6735 39491 6756
rect 39050 6619 39066 6653
rect 39100 6642 39116 6653
rect 39050 6608 39068 6619
rect 39102 6608 39116 6642
rect 39267 6638 39303 6710
rect 39358 6701 39491 6735
rect 39662 6797 39728 6809
rect 39662 6763 39678 6797
rect 39712 6763 39728 6797
rect 39662 6746 39728 6763
rect 39358 6650 39392 6701
rect 39662 6695 39678 6746
rect 39712 6695 39728 6746
rect 39662 6683 39728 6695
rect 39762 6797 39808 6843
rect 39796 6763 39808 6797
rect 39762 6729 39808 6763
rect 39796 6695 39808 6729
rect 40032 6828 40038 6862
rect 40072 6828 40080 6862
rect 40664 6856 40670 6876
rect 40704 6856 40710 6890
rect 40664 6846 40710 6856
rect 40792 6851 40821 6885
rect 40855 6851 40913 6885
rect 40947 6851 41005 6885
rect 41039 6851 41068 6885
rect 40032 6740 40080 6828
rect 40406 6785 40422 6819
rect 40456 6818 40472 6819
rect 40456 6786 40618 6818
rect 40858 6810 40924 6817
rect 40852 6805 40924 6810
rect 40852 6786 40874 6805
rect 40456 6785 40874 6786
rect 40406 6782 40874 6785
rect 40582 6771 40874 6782
rect 40908 6771 40924 6805
rect 40582 6750 40924 6771
rect 40278 6740 40312 6742
rect 40032 6723 40312 6740
rect 40032 6706 40278 6723
rect 39050 6605 39116 6608
rect 39262 6636 39303 6638
rect 39262 6602 39264 6636
rect 39298 6602 39303 6636
rect 39262 6600 39303 6602
rect 38970 6553 39036 6571
rect 38970 6519 38986 6553
rect 39020 6519 39036 6553
rect 38970 6485 39036 6519
rect 38970 6451 38986 6485
rect 39020 6451 39036 6485
rect 38970 6417 39036 6451
rect 38970 6383 38986 6417
rect 39020 6383 39036 6417
rect 38970 6375 39036 6383
rect 39070 6553 39112 6569
rect 39104 6519 39112 6553
rect 39070 6485 39112 6519
rect 39104 6451 39112 6485
rect 39070 6417 39112 6451
rect 39104 6383 39112 6417
rect 38541 6349 38580 6374
rect 38092 6297 38108 6331
rect 38142 6297 38158 6331
rect 38298 6310 38580 6349
rect 39070 6341 39112 6383
rect 39267 6550 39303 6600
rect 39337 6634 39392 6650
rect 39371 6600 39392 6634
rect 39337 6584 39392 6600
rect 39437 6648 39505 6665
rect 39437 6647 39457 6648
rect 39437 6613 39455 6647
rect 39491 6614 39505 6648
rect 39489 6613 39505 6614
rect 39437 6591 39505 6613
rect 39358 6555 39392 6584
rect 39662 6563 39708 6683
rect 39762 6679 39808 6695
rect 39980 6658 39996 6659
rect 39742 6611 39758 6645
rect 39792 6638 39808 6645
rect 39860 6638 39996 6658
rect 39792 6625 39996 6638
rect 40030 6625 40046 6659
rect 39792 6624 40046 6625
rect 39792 6611 39900 6624
rect 39980 6622 40046 6624
rect 40278 6655 40312 6657
rect 39742 6597 39900 6611
rect 39756 6596 39900 6597
rect 40278 6619 40312 6621
rect 39952 6563 39986 6582
rect 39267 6500 39321 6550
rect 39358 6521 39493 6555
rect 39267 6466 39285 6500
rect 39319 6466 39321 6500
rect 39457 6487 39493 6521
rect 39267 6419 39321 6466
rect 39267 6385 39285 6419
rect 39319 6385 39321 6419
rect 39267 6369 39321 6385
rect 39355 6453 39371 6487
rect 39405 6453 39421 6487
rect 39355 6419 39421 6453
rect 39355 6385 39371 6419
rect 39405 6385 39421 6419
rect 38466 6308 38580 6310
rect 38738 6297 38754 6331
rect 38788 6297 38804 6331
rect 38904 6307 38933 6341
rect 38967 6307 39025 6341
rect 39059 6307 39117 6341
rect 39151 6307 39180 6341
rect 39355 6335 39421 6385
rect 39491 6453 39493 6487
rect 39457 6419 39493 6453
rect 39491 6385 39493 6419
rect 39457 6369 39493 6385
rect 39662 6545 39728 6563
rect 39662 6511 39678 6545
rect 39712 6511 39728 6545
rect 39662 6477 39728 6511
rect 39662 6443 39678 6477
rect 39712 6443 39728 6477
rect 39662 6409 39728 6443
rect 39662 6375 39678 6409
rect 39712 6375 39728 6409
rect 39662 6367 39728 6375
rect 39762 6545 39804 6561
rect 39796 6511 39804 6545
rect 39762 6477 39804 6511
rect 39796 6443 39804 6477
rect 39762 6409 39804 6443
rect 39952 6495 39986 6497
rect 39952 6459 39986 6461
rect 39796 6375 39804 6409
rect 39071 6300 39105 6307
rect 39250 6301 39279 6335
rect 39313 6301 39371 6335
rect 39405 6301 39463 6335
rect 39497 6301 39526 6335
rect 39762 6333 39804 6375
rect 39912 6393 39952 6414
rect 40040 6563 40074 6582
rect 40278 6534 40312 6553
rect 40374 6723 40408 6742
rect 40374 6655 40408 6657
rect 40374 6619 40408 6621
rect 40374 6534 40408 6553
rect 40470 6723 40504 6742
rect 40858 6737 40924 6750
rect 40858 6703 40874 6737
rect 40908 6703 40924 6737
rect 40858 6691 40924 6703
rect 40958 6805 41004 6851
rect 41138 6845 41167 6879
rect 41201 6845 41259 6879
rect 41293 6845 41351 6879
rect 41385 6845 41414 6879
rect 40992 6771 41004 6805
rect 40958 6737 41004 6771
rect 40992 6703 41004 6737
rect 40470 6655 40504 6657
rect 40626 6625 40642 6659
rect 40676 6625 40692 6659
rect 40470 6619 40504 6621
rect 40470 6534 40504 6553
rect 40598 6563 40632 6582
rect 40040 6495 40074 6497
rect 40598 6495 40632 6497
rect 40040 6459 40074 6461
rect 40310 6457 40326 6491
rect 40360 6457 40376 6491
rect 40598 6459 40632 6461
rect 39986 6393 39988 6414
rect 39912 6374 39988 6393
rect 40074 6393 40598 6418
rect 40686 6563 40720 6582
rect 40686 6495 40720 6497
rect 40686 6459 40720 6461
rect 40632 6393 40634 6418
rect 40040 6385 40634 6393
rect 40040 6374 40276 6385
rect 39596 6299 39625 6333
rect 39659 6299 39717 6333
rect 39751 6299 39809 6333
rect 39843 6299 39872 6333
rect 38158 6212 38204 6218
rect 38158 6210 38646 6212
rect 38158 6176 38166 6210
rect 38200 6193 38646 6210
rect 38200 6188 38596 6193
rect 38200 6178 38475 6188
rect 38200 6176 38204 6178
rect 38158 6174 38204 6176
rect 38376 6154 38475 6178
rect 38509 6159 38596 6188
rect 38630 6168 38646 6193
rect 38630 6159 38771 6168
rect 38509 6154 38771 6159
rect 38376 6134 38771 6154
rect 38500 6050 38516 6084
rect 38550 6050 38686 6084
rect 38024 6000 38406 6016
rect 38024 5976 38372 6000
rect 38372 5930 38406 5964
rect 38372 5878 38406 5894
rect 38468 6000 38502 6016
rect 38468 5930 38502 5964
rect 38468 5878 38502 5894
rect 38564 6000 38598 6016
rect 38564 5930 38598 5964
rect 38564 5878 38598 5894
rect 36838 5797 36867 5831
rect 36901 5797 36959 5831
rect 36993 5797 37051 5831
rect 37085 5797 37114 5831
rect 37912 5797 37941 5831
rect 37975 5797 38033 5831
rect 38067 5797 38125 5831
rect 38159 5797 38188 5831
rect 38404 5810 38420 5844
rect 38454 5810 38470 5844
rect 36857 5753 36911 5797
rect 36857 5719 36877 5753
rect 36857 5685 36911 5719
rect 36857 5651 36877 5685
rect 36857 5635 36911 5651
rect 36945 5753 37011 5763
rect 36945 5719 36961 5753
rect 36995 5719 37011 5753
rect 36945 5710 37011 5719
rect 36945 5685 36963 5710
rect 36945 5651 36961 5685
rect 36997 5676 37011 5710
rect 36995 5651 37011 5676
rect 36945 5635 37011 5651
rect 37045 5753 37093 5797
rect 37079 5719 37093 5753
rect 37045 5685 37093 5719
rect 37079 5651 37093 5685
rect 37045 5635 37093 5651
rect 37931 5753 37985 5797
rect 37931 5719 37951 5753
rect 37931 5685 37985 5719
rect 37931 5651 37951 5685
rect 37931 5635 37985 5651
rect 38019 5753 38085 5763
rect 38019 5719 38035 5753
rect 38069 5719 38085 5753
rect 38019 5715 38085 5719
rect 38019 5681 38033 5715
rect 38067 5685 38085 5715
rect 38019 5651 38035 5681
rect 38069 5651 38085 5685
rect 38019 5635 38085 5651
rect 38119 5753 38167 5797
rect 38153 5719 38167 5753
rect 38516 5729 38532 5763
rect 38566 5729 38582 5763
rect 38119 5685 38167 5719
rect 38153 5651 38167 5685
rect 38119 5635 38167 5651
rect 38388 5667 38422 5686
rect 36855 5594 36875 5599
rect 36855 5560 36872 5594
rect 36909 5565 36925 5599
rect 36906 5560 36925 5565
rect 36855 5549 36925 5560
rect 36959 5515 36993 5635
rect 37027 5565 37043 5599
rect 37077 5590 37097 5599
rect 37027 5556 37045 5565
rect 37079 5556 37097 5590
rect 37027 5549 37097 5556
rect 37929 5592 37949 5599
rect 37929 5558 37947 5592
rect 37983 5565 37999 5599
rect 37981 5558 37999 5565
rect 37929 5549 37999 5558
rect 38033 5515 38067 5635
rect 38388 5599 38422 5601
rect 38101 5565 38117 5599
rect 38151 5592 38171 5599
rect 38101 5558 38121 5565
rect 38155 5558 38171 5592
rect 38101 5549 38171 5558
rect 38388 5563 38422 5565
rect 36532 5435 36798 5436
rect 36532 5401 36548 5435
rect 36582 5401 36798 5435
rect 36532 5400 36798 5401
rect 36857 5499 36923 5515
rect 36857 5465 36889 5499
rect 36959 5499 37095 5515
rect 36959 5481 37045 5499
rect 36857 5431 36923 5465
rect 36215 5363 36281 5397
rect 36215 5329 36231 5363
rect 36265 5329 36281 5363
rect 36857 5397 36889 5431
rect 36857 5363 36923 5397
rect 36215 5324 36281 5329
rect 36408 5329 36690 5362
rect 36408 5295 36498 5329
rect 36532 5327 36690 5329
rect 36532 5295 36617 5327
rect 36408 5293 36617 5295
rect 36651 5293 36690 5327
rect 36408 5287 36690 5293
rect 36857 5329 36889 5363
rect 36857 5287 36923 5329
rect 37029 5465 37045 5481
rect 37079 5465 37095 5499
rect 37029 5431 37095 5465
rect 37029 5397 37045 5431
rect 37079 5397 37095 5431
rect 37029 5363 37095 5397
rect 37029 5329 37045 5363
rect 37079 5329 37095 5363
rect 37029 5324 37095 5329
rect 37931 5499 37997 5515
rect 37931 5465 37963 5499
rect 38033 5499 38169 5515
rect 38033 5481 38119 5499
rect 37931 5431 37997 5465
rect 37931 5397 37963 5431
rect 37931 5363 37997 5397
rect 37931 5329 37963 5363
rect 37931 5287 37997 5329
rect 38103 5465 38119 5481
rect 38153 5465 38169 5499
rect 38388 5478 38422 5497
rect 38484 5667 38518 5686
rect 38484 5599 38518 5601
rect 38484 5563 38518 5565
rect 38484 5478 38518 5497
rect 38580 5667 38614 5686
rect 38580 5599 38614 5601
rect 38580 5563 38614 5565
rect 38580 5478 38614 5497
rect 38103 5431 38169 5465
rect 38103 5397 38119 5431
rect 38153 5397 38169 5431
rect 38420 5436 38486 5438
rect 38652 5436 38686 6050
rect 38737 5831 38771 6134
rect 38968 5831 39002 6042
rect 39912 6016 39946 6374
rect 40186 6351 40276 6374
rect 40310 6383 40634 6385
rect 40310 6351 40395 6383
rect 40186 6349 40395 6351
rect 40429 6374 40634 6383
rect 40686 6374 40720 6393
rect 40858 6571 40904 6691
rect 40958 6687 41004 6703
rect 41155 6773 41207 6811
rect 41155 6739 41173 6773
rect 41243 6803 41309 6845
rect 41484 6843 41513 6877
rect 41547 6843 41605 6877
rect 41639 6843 41697 6877
rect 41731 6843 41760 6877
rect 41920 6862 41968 6874
rect 42182 6866 42198 6900
rect 42232 6866 42248 6900
rect 42548 6890 42598 6960
rect 44038 6934 44072 6950
rect 44134 7056 44168 7072
rect 44230 7058 44264 7072
rect 44348 7058 44568 7080
rect 44228 7056 44568 7058
rect 44228 7022 44230 7056
rect 44264 7044 44568 7056
rect 44264 7022 44384 7044
rect 44134 6986 44168 7020
rect 44229 7020 44230 7022
rect 44229 6986 44264 7020
rect 44532 6996 44568 7044
rect 44229 6985 44230 6986
rect 44134 6934 44168 6950
rect 44230 6934 44264 6950
rect 44436 6960 44568 6996
rect 45920 7056 45954 7072
rect 45920 6986 45954 7020
rect 42548 6876 42558 6890
rect 41243 6769 41259 6803
rect 41293 6769 41309 6803
rect 41345 6790 41379 6811
rect 41155 6710 41207 6739
rect 41345 6735 41379 6756
rect 40938 6619 40954 6653
rect 40988 6642 41004 6653
rect 40938 6608 40956 6619
rect 40990 6608 41004 6642
rect 41155 6638 41191 6710
rect 41246 6701 41379 6735
rect 41550 6797 41616 6809
rect 41550 6763 41566 6797
rect 41600 6763 41616 6797
rect 41550 6746 41616 6763
rect 41246 6650 41280 6701
rect 41550 6695 41566 6746
rect 41600 6695 41616 6746
rect 41550 6683 41616 6695
rect 41650 6797 41696 6843
rect 41684 6763 41696 6797
rect 41650 6729 41696 6763
rect 41684 6695 41696 6729
rect 41920 6828 41926 6862
rect 41960 6828 41968 6862
rect 42552 6856 42558 6876
rect 42592 6856 42598 6890
rect 42552 6846 42598 6856
rect 42680 6851 42709 6885
rect 42743 6851 42801 6885
rect 42835 6851 42893 6885
rect 42927 6851 42956 6885
rect 41920 6740 41968 6828
rect 42294 6785 42310 6819
rect 42344 6818 42360 6819
rect 42344 6786 42506 6818
rect 42746 6810 42812 6817
rect 42740 6805 42812 6810
rect 42740 6786 42762 6805
rect 42344 6785 42762 6786
rect 42294 6782 42762 6785
rect 42470 6771 42762 6782
rect 42796 6771 42812 6805
rect 42470 6750 42812 6771
rect 42166 6740 42200 6742
rect 41920 6723 42200 6740
rect 41920 6706 42166 6723
rect 40938 6605 41004 6608
rect 41150 6636 41191 6638
rect 41150 6602 41152 6636
rect 41186 6602 41191 6636
rect 41150 6600 41191 6602
rect 40858 6553 40924 6571
rect 40858 6519 40874 6553
rect 40908 6519 40924 6553
rect 40858 6485 40924 6519
rect 40858 6451 40874 6485
rect 40908 6451 40924 6485
rect 40858 6417 40924 6451
rect 40858 6383 40874 6417
rect 40908 6383 40924 6417
rect 40858 6375 40924 6383
rect 40958 6553 41000 6569
rect 40992 6519 41000 6553
rect 40958 6485 41000 6519
rect 40992 6451 41000 6485
rect 40958 6417 41000 6451
rect 40992 6383 41000 6417
rect 40429 6349 40468 6374
rect 39980 6297 39996 6331
rect 40030 6297 40046 6331
rect 40186 6310 40468 6349
rect 40958 6341 41000 6383
rect 41155 6550 41191 6600
rect 41225 6634 41280 6650
rect 41259 6600 41280 6634
rect 41225 6584 41280 6600
rect 41325 6648 41393 6665
rect 41325 6647 41345 6648
rect 41325 6613 41343 6647
rect 41379 6614 41393 6648
rect 41377 6613 41393 6614
rect 41325 6591 41393 6613
rect 41246 6555 41280 6584
rect 41550 6563 41596 6683
rect 41650 6679 41696 6695
rect 41868 6658 41884 6659
rect 41630 6611 41646 6645
rect 41680 6638 41696 6645
rect 41748 6638 41884 6658
rect 41680 6625 41884 6638
rect 41918 6625 41934 6659
rect 41680 6624 41934 6625
rect 41680 6611 41788 6624
rect 41868 6622 41934 6624
rect 42166 6655 42200 6657
rect 41630 6597 41788 6611
rect 41644 6596 41788 6597
rect 42166 6619 42200 6621
rect 41840 6563 41874 6582
rect 41155 6500 41209 6550
rect 41246 6521 41381 6555
rect 41155 6466 41173 6500
rect 41207 6466 41209 6500
rect 41345 6487 41381 6521
rect 41155 6419 41209 6466
rect 41155 6385 41173 6419
rect 41207 6385 41209 6419
rect 41155 6369 41209 6385
rect 41243 6453 41259 6487
rect 41293 6453 41309 6487
rect 41243 6419 41309 6453
rect 41243 6385 41259 6419
rect 41293 6385 41309 6419
rect 40354 6308 40468 6310
rect 40626 6297 40642 6331
rect 40676 6297 40692 6331
rect 40792 6307 40821 6341
rect 40855 6307 40913 6341
rect 40947 6307 41005 6341
rect 41039 6307 41068 6341
rect 41243 6335 41309 6385
rect 41379 6453 41381 6487
rect 41345 6419 41381 6453
rect 41379 6385 41381 6419
rect 41345 6369 41381 6385
rect 41550 6545 41616 6563
rect 41550 6511 41566 6545
rect 41600 6511 41616 6545
rect 41550 6477 41616 6511
rect 41550 6443 41566 6477
rect 41600 6443 41616 6477
rect 41550 6409 41616 6443
rect 41550 6375 41566 6409
rect 41600 6375 41616 6409
rect 41550 6367 41616 6375
rect 41650 6545 41692 6561
rect 41684 6511 41692 6545
rect 41650 6477 41692 6511
rect 41684 6443 41692 6477
rect 41650 6409 41692 6443
rect 41840 6495 41874 6497
rect 41840 6459 41874 6461
rect 41684 6375 41692 6409
rect 40959 6300 40993 6307
rect 41138 6301 41167 6335
rect 41201 6301 41259 6335
rect 41293 6301 41351 6335
rect 41385 6301 41414 6335
rect 41650 6333 41692 6375
rect 41800 6393 41840 6414
rect 41928 6563 41962 6582
rect 42166 6534 42200 6553
rect 42262 6723 42296 6742
rect 42262 6655 42296 6657
rect 42262 6619 42296 6621
rect 42262 6534 42296 6553
rect 42358 6723 42392 6742
rect 42746 6737 42812 6750
rect 42746 6703 42762 6737
rect 42796 6703 42812 6737
rect 42746 6691 42812 6703
rect 42846 6805 42892 6851
rect 43026 6845 43055 6879
rect 43089 6845 43147 6879
rect 43181 6845 43239 6879
rect 43273 6845 43302 6879
rect 42880 6771 42892 6805
rect 42846 6737 42892 6771
rect 42880 6703 42892 6737
rect 42358 6655 42392 6657
rect 42514 6625 42530 6659
rect 42564 6625 42580 6659
rect 42358 6619 42392 6621
rect 42358 6534 42392 6553
rect 42486 6563 42520 6582
rect 41928 6495 41962 6497
rect 42486 6495 42520 6497
rect 41928 6459 41962 6461
rect 42198 6457 42214 6491
rect 42248 6457 42264 6491
rect 42486 6459 42520 6461
rect 41874 6393 41876 6414
rect 41800 6374 41876 6393
rect 41962 6393 42486 6418
rect 42574 6563 42608 6582
rect 42574 6495 42608 6497
rect 42574 6459 42608 6461
rect 42520 6393 42522 6418
rect 41928 6385 42522 6393
rect 41928 6374 42164 6385
rect 41484 6299 41513 6333
rect 41547 6299 41605 6333
rect 41639 6299 41697 6333
rect 41731 6299 41760 6333
rect 40046 6212 40092 6218
rect 40046 6210 40534 6212
rect 40046 6176 40054 6210
rect 40088 6193 40534 6210
rect 40088 6188 40484 6193
rect 40088 6178 40363 6188
rect 40088 6176 40092 6178
rect 40046 6174 40092 6176
rect 40264 6154 40363 6178
rect 40397 6159 40484 6188
rect 40518 6168 40534 6193
rect 40518 6159 40659 6168
rect 40397 6154 40659 6159
rect 40264 6134 40659 6154
rect 40388 6050 40404 6084
rect 40438 6050 40574 6084
rect 39912 6000 40294 6016
rect 39912 5976 40260 6000
rect 40260 5930 40294 5964
rect 40260 5878 40294 5894
rect 40356 6000 40390 6016
rect 40356 5930 40390 5964
rect 40356 5878 40390 5894
rect 40452 6000 40486 6016
rect 40452 5930 40486 5964
rect 40452 5878 40486 5894
rect 38726 5797 38755 5831
rect 38789 5797 38847 5831
rect 38881 5797 38939 5831
rect 38973 5797 39002 5831
rect 39800 5797 39829 5831
rect 39863 5797 39921 5831
rect 39955 5797 40013 5831
rect 40047 5797 40076 5831
rect 40292 5810 40308 5844
rect 40342 5810 40358 5844
rect 38745 5753 38799 5797
rect 38745 5719 38765 5753
rect 38745 5685 38799 5719
rect 38745 5651 38765 5685
rect 38745 5635 38799 5651
rect 38833 5753 38899 5763
rect 38833 5719 38849 5753
rect 38883 5719 38899 5753
rect 38833 5710 38899 5719
rect 38833 5685 38851 5710
rect 38833 5651 38849 5685
rect 38885 5676 38899 5710
rect 38883 5651 38899 5676
rect 38833 5635 38899 5651
rect 38933 5753 38981 5797
rect 38967 5719 38981 5753
rect 38933 5685 38981 5719
rect 38967 5651 38981 5685
rect 38933 5635 38981 5651
rect 39819 5753 39873 5797
rect 39819 5719 39839 5753
rect 39819 5685 39873 5719
rect 39819 5651 39839 5685
rect 39819 5635 39873 5651
rect 39907 5753 39973 5763
rect 39907 5719 39923 5753
rect 39957 5719 39973 5753
rect 39907 5715 39973 5719
rect 39907 5681 39921 5715
rect 39955 5685 39973 5715
rect 39907 5651 39923 5681
rect 39957 5651 39973 5685
rect 39907 5635 39973 5651
rect 40007 5753 40055 5797
rect 40041 5719 40055 5753
rect 40404 5729 40420 5763
rect 40454 5729 40470 5763
rect 40007 5685 40055 5719
rect 40041 5651 40055 5685
rect 40007 5635 40055 5651
rect 40276 5667 40310 5686
rect 38743 5594 38763 5599
rect 38743 5560 38760 5594
rect 38797 5565 38813 5599
rect 38794 5560 38813 5565
rect 38743 5549 38813 5560
rect 38847 5515 38881 5635
rect 38915 5565 38931 5599
rect 38965 5590 38985 5599
rect 38915 5556 38933 5565
rect 38967 5556 38985 5590
rect 38915 5549 38985 5556
rect 39817 5592 39837 5599
rect 39817 5558 39835 5592
rect 39871 5565 39887 5599
rect 39869 5558 39887 5565
rect 39817 5549 39887 5558
rect 39921 5515 39955 5635
rect 40276 5599 40310 5601
rect 39989 5565 40005 5599
rect 40039 5592 40059 5599
rect 39989 5558 40009 5565
rect 40043 5558 40059 5592
rect 39989 5549 40059 5558
rect 40276 5563 40310 5565
rect 38420 5435 38686 5436
rect 38420 5401 38436 5435
rect 38470 5401 38686 5435
rect 38420 5400 38686 5401
rect 38745 5499 38811 5515
rect 38745 5465 38777 5499
rect 38847 5499 38983 5515
rect 38847 5481 38933 5499
rect 38745 5431 38811 5465
rect 38103 5363 38169 5397
rect 38103 5329 38119 5363
rect 38153 5329 38169 5363
rect 38745 5397 38777 5431
rect 38745 5363 38811 5397
rect 38103 5324 38169 5329
rect 38296 5329 38578 5362
rect 38296 5295 38386 5329
rect 38420 5327 38578 5329
rect 38420 5295 38505 5327
rect 38296 5293 38505 5295
rect 38539 5293 38578 5327
rect 38296 5287 38578 5293
rect 38745 5329 38777 5363
rect 38745 5287 38811 5329
rect 38917 5465 38933 5481
rect 38967 5465 38983 5499
rect 38917 5431 38983 5465
rect 38917 5397 38933 5431
rect 38967 5397 38983 5431
rect 38917 5363 38983 5397
rect 38917 5329 38933 5363
rect 38967 5329 38983 5363
rect 38917 5324 38983 5329
rect 39819 5499 39885 5515
rect 39819 5465 39851 5499
rect 39921 5499 40057 5515
rect 39921 5481 40007 5499
rect 39819 5431 39885 5465
rect 39819 5397 39851 5431
rect 39819 5363 39885 5397
rect 39819 5329 39851 5363
rect 39819 5287 39885 5329
rect 39991 5465 40007 5481
rect 40041 5465 40057 5499
rect 40276 5478 40310 5497
rect 40372 5667 40406 5686
rect 40372 5599 40406 5601
rect 40372 5563 40406 5565
rect 40372 5478 40406 5497
rect 40468 5667 40502 5686
rect 40468 5599 40502 5601
rect 40468 5563 40502 5565
rect 40468 5478 40502 5497
rect 39991 5431 40057 5465
rect 39991 5397 40007 5431
rect 40041 5397 40057 5431
rect 40308 5436 40374 5438
rect 40540 5436 40574 6050
rect 40625 5831 40659 6134
rect 40856 5831 40890 6042
rect 41800 6016 41834 6374
rect 42074 6351 42164 6374
rect 42198 6383 42522 6385
rect 42198 6351 42283 6383
rect 42074 6349 42283 6351
rect 42317 6374 42522 6383
rect 42574 6374 42608 6393
rect 42746 6571 42792 6691
rect 42846 6687 42892 6703
rect 43043 6773 43095 6811
rect 43043 6739 43061 6773
rect 43131 6803 43197 6845
rect 43372 6843 43401 6877
rect 43435 6843 43493 6877
rect 43527 6843 43585 6877
rect 43619 6843 43648 6877
rect 43808 6862 43856 6874
rect 44070 6866 44086 6900
rect 44120 6866 44136 6900
rect 44436 6890 44486 6960
rect 45920 6934 45954 6950
rect 46016 7056 46050 7072
rect 46112 7058 46146 7072
rect 46230 7058 46450 7080
rect 46110 7056 46450 7058
rect 46110 7022 46112 7056
rect 46146 7044 46450 7056
rect 46146 7022 46266 7044
rect 46016 6986 46050 7020
rect 46111 7020 46112 7022
rect 46111 6986 46146 7020
rect 46414 6996 46450 7044
rect 46111 6985 46112 6986
rect 46016 6934 46050 6950
rect 46112 6934 46146 6950
rect 46318 6960 46450 6996
rect 47808 7056 47842 7072
rect 47808 6986 47842 7020
rect 44436 6876 44446 6890
rect 43131 6769 43147 6803
rect 43181 6769 43197 6803
rect 43233 6790 43267 6811
rect 43043 6710 43095 6739
rect 43233 6735 43267 6756
rect 42826 6619 42842 6653
rect 42876 6642 42892 6653
rect 42826 6608 42844 6619
rect 42878 6608 42892 6642
rect 43043 6638 43079 6710
rect 43134 6701 43267 6735
rect 43438 6797 43504 6809
rect 43438 6763 43454 6797
rect 43488 6763 43504 6797
rect 43438 6746 43504 6763
rect 43134 6650 43168 6701
rect 43438 6695 43454 6746
rect 43488 6695 43504 6746
rect 43438 6683 43504 6695
rect 43538 6797 43584 6843
rect 43572 6763 43584 6797
rect 43538 6729 43584 6763
rect 43572 6695 43584 6729
rect 43808 6828 43814 6862
rect 43848 6828 43856 6862
rect 44440 6856 44446 6876
rect 44480 6856 44486 6890
rect 44440 6846 44486 6856
rect 44568 6851 44597 6885
rect 44631 6851 44689 6885
rect 44723 6851 44781 6885
rect 44815 6851 44844 6885
rect 43808 6740 43856 6828
rect 44182 6785 44198 6819
rect 44232 6818 44248 6819
rect 44232 6786 44394 6818
rect 44634 6810 44700 6817
rect 44628 6805 44700 6810
rect 44628 6786 44650 6805
rect 44232 6785 44650 6786
rect 44182 6782 44650 6785
rect 44358 6771 44650 6782
rect 44684 6771 44700 6805
rect 44358 6750 44700 6771
rect 44054 6740 44088 6742
rect 43808 6723 44088 6740
rect 43808 6706 44054 6723
rect 42826 6605 42892 6608
rect 43038 6636 43079 6638
rect 43038 6602 43040 6636
rect 43074 6602 43079 6636
rect 43038 6600 43079 6602
rect 42746 6553 42812 6571
rect 42746 6519 42762 6553
rect 42796 6519 42812 6553
rect 42746 6485 42812 6519
rect 42746 6451 42762 6485
rect 42796 6451 42812 6485
rect 42746 6417 42812 6451
rect 42746 6383 42762 6417
rect 42796 6383 42812 6417
rect 42746 6375 42812 6383
rect 42846 6553 42888 6569
rect 42880 6519 42888 6553
rect 42846 6485 42888 6519
rect 42880 6451 42888 6485
rect 42846 6417 42888 6451
rect 42880 6383 42888 6417
rect 42317 6349 42356 6374
rect 41868 6297 41884 6331
rect 41918 6297 41934 6331
rect 42074 6310 42356 6349
rect 42846 6341 42888 6383
rect 43043 6550 43079 6600
rect 43113 6634 43168 6650
rect 43147 6600 43168 6634
rect 43113 6584 43168 6600
rect 43213 6648 43281 6665
rect 43213 6647 43233 6648
rect 43213 6613 43231 6647
rect 43267 6614 43281 6648
rect 43265 6613 43281 6614
rect 43213 6591 43281 6613
rect 43134 6555 43168 6584
rect 43438 6563 43484 6683
rect 43538 6679 43584 6695
rect 43756 6658 43772 6659
rect 43518 6611 43534 6645
rect 43568 6638 43584 6645
rect 43636 6638 43772 6658
rect 43568 6625 43772 6638
rect 43806 6625 43822 6659
rect 43568 6624 43822 6625
rect 43568 6611 43676 6624
rect 43756 6622 43822 6624
rect 44054 6655 44088 6657
rect 43518 6597 43676 6611
rect 43532 6596 43676 6597
rect 44054 6619 44088 6621
rect 43728 6563 43762 6582
rect 43043 6500 43097 6550
rect 43134 6521 43269 6555
rect 43043 6466 43061 6500
rect 43095 6466 43097 6500
rect 43233 6487 43269 6521
rect 43043 6419 43097 6466
rect 43043 6385 43061 6419
rect 43095 6385 43097 6419
rect 43043 6369 43097 6385
rect 43131 6453 43147 6487
rect 43181 6453 43197 6487
rect 43131 6419 43197 6453
rect 43131 6385 43147 6419
rect 43181 6385 43197 6419
rect 42242 6308 42356 6310
rect 42514 6297 42530 6331
rect 42564 6297 42580 6331
rect 42680 6307 42709 6341
rect 42743 6307 42801 6341
rect 42835 6307 42893 6341
rect 42927 6307 42956 6341
rect 43131 6335 43197 6385
rect 43267 6453 43269 6487
rect 43233 6419 43269 6453
rect 43267 6385 43269 6419
rect 43233 6369 43269 6385
rect 43438 6545 43504 6563
rect 43438 6511 43454 6545
rect 43488 6511 43504 6545
rect 43438 6477 43504 6511
rect 43438 6443 43454 6477
rect 43488 6443 43504 6477
rect 43438 6409 43504 6443
rect 43438 6375 43454 6409
rect 43488 6375 43504 6409
rect 43438 6367 43504 6375
rect 43538 6545 43580 6561
rect 43572 6511 43580 6545
rect 43538 6477 43580 6511
rect 43572 6443 43580 6477
rect 43538 6409 43580 6443
rect 43728 6495 43762 6497
rect 43728 6459 43762 6461
rect 43572 6375 43580 6409
rect 42847 6300 42881 6307
rect 43026 6301 43055 6335
rect 43089 6301 43147 6335
rect 43181 6301 43239 6335
rect 43273 6301 43302 6335
rect 43538 6333 43580 6375
rect 43688 6393 43728 6414
rect 43816 6563 43850 6582
rect 44054 6534 44088 6553
rect 44150 6723 44184 6742
rect 44150 6655 44184 6657
rect 44150 6619 44184 6621
rect 44150 6534 44184 6553
rect 44246 6723 44280 6742
rect 44634 6737 44700 6750
rect 44634 6703 44650 6737
rect 44684 6703 44700 6737
rect 44634 6691 44700 6703
rect 44734 6805 44780 6851
rect 44908 6845 44937 6879
rect 44971 6845 45029 6879
rect 45063 6845 45121 6879
rect 45155 6845 45184 6879
rect 44768 6771 44780 6805
rect 44734 6737 44780 6771
rect 44768 6703 44780 6737
rect 44246 6655 44280 6657
rect 44402 6625 44418 6659
rect 44452 6625 44468 6659
rect 44246 6619 44280 6621
rect 44246 6534 44280 6553
rect 44374 6563 44408 6582
rect 43816 6495 43850 6497
rect 44374 6495 44408 6497
rect 43816 6459 43850 6461
rect 44086 6457 44102 6491
rect 44136 6457 44152 6491
rect 44374 6459 44408 6461
rect 43762 6393 43764 6414
rect 43688 6374 43764 6393
rect 43850 6393 44374 6418
rect 44462 6563 44496 6582
rect 44462 6495 44496 6497
rect 44462 6459 44496 6461
rect 44408 6393 44410 6418
rect 43816 6385 44410 6393
rect 43816 6374 44052 6385
rect 43372 6299 43401 6333
rect 43435 6299 43493 6333
rect 43527 6299 43585 6333
rect 43619 6299 43648 6333
rect 41934 6212 41980 6218
rect 41934 6210 42422 6212
rect 41934 6176 41942 6210
rect 41976 6193 42422 6210
rect 41976 6188 42372 6193
rect 41976 6178 42251 6188
rect 41976 6176 41980 6178
rect 41934 6174 41980 6176
rect 42152 6154 42251 6178
rect 42285 6159 42372 6188
rect 42406 6168 42422 6193
rect 42406 6159 42547 6168
rect 42285 6154 42547 6159
rect 42152 6134 42547 6154
rect 42276 6050 42292 6084
rect 42326 6050 42462 6084
rect 41800 6000 42182 6016
rect 41800 5976 42148 6000
rect 42148 5930 42182 5964
rect 42148 5878 42182 5894
rect 42244 6000 42278 6016
rect 42244 5930 42278 5964
rect 42244 5878 42278 5894
rect 42340 6000 42374 6016
rect 42340 5930 42374 5964
rect 42340 5878 42374 5894
rect 40614 5797 40643 5831
rect 40677 5797 40735 5831
rect 40769 5797 40827 5831
rect 40861 5797 40890 5831
rect 41688 5797 41717 5831
rect 41751 5797 41809 5831
rect 41843 5797 41901 5831
rect 41935 5797 41964 5831
rect 42180 5810 42196 5844
rect 42230 5810 42246 5844
rect 40633 5753 40687 5797
rect 40633 5719 40653 5753
rect 40633 5685 40687 5719
rect 40633 5651 40653 5685
rect 40633 5635 40687 5651
rect 40721 5753 40787 5763
rect 40721 5719 40737 5753
rect 40771 5719 40787 5753
rect 40721 5710 40787 5719
rect 40721 5685 40739 5710
rect 40721 5651 40737 5685
rect 40773 5676 40787 5710
rect 40771 5651 40787 5676
rect 40721 5635 40787 5651
rect 40821 5753 40869 5797
rect 40855 5719 40869 5753
rect 40821 5685 40869 5719
rect 40855 5651 40869 5685
rect 40821 5635 40869 5651
rect 41707 5753 41761 5797
rect 41707 5719 41727 5753
rect 41707 5685 41761 5719
rect 41707 5651 41727 5685
rect 41707 5635 41761 5651
rect 41795 5753 41861 5763
rect 41795 5719 41811 5753
rect 41845 5719 41861 5753
rect 41795 5715 41861 5719
rect 41795 5681 41809 5715
rect 41843 5685 41861 5715
rect 41795 5651 41811 5681
rect 41845 5651 41861 5685
rect 41795 5635 41861 5651
rect 41895 5753 41943 5797
rect 41929 5719 41943 5753
rect 42292 5729 42308 5763
rect 42342 5729 42358 5763
rect 41895 5685 41943 5719
rect 41929 5651 41943 5685
rect 41895 5635 41943 5651
rect 42164 5667 42198 5686
rect 40631 5594 40651 5599
rect 40631 5560 40648 5594
rect 40685 5565 40701 5599
rect 40682 5560 40701 5565
rect 40631 5549 40701 5560
rect 40735 5515 40769 5635
rect 40803 5565 40819 5599
rect 40853 5590 40873 5599
rect 40803 5556 40821 5565
rect 40855 5556 40873 5590
rect 40803 5549 40873 5556
rect 41705 5592 41725 5599
rect 41705 5558 41723 5592
rect 41759 5565 41775 5599
rect 41757 5558 41775 5565
rect 41705 5549 41775 5558
rect 41809 5515 41843 5635
rect 42164 5599 42198 5601
rect 41877 5565 41893 5599
rect 41927 5592 41947 5599
rect 41877 5558 41897 5565
rect 41931 5558 41947 5592
rect 41877 5549 41947 5558
rect 42164 5563 42198 5565
rect 40308 5435 40574 5436
rect 40308 5401 40324 5435
rect 40358 5401 40574 5435
rect 40308 5400 40574 5401
rect 40633 5499 40699 5515
rect 40633 5465 40665 5499
rect 40735 5499 40871 5515
rect 40735 5481 40821 5499
rect 40633 5431 40699 5465
rect 39991 5363 40057 5397
rect 39991 5329 40007 5363
rect 40041 5329 40057 5363
rect 40633 5397 40665 5431
rect 40633 5363 40699 5397
rect 39991 5324 40057 5329
rect 40184 5329 40466 5362
rect 40184 5295 40274 5329
rect 40308 5327 40466 5329
rect 40308 5295 40393 5327
rect 40184 5293 40393 5295
rect 40427 5293 40466 5327
rect 40184 5287 40466 5293
rect 40633 5329 40665 5363
rect 40633 5287 40699 5329
rect 40805 5465 40821 5481
rect 40855 5465 40871 5499
rect 40805 5431 40871 5465
rect 40805 5397 40821 5431
rect 40855 5397 40871 5431
rect 40805 5363 40871 5397
rect 40805 5329 40821 5363
rect 40855 5329 40871 5363
rect 40805 5324 40871 5329
rect 41707 5499 41773 5515
rect 41707 5465 41739 5499
rect 41809 5499 41945 5515
rect 41809 5481 41895 5499
rect 41707 5431 41773 5465
rect 41707 5397 41739 5431
rect 41707 5363 41773 5397
rect 41707 5329 41739 5363
rect 41707 5287 41773 5329
rect 41879 5465 41895 5481
rect 41929 5465 41945 5499
rect 42164 5478 42198 5497
rect 42260 5667 42294 5686
rect 42260 5599 42294 5601
rect 42260 5563 42294 5565
rect 42260 5478 42294 5497
rect 42356 5667 42390 5686
rect 42356 5599 42390 5601
rect 42356 5563 42390 5565
rect 42356 5478 42390 5497
rect 41879 5431 41945 5465
rect 41879 5397 41895 5431
rect 41929 5397 41945 5431
rect 42196 5436 42262 5438
rect 42428 5436 42462 6050
rect 42513 5831 42547 6134
rect 42744 5831 42778 6042
rect 43688 6016 43722 6374
rect 43962 6351 44052 6374
rect 44086 6383 44410 6385
rect 44086 6351 44171 6383
rect 43962 6349 44171 6351
rect 44205 6374 44410 6383
rect 44462 6374 44496 6393
rect 44634 6571 44680 6691
rect 44734 6687 44780 6703
rect 44925 6773 44977 6811
rect 44925 6739 44943 6773
rect 45013 6803 45079 6845
rect 45254 6843 45283 6877
rect 45317 6843 45375 6877
rect 45409 6843 45467 6877
rect 45501 6843 45530 6877
rect 45690 6862 45738 6874
rect 45952 6866 45968 6900
rect 46002 6866 46018 6900
rect 46318 6890 46368 6960
rect 47808 6934 47842 6950
rect 47904 7056 47938 7072
rect 48000 7058 48034 7072
rect 48118 7058 48338 7080
rect 47998 7056 48338 7058
rect 47998 7022 48000 7056
rect 48034 7044 48338 7056
rect 48034 7022 48154 7044
rect 47904 6986 47938 7020
rect 47999 7020 48000 7022
rect 47999 6986 48034 7020
rect 48302 6996 48338 7044
rect 47999 6985 48000 6986
rect 47904 6934 47938 6950
rect 48000 6934 48034 6950
rect 48206 6960 48338 6996
rect 49696 7056 49730 7072
rect 49696 6986 49730 7020
rect 46318 6876 46328 6890
rect 45013 6769 45029 6803
rect 45063 6769 45079 6803
rect 45115 6790 45149 6811
rect 44925 6710 44977 6739
rect 45115 6735 45149 6756
rect 44714 6619 44730 6653
rect 44764 6642 44780 6653
rect 44714 6608 44732 6619
rect 44766 6608 44780 6642
rect 44925 6638 44961 6710
rect 45016 6701 45149 6735
rect 45320 6797 45386 6809
rect 45320 6763 45336 6797
rect 45370 6763 45386 6797
rect 45320 6746 45386 6763
rect 45016 6650 45050 6701
rect 45320 6695 45336 6746
rect 45370 6695 45386 6746
rect 45320 6683 45386 6695
rect 45420 6797 45466 6843
rect 45454 6763 45466 6797
rect 45420 6729 45466 6763
rect 45454 6695 45466 6729
rect 45690 6828 45696 6862
rect 45730 6828 45738 6862
rect 46322 6856 46328 6876
rect 46362 6856 46368 6890
rect 46322 6846 46368 6856
rect 46450 6851 46479 6885
rect 46513 6851 46571 6885
rect 46605 6851 46663 6885
rect 46697 6851 46726 6885
rect 45690 6740 45738 6828
rect 46064 6785 46080 6819
rect 46114 6818 46130 6819
rect 46114 6786 46276 6818
rect 46516 6810 46582 6817
rect 46510 6805 46582 6810
rect 46510 6786 46532 6805
rect 46114 6785 46532 6786
rect 46064 6782 46532 6785
rect 46240 6771 46532 6782
rect 46566 6771 46582 6805
rect 46240 6750 46582 6771
rect 45936 6740 45970 6742
rect 45690 6723 45970 6740
rect 45690 6706 45936 6723
rect 44714 6605 44780 6608
rect 44920 6636 44961 6638
rect 44920 6602 44922 6636
rect 44956 6602 44961 6636
rect 44920 6600 44961 6602
rect 44634 6553 44700 6571
rect 44634 6519 44650 6553
rect 44684 6519 44700 6553
rect 44634 6485 44700 6519
rect 44634 6451 44650 6485
rect 44684 6451 44700 6485
rect 44634 6417 44700 6451
rect 44634 6383 44650 6417
rect 44684 6383 44700 6417
rect 44634 6375 44700 6383
rect 44734 6553 44776 6569
rect 44768 6519 44776 6553
rect 44734 6485 44776 6519
rect 44768 6451 44776 6485
rect 44734 6417 44776 6451
rect 44768 6383 44776 6417
rect 44205 6349 44244 6374
rect 43756 6297 43772 6331
rect 43806 6297 43822 6331
rect 43962 6310 44244 6349
rect 44734 6341 44776 6383
rect 44925 6550 44961 6600
rect 44995 6634 45050 6650
rect 45029 6600 45050 6634
rect 44995 6584 45050 6600
rect 45095 6648 45163 6665
rect 45095 6647 45115 6648
rect 45095 6613 45113 6647
rect 45149 6614 45163 6648
rect 45147 6613 45163 6614
rect 45095 6591 45163 6613
rect 45016 6555 45050 6584
rect 45320 6563 45366 6683
rect 45420 6679 45466 6695
rect 45638 6658 45654 6659
rect 45400 6611 45416 6645
rect 45450 6638 45466 6645
rect 45518 6638 45654 6658
rect 45450 6625 45654 6638
rect 45688 6625 45704 6659
rect 45450 6624 45704 6625
rect 45450 6611 45558 6624
rect 45638 6622 45704 6624
rect 45936 6655 45970 6657
rect 45400 6597 45558 6611
rect 45414 6596 45558 6597
rect 45936 6619 45970 6621
rect 45610 6563 45644 6582
rect 44925 6500 44979 6550
rect 45016 6521 45151 6555
rect 44925 6466 44943 6500
rect 44977 6466 44979 6500
rect 45115 6487 45151 6521
rect 44925 6419 44979 6466
rect 44925 6385 44943 6419
rect 44977 6385 44979 6419
rect 44925 6369 44979 6385
rect 45013 6453 45029 6487
rect 45063 6453 45079 6487
rect 45013 6419 45079 6453
rect 45013 6385 45029 6419
rect 45063 6385 45079 6419
rect 44130 6308 44244 6310
rect 44402 6297 44418 6331
rect 44452 6297 44468 6331
rect 44568 6307 44597 6341
rect 44631 6307 44689 6341
rect 44723 6307 44781 6341
rect 44815 6307 44844 6341
rect 45013 6335 45079 6385
rect 45149 6453 45151 6487
rect 45115 6419 45151 6453
rect 45149 6385 45151 6419
rect 45115 6369 45151 6385
rect 45320 6545 45386 6563
rect 45320 6511 45336 6545
rect 45370 6511 45386 6545
rect 45320 6477 45386 6511
rect 45320 6443 45336 6477
rect 45370 6443 45386 6477
rect 45320 6409 45386 6443
rect 45320 6375 45336 6409
rect 45370 6375 45386 6409
rect 45320 6367 45386 6375
rect 45420 6545 45462 6561
rect 45454 6511 45462 6545
rect 45420 6477 45462 6511
rect 45454 6443 45462 6477
rect 45420 6409 45462 6443
rect 45610 6495 45644 6497
rect 45610 6459 45644 6461
rect 45454 6375 45462 6409
rect 44735 6300 44769 6307
rect 44908 6301 44937 6335
rect 44971 6301 45029 6335
rect 45063 6301 45121 6335
rect 45155 6301 45184 6335
rect 45420 6333 45462 6375
rect 45570 6393 45610 6414
rect 45698 6563 45732 6582
rect 45936 6534 45970 6553
rect 46032 6723 46066 6742
rect 46032 6655 46066 6657
rect 46032 6619 46066 6621
rect 46032 6534 46066 6553
rect 46128 6723 46162 6742
rect 46516 6737 46582 6750
rect 46516 6703 46532 6737
rect 46566 6703 46582 6737
rect 46516 6691 46582 6703
rect 46616 6805 46662 6851
rect 46796 6845 46825 6879
rect 46859 6845 46917 6879
rect 46951 6845 47009 6879
rect 47043 6845 47072 6879
rect 46650 6771 46662 6805
rect 46616 6737 46662 6771
rect 46650 6703 46662 6737
rect 46128 6655 46162 6657
rect 46284 6625 46300 6659
rect 46334 6625 46350 6659
rect 46128 6619 46162 6621
rect 46128 6534 46162 6553
rect 46256 6563 46290 6582
rect 45698 6495 45732 6497
rect 46256 6495 46290 6497
rect 45698 6459 45732 6461
rect 45968 6457 45984 6491
rect 46018 6457 46034 6491
rect 46256 6459 46290 6461
rect 45644 6393 45646 6414
rect 45570 6374 45646 6393
rect 45732 6393 46256 6418
rect 46344 6563 46378 6582
rect 46344 6495 46378 6497
rect 46344 6459 46378 6461
rect 46290 6393 46292 6418
rect 45698 6385 46292 6393
rect 45698 6374 45934 6385
rect 45254 6299 45283 6333
rect 45317 6299 45375 6333
rect 45409 6299 45467 6333
rect 45501 6299 45530 6333
rect 43822 6212 43868 6218
rect 43822 6210 44310 6212
rect 43822 6176 43830 6210
rect 43864 6193 44310 6210
rect 43864 6188 44260 6193
rect 43864 6178 44139 6188
rect 43864 6176 43868 6178
rect 43822 6174 43868 6176
rect 44040 6154 44139 6178
rect 44173 6159 44260 6188
rect 44294 6168 44310 6193
rect 44294 6159 44435 6168
rect 44173 6154 44435 6159
rect 44040 6134 44435 6154
rect 44164 6050 44180 6084
rect 44214 6050 44350 6084
rect 43688 6000 44070 6016
rect 43688 5976 44036 6000
rect 44036 5930 44070 5964
rect 44036 5878 44070 5894
rect 44132 6000 44166 6016
rect 44132 5930 44166 5964
rect 44132 5878 44166 5894
rect 44228 6000 44262 6016
rect 44228 5930 44262 5964
rect 44228 5878 44262 5894
rect 42502 5797 42531 5831
rect 42565 5797 42623 5831
rect 42657 5797 42715 5831
rect 42749 5797 42778 5831
rect 43576 5797 43605 5831
rect 43639 5797 43697 5831
rect 43731 5797 43789 5831
rect 43823 5797 43852 5831
rect 44068 5810 44084 5844
rect 44118 5810 44134 5844
rect 42521 5753 42575 5797
rect 42521 5719 42541 5753
rect 42521 5685 42575 5719
rect 42521 5651 42541 5685
rect 42521 5635 42575 5651
rect 42609 5753 42675 5763
rect 42609 5719 42625 5753
rect 42659 5719 42675 5753
rect 42609 5710 42675 5719
rect 42609 5685 42627 5710
rect 42609 5651 42625 5685
rect 42661 5676 42675 5710
rect 42659 5651 42675 5676
rect 42609 5635 42675 5651
rect 42709 5753 42757 5797
rect 42743 5719 42757 5753
rect 42709 5685 42757 5719
rect 42743 5651 42757 5685
rect 42709 5635 42757 5651
rect 43595 5753 43649 5797
rect 43595 5719 43615 5753
rect 43595 5685 43649 5719
rect 43595 5651 43615 5685
rect 43595 5635 43649 5651
rect 43683 5753 43749 5763
rect 43683 5719 43699 5753
rect 43733 5719 43749 5753
rect 43683 5715 43749 5719
rect 43683 5681 43697 5715
rect 43731 5685 43749 5715
rect 43683 5651 43699 5681
rect 43733 5651 43749 5685
rect 43683 5635 43749 5651
rect 43783 5753 43831 5797
rect 43817 5719 43831 5753
rect 44180 5729 44196 5763
rect 44230 5729 44246 5763
rect 43783 5685 43831 5719
rect 43817 5651 43831 5685
rect 43783 5635 43831 5651
rect 44052 5667 44086 5686
rect 42519 5594 42539 5599
rect 42519 5560 42536 5594
rect 42573 5565 42589 5599
rect 42570 5560 42589 5565
rect 42519 5549 42589 5560
rect 42623 5515 42657 5635
rect 42691 5565 42707 5599
rect 42741 5590 42761 5599
rect 42691 5556 42709 5565
rect 42743 5556 42761 5590
rect 42691 5549 42761 5556
rect 43593 5592 43613 5599
rect 43593 5558 43611 5592
rect 43647 5565 43663 5599
rect 43645 5558 43663 5565
rect 43593 5549 43663 5558
rect 43697 5515 43731 5635
rect 44052 5599 44086 5601
rect 43765 5565 43781 5599
rect 43815 5592 43835 5599
rect 43765 5558 43785 5565
rect 43819 5558 43835 5592
rect 43765 5549 43835 5558
rect 44052 5563 44086 5565
rect 42196 5435 42462 5436
rect 42196 5401 42212 5435
rect 42246 5401 42462 5435
rect 42196 5400 42462 5401
rect 42521 5499 42587 5515
rect 42521 5465 42553 5499
rect 42623 5499 42759 5515
rect 42623 5481 42709 5499
rect 42521 5431 42587 5465
rect 41879 5363 41945 5397
rect 41879 5329 41895 5363
rect 41929 5329 41945 5363
rect 42521 5397 42553 5431
rect 42521 5363 42587 5397
rect 41879 5324 41945 5329
rect 42072 5329 42354 5362
rect 42072 5295 42162 5329
rect 42196 5327 42354 5329
rect 42196 5295 42281 5327
rect 42072 5293 42281 5295
rect 42315 5293 42354 5327
rect 42072 5287 42354 5293
rect 42521 5329 42553 5363
rect 42521 5287 42587 5329
rect 42693 5465 42709 5481
rect 42743 5465 42759 5499
rect 42693 5431 42759 5465
rect 42693 5397 42709 5431
rect 42743 5397 42759 5431
rect 42693 5363 42759 5397
rect 42693 5329 42709 5363
rect 42743 5329 42759 5363
rect 42693 5324 42759 5329
rect 43595 5499 43661 5515
rect 43595 5465 43627 5499
rect 43697 5499 43833 5515
rect 43697 5481 43783 5499
rect 43595 5431 43661 5465
rect 43595 5397 43627 5431
rect 43595 5363 43661 5397
rect 43595 5329 43627 5363
rect 43595 5287 43661 5329
rect 43767 5465 43783 5481
rect 43817 5465 43833 5499
rect 44052 5478 44086 5497
rect 44148 5667 44182 5686
rect 44148 5599 44182 5601
rect 44148 5563 44182 5565
rect 44148 5478 44182 5497
rect 44244 5667 44278 5686
rect 44244 5599 44278 5601
rect 44244 5563 44278 5565
rect 44244 5478 44278 5497
rect 43767 5431 43833 5465
rect 43767 5397 43783 5431
rect 43817 5397 43833 5431
rect 44084 5436 44150 5438
rect 44316 5436 44350 6050
rect 44401 5831 44435 6134
rect 44632 5831 44666 6042
rect 45570 6016 45604 6374
rect 45844 6351 45934 6374
rect 45968 6383 46292 6385
rect 45968 6351 46053 6383
rect 45844 6349 46053 6351
rect 46087 6374 46292 6383
rect 46344 6374 46378 6393
rect 46516 6571 46562 6691
rect 46616 6687 46662 6703
rect 46813 6773 46865 6811
rect 46813 6739 46831 6773
rect 46901 6803 46967 6845
rect 47142 6843 47171 6877
rect 47205 6843 47263 6877
rect 47297 6843 47355 6877
rect 47389 6843 47418 6877
rect 47578 6862 47626 6874
rect 47840 6866 47856 6900
rect 47890 6866 47906 6900
rect 48206 6890 48256 6960
rect 49696 6934 49730 6950
rect 49792 7056 49826 7072
rect 49888 7058 49922 7072
rect 50006 7058 50226 7080
rect 49886 7056 50226 7058
rect 49886 7022 49888 7056
rect 49922 7044 50226 7056
rect 49922 7022 50042 7044
rect 49792 6986 49826 7020
rect 49887 7020 49888 7022
rect 49887 6986 49922 7020
rect 50190 6996 50226 7044
rect 49887 6985 49888 6986
rect 49792 6934 49826 6950
rect 49888 6934 49922 6950
rect 50094 6960 50226 6996
rect 51584 7056 51618 7072
rect 51584 6986 51618 7020
rect 48206 6876 48216 6890
rect 46901 6769 46917 6803
rect 46951 6769 46967 6803
rect 47003 6790 47037 6811
rect 46813 6710 46865 6739
rect 47003 6735 47037 6756
rect 46596 6619 46612 6653
rect 46646 6642 46662 6653
rect 46596 6608 46614 6619
rect 46648 6608 46662 6642
rect 46813 6638 46849 6710
rect 46904 6701 47037 6735
rect 47208 6797 47274 6809
rect 47208 6763 47224 6797
rect 47258 6763 47274 6797
rect 47208 6746 47274 6763
rect 46904 6650 46938 6701
rect 47208 6695 47224 6746
rect 47258 6695 47274 6746
rect 47208 6683 47274 6695
rect 47308 6797 47354 6843
rect 47342 6763 47354 6797
rect 47308 6729 47354 6763
rect 47342 6695 47354 6729
rect 47578 6828 47584 6862
rect 47618 6828 47626 6862
rect 48210 6856 48216 6876
rect 48250 6856 48256 6890
rect 48210 6846 48256 6856
rect 48338 6851 48367 6885
rect 48401 6851 48459 6885
rect 48493 6851 48551 6885
rect 48585 6851 48614 6885
rect 47578 6740 47626 6828
rect 47952 6785 47968 6819
rect 48002 6818 48018 6819
rect 48002 6786 48164 6818
rect 48404 6810 48470 6817
rect 48398 6805 48470 6810
rect 48398 6786 48420 6805
rect 48002 6785 48420 6786
rect 47952 6782 48420 6785
rect 48128 6771 48420 6782
rect 48454 6771 48470 6805
rect 48128 6750 48470 6771
rect 47824 6740 47858 6742
rect 47578 6723 47858 6740
rect 47578 6706 47824 6723
rect 46596 6605 46662 6608
rect 46808 6636 46849 6638
rect 46808 6602 46810 6636
rect 46844 6602 46849 6636
rect 46808 6600 46849 6602
rect 46516 6553 46582 6571
rect 46516 6519 46532 6553
rect 46566 6519 46582 6553
rect 46516 6485 46582 6519
rect 46516 6451 46532 6485
rect 46566 6451 46582 6485
rect 46516 6417 46582 6451
rect 46516 6383 46532 6417
rect 46566 6383 46582 6417
rect 46516 6375 46582 6383
rect 46616 6553 46658 6569
rect 46650 6519 46658 6553
rect 46616 6485 46658 6519
rect 46650 6451 46658 6485
rect 46616 6417 46658 6451
rect 46650 6383 46658 6417
rect 46087 6349 46126 6374
rect 45638 6297 45654 6331
rect 45688 6297 45704 6331
rect 45844 6310 46126 6349
rect 46616 6341 46658 6383
rect 46813 6550 46849 6600
rect 46883 6634 46938 6650
rect 46917 6600 46938 6634
rect 46883 6584 46938 6600
rect 46983 6648 47051 6665
rect 46983 6647 47003 6648
rect 46983 6613 47001 6647
rect 47037 6614 47051 6648
rect 47035 6613 47051 6614
rect 46983 6591 47051 6613
rect 46904 6555 46938 6584
rect 47208 6563 47254 6683
rect 47308 6679 47354 6695
rect 47526 6658 47542 6659
rect 47288 6611 47304 6645
rect 47338 6638 47354 6645
rect 47406 6638 47542 6658
rect 47338 6625 47542 6638
rect 47576 6625 47592 6659
rect 47338 6624 47592 6625
rect 47338 6611 47446 6624
rect 47526 6622 47592 6624
rect 47824 6655 47858 6657
rect 47288 6597 47446 6611
rect 47302 6596 47446 6597
rect 47824 6619 47858 6621
rect 47498 6563 47532 6582
rect 46813 6500 46867 6550
rect 46904 6521 47039 6555
rect 46813 6466 46831 6500
rect 46865 6466 46867 6500
rect 47003 6487 47039 6521
rect 46813 6419 46867 6466
rect 46813 6385 46831 6419
rect 46865 6385 46867 6419
rect 46813 6369 46867 6385
rect 46901 6453 46917 6487
rect 46951 6453 46967 6487
rect 46901 6419 46967 6453
rect 46901 6385 46917 6419
rect 46951 6385 46967 6419
rect 46012 6308 46126 6310
rect 46284 6297 46300 6331
rect 46334 6297 46350 6331
rect 46450 6307 46479 6341
rect 46513 6307 46571 6341
rect 46605 6307 46663 6341
rect 46697 6307 46726 6341
rect 46901 6335 46967 6385
rect 47037 6453 47039 6487
rect 47003 6419 47039 6453
rect 47037 6385 47039 6419
rect 47003 6369 47039 6385
rect 47208 6545 47274 6563
rect 47208 6511 47224 6545
rect 47258 6511 47274 6545
rect 47208 6477 47274 6511
rect 47208 6443 47224 6477
rect 47258 6443 47274 6477
rect 47208 6409 47274 6443
rect 47208 6375 47224 6409
rect 47258 6375 47274 6409
rect 47208 6367 47274 6375
rect 47308 6545 47350 6561
rect 47342 6511 47350 6545
rect 47308 6477 47350 6511
rect 47342 6443 47350 6477
rect 47308 6409 47350 6443
rect 47498 6495 47532 6497
rect 47498 6459 47532 6461
rect 47342 6375 47350 6409
rect 46617 6300 46651 6307
rect 46796 6301 46825 6335
rect 46859 6301 46917 6335
rect 46951 6301 47009 6335
rect 47043 6301 47072 6335
rect 47308 6333 47350 6375
rect 47458 6393 47498 6414
rect 47586 6563 47620 6582
rect 47824 6534 47858 6553
rect 47920 6723 47954 6742
rect 47920 6655 47954 6657
rect 47920 6619 47954 6621
rect 47920 6534 47954 6553
rect 48016 6723 48050 6742
rect 48404 6737 48470 6750
rect 48404 6703 48420 6737
rect 48454 6703 48470 6737
rect 48404 6691 48470 6703
rect 48504 6805 48550 6851
rect 48684 6845 48713 6879
rect 48747 6845 48805 6879
rect 48839 6845 48897 6879
rect 48931 6845 48960 6879
rect 48538 6771 48550 6805
rect 48504 6737 48550 6771
rect 48538 6703 48550 6737
rect 48016 6655 48050 6657
rect 48172 6625 48188 6659
rect 48222 6625 48238 6659
rect 48016 6619 48050 6621
rect 48016 6534 48050 6553
rect 48144 6563 48178 6582
rect 47586 6495 47620 6497
rect 48144 6495 48178 6497
rect 47586 6459 47620 6461
rect 47856 6457 47872 6491
rect 47906 6457 47922 6491
rect 48144 6459 48178 6461
rect 47532 6393 47534 6414
rect 47458 6374 47534 6393
rect 47620 6393 48144 6418
rect 48232 6563 48266 6582
rect 48232 6495 48266 6497
rect 48232 6459 48266 6461
rect 48178 6393 48180 6418
rect 47586 6385 48180 6393
rect 47586 6374 47822 6385
rect 47142 6299 47171 6333
rect 47205 6299 47263 6333
rect 47297 6299 47355 6333
rect 47389 6299 47418 6333
rect 45704 6212 45750 6218
rect 45704 6210 46192 6212
rect 45704 6176 45712 6210
rect 45746 6193 46192 6210
rect 45746 6188 46142 6193
rect 45746 6178 46021 6188
rect 45746 6176 45750 6178
rect 45704 6174 45750 6176
rect 45922 6154 46021 6178
rect 46055 6159 46142 6188
rect 46176 6168 46192 6193
rect 46176 6159 46317 6168
rect 46055 6154 46317 6159
rect 45922 6134 46317 6154
rect 46046 6050 46062 6084
rect 46096 6050 46232 6084
rect 45570 6000 45952 6016
rect 45570 5976 45918 6000
rect 45918 5930 45952 5964
rect 45918 5878 45952 5894
rect 46014 6000 46048 6016
rect 46014 5930 46048 5964
rect 46014 5878 46048 5894
rect 46110 6000 46144 6016
rect 46110 5930 46144 5964
rect 46110 5878 46144 5894
rect 44390 5797 44419 5831
rect 44453 5797 44511 5831
rect 44545 5797 44603 5831
rect 44637 5797 44666 5831
rect 45458 5797 45487 5831
rect 45521 5797 45579 5831
rect 45613 5797 45671 5831
rect 45705 5797 45734 5831
rect 45950 5810 45966 5844
rect 46000 5810 46016 5844
rect 44409 5753 44463 5797
rect 44409 5719 44429 5753
rect 44409 5685 44463 5719
rect 44409 5651 44429 5685
rect 44409 5635 44463 5651
rect 44497 5753 44563 5763
rect 44497 5719 44513 5753
rect 44547 5719 44563 5753
rect 44497 5710 44563 5719
rect 44497 5685 44515 5710
rect 44497 5651 44513 5685
rect 44549 5676 44563 5710
rect 44547 5651 44563 5676
rect 44497 5635 44563 5651
rect 44597 5753 44645 5797
rect 44631 5719 44645 5753
rect 44597 5685 44645 5719
rect 44631 5651 44645 5685
rect 44597 5635 44645 5651
rect 45477 5753 45531 5797
rect 45477 5719 45497 5753
rect 45477 5685 45531 5719
rect 45477 5651 45497 5685
rect 45477 5635 45531 5651
rect 45565 5753 45631 5763
rect 45565 5719 45581 5753
rect 45615 5719 45631 5753
rect 45565 5715 45631 5719
rect 45565 5681 45579 5715
rect 45613 5685 45631 5715
rect 45565 5651 45581 5681
rect 45615 5651 45631 5685
rect 45565 5635 45631 5651
rect 45665 5753 45713 5797
rect 45699 5719 45713 5753
rect 46062 5729 46078 5763
rect 46112 5729 46128 5763
rect 45665 5685 45713 5719
rect 45699 5651 45713 5685
rect 45665 5635 45713 5651
rect 45934 5667 45968 5686
rect 44407 5594 44427 5599
rect 44407 5560 44424 5594
rect 44461 5565 44477 5599
rect 44458 5560 44477 5565
rect 44407 5549 44477 5560
rect 44511 5515 44545 5635
rect 44579 5565 44595 5599
rect 44629 5590 44649 5599
rect 44579 5556 44597 5565
rect 44631 5556 44649 5590
rect 44579 5549 44649 5556
rect 45475 5592 45495 5599
rect 45475 5558 45493 5592
rect 45529 5565 45545 5599
rect 45527 5558 45545 5565
rect 45475 5549 45545 5558
rect 45579 5515 45613 5635
rect 45934 5599 45968 5601
rect 45647 5565 45663 5599
rect 45697 5592 45717 5599
rect 45647 5558 45667 5565
rect 45701 5558 45717 5592
rect 45647 5549 45717 5558
rect 45934 5563 45968 5565
rect 44084 5435 44350 5436
rect 44084 5401 44100 5435
rect 44134 5401 44350 5435
rect 44084 5400 44350 5401
rect 44409 5499 44475 5515
rect 44409 5465 44441 5499
rect 44511 5499 44647 5515
rect 44511 5481 44597 5499
rect 44409 5431 44475 5465
rect 43767 5363 43833 5397
rect 43767 5329 43783 5363
rect 43817 5329 43833 5363
rect 44409 5397 44441 5431
rect 44409 5363 44475 5397
rect 43767 5324 43833 5329
rect 43960 5329 44242 5362
rect 43960 5295 44050 5329
rect 44084 5327 44242 5329
rect 44084 5295 44169 5327
rect 43960 5293 44169 5295
rect 44203 5293 44242 5327
rect 43960 5287 44242 5293
rect 44409 5329 44441 5363
rect 44409 5287 44475 5329
rect 44581 5465 44597 5481
rect 44631 5465 44647 5499
rect 44581 5431 44647 5465
rect 44581 5397 44597 5431
rect 44631 5397 44647 5431
rect 44581 5363 44647 5397
rect 44581 5329 44597 5363
rect 44631 5329 44647 5363
rect 44581 5324 44647 5329
rect 45477 5499 45543 5515
rect 45477 5465 45509 5499
rect 45579 5499 45715 5515
rect 45579 5481 45665 5499
rect 45477 5431 45543 5465
rect 45477 5397 45509 5431
rect 45477 5363 45543 5397
rect 45477 5329 45509 5363
rect 45477 5287 45543 5329
rect 45649 5465 45665 5481
rect 45699 5465 45715 5499
rect 45934 5478 45968 5497
rect 46030 5667 46064 5686
rect 46030 5599 46064 5601
rect 46030 5563 46064 5565
rect 46030 5478 46064 5497
rect 46126 5667 46160 5686
rect 46126 5599 46160 5601
rect 46126 5563 46160 5565
rect 46126 5478 46160 5497
rect 45649 5431 45715 5465
rect 45649 5397 45665 5431
rect 45699 5397 45715 5431
rect 45966 5436 46032 5438
rect 46198 5436 46232 6050
rect 46283 5831 46317 6134
rect 46514 5831 46548 6042
rect 47458 6016 47492 6374
rect 47732 6351 47822 6374
rect 47856 6383 48180 6385
rect 47856 6351 47941 6383
rect 47732 6349 47941 6351
rect 47975 6374 48180 6383
rect 48232 6374 48266 6393
rect 48404 6571 48450 6691
rect 48504 6687 48550 6703
rect 48701 6773 48753 6811
rect 48701 6739 48719 6773
rect 48789 6803 48855 6845
rect 49030 6843 49059 6877
rect 49093 6843 49151 6877
rect 49185 6843 49243 6877
rect 49277 6843 49306 6877
rect 49466 6862 49514 6874
rect 49728 6866 49744 6900
rect 49778 6866 49794 6900
rect 50094 6890 50144 6960
rect 51584 6934 51618 6950
rect 51680 7056 51714 7072
rect 51776 7058 51810 7072
rect 51894 7058 52114 7080
rect 51774 7056 52114 7058
rect 51774 7022 51776 7056
rect 51810 7044 52114 7056
rect 51810 7022 51930 7044
rect 51680 6986 51714 7020
rect 51775 7020 51776 7022
rect 51775 6986 51810 7020
rect 52078 6996 52114 7044
rect 51775 6985 51776 6986
rect 51680 6934 51714 6950
rect 51776 6934 51810 6950
rect 51982 6960 52114 6996
rect 53472 7056 53506 7072
rect 53472 6986 53506 7020
rect 50094 6876 50104 6890
rect 48789 6769 48805 6803
rect 48839 6769 48855 6803
rect 48891 6790 48925 6811
rect 48701 6710 48753 6739
rect 48891 6735 48925 6756
rect 48484 6619 48500 6653
rect 48534 6642 48550 6653
rect 48484 6608 48502 6619
rect 48536 6608 48550 6642
rect 48701 6638 48737 6710
rect 48792 6701 48925 6735
rect 49096 6797 49162 6809
rect 49096 6763 49112 6797
rect 49146 6763 49162 6797
rect 49096 6746 49162 6763
rect 48792 6650 48826 6701
rect 49096 6695 49112 6746
rect 49146 6695 49162 6746
rect 49096 6683 49162 6695
rect 49196 6797 49242 6843
rect 49230 6763 49242 6797
rect 49196 6729 49242 6763
rect 49230 6695 49242 6729
rect 49466 6828 49472 6862
rect 49506 6828 49514 6862
rect 50098 6856 50104 6876
rect 50138 6856 50144 6890
rect 50098 6846 50144 6856
rect 50226 6851 50255 6885
rect 50289 6851 50347 6885
rect 50381 6851 50439 6885
rect 50473 6851 50502 6885
rect 49466 6740 49514 6828
rect 49840 6785 49856 6819
rect 49890 6818 49906 6819
rect 49890 6786 50052 6818
rect 50292 6810 50358 6817
rect 50286 6805 50358 6810
rect 50286 6786 50308 6805
rect 49890 6785 50308 6786
rect 49840 6782 50308 6785
rect 50016 6771 50308 6782
rect 50342 6771 50358 6805
rect 50016 6750 50358 6771
rect 49712 6740 49746 6742
rect 49466 6723 49746 6740
rect 49466 6706 49712 6723
rect 48484 6605 48550 6608
rect 48696 6636 48737 6638
rect 48696 6602 48698 6636
rect 48732 6602 48737 6636
rect 48696 6600 48737 6602
rect 48404 6553 48470 6571
rect 48404 6519 48420 6553
rect 48454 6519 48470 6553
rect 48404 6485 48470 6519
rect 48404 6451 48420 6485
rect 48454 6451 48470 6485
rect 48404 6417 48470 6451
rect 48404 6383 48420 6417
rect 48454 6383 48470 6417
rect 48404 6375 48470 6383
rect 48504 6553 48546 6569
rect 48538 6519 48546 6553
rect 48504 6485 48546 6519
rect 48538 6451 48546 6485
rect 48504 6417 48546 6451
rect 48538 6383 48546 6417
rect 47975 6349 48014 6374
rect 47526 6297 47542 6331
rect 47576 6297 47592 6331
rect 47732 6310 48014 6349
rect 48504 6341 48546 6383
rect 48701 6550 48737 6600
rect 48771 6634 48826 6650
rect 48805 6600 48826 6634
rect 48771 6584 48826 6600
rect 48871 6648 48939 6665
rect 48871 6647 48891 6648
rect 48871 6613 48889 6647
rect 48925 6614 48939 6648
rect 48923 6613 48939 6614
rect 48871 6591 48939 6613
rect 48792 6555 48826 6584
rect 49096 6563 49142 6683
rect 49196 6679 49242 6695
rect 49414 6658 49430 6659
rect 49176 6611 49192 6645
rect 49226 6638 49242 6645
rect 49294 6638 49430 6658
rect 49226 6625 49430 6638
rect 49464 6625 49480 6659
rect 49226 6624 49480 6625
rect 49226 6611 49334 6624
rect 49414 6622 49480 6624
rect 49712 6655 49746 6657
rect 49176 6597 49334 6611
rect 49190 6596 49334 6597
rect 49712 6619 49746 6621
rect 49386 6563 49420 6582
rect 48701 6500 48755 6550
rect 48792 6521 48927 6555
rect 48701 6466 48719 6500
rect 48753 6466 48755 6500
rect 48891 6487 48927 6521
rect 48701 6419 48755 6466
rect 48701 6385 48719 6419
rect 48753 6385 48755 6419
rect 48701 6369 48755 6385
rect 48789 6453 48805 6487
rect 48839 6453 48855 6487
rect 48789 6419 48855 6453
rect 48789 6385 48805 6419
rect 48839 6385 48855 6419
rect 47900 6308 48014 6310
rect 48172 6297 48188 6331
rect 48222 6297 48238 6331
rect 48338 6307 48367 6341
rect 48401 6307 48459 6341
rect 48493 6307 48551 6341
rect 48585 6307 48614 6341
rect 48789 6335 48855 6385
rect 48925 6453 48927 6487
rect 48891 6419 48927 6453
rect 48925 6385 48927 6419
rect 48891 6369 48927 6385
rect 49096 6545 49162 6563
rect 49096 6511 49112 6545
rect 49146 6511 49162 6545
rect 49096 6477 49162 6511
rect 49096 6443 49112 6477
rect 49146 6443 49162 6477
rect 49096 6409 49162 6443
rect 49096 6375 49112 6409
rect 49146 6375 49162 6409
rect 49096 6367 49162 6375
rect 49196 6545 49238 6561
rect 49230 6511 49238 6545
rect 49196 6477 49238 6511
rect 49230 6443 49238 6477
rect 49196 6409 49238 6443
rect 49386 6495 49420 6497
rect 49386 6459 49420 6461
rect 49230 6375 49238 6409
rect 48505 6300 48539 6307
rect 48684 6301 48713 6335
rect 48747 6301 48805 6335
rect 48839 6301 48897 6335
rect 48931 6301 48960 6335
rect 49196 6333 49238 6375
rect 49346 6393 49386 6414
rect 49474 6563 49508 6582
rect 49712 6534 49746 6553
rect 49808 6723 49842 6742
rect 49808 6655 49842 6657
rect 49808 6619 49842 6621
rect 49808 6534 49842 6553
rect 49904 6723 49938 6742
rect 50292 6737 50358 6750
rect 50292 6703 50308 6737
rect 50342 6703 50358 6737
rect 50292 6691 50358 6703
rect 50392 6805 50438 6851
rect 50572 6845 50601 6879
rect 50635 6845 50693 6879
rect 50727 6845 50785 6879
rect 50819 6845 50848 6879
rect 50426 6771 50438 6805
rect 50392 6737 50438 6771
rect 50426 6703 50438 6737
rect 49904 6655 49938 6657
rect 50060 6625 50076 6659
rect 50110 6625 50126 6659
rect 49904 6619 49938 6621
rect 49904 6534 49938 6553
rect 50032 6563 50066 6582
rect 49474 6495 49508 6497
rect 50032 6495 50066 6497
rect 49474 6459 49508 6461
rect 49744 6457 49760 6491
rect 49794 6457 49810 6491
rect 50032 6459 50066 6461
rect 49420 6393 49422 6414
rect 49346 6374 49422 6393
rect 49508 6393 50032 6418
rect 50120 6563 50154 6582
rect 50120 6495 50154 6497
rect 50120 6459 50154 6461
rect 50066 6393 50068 6418
rect 49474 6385 50068 6393
rect 49474 6374 49710 6385
rect 49030 6299 49059 6333
rect 49093 6299 49151 6333
rect 49185 6299 49243 6333
rect 49277 6299 49306 6333
rect 47592 6212 47638 6218
rect 47592 6210 48080 6212
rect 47592 6176 47600 6210
rect 47634 6193 48080 6210
rect 47634 6188 48030 6193
rect 47634 6178 47909 6188
rect 47634 6176 47638 6178
rect 47592 6174 47638 6176
rect 47810 6154 47909 6178
rect 47943 6159 48030 6188
rect 48064 6168 48080 6193
rect 48064 6159 48205 6168
rect 47943 6154 48205 6159
rect 47810 6134 48205 6154
rect 47934 6050 47950 6084
rect 47984 6050 48120 6084
rect 47458 6000 47840 6016
rect 47458 5976 47806 6000
rect 47806 5930 47840 5964
rect 47806 5878 47840 5894
rect 47902 6000 47936 6016
rect 47902 5930 47936 5964
rect 47902 5878 47936 5894
rect 47998 6000 48032 6016
rect 47998 5930 48032 5964
rect 47998 5878 48032 5894
rect 46272 5797 46301 5831
rect 46335 5797 46393 5831
rect 46427 5797 46485 5831
rect 46519 5797 46548 5831
rect 47346 5797 47375 5831
rect 47409 5797 47467 5831
rect 47501 5797 47559 5831
rect 47593 5797 47622 5831
rect 47838 5810 47854 5844
rect 47888 5810 47904 5844
rect 46291 5753 46345 5797
rect 46291 5719 46311 5753
rect 46291 5685 46345 5719
rect 46291 5651 46311 5685
rect 46291 5635 46345 5651
rect 46379 5753 46445 5763
rect 46379 5719 46395 5753
rect 46429 5719 46445 5753
rect 46379 5710 46445 5719
rect 46379 5685 46397 5710
rect 46379 5651 46395 5685
rect 46431 5676 46445 5710
rect 46429 5651 46445 5676
rect 46379 5635 46445 5651
rect 46479 5753 46527 5797
rect 46513 5719 46527 5753
rect 46479 5685 46527 5719
rect 46513 5651 46527 5685
rect 46479 5635 46527 5651
rect 47365 5753 47419 5797
rect 47365 5719 47385 5753
rect 47365 5685 47419 5719
rect 47365 5651 47385 5685
rect 47365 5635 47419 5651
rect 47453 5753 47519 5763
rect 47453 5719 47469 5753
rect 47503 5719 47519 5753
rect 47453 5715 47519 5719
rect 47453 5681 47467 5715
rect 47501 5685 47519 5715
rect 47453 5651 47469 5681
rect 47503 5651 47519 5685
rect 47453 5635 47519 5651
rect 47553 5753 47601 5797
rect 47587 5719 47601 5753
rect 47950 5729 47966 5763
rect 48000 5729 48016 5763
rect 47553 5685 47601 5719
rect 47587 5651 47601 5685
rect 47553 5635 47601 5651
rect 47822 5667 47856 5686
rect 46289 5594 46309 5599
rect 46289 5560 46306 5594
rect 46343 5565 46359 5599
rect 46340 5560 46359 5565
rect 46289 5549 46359 5560
rect 46393 5515 46427 5635
rect 46461 5565 46477 5599
rect 46511 5590 46531 5599
rect 46461 5556 46479 5565
rect 46513 5556 46531 5590
rect 46461 5549 46531 5556
rect 47363 5592 47383 5599
rect 47363 5558 47381 5592
rect 47417 5565 47433 5599
rect 47415 5558 47433 5565
rect 47363 5549 47433 5558
rect 47467 5515 47501 5635
rect 47822 5599 47856 5601
rect 47535 5565 47551 5599
rect 47585 5592 47605 5599
rect 47535 5558 47555 5565
rect 47589 5558 47605 5592
rect 47535 5549 47605 5558
rect 47822 5563 47856 5565
rect 45966 5435 46232 5436
rect 45966 5401 45982 5435
rect 46016 5401 46232 5435
rect 45966 5400 46232 5401
rect 46291 5499 46357 5515
rect 46291 5465 46323 5499
rect 46393 5499 46529 5515
rect 46393 5481 46479 5499
rect 46291 5431 46357 5465
rect 45649 5363 45715 5397
rect 45649 5329 45665 5363
rect 45699 5329 45715 5363
rect 46291 5397 46323 5431
rect 46291 5363 46357 5397
rect 45649 5324 45715 5329
rect 45842 5329 46124 5362
rect 45842 5295 45932 5329
rect 45966 5327 46124 5329
rect 45966 5295 46051 5327
rect 45842 5293 46051 5295
rect 46085 5293 46124 5327
rect 45842 5287 46124 5293
rect 46291 5329 46323 5363
rect 46291 5287 46357 5329
rect 46463 5465 46479 5481
rect 46513 5465 46529 5499
rect 46463 5431 46529 5465
rect 46463 5397 46479 5431
rect 46513 5397 46529 5431
rect 46463 5363 46529 5397
rect 46463 5329 46479 5363
rect 46513 5329 46529 5363
rect 46463 5324 46529 5329
rect 47365 5499 47431 5515
rect 47365 5465 47397 5499
rect 47467 5499 47603 5515
rect 47467 5481 47553 5499
rect 47365 5431 47431 5465
rect 47365 5397 47397 5431
rect 47365 5363 47431 5397
rect 47365 5329 47397 5363
rect 47365 5287 47431 5329
rect 47537 5465 47553 5481
rect 47587 5465 47603 5499
rect 47822 5478 47856 5497
rect 47918 5667 47952 5686
rect 47918 5599 47952 5601
rect 47918 5563 47952 5565
rect 47918 5478 47952 5497
rect 48014 5667 48048 5686
rect 48014 5599 48048 5601
rect 48014 5563 48048 5565
rect 48014 5478 48048 5497
rect 47537 5431 47603 5465
rect 47537 5397 47553 5431
rect 47587 5397 47603 5431
rect 47854 5436 47920 5438
rect 48086 5436 48120 6050
rect 48171 5831 48205 6134
rect 48402 5831 48436 6042
rect 49346 6016 49380 6374
rect 49620 6351 49710 6374
rect 49744 6383 50068 6385
rect 49744 6351 49829 6383
rect 49620 6349 49829 6351
rect 49863 6374 50068 6383
rect 50120 6374 50154 6393
rect 50292 6571 50338 6691
rect 50392 6687 50438 6703
rect 50589 6773 50641 6811
rect 50589 6739 50607 6773
rect 50677 6803 50743 6845
rect 50918 6843 50947 6877
rect 50981 6843 51039 6877
rect 51073 6843 51131 6877
rect 51165 6843 51194 6877
rect 51354 6862 51402 6874
rect 51616 6866 51632 6900
rect 51666 6866 51682 6900
rect 51982 6890 52032 6960
rect 53472 6934 53506 6950
rect 53568 7056 53602 7072
rect 53664 7058 53698 7072
rect 53782 7058 54002 7080
rect 53662 7056 54002 7058
rect 53662 7022 53664 7056
rect 53698 7044 54002 7056
rect 53698 7022 53818 7044
rect 53568 6986 53602 7020
rect 53663 7020 53664 7022
rect 53663 6986 53698 7020
rect 53966 6996 54002 7044
rect 53663 6985 53664 6986
rect 53568 6934 53602 6950
rect 53664 6934 53698 6950
rect 53870 6960 54002 6996
rect 55360 7056 55394 7072
rect 55360 6986 55394 7020
rect 51982 6876 51992 6890
rect 50677 6769 50693 6803
rect 50727 6769 50743 6803
rect 50779 6790 50813 6811
rect 50589 6710 50641 6739
rect 50779 6735 50813 6756
rect 50372 6619 50388 6653
rect 50422 6642 50438 6653
rect 50372 6608 50390 6619
rect 50424 6608 50438 6642
rect 50589 6638 50625 6710
rect 50680 6701 50813 6735
rect 50984 6797 51050 6809
rect 50984 6763 51000 6797
rect 51034 6763 51050 6797
rect 50984 6746 51050 6763
rect 50680 6650 50714 6701
rect 50984 6695 51000 6746
rect 51034 6695 51050 6746
rect 50984 6683 51050 6695
rect 51084 6797 51130 6843
rect 51118 6763 51130 6797
rect 51084 6729 51130 6763
rect 51118 6695 51130 6729
rect 51354 6828 51360 6862
rect 51394 6828 51402 6862
rect 51986 6856 51992 6876
rect 52026 6856 52032 6890
rect 51986 6846 52032 6856
rect 52114 6851 52143 6885
rect 52177 6851 52235 6885
rect 52269 6851 52327 6885
rect 52361 6851 52390 6885
rect 51354 6740 51402 6828
rect 51728 6785 51744 6819
rect 51778 6818 51794 6819
rect 51778 6786 51940 6818
rect 52180 6810 52246 6817
rect 52174 6805 52246 6810
rect 52174 6786 52196 6805
rect 51778 6785 52196 6786
rect 51728 6782 52196 6785
rect 51904 6771 52196 6782
rect 52230 6771 52246 6805
rect 51904 6750 52246 6771
rect 51600 6740 51634 6742
rect 51354 6723 51634 6740
rect 51354 6706 51600 6723
rect 50372 6605 50438 6608
rect 50584 6636 50625 6638
rect 50584 6602 50586 6636
rect 50620 6602 50625 6636
rect 50584 6600 50625 6602
rect 50292 6553 50358 6571
rect 50292 6519 50308 6553
rect 50342 6519 50358 6553
rect 50292 6485 50358 6519
rect 50292 6451 50308 6485
rect 50342 6451 50358 6485
rect 50292 6417 50358 6451
rect 50292 6383 50308 6417
rect 50342 6383 50358 6417
rect 50292 6375 50358 6383
rect 50392 6553 50434 6569
rect 50426 6519 50434 6553
rect 50392 6485 50434 6519
rect 50426 6451 50434 6485
rect 50392 6417 50434 6451
rect 50426 6383 50434 6417
rect 49863 6349 49902 6374
rect 49414 6297 49430 6331
rect 49464 6297 49480 6331
rect 49620 6310 49902 6349
rect 50392 6341 50434 6383
rect 50589 6550 50625 6600
rect 50659 6634 50714 6650
rect 50693 6600 50714 6634
rect 50659 6584 50714 6600
rect 50759 6648 50827 6665
rect 50759 6647 50779 6648
rect 50759 6613 50777 6647
rect 50813 6614 50827 6648
rect 50811 6613 50827 6614
rect 50759 6591 50827 6613
rect 50680 6555 50714 6584
rect 50984 6563 51030 6683
rect 51084 6679 51130 6695
rect 51302 6658 51318 6659
rect 51064 6611 51080 6645
rect 51114 6638 51130 6645
rect 51182 6638 51318 6658
rect 51114 6625 51318 6638
rect 51352 6625 51368 6659
rect 51114 6624 51368 6625
rect 51114 6611 51222 6624
rect 51302 6622 51368 6624
rect 51600 6655 51634 6657
rect 51064 6597 51222 6611
rect 51078 6596 51222 6597
rect 51600 6619 51634 6621
rect 51274 6563 51308 6582
rect 50589 6500 50643 6550
rect 50680 6521 50815 6555
rect 50589 6466 50607 6500
rect 50641 6466 50643 6500
rect 50779 6487 50815 6521
rect 50589 6419 50643 6466
rect 50589 6385 50607 6419
rect 50641 6385 50643 6419
rect 50589 6369 50643 6385
rect 50677 6453 50693 6487
rect 50727 6453 50743 6487
rect 50677 6419 50743 6453
rect 50677 6385 50693 6419
rect 50727 6385 50743 6419
rect 49788 6308 49902 6310
rect 50060 6297 50076 6331
rect 50110 6297 50126 6331
rect 50226 6307 50255 6341
rect 50289 6307 50347 6341
rect 50381 6307 50439 6341
rect 50473 6307 50502 6341
rect 50677 6335 50743 6385
rect 50813 6453 50815 6487
rect 50779 6419 50815 6453
rect 50813 6385 50815 6419
rect 50779 6369 50815 6385
rect 50984 6545 51050 6563
rect 50984 6511 51000 6545
rect 51034 6511 51050 6545
rect 50984 6477 51050 6511
rect 50984 6443 51000 6477
rect 51034 6443 51050 6477
rect 50984 6409 51050 6443
rect 50984 6375 51000 6409
rect 51034 6375 51050 6409
rect 50984 6367 51050 6375
rect 51084 6545 51126 6561
rect 51118 6511 51126 6545
rect 51084 6477 51126 6511
rect 51118 6443 51126 6477
rect 51084 6409 51126 6443
rect 51274 6495 51308 6497
rect 51274 6459 51308 6461
rect 51118 6375 51126 6409
rect 50393 6300 50427 6307
rect 50572 6301 50601 6335
rect 50635 6301 50693 6335
rect 50727 6301 50785 6335
rect 50819 6301 50848 6335
rect 51084 6333 51126 6375
rect 51234 6393 51274 6414
rect 51362 6563 51396 6582
rect 51600 6534 51634 6553
rect 51696 6723 51730 6742
rect 51696 6655 51730 6657
rect 51696 6619 51730 6621
rect 51696 6534 51730 6553
rect 51792 6723 51826 6742
rect 52180 6737 52246 6750
rect 52180 6703 52196 6737
rect 52230 6703 52246 6737
rect 52180 6691 52246 6703
rect 52280 6805 52326 6851
rect 52460 6845 52489 6879
rect 52523 6845 52581 6879
rect 52615 6845 52673 6879
rect 52707 6845 52736 6879
rect 52314 6771 52326 6805
rect 52280 6737 52326 6771
rect 52314 6703 52326 6737
rect 51792 6655 51826 6657
rect 51948 6625 51964 6659
rect 51998 6625 52014 6659
rect 51792 6619 51826 6621
rect 51792 6534 51826 6553
rect 51920 6563 51954 6582
rect 51362 6495 51396 6497
rect 51920 6495 51954 6497
rect 51362 6459 51396 6461
rect 51632 6457 51648 6491
rect 51682 6457 51698 6491
rect 51920 6459 51954 6461
rect 51308 6393 51310 6414
rect 51234 6374 51310 6393
rect 51396 6393 51920 6418
rect 52008 6563 52042 6582
rect 52008 6495 52042 6497
rect 52008 6459 52042 6461
rect 51954 6393 51956 6418
rect 51362 6385 51956 6393
rect 51362 6374 51598 6385
rect 50918 6299 50947 6333
rect 50981 6299 51039 6333
rect 51073 6299 51131 6333
rect 51165 6299 51194 6333
rect 49480 6212 49526 6218
rect 49480 6210 49968 6212
rect 49480 6176 49488 6210
rect 49522 6193 49968 6210
rect 49522 6188 49918 6193
rect 49522 6178 49797 6188
rect 49522 6176 49526 6178
rect 49480 6174 49526 6176
rect 49698 6154 49797 6178
rect 49831 6159 49918 6188
rect 49952 6168 49968 6193
rect 49952 6159 50093 6168
rect 49831 6154 50093 6159
rect 49698 6134 50093 6154
rect 49822 6050 49838 6084
rect 49872 6050 50008 6084
rect 49346 6000 49728 6016
rect 49346 5976 49694 6000
rect 49694 5930 49728 5964
rect 49694 5878 49728 5894
rect 49790 6000 49824 6016
rect 49790 5930 49824 5964
rect 49790 5878 49824 5894
rect 49886 6000 49920 6016
rect 49886 5930 49920 5964
rect 49886 5878 49920 5894
rect 48160 5797 48189 5831
rect 48223 5797 48281 5831
rect 48315 5797 48373 5831
rect 48407 5797 48436 5831
rect 49234 5797 49263 5831
rect 49297 5797 49355 5831
rect 49389 5797 49447 5831
rect 49481 5797 49510 5831
rect 49726 5810 49742 5844
rect 49776 5810 49792 5844
rect 48179 5753 48233 5797
rect 48179 5719 48199 5753
rect 48179 5685 48233 5719
rect 48179 5651 48199 5685
rect 48179 5635 48233 5651
rect 48267 5753 48333 5763
rect 48267 5719 48283 5753
rect 48317 5719 48333 5753
rect 48267 5710 48333 5719
rect 48267 5685 48285 5710
rect 48267 5651 48283 5685
rect 48319 5676 48333 5710
rect 48317 5651 48333 5676
rect 48267 5635 48333 5651
rect 48367 5753 48415 5797
rect 48401 5719 48415 5753
rect 48367 5685 48415 5719
rect 48401 5651 48415 5685
rect 48367 5635 48415 5651
rect 49253 5753 49307 5797
rect 49253 5719 49273 5753
rect 49253 5685 49307 5719
rect 49253 5651 49273 5685
rect 49253 5635 49307 5651
rect 49341 5753 49407 5763
rect 49341 5719 49357 5753
rect 49391 5719 49407 5753
rect 49341 5715 49407 5719
rect 49341 5681 49355 5715
rect 49389 5685 49407 5715
rect 49341 5651 49357 5681
rect 49391 5651 49407 5685
rect 49341 5635 49407 5651
rect 49441 5753 49489 5797
rect 49475 5719 49489 5753
rect 49838 5729 49854 5763
rect 49888 5729 49904 5763
rect 49441 5685 49489 5719
rect 49475 5651 49489 5685
rect 49441 5635 49489 5651
rect 49710 5667 49744 5686
rect 48177 5594 48197 5599
rect 48177 5560 48194 5594
rect 48231 5565 48247 5599
rect 48228 5560 48247 5565
rect 48177 5549 48247 5560
rect 48281 5515 48315 5635
rect 48349 5565 48365 5599
rect 48399 5590 48419 5599
rect 48349 5556 48367 5565
rect 48401 5556 48419 5590
rect 48349 5549 48419 5556
rect 49251 5592 49271 5599
rect 49251 5558 49269 5592
rect 49305 5565 49321 5599
rect 49303 5558 49321 5565
rect 49251 5549 49321 5558
rect 49355 5515 49389 5635
rect 49710 5599 49744 5601
rect 49423 5565 49439 5599
rect 49473 5592 49493 5599
rect 49423 5558 49443 5565
rect 49477 5558 49493 5592
rect 49423 5549 49493 5558
rect 49710 5563 49744 5565
rect 47854 5435 48120 5436
rect 47854 5401 47870 5435
rect 47904 5401 48120 5435
rect 47854 5400 48120 5401
rect 48179 5499 48245 5515
rect 48179 5465 48211 5499
rect 48281 5499 48417 5515
rect 48281 5481 48367 5499
rect 48179 5431 48245 5465
rect 47537 5363 47603 5397
rect 47537 5329 47553 5363
rect 47587 5329 47603 5363
rect 48179 5397 48211 5431
rect 48179 5363 48245 5397
rect 47537 5324 47603 5329
rect 47730 5329 48012 5362
rect 47730 5295 47820 5329
rect 47854 5327 48012 5329
rect 47854 5295 47939 5327
rect 47730 5293 47939 5295
rect 47973 5293 48012 5327
rect 47730 5287 48012 5293
rect 48179 5329 48211 5363
rect 48179 5287 48245 5329
rect 48351 5465 48367 5481
rect 48401 5465 48417 5499
rect 48351 5431 48417 5465
rect 48351 5397 48367 5431
rect 48401 5397 48417 5431
rect 48351 5363 48417 5397
rect 48351 5329 48367 5363
rect 48401 5329 48417 5363
rect 48351 5324 48417 5329
rect 49253 5499 49319 5515
rect 49253 5465 49285 5499
rect 49355 5499 49491 5515
rect 49355 5481 49441 5499
rect 49253 5431 49319 5465
rect 49253 5397 49285 5431
rect 49253 5363 49319 5397
rect 49253 5329 49285 5363
rect 49253 5287 49319 5329
rect 49425 5465 49441 5481
rect 49475 5465 49491 5499
rect 49710 5478 49744 5497
rect 49806 5667 49840 5686
rect 49806 5599 49840 5601
rect 49806 5563 49840 5565
rect 49806 5478 49840 5497
rect 49902 5667 49936 5686
rect 49902 5599 49936 5601
rect 49902 5563 49936 5565
rect 49902 5478 49936 5497
rect 49425 5431 49491 5465
rect 49425 5397 49441 5431
rect 49475 5397 49491 5431
rect 49742 5436 49808 5438
rect 49974 5436 50008 6050
rect 50059 5831 50093 6134
rect 50290 5831 50324 6042
rect 51234 6016 51268 6374
rect 51508 6351 51598 6374
rect 51632 6383 51956 6385
rect 51632 6351 51717 6383
rect 51508 6349 51717 6351
rect 51751 6374 51956 6383
rect 52008 6374 52042 6393
rect 52180 6571 52226 6691
rect 52280 6687 52326 6703
rect 52477 6773 52529 6811
rect 52477 6739 52495 6773
rect 52565 6803 52631 6845
rect 52806 6843 52835 6877
rect 52869 6843 52927 6877
rect 52961 6843 53019 6877
rect 53053 6843 53082 6877
rect 53242 6862 53290 6874
rect 53504 6866 53520 6900
rect 53554 6866 53570 6900
rect 53870 6890 53920 6960
rect 55360 6934 55394 6950
rect 55456 7056 55490 7072
rect 55552 7058 55586 7072
rect 55670 7058 55890 7080
rect 55550 7056 55890 7058
rect 55550 7022 55552 7056
rect 55586 7044 55890 7056
rect 55586 7022 55706 7044
rect 55456 6986 55490 7020
rect 55551 7020 55552 7022
rect 55551 6986 55586 7020
rect 55854 6996 55890 7044
rect 55551 6985 55552 6986
rect 55456 6934 55490 6950
rect 55552 6934 55586 6950
rect 55758 6960 55890 6996
rect 57248 7056 57282 7072
rect 57248 6986 57282 7020
rect 53870 6876 53880 6890
rect 52565 6769 52581 6803
rect 52615 6769 52631 6803
rect 52667 6790 52701 6811
rect 52477 6710 52529 6739
rect 52667 6735 52701 6756
rect 52260 6619 52276 6653
rect 52310 6642 52326 6653
rect 52260 6608 52278 6619
rect 52312 6608 52326 6642
rect 52477 6638 52513 6710
rect 52568 6701 52701 6735
rect 52872 6797 52938 6809
rect 52872 6763 52888 6797
rect 52922 6763 52938 6797
rect 52872 6746 52938 6763
rect 52568 6650 52602 6701
rect 52872 6695 52888 6746
rect 52922 6695 52938 6746
rect 52872 6683 52938 6695
rect 52972 6797 53018 6843
rect 53006 6763 53018 6797
rect 52972 6729 53018 6763
rect 53006 6695 53018 6729
rect 53242 6828 53248 6862
rect 53282 6828 53290 6862
rect 53874 6856 53880 6876
rect 53914 6856 53920 6890
rect 53874 6846 53920 6856
rect 54002 6851 54031 6885
rect 54065 6851 54123 6885
rect 54157 6851 54215 6885
rect 54249 6851 54278 6885
rect 53242 6740 53290 6828
rect 53616 6785 53632 6819
rect 53666 6818 53682 6819
rect 53666 6786 53828 6818
rect 54068 6810 54134 6817
rect 54062 6805 54134 6810
rect 54062 6786 54084 6805
rect 53666 6785 54084 6786
rect 53616 6782 54084 6785
rect 53792 6771 54084 6782
rect 54118 6771 54134 6805
rect 53792 6750 54134 6771
rect 53488 6740 53522 6742
rect 53242 6723 53522 6740
rect 53242 6706 53488 6723
rect 52260 6605 52326 6608
rect 52472 6636 52513 6638
rect 52472 6602 52474 6636
rect 52508 6602 52513 6636
rect 52472 6600 52513 6602
rect 52180 6553 52246 6571
rect 52180 6519 52196 6553
rect 52230 6519 52246 6553
rect 52180 6485 52246 6519
rect 52180 6451 52196 6485
rect 52230 6451 52246 6485
rect 52180 6417 52246 6451
rect 52180 6383 52196 6417
rect 52230 6383 52246 6417
rect 52180 6375 52246 6383
rect 52280 6553 52322 6569
rect 52314 6519 52322 6553
rect 52280 6485 52322 6519
rect 52314 6451 52322 6485
rect 52280 6417 52322 6451
rect 52314 6383 52322 6417
rect 51751 6349 51790 6374
rect 51302 6297 51318 6331
rect 51352 6297 51368 6331
rect 51508 6310 51790 6349
rect 52280 6341 52322 6383
rect 52477 6550 52513 6600
rect 52547 6634 52602 6650
rect 52581 6600 52602 6634
rect 52547 6584 52602 6600
rect 52647 6648 52715 6665
rect 52647 6647 52667 6648
rect 52647 6613 52665 6647
rect 52701 6614 52715 6648
rect 52699 6613 52715 6614
rect 52647 6591 52715 6613
rect 52568 6555 52602 6584
rect 52872 6563 52918 6683
rect 52972 6679 53018 6695
rect 53190 6658 53206 6659
rect 52952 6611 52968 6645
rect 53002 6638 53018 6645
rect 53070 6638 53206 6658
rect 53002 6625 53206 6638
rect 53240 6625 53256 6659
rect 53002 6624 53256 6625
rect 53002 6611 53110 6624
rect 53190 6622 53256 6624
rect 53488 6655 53522 6657
rect 52952 6597 53110 6611
rect 52966 6596 53110 6597
rect 53488 6619 53522 6621
rect 53162 6563 53196 6582
rect 52477 6500 52531 6550
rect 52568 6521 52703 6555
rect 52477 6466 52495 6500
rect 52529 6466 52531 6500
rect 52667 6487 52703 6521
rect 52477 6419 52531 6466
rect 52477 6385 52495 6419
rect 52529 6385 52531 6419
rect 52477 6369 52531 6385
rect 52565 6453 52581 6487
rect 52615 6453 52631 6487
rect 52565 6419 52631 6453
rect 52565 6385 52581 6419
rect 52615 6385 52631 6419
rect 51676 6308 51790 6310
rect 51948 6297 51964 6331
rect 51998 6297 52014 6331
rect 52114 6307 52143 6341
rect 52177 6307 52235 6341
rect 52269 6307 52327 6341
rect 52361 6307 52390 6341
rect 52565 6335 52631 6385
rect 52701 6453 52703 6487
rect 52667 6419 52703 6453
rect 52701 6385 52703 6419
rect 52667 6369 52703 6385
rect 52872 6545 52938 6563
rect 52872 6511 52888 6545
rect 52922 6511 52938 6545
rect 52872 6477 52938 6511
rect 52872 6443 52888 6477
rect 52922 6443 52938 6477
rect 52872 6409 52938 6443
rect 52872 6375 52888 6409
rect 52922 6375 52938 6409
rect 52872 6367 52938 6375
rect 52972 6545 53014 6561
rect 53006 6511 53014 6545
rect 52972 6477 53014 6511
rect 53006 6443 53014 6477
rect 52972 6409 53014 6443
rect 53162 6495 53196 6497
rect 53162 6459 53196 6461
rect 53006 6375 53014 6409
rect 52281 6300 52315 6307
rect 52460 6301 52489 6335
rect 52523 6301 52581 6335
rect 52615 6301 52673 6335
rect 52707 6301 52736 6335
rect 52972 6333 53014 6375
rect 53122 6393 53162 6414
rect 53250 6563 53284 6582
rect 53488 6534 53522 6553
rect 53584 6723 53618 6742
rect 53584 6655 53618 6657
rect 53584 6619 53618 6621
rect 53584 6534 53618 6553
rect 53680 6723 53714 6742
rect 54068 6737 54134 6750
rect 54068 6703 54084 6737
rect 54118 6703 54134 6737
rect 54068 6691 54134 6703
rect 54168 6805 54214 6851
rect 54348 6845 54377 6879
rect 54411 6845 54469 6879
rect 54503 6845 54561 6879
rect 54595 6845 54624 6879
rect 54202 6771 54214 6805
rect 54168 6737 54214 6771
rect 54202 6703 54214 6737
rect 53680 6655 53714 6657
rect 53836 6625 53852 6659
rect 53886 6625 53902 6659
rect 53680 6619 53714 6621
rect 53680 6534 53714 6553
rect 53808 6563 53842 6582
rect 53250 6495 53284 6497
rect 53808 6495 53842 6497
rect 53250 6459 53284 6461
rect 53520 6457 53536 6491
rect 53570 6457 53586 6491
rect 53808 6459 53842 6461
rect 53196 6393 53198 6414
rect 53122 6374 53198 6393
rect 53284 6393 53808 6418
rect 53896 6563 53930 6582
rect 53896 6495 53930 6497
rect 53896 6459 53930 6461
rect 53842 6393 53844 6418
rect 53250 6385 53844 6393
rect 53250 6374 53486 6385
rect 52806 6299 52835 6333
rect 52869 6299 52927 6333
rect 52961 6299 53019 6333
rect 53053 6299 53082 6333
rect 51368 6212 51414 6218
rect 51368 6210 51856 6212
rect 51368 6176 51376 6210
rect 51410 6193 51856 6210
rect 51410 6188 51806 6193
rect 51410 6178 51685 6188
rect 51410 6176 51414 6178
rect 51368 6174 51414 6176
rect 51586 6154 51685 6178
rect 51719 6159 51806 6188
rect 51840 6168 51856 6193
rect 51840 6159 51981 6168
rect 51719 6154 51981 6159
rect 51586 6134 51981 6154
rect 51710 6050 51726 6084
rect 51760 6050 51896 6084
rect 51234 6000 51616 6016
rect 51234 5976 51582 6000
rect 51582 5930 51616 5964
rect 51582 5878 51616 5894
rect 51678 6000 51712 6016
rect 51678 5930 51712 5964
rect 51678 5878 51712 5894
rect 51774 6000 51808 6016
rect 51774 5930 51808 5964
rect 51774 5878 51808 5894
rect 50048 5797 50077 5831
rect 50111 5797 50169 5831
rect 50203 5797 50261 5831
rect 50295 5797 50324 5831
rect 51122 5797 51151 5831
rect 51185 5797 51243 5831
rect 51277 5797 51335 5831
rect 51369 5797 51398 5831
rect 51614 5810 51630 5844
rect 51664 5810 51680 5844
rect 50067 5753 50121 5797
rect 50067 5719 50087 5753
rect 50067 5685 50121 5719
rect 50067 5651 50087 5685
rect 50067 5635 50121 5651
rect 50155 5753 50221 5763
rect 50155 5719 50171 5753
rect 50205 5719 50221 5753
rect 50155 5710 50221 5719
rect 50155 5685 50173 5710
rect 50155 5651 50171 5685
rect 50207 5676 50221 5710
rect 50205 5651 50221 5676
rect 50155 5635 50221 5651
rect 50255 5753 50303 5797
rect 50289 5719 50303 5753
rect 50255 5685 50303 5719
rect 50289 5651 50303 5685
rect 50255 5635 50303 5651
rect 51141 5753 51195 5797
rect 51141 5719 51161 5753
rect 51141 5685 51195 5719
rect 51141 5651 51161 5685
rect 51141 5635 51195 5651
rect 51229 5753 51295 5763
rect 51229 5719 51245 5753
rect 51279 5719 51295 5753
rect 51229 5715 51295 5719
rect 51229 5681 51243 5715
rect 51277 5685 51295 5715
rect 51229 5651 51245 5681
rect 51279 5651 51295 5685
rect 51229 5635 51295 5651
rect 51329 5753 51377 5797
rect 51363 5719 51377 5753
rect 51726 5729 51742 5763
rect 51776 5729 51792 5763
rect 51329 5685 51377 5719
rect 51363 5651 51377 5685
rect 51329 5635 51377 5651
rect 51598 5667 51632 5686
rect 50065 5594 50085 5599
rect 50065 5560 50082 5594
rect 50119 5565 50135 5599
rect 50116 5560 50135 5565
rect 50065 5549 50135 5560
rect 50169 5515 50203 5635
rect 50237 5565 50253 5599
rect 50287 5590 50307 5599
rect 50237 5556 50255 5565
rect 50289 5556 50307 5590
rect 50237 5549 50307 5556
rect 51139 5592 51159 5599
rect 51139 5558 51157 5592
rect 51193 5565 51209 5599
rect 51191 5558 51209 5565
rect 51139 5549 51209 5558
rect 51243 5515 51277 5635
rect 51598 5599 51632 5601
rect 51311 5565 51327 5599
rect 51361 5592 51381 5599
rect 51311 5558 51331 5565
rect 51365 5558 51381 5592
rect 51311 5549 51381 5558
rect 51598 5563 51632 5565
rect 49742 5435 50008 5436
rect 49742 5401 49758 5435
rect 49792 5401 50008 5435
rect 49742 5400 50008 5401
rect 50067 5499 50133 5515
rect 50067 5465 50099 5499
rect 50169 5499 50305 5515
rect 50169 5481 50255 5499
rect 50067 5431 50133 5465
rect 49425 5363 49491 5397
rect 49425 5329 49441 5363
rect 49475 5329 49491 5363
rect 50067 5397 50099 5431
rect 50067 5363 50133 5397
rect 49425 5324 49491 5329
rect 49618 5329 49900 5362
rect 49618 5295 49708 5329
rect 49742 5327 49900 5329
rect 49742 5295 49827 5327
rect 49618 5293 49827 5295
rect 49861 5293 49900 5327
rect 49618 5287 49900 5293
rect 50067 5329 50099 5363
rect 50067 5287 50133 5329
rect 50239 5465 50255 5481
rect 50289 5465 50305 5499
rect 50239 5431 50305 5465
rect 50239 5397 50255 5431
rect 50289 5397 50305 5431
rect 50239 5363 50305 5397
rect 50239 5329 50255 5363
rect 50289 5329 50305 5363
rect 50239 5324 50305 5329
rect 51141 5499 51207 5515
rect 51141 5465 51173 5499
rect 51243 5499 51379 5515
rect 51243 5481 51329 5499
rect 51141 5431 51207 5465
rect 51141 5397 51173 5431
rect 51141 5363 51207 5397
rect 51141 5329 51173 5363
rect 51141 5287 51207 5329
rect 51313 5465 51329 5481
rect 51363 5465 51379 5499
rect 51598 5478 51632 5497
rect 51694 5667 51728 5686
rect 51694 5599 51728 5601
rect 51694 5563 51728 5565
rect 51694 5478 51728 5497
rect 51790 5667 51824 5686
rect 51790 5599 51824 5601
rect 51790 5563 51824 5565
rect 51790 5478 51824 5497
rect 51313 5431 51379 5465
rect 51313 5397 51329 5431
rect 51363 5397 51379 5431
rect 51630 5436 51696 5438
rect 51862 5436 51896 6050
rect 51947 5831 51981 6134
rect 52178 5831 52212 6042
rect 53122 6016 53156 6374
rect 53396 6351 53486 6374
rect 53520 6383 53844 6385
rect 53520 6351 53605 6383
rect 53396 6349 53605 6351
rect 53639 6374 53844 6383
rect 53896 6374 53930 6393
rect 54068 6571 54114 6691
rect 54168 6687 54214 6703
rect 54365 6773 54417 6811
rect 54365 6739 54383 6773
rect 54453 6803 54519 6845
rect 54694 6843 54723 6877
rect 54757 6843 54815 6877
rect 54849 6843 54907 6877
rect 54941 6843 54970 6877
rect 55130 6862 55178 6874
rect 55392 6866 55408 6900
rect 55442 6866 55458 6900
rect 55758 6890 55808 6960
rect 57248 6934 57282 6950
rect 57344 7056 57378 7072
rect 57440 7058 57474 7072
rect 57558 7058 57778 7080
rect 57438 7056 57778 7058
rect 57438 7022 57440 7056
rect 57474 7044 57778 7056
rect 57474 7022 57594 7044
rect 57344 6986 57378 7020
rect 57439 7020 57440 7022
rect 57439 6986 57474 7020
rect 57742 6996 57778 7044
rect 57439 6985 57440 6986
rect 57344 6934 57378 6950
rect 57440 6934 57474 6950
rect 57646 6960 57778 6996
rect 59136 7056 59170 7072
rect 59136 6986 59170 7020
rect 55758 6876 55768 6890
rect 54453 6769 54469 6803
rect 54503 6769 54519 6803
rect 54555 6790 54589 6811
rect 54365 6710 54417 6739
rect 54555 6735 54589 6756
rect 54148 6619 54164 6653
rect 54198 6642 54214 6653
rect 54148 6608 54166 6619
rect 54200 6608 54214 6642
rect 54365 6638 54401 6710
rect 54456 6701 54589 6735
rect 54760 6797 54826 6809
rect 54760 6763 54776 6797
rect 54810 6763 54826 6797
rect 54760 6746 54826 6763
rect 54456 6650 54490 6701
rect 54760 6695 54776 6746
rect 54810 6695 54826 6746
rect 54760 6683 54826 6695
rect 54860 6797 54906 6843
rect 54894 6763 54906 6797
rect 54860 6729 54906 6763
rect 54894 6695 54906 6729
rect 55130 6828 55136 6862
rect 55170 6828 55178 6862
rect 55762 6856 55768 6876
rect 55802 6856 55808 6890
rect 55762 6846 55808 6856
rect 55890 6851 55919 6885
rect 55953 6851 56011 6885
rect 56045 6851 56103 6885
rect 56137 6851 56166 6885
rect 55130 6740 55178 6828
rect 55504 6785 55520 6819
rect 55554 6818 55570 6819
rect 55554 6786 55716 6818
rect 55956 6810 56022 6817
rect 55950 6805 56022 6810
rect 55950 6786 55972 6805
rect 55554 6785 55972 6786
rect 55504 6782 55972 6785
rect 55680 6771 55972 6782
rect 56006 6771 56022 6805
rect 55680 6750 56022 6771
rect 55376 6740 55410 6742
rect 55130 6723 55410 6740
rect 55130 6706 55376 6723
rect 54148 6605 54214 6608
rect 54360 6636 54401 6638
rect 54360 6602 54362 6636
rect 54396 6602 54401 6636
rect 54360 6600 54401 6602
rect 54068 6553 54134 6571
rect 54068 6519 54084 6553
rect 54118 6519 54134 6553
rect 54068 6485 54134 6519
rect 54068 6451 54084 6485
rect 54118 6451 54134 6485
rect 54068 6417 54134 6451
rect 54068 6383 54084 6417
rect 54118 6383 54134 6417
rect 54068 6375 54134 6383
rect 54168 6553 54210 6569
rect 54202 6519 54210 6553
rect 54168 6485 54210 6519
rect 54202 6451 54210 6485
rect 54168 6417 54210 6451
rect 54202 6383 54210 6417
rect 53639 6349 53678 6374
rect 53190 6297 53206 6331
rect 53240 6297 53256 6331
rect 53396 6310 53678 6349
rect 54168 6341 54210 6383
rect 54365 6550 54401 6600
rect 54435 6634 54490 6650
rect 54469 6600 54490 6634
rect 54435 6584 54490 6600
rect 54535 6648 54603 6665
rect 54535 6647 54555 6648
rect 54535 6613 54553 6647
rect 54589 6614 54603 6648
rect 54587 6613 54603 6614
rect 54535 6591 54603 6613
rect 54456 6555 54490 6584
rect 54760 6563 54806 6683
rect 54860 6679 54906 6695
rect 55078 6658 55094 6659
rect 54840 6611 54856 6645
rect 54890 6638 54906 6645
rect 54958 6638 55094 6658
rect 54890 6625 55094 6638
rect 55128 6625 55144 6659
rect 54890 6624 55144 6625
rect 54890 6611 54998 6624
rect 55078 6622 55144 6624
rect 55376 6655 55410 6657
rect 54840 6597 54998 6611
rect 54854 6596 54998 6597
rect 55376 6619 55410 6621
rect 55050 6563 55084 6582
rect 54365 6500 54419 6550
rect 54456 6521 54591 6555
rect 54365 6466 54383 6500
rect 54417 6466 54419 6500
rect 54555 6487 54591 6521
rect 54365 6419 54419 6466
rect 54365 6385 54383 6419
rect 54417 6385 54419 6419
rect 54365 6369 54419 6385
rect 54453 6453 54469 6487
rect 54503 6453 54519 6487
rect 54453 6419 54519 6453
rect 54453 6385 54469 6419
rect 54503 6385 54519 6419
rect 53564 6308 53678 6310
rect 53836 6297 53852 6331
rect 53886 6297 53902 6331
rect 54002 6307 54031 6341
rect 54065 6307 54123 6341
rect 54157 6307 54215 6341
rect 54249 6307 54278 6341
rect 54453 6335 54519 6385
rect 54589 6453 54591 6487
rect 54555 6419 54591 6453
rect 54589 6385 54591 6419
rect 54555 6369 54591 6385
rect 54760 6545 54826 6563
rect 54760 6511 54776 6545
rect 54810 6511 54826 6545
rect 54760 6477 54826 6511
rect 54760 6443 54776 6477
rect 54810 6443 54826 6477
rect 54760 6409 54826 6443
rect 54760 6375 54776 6409
rect 54810 6375 54826 6409
rect 54760 6367 54826 6375
rect 54860 6545 54902 6561
rect 54894 6511 54902 6545
rect 54860 6477 54902 6511
rect 54894 6443 54902 6477
rect 54860 6409 54902 6443
rect 55050 6495 55084 6497
rect 55050 6459 55084 6461
rect 54894 6375 54902 6409
rect 54169 6300 54203 6307
rect 54348 6301 54377 6335
rect 54411 6301 54469 6335
rect 54503 6301 54561 6335
rect 54595 6301 54624 6335
rect 54860 6333 54902 6375
rect 55010 6393 55050 6414
rect 55138 6563 55172 6582
rect 55376 6534 55410 6553
rect 55472 6723 55506 6742
rect 55472 6655 55506 6657
rect 55472 6619 55506 6621
rect 55472 6534 55506 6553
rect 55568 6723 55602 6742
rect 55956 6737 56022 6750
rect 55956 6703 55972 6737
rect 56006 6703 56022 6737
rect 55956 6691 56022 6703
rect 56056 6805 56102 6851
rect 56236 6845 56265 6879
rect 56299 6845 56357 6879
rect 56391 6845 56449 6879
rect 56483 6845 56512 6879
rect 56090 6771 56102 6805
rect 56056 6737 56102 6771
rect 56090 6703 56102 6737
rect 55568 6655 55602 6657
rect 55724 6625 55740 6659
rect 55774 6625 55790 6659
rect 55568 6619 55602 6621
rect 55568 6534 55602 6553
rect 55696 6563 55730 6582
rect 55138 6495 55172 6497
rect 55696 6495 55730 6497
rect 55138 6459 55172 6461
rect 55408 6457 55424 6491
rect 55458 6457 55474 6491
rect 55696 6459 55730 6461
rect 55084 6393 55086 6414
rect 55010 6374 55086 6393
rect 55172 6393 55696 6418
rect 55784 6563 55818 6582
rect 55784 6495 55818 6497
rect 55784 6459 55818 6461
rect 55730 6393 55732 6418
rect 55138 6385 55732 6393
rect 55138 6374 55374 6385
rect 54694 6299 54723 6333
rect 54757 6299 54815 6333
rect 54849 6299 54907 6333
rect 54941 6299 54970 6333
rect 53256 6212 53302 6218
rect 53256 6210 53744 6212
rect 53256 6176 53264 6210
rect 53298 6193 53744 6210
rect 53298 6188 53694 6193
rect 53298 6178 53573 6188
rect 53298 6176 53302 6178
rect 53256 6174 53302 6176
rect 53474 6154 53573 6178
rect 53607 6159 53694 6188
rect 53728 6168 53744 6193
rect 53728 6159 53869 6168
rect 53607 6154 53869 6159
rect 53474 6134 53869 6154
rect 53598 6050 53614 6084
rect 53648 6050 53784 6084
rect 53122 6000 53504 6016
rect 53122 5976 53470 6000
rect 53470 5930 53504 5964
rect 53470 5878 53504 5894
rect 53566 6000 53600 6016
rect 53566 5930 53600 5964
rect 53566 5878 53600 5894
rect 53662 6000 53696 6016
rect 53662 5930 53696 5964
rect 53662 5878 53696 5894
rect 51936 5797 51965 5831
rect 51999 5797 52057 5831
rect 52091 5797 52149 5831
rect 52183 5797 52212 5831
rect 53010 5797 53039 5831
rect 53073 5797 53131 5831
rect 53165 5797 53223 5831
rect 53257 5797 53286 5831
rect 53502 5810 53518 5844
rect 53552 5810 53568 5844
rect 51955 5753 52009 5797
rect 51955 5719 51975 5753
rect 51955 5685 52009 5719
rect 51955 5651 51975 5685
rect 51955 5635 52009 5651
rect 52043 5753 52109 5763
rect 52043 5719 52059 5753
rect 52093 5719 52109 5753
rect 52043 5710 52109 5719
rect 52043 5685 52061 5710
rect 52043 5651 52059 5685
rect 52095 5676 52109 5710
rect 52093 5651 52109 5676
rect 52043 5635 52109 5651
rect 52143 5753 52191 5797
rect 52177 5719 52191 5753
rect 52143 5685 52191 5719
rect 52177 5651 52191 5685
rect 52143 5635 52191 5651
rect 53029 5753 53083 5797
rect 53029 5719 53049 5753
rect 53029 5685 53083 5719
rect 53029 5651 53049 5685
rect 53029 5635 53083 5651
rect 53117 5753 53183 5763
rect 53117 5719 53133 5753
rect 53167 5719 53183 5753
rect 53117 5715 53183 5719
rect 53117 5681 53131 5715
rect 53165 5685 53183 5715
rect 53117 5651 53133 5681
rect 53167 5651 53183 5685
rect 53117 5635 53183 5651
rect 53217 5753 53265 5797
rect 53251 5719 53265 5753
rect 53614 5729 53630 5763
rect 53664 5729 53680 5763
rect 53217 5685 53265 5719
rect 53251 5651 53265 5685
rect 53217 5635 53265 5651
rect 53486 5667 53520 5686
rect 51953 5594 51973 5599
rect 51953 5560 51970 5594
rect 52007 5565 52023 5599
rect 52004 5560 52023 5565
rect 51953 5549 52023 5560
rect 52057 5515 52091 5635
rect 52125 5565 52141 5599
rect 52175 5590 52195 5599
rect 52125 5556 52143 5565
rect 52177 5556 52195 5590
rect 52125 5549 52195 5556
rect 53027 5592 53047 5599
rect 53027 5558 53045 5592
rect 53081 5565 53097 5599
rect 53079 5558 53097 5565
rect 53027 5549 53097 5558
rect 53131 5515 53165 5635
rect 53486 5599 53520 5601
rect 53199 5565 53215 5599
rect 53249 5592 53269 5599
rect 53199 5558 53219 5565
rect 53253 5558 53269 5592
rect 53199 5549 53269 5558
rect 53486 5563 53520 5565
rect 51630 5435 51896 5436
rect 51630 5401 51646 5435
rect 51680 5401 51896 5435
rect 51630 5400 51896 5401
rect 51955 5499 52021 5515
rect 51955 5465 51987 5499
rect 52057 5499 52193 5515
rect 52057 5481 52143 5499
rect 51955 5431 52021 5465
rect 51313 5363 51379 5397
rect 51313 5329 51329 5363
rect 51363 5329 51379 5363
rect 51955 5397 51987 5431
rect 51955 5363 52021 5397
rect 51313 5324 51379 5329
rect 51506 5329 51788 5362
rect 51506 5295 51596 5329
rect 51630 5327 51788 5329
rect 51630 5295 51715 5327
rect 51506 5293 51715 5295
rect 51749 5293 51788 5327
rect 51506 5287 51788 5293
rect 51955 5329 51987 5363
rect 51955 5287 52021 5329
rect 52127 5465 52143 5481
rect 52177 5465 52193 5499
rect 52127 5431 52193 5465
rect 52127 5397 52143 5431
rect 52177 5397 52193 5431
rect 52127 5363 52193 5397
rect 52127 5329 52143 5363
rect 52177 5329 52193 5363
rect 52127 5324 52193 5329
rect 53029 5499 53095 5515
rect 53029 5465 53061 5499
rect 53131 5499 53267 5515
rect 53131 5481 53217 5499
rect 53029 5431 53095 5465
rect 53029 5397 53061 5431
rect 53029 5363 53095 5397
rect 53029 5329 53061 5363
rect 53029 5287 53095 5329
rect 53201 5465 53217 5481
rect 53251 5465 53267 5499
rect 53486 5478 53520 5497
rect 53582 5667 53616 5686
rect 53582 5599 53616 5601
rect 53582 5563 53616 5565
rect 53582 5478 53616 5497
rect 53678 5667 53712 5686
rect 53678 5599 53712 5601
rect 53678 5563 53712 5565
rect 53678 5478 53712 5497
rect 53201 5431 53267 5465
rect 53201 5397 53217 5431
rect 53251 5397 53267 5431
rect 53518 5436 53584 5438
rect 53750 5436 53784 6050
rect 53835 5831 53869 6134
rect 54066 5831 54100 6042
rect 55010 6016 55044 6374
rect 55284 6351 55374 6374
rect 55408 6383 55732 6385
rect 55408 6351 55493 6383
rect 55284 6349 55493 6351
rect 55527 6374 55732 6383
rect 55784 6374 55818 6393
rect 55956 6571 56002 6691
rect 56056 6687 56102 6703
rect 56253 6773 56305 6811
rect 56253 6739 56271 6773
rect 56341 6803 56407 6845
rect 56582 6843 56611 6877
rect 56645 6843 56703 6877
rect 56737 6843 56795 6877
rect 56829 6843 56858 6877
rect 57018 6862 57066 6874
rect 57280 6866 57296 6900
rect 57330 6866 57346 6900
rect 57646 6890 57696 6960
rect 59136 6934 59170 6950
rect 59232 7056 59266 7072
rect 59328 7058 59362 7072
rect 59446 7058 59666 7080
rect 59326 7056 59666 7058
rect 59326 7022 59328 7056
rect 59362 7044 59666 7056
rect 59362 7022 59482 7044
rect 59232 6986 59266 7020
rect 59327 7020 59328 7022
rect 59327 6986 59362 7020
rect 59630 6996 59666 7044
rect 59327 6985 59328 6986
rect 59232 6934 59266 6950
rect 59328 6934 59362 6950
rect 59534 6960 59666 6996
rect 57646 6876 57656 6890
rect 56341 6769 56357 6803
rect 56391 6769 56407 6803
rect 56443 6790 56477 6811
rect 56253 6710 56305 6739
rect 56443 6735 56477 6756
rect 56036 6619 56052 6653
rect 56086 6642 56102 6653
rect 56036 6608 56054 6619
rect 56088 6608 56102 6642
rect 56253 6638 56289 6710
rect 56344 6701 56477 6735
rect 56648 6797 56714 6809
rect 56648 6763 56664 6797
rect 56698 6763 56714 6797
rect 56648 6746 56714 6763
rect 56344 6650 56378 6701
rect 56648 6695 56664 6746
rect 56698 6695 56714 6746
rect 56648 6683 56714 6695
rect 56748 6797 56794 6843
rect 56782 6763 56794 6797
rect 56748 6729 56794 6763
rect 56782 6695 56794 6729
rect 57018 6828 57024 6862
rect 57058 6828 57066 6862
rect 57650 6856 57656 6876
rect 57690 6856 57696 6890
rect 57650 6846 57696 6856
rect 57778 6851 57807 6885
rect 57841 6851 57899 6885
rect 57933 6851 57991 6885
rect 58025 6851 58054 6885
rect 57018 6740 57066 6828
rect 57392 6785 57408 6819
rect 57442 6818 57458 6819
rect 57442 6786 57604 6818
rect 57844 6810 57910 6817
rect 57838 6805 57910 6810
rect 57838 6786 57860 6805
rect 57442 6785 57860 6786
rect 57392 6782 57860 6785
rect 57568 6771 57860 6782
rect 57894 6771 57910 6805
rect 57568 6750 57910 6771
rect 57264 6740 57298 6742
rect 57018 6723 57298 6740
rect 57018 6706 57264 6723
rect 56036 6605 56102 6608
rect 56248 6636 56289 6638
rect 56248 6602 56250 6636
rect 56284 6602 56289 6636
rect 56248 6600 56289 6602
rect 55956 6553 56022 6571
rect 55956 6519 55972 6553
rect 56006 6519 56022 6553
rect 55956 6485 56022 6519
rect 55956 6451 55972 6485
rect 56006 6451 56022 6485
rect 55956 6417 56022 6451
rect 55956 6383 55972 6417
rect 56006 6383 56022 6417
rect 55956 6375 56022 6383
rect 56056 6553 56098 6569
rect 56090 6519 56098 6553
rect 56056 6485 56098 6519
rect 56090 6451 56098 6485
rect 56056 6417 56098 6451
rect 56090 6383 56098 6417
rect 55527 6349 55566 6374
rect 55078 6297 55094 6331
rect 55128 6297 55144 6331
rect 55284 6310 55566 6349
rect 56056 6341 56098 6383
rect 56253 6550 56289 6600
rect 56323 6634 56378 6650
rect 56357 6600 56378 6634
rect 56323 6584 56378 6600
rect 56423 6648 56491 6665
rect 56423 6647 56443 6648
rect 56423 6613 56441 6647
rect 56477 6614 56491 6648
rect 56475 6613 56491 6614
rect 56423 6591 56491 6613
rect 56344 6555 56378 6584
rect 56648 6563 56694 6683
rect 56748 6679 56794 6695
rect 56966 6658 56982 6659
rect 56728 6611 56744 6645
rect 56778 6638 56794 6645
rect 56846 6638 56982 6658
rect 56778 6625 56982 6638
rect 57016 6625 57032 6659
rect 56778 6624 57032 6625
rect 56778 6611 56886 6624
rect 56966 6622 57032 6624
rect 57264 6655 57298 6657
rect 56728 6597 56886 6611
rect 56742 6596 56886 6597
rect 57264 6619 57298 6621
rect 56938 6563 56972 6582
rect 56253 6500 56307 6550
rect 56344 6521 56479 6555
rect 56253 6466 56271 6500
rect 56305 6466 56307 6500
rect 56443 6487 56479 6521
rect 56253 6419 56307 6466
rect 56253 6385 56271 6419
rect 56305 6385 56307 6419
rect 56253 6369 56307 6385
rect 56341 6453 56357 6487
rect 56391 6453 56407 6487
rect 56341 6419 56407 6453
rect 56341 6385 56357 6419
rect 56391 6385 56407 6419
rect 55452 6308 55566 6310
rect 55724 6297 55740 6331
rect 55774 6297 55790 6331
rect 55890 6307 55919 6341
rect 55953 6307 56011 6341
rect 56045 6307 56103 6341
rect 56137 6307 56166 6341
rect 56341 6335 56407 6385
rect 56477 6453 56479 6487
rect 56443 6419 56479 6453
rect 56477 6385 56479 6419
rect 56443 6369 56479 6385
rect 56648 6545 56714 6563
rect 56648 6511 56664 6545
rect 56698 6511 56714 6545
rect 56648 6477 56714 6511
rect 56648 6443 56664 6477
rect 56698 6443 56714 6477
rect 56648 6409 56714 6443
rect 56648 6375 56664 6409
rect 56698 6375 56714 6409
rect 56648 6367 56714 6375
rect 56748 6545 56790 6561
rect 56782 6511 56790 6545
rect 56748 6477 56790 6511
rect 56782 6443 56790 6477
rect 56748 6409 56790 6443
rect 56938 6495 56972 6497
rect 56938 6459 56972 6461
rect 56782 6375 56790 6409
rect 56057 6300 56091 6307
rect 56236 6301 56265 6335
rect 56299 6301 56357 6335
rect 56391 6301 56449 6335
rect 56483 6301 56512 6335
rect 56748 6333 56790 6375
rect 56898 6393 56938 6414
rect 57026 6563 57060 6582
rect 57264 6534 57298 6553
rect 57360 6723 57394 6742
rect 57360 6655 57394 6657
rect 57360 6619 57394 6621
rect 57360 6534 57394 6553
rect 57456 6723 57490 6742
rect 57844 6737 57910 6750
rect 57844 6703 57860 6737
rect 57894 6703 57910 6737
rect 57844 6691 57910 6703
rect 57944 6805 57990 6851
rect 58124 6845 58153 6879
rect 58187 6845 58245 6879
rect 58279 6845 58337 6879
rect 58371 6845 58400 6879
rect 57978 6771 57990 6805
rect 57944 6737 57990 6771
rect 57978 6703 57990 6737
rect 57456 6655 57490 6657
rect 57612 6625 57628 6659
rect 57662 6625 57678 6659
rect 57456 6619 57490 6621
rect 57456 6534 57490 6553
rect 57584 6563 57618 6582
rect 57026 6495 57060 6497
rect 57584 6495 57618 6497
rect 57026 6459 57060 6461
rect 57296 6457 57312 6491
rect 57346 6457 57362 6491
rect 57584 6459 57618 6461
rect 56972 6393 56974 6414
rect 56898 6374 56974 6393
rect 57060 6393 57584 6418
rect 57672 6563 57706 6582
rect 57672 6495 57706 6497
rect 57672 6459 57706 6461
rect 57618 6393 57620 6418
rect 57026 6385 57620 6393
rect 57026 6374 57262 6385
rect 56582 6299 56611 6333
rect 56645 6299 56703 6333
rect 56737 6299 56795 6333
rect 56829 6299 56858 6333
rect 55144 6212 55190 6218
rect 55144 6210 55632 6212
rect 55144 6176 55152 6210
rect 55186 6193 55632 6210
rect 55186 6188 55582 6193
rect 55186 6178 55461 6188
rect 55186 6176 55190 6178
rect 55144 6174 55190 6176
rect 55362 6154 55461 6178
rect 55495 6159 55582 6188
rect 55616 6168 55632 6193
rect 55616 6159 55757 6168
rect 55495 6154 55757 6159
rect 55362 6134 55757 6154
rect 55486 6050 55502 6084
rect 55536 6050 55672 6084
rect 55010 6000 55392 6016
rect 55010 5976 55358 6000
rect 55358 5930 55392 5964
rect 55358 5878 55392 5894
rect 55454 6000 55488 6016
rect 55454 5930 55488 5964
rect 55454 5878 55488 5894
rect 55550 6000 55584 6016
rect 55550 5930 55584 5964
rect 55550 5878 55584 5894
rect 53824 5797 53853 5831
rect 53887 5797 53945 5831
rect 53979 5797 54037 5831
rect 54071 5797 54100 5831
rect 54898 5797 54927 5831
rect 54961 5797 55019 5831
rect 55053 5797 55111 5831
rect 55145 5797 55174 5831
rect 55390 5810 55406 5844
rect 55440 5810 55456 5844
rect 53843 5753 53897 5797
rect 53843 5719 53863 5753
rect 53843 5685 53897 5719
rect 53843 5651 53863 5685
rect 53843 5635 53897 5651
rect 53931 5753 53997 5763
rect 53931 5719 53947 5753
rect 53981 5719 53997 5753
rect 53931 5710 53997 5719
rect 53931 5685 53949 5710
rect 53931 5651 53947 5685
rect 53983 5676 53997 5710
rect 53981 5651 53997 5676
rect 53931 5635 53997 5651
rect 54031 5753 54079 5797
rect 54065 5719 54079 5753
rect 54031 5685 54079 5719
rect 54065 5651 54079 5685
rect 54031 5635 54079 5651
rect 54917 5753 54971 5797
rect 54917 5719 54937 5753
rect 54917 5685 54971 5719
rect 54917 5651 54937 5685
rect 54917 5635 54971 5651
rect 55005 5753 55071 5763
rect 55005 5719 55021 5753
rect 55055 5719 55071 5753
rect 55005 5715 55071 5719
rect 55005 5681 55019 5715
rect 55053 5685 55071 5715
rect 55005 5651 55021 5681
rect 55055 5651 55071 5685
rect 55005 5635 55071 5651
rect 55105 5753 55153 5797
rect 55139 5719 55153 5753
rect 55502 5729 55518 5763
rect 55552 5729 55568 5763
rect 55105 5685 55153 5719
rect 55139 5651 55153 5685
rect 55105 5635 55153 5651
rect 55374 5667 55408 5686
rect 53841 5594 53861 5599
rect 53841 5560 53858 5594
rect 53895 5565 53911 5599
rect 53892 5560 53911 5565
rect 53841 5549 53911 5560
rect 53945 5515 53979 5635
rect 54013 5565 54029 5599
rect 54063 5590 54083 5599
rect 54013 5556 54031 5565
rect 54065 5556 54083 5590
rect 54013 5549 54083 5556
rect 54915 5592 54935 5599
rect 54915 5558 54933 5592
rect 54969 5565 54985 5599
rect 54967 5558 54985 5565
rect 54915 5549 54985 5558
rect 55019 5515 55053 5635
rect 55374 5599 55408 5601
rect 55087 5565 55103 5599
rect 55137 5592 55157 5599
rect 55087 5558 55107 5565
rect 55141 5558 55157 5592
rect 55087 5549 55157 5558
rect 55374 5563 55408 5565
rect 53518 5435 53784 5436
rect 53518 5401 53534 5435
rect 53568 5401 53784 5435
rect 53518 5400 53784 5401
rect 53843 5499 53909 5515
rect 53843 5465 53875 5499
rect 53945 5499 54081 5515
rect 53945 5481 54031 5499
rect 53843 5431 53909 5465
rect 53201 5363 53267 5397
rect 53201 5329 53217 5363
rect 53251 5329 53267 5363
rect 53843 5397 53875 5431
rect 53843 5363 53909 5397
rect 53201 5324 53267 5329
rect 53394 5329 53676 5362
rect 53394 5295 53484 5329
rect 53518 5327 53676 5329
rect 53518 5295 53603 5327
rect 53394 5293 53603 5295
rect 53637 5293 53676 5327
rect 53394 5287 53676 5293
rect 53843 5329 53875 5363
rect 53843 5287 53909 5329
rect 54015 5465 54031 5481
rect 54065 5465 54081 5499
rect 54015 5431 54081 5465
rect 54015 5397 54031 5431
rect 54065 5397 54081 5431
rect 54015 5363 54081 5397
rect 54015 5329 54031 5363
rect 54065 5329 54081 5363
rect 54015 5324 54081 5329
rect 54917 5499 54983 5515
rect 54917 5465 54949 5499
rect 55019 5499 55155 5515
rect 55019 5481 55105 5499
rect 54917 5431 54983 5465
rect 54917 5397 54949 5431
rect 54917 5363 54983 5397
rect 54917 5329 54949 5363
rect 54917 5287 54983 5329
rect 55089 5465 55105 5481
rect 55139 5465 55155 5499
rect 55374 5478 55408 5497
rect 55470 5667 55504 5686
rect 55470 5599 55504 5601
rect 55470 5563 55504 5565
rect 55470 5478 55504 5497
rect 55566 5667 55600 5686
rect 55566 5599 55600 5601
rect 55566 5563 55600 5565
rect 55566 5478 55600 5497
rect 55089 5431 55155 5465
rect 55089 5397 55105 5431
rect 55139 5397 55155 5431
rect 55406 5436 55472 5438
rect 55638 5436 55672 6050
rect 55723 5831 55757 6134
rect 55954 5831 55988 6042
rect 56898 6016 56932 6374
rect 57172 6351 57262 6374
rect 57296 6383 57620 6385
rect 57296 6351 57381 6383
rect 57172 6349 57381 6351
rect 57415 6374 57620 6383
rect 57672 6374 57706 6393
rect 57844 6571 57890 6691
rect 57944 6687 57990 6703
rect 58141 6773 58193 6811
rect 58141 6739 58159 6773
rect 58229 6803 58295 6845
rect 58470 6843 58499 6877
rect 58533 6843 58591 6877
rect 58625 6843 58683 6877
rect 58717 6843 58746 6877
rect 58906 6862 58954 6874
rect 59168 6866 59184 6900
rect 59218 6866 59234 6900
rect 59534 6890 59584 6960
rect 59534 6876 59544 6890
rect 58229 6769 58245 6803
rect 58279 6769 58295 6803
rect 58331 6790 58365 6811
rect 58141 6710 58193 6739
rect 58331 6735 58365 6756
rect 57924 6619 57940 6653
rect 57974 6642 57990 6653
rect 57924 6608 57942 6619
rect 57976 6608 57990 6642
rect 58141 6638 58177 6710
rect 58232 6701 58365 6735
rect 58536 6797 58602 6809
rect 58536 6763 58552 6797
rect 58586 6763 58602 6797
rect 58536 6746 58602 6763
rect 58232 6650 58266 6701
rect 58536 6695 58552 6746
rect 58586 6695 58602 6746
rect 58536 6683 58602 6695
rect 58636 6797 58682 6843
rect 58670 6763 58682 6797
rect 58636 6729 58682 6763
rect 58670 6695 58682 6729
rect 58906 6828 58912 6862
rect 58946 6828 58954 6862
rect 59538 6856 59544 6876
rect 59578 6856 59584 6890
rect 59538 6846 59584 6856
rect 59666 6851 59695 6885
rect 59729 6851 59787 6885
rect 59821 6851 59879 6885
rect 59913 6851 59942 6885
rect 58906 6740 58954 6828
rect 59280 6785 59296 6819
rect 59330 6818 59346 6819
rect 59330 6786 59492 6818
rect 59732 6810 59798 6817
rect 59726 6805 59798 6810
rect 59726 6786 59748 6805
rect 59330 6785 59748 6786
rect 59280 6782 59748 6785
rect 59456 6771 59748 6782
rect 59782 6771 59798 6805
rect 59456 6750 59798 6771
rect 59152 6740 59186 6742
rect 58906 6723 59186 6740
rect 58906 6706 59152 6723
rect 57924 6605 57990 6608
rect 58136 6636 58177 6638
rect 58136 6602 58138 6636
rect 58172 6602 58177 6636
rect 58136 6600 58177 6602
rect 57844 6553 57910 6571
rect 57844 6519 57860 6553
rect 57894 6519 57910 6553
rect 57844 6485 57910 6519
rect 57844 6451 57860 6485
rect 57894 6451 57910 6485
rect 57844 6417 57910 6451
rect 57844 6383 57860 6417
rect 57894 6383 57910 6417
rect 57844 6375 57910 6383
rect 57944 6553 57986 6569
rect 57978 6519 57986 6553
rect 57944 6485 57986 6519
rect 57978 6451 57986 6485
rect 57944 6417 57986 6451
rect 57978 6383 57986 6417
rect 57415 6349 57454 6374
rect 56966 6297 56982 6331
rect 57016 6297 57032 6331
rect 57172 6310 57454 6349
rect 57944 6341 57986 6383
rect 58141 6550 58177 6600
rect 58211 6634 58266 6650
rect 58245 6600 58266 6634
rect 58211 6584 58266 6600
rect 58311 6648 58379 6665
rect 58311 6647 58331 6648
rect 58311 6613 58329 6647
rect 58365 6614 58379 6648
rect 58363 6613 58379 6614
rect 58311 6591 58379 6613
rect 58232 6555 58266 6584
rect 58536 6563 58582 6683
rect 58636 6679 58682 6695
rect 58854 6658 58870 6659
rect 58616 6611 58632 6645
rect 58666 6638 58682 6645
rect 58734 6638 58870 6658
rect 58666 6625 58870 6638
rect 58904 6625 58920 6659
rect 58666 6624 58920 6625
rect 58666 6611 58774 6624
rect 58854 6622 58920 6624
rect 59152 6655 59186 6657
rect 58616 6597 58774 6611
rect 58630 6596 58774 6597
rect 59152 6619 59186 6621
rect 58826 6563 58860 6582
rect 58141 6500 58195 6550
rect 58232 6521 58367 6555
rect 58141 6466 58159 6500
rect 58193 6466 58195 6500
rect 58331 6487 58367 6521
rect 58141 6419 58195 6466
rect 58141 6385 58159 6419
rect 58193 6385 58195 6419
rect 58141 6369 58195 6385
rect 58229 6453 58245 6487
rect 58279 6453 58295 6487
rect 58229 6419 58295 6453
rect 58229 6385 58245 6419
rect 58279 6385 58295 6419
rect 57340 6308 57454 6310
rect 57612 6297 57628 6331
rect 57662 6297 57678 6331
rect 57778 6307 57807 6341
rect 57841 6307 57899 6341
rect 57933 6307 57991 6341
rect 58025 6307 58054 6341
rect 58229 6335 58295 6385
rect 58365 6453 58367 6487
rect 58331 6419 58367 6453
rect 58365 6385 58367 6419
rect 58331 6369 58367 6385
rect 58536 6545 58602 6563
rect 58536 6511 58552 6545
rect 58586 6511 58602 6545
rect 58536 6477 58602 6511
rect 58536 6443 58552 6477
rect 58586 6443 58602 6477
rect 58536 6409 58602 6443
rect 58536 6375 58552 6409
rect 58586 6375 58602 6409
rect 58536 6367 58602 6375
rect 58636 6545 58678 6561
rect 58670 6511 58678 6545
rect 58636 6477 58678 6511
rect 58670 6443 58678 6477
rect 58636 6409 58678 6443
rect 58826 6495 58860 6497
rect 58826 6459 58860 6461
rect 58670 6375 58678 6409
rect 57945 6300 57979 6307
rect 58124 6301 58153 6335
rect 58187 6301 58245 6335
rect 58279 6301 58337 6335
rect 58371 6301 58400 6335
rect 58636 6333 58678 6375
rect 58786 6393 58826 6414
rect 58914 6563 58948 6582
rect 59152 6534 59186 6553
rect 59248 6723 59282 6742
rect 59248 6655 59282 6657
rect 59248 6619 59282 6621
rect 59248 6534 59282 6553
rect 59344 6723 59378 6742
rect 59732 6737 59798 6750
rect 59732 6703 59748 6737
rect 59782 6703 59798 6737
rect 59732 6691 59798 6703
rect 59832 6805 59878 6851
rect 59866 6771 59878 6805
rect 59832 6737 59878 6771
rect 59866 6703 59878 6737
rect 59344 6655 59378 6657
rect 59500 6625 59516 6659
rect 59550 6625 59566 6659
rect 59344 6619 59378 6621
rect 59344 6534 59378 6553
rect 59472 6563 59506 6582
rect 58914 6495 58948 6497
rect 59472 6495 59506 6497
rect 58914 6459 58948 6461
rect 59184 6457 59200 6491
rect 59234 6457 59250 6491
rect 59472 6459 59506 6461
rect 58860 6393 58862 6414
rect 58786 6374 58862 6393
rect 58948 6393 59472 6418
rect 59560 6563 59594 6582
rect 59560 6495 59594 6497
rect 59560 6459 59594 6461
rect 59506 6393 59508 6418
rect 58914 6385 59508 6393
rect 58914 6374 59150 6385
rect 58470 6299 58499 6333
rect 58533 6299 58591 6333
rect 58625 6299 58683 6333
rect 58717 6299 58746 6333
rect 57032 6212 57078 6218
rect 57032 6210 57520 6212
rect 57032 6176 57040 6210
rect 57074 6193 57520 6210
rect 57074 6188 57470 6193
rect 57074 6178 57349 6188
rect 57074 6176 57078 6178
rect 57032 6174 57078 6176
rect 57250 6154 57349 6178
rect 57383 6159 57470 6188
rect 57504 6168 57520 6193
rect 57504 6159 57645 6168
rect 57383 6154 57645 6159
rect 57250 6134 57645 6154
rect 57374 6050 57390 6084
rect 57424 6050 57560 6084
rect 56898 6000 57280 6016
rect 56898 5976 57246 6000
rect 57246 5930 57280 5964
rect 57246 5878 57280 5894
rect 57342 6000 57376 6016
rect 57342 5930 57376 5964
rect 57342 5878 57376 5894
rect 57438 6000 57472 6016
rect 57438 5930 57472 5964
rect 57438 5878 57472 5894
rect 55712 5797 55741 5831
rect 55775 5797 55833 5831
rect 55867 5797 55925 5831
rect 55959 5797 55988 5831
rect 56786 5797 56815 5831
rect 56849 5797 56907 5831
rect 56941 5797 56999 5831
rect 57033 5797 57062 5831
rect 57278 5810 57294 5844
rect 57328 5810 57344 5844
rect 55731 5753 55785 5797
rect 55731 5719 55751 5753
rect 55731 5685 55785 5719
rect 55731 5651 55751 5685
rect 55731 5635 55785 5651
rect 55819 5753 55885 5763
rect 55819 5719 55835 5753
rect 55869 5719 55885 5753
rect 55819 5710 55885 5719
rect 55819 5685 55837 5710
rect 55819 5651 55835 5685
rect 55871 5676 55885 5710
rect 55869 5651 55885 5676
rect 55819 5635 55885 5651
rect 55919 5753 55967 5797
rect 55953 5719 55967 5753
rect 55919 5685 55967 5719
rect 55953 5651 55967 5685
rect 55919 5635 55967 5651
rect 56805 5753 56859 5797
rect 56805 5719 56825 5753
rect 56805 5685 56859 5719
rect 56805 5651 56825 5685
rect 56805 5635 56859 5651
rect 56893 5753 56959 5763
rect 56893 5719 56909 5753
rect 56943 5719 56959 5753
rect 56893 5715 56959 5719
rect 56893 5681 56907 5715
rect 56941 5685 56959 5715
rect 56893 5651 56909 5681
rect 56943 5651 56959 5685
rect 56893 5635 56959 5651
rect 56993 5753 57041 5797
rect 57027 5719 57041 5753
rect 57390 5729 57406 5763
rect 57440 5729 57456 5763
rect 56993 5685 57041 5719
rect 57027 5651 57041 5685
rect 56993 5635 57041 5651
rect 57262 5667 57296 5686
rect 55729 5594 55749 5599
rect 55729 5560 55746 5594
rect 55783 5565 55799 5599
rect 55780 5560 55799 5565
rect 55729 5549 55799 5560
rect 55833 5515 55867 5635
rect 55901 5565 55917 5599
rect 55951 5590 55971 5599
rect 55901 5556 55919 5565
rect 55953 5556 55971 5590
rect 55901 5549 55971 5556
rect 56803 5592 56823 5599
rect 56803 5558 56821 5592
rect 56857 5565 56873 5599
rect 56855 5558 56873 5565
rect 56803 5549 56873 5558
rect 56907 5515 56941 5635
rect 57262 5599 57296 5601
rect 56975 5565 56991 5599
rect 57025 5592 57045 5599
rect 56975 5558 56995 5565
rect 57029 5558 57045 5592
rect 56975 5549 57045 5558
rect 57262 5563 57296 5565
rect 55406 5435 55672 5436
rect 55406 5401 55422 5435
rect 55456 5401 55672 5435
rect 55406 5400 55672 5401
rect 55731 5499 55797 5515
rect 55731 5465 55763 5499
rect 55833 5499 55969 5515
rect 55833 5481 55919 5499
rect 55731 5431 55797 5465
rect 55089 5363 55155 5397
rect 55089 5329 55105 5363
rect 55139 5329 55155 5363
rect 55731 5397 55763 5431
rect 55731 5363 55797 5397
rect 55089 5324 55155 5329
rect 55282 5329 55564 5362
rect 55282 5295 55372 5329
rect 55406 5327 55564 5329
rect 55406 5295 55491 5327
rect 55282 5293 55491 5295
rect 55525 5293 55564 5327
rect 55282 5287 55564 5293
rect 55731 5329 55763 5363
rect 55731 5287 55797 5329
rect 55903 5465 55919 5481
rect 55953 5465 55969 5499
rect 55903 5431 55969 5465
rect 55903 5397 55919 5431
rect 55953 5397 55969 5431
rect 55903 5363 55969 5397
rect 55903 5329 55919 5363
rect 55953 5329 55969 5363
rect 55903 5324 55969 5329
rect 56805 5499 56871 5515
rect 56805 5465 56837 5499
rect 56907 5499 57043 5515
rect 56907 5481 56993 5499
rect 56805 5431 56871 5465
rect 56805 5397 56837 5431
rect 56805 5363 56871 5397
rect 56805 5329 56837 5363
rect 56805 5287 56871 5329
rect 56977 5465 56993 5481
rect 57027 5465 57043 5499
rect 57262 5478 57296 5497
rect 57358 5667 57392 5686
rect 57358 5599 57392 5601
rect 57358 5563 57392 5565
rect 57358 5478 57392 5497
rect 57454 5667 57488 5686
rect 57454 5599 57488 5601
rect 57454 5563 57488 5565
rect 57454 5478 57488 5497
rect 56977 5431 57043 5465
rect 56977 5397 56993 5431
rect 57027 5397 57043 5431
rect 57294 5436 57360 5438
rect 57526 5436 57560 6050
rect 57611 5831 57645 6134
rect 57842 5831 57876 6042
rect 58786 6016 58820 6374
rect 59060 6351 59150 6374
rect 59184 6383 59508 6385
rect 59184 6351 59269 6383
rect 59060 6349 59269 6351
rect 59303 6374 59508 6383
rect 59560 6374 59594 6393
rect 59732 6571 59778 6691
rect 59832 6687 59878 6703
rect 59812 6619 59828 6653
rect 59862 6642 59878 6653
rect 59812 6608 59830 6619
rect 59864 6608 59878 6642
rect 59812 6605 59878 6608
rect 59732 6553 59798 6571
rect 59732 6519 59748 6553
rect 59782 6519 59798 6553
rect 59732 6485 59798 6519
rect 59732 6451 59748 6485
rect 59782 6451 59798 6485
rect 59732 6417 59798 6451
rect 59732 6383 59748 6417
rect 59782 6383 59798 6417
rect 59732 6375 59798 6383
rect 59832 6553 59874 6569
rect 59866 6519 59874 6553
rect 59832 6485 59874 6519
rect 59866 6451 59874 6485
rect 59832 6417 59874 6451
rect 59866 6383 59874 6417
rect 59303 6349 59342 6374
rect 58854 6297 58870 6331
rect 58904 6297 58920 6331
rect 59060 6310 59342 6349
rect 59832 6341 59874 6383
rect 59228 6308 59342 6310
rect 59500 6297 59516 6331
rect 59550 6297 59566 6331
rect 59666 6307 59695 6341
rect 59729 6307 59787 6341
rect 59821 6307 59879 6341
rect 59913 6307 59942 6341
rect 59833 6300 59867 6307
rect 58920 6212 58966 6218
rect 58920 6210 59408 6212
rect 58920 6176 58928 6210
rect 58962 6193 59408 6210
rect 58962 6188 59358 6193
rect 58962 6178 59237 6188
rect 58962 6176 58966 6178
rect 58920 6174 58966 6176
rect 59138 6154 59237 6178
rect 59271 6159 59358 6188
rect 59392 6168 59408 6193
rect 59392 6159 59533 6168
rect 59271 6154 59533 6159
rect 59138 6134 59533 6154
rect 59262 6050 59278 6084
rect 59312 6050 59448 6084
rect 58786 6000 59168 6016
rect 58786 5976 59134 6000
rect 59134 5930 59168 5964
rect 59134 5878 59168 5894
rect 59230 6000 59264 6016
rect 59230 5930 59264 5964
rect 59230 5878 59264 5894
rect 59326 6000 59360 6016
rect 59326 5930 59360 5964
rect 59326 5878 59360 5894
rect 57600 5797 57629 5831
rect 57663 5797 57721 5831
rect 57755 5797 57813 5831
rect 57847 5797 57876 5831
rect 58674 5797 58703 5831
rect 58737 5797 58795 5831
rect 58829 5797 58887 5831
rect 58921 5797 58950 5831
rect 59166 5810 59182 5844
rect 59216 5810 59232 5844
rect 57619 5753 57673 5797
rect 57619 5719 57639 5753
rect 57619 5685 57673 5719
rect 57619 5651 57639 5685
rect 57619 5635 57673 5651
rect 57707 5753 57773 5763
rect 57707 5719 57723 5753
rect 57757 5719 57773 5753
rect 57707 5710 57773 5719
rect 57707 5685 57725 5710
rect 57707 5651 57723 5685
rect 57759 5676 57773 5710
rect 57757 5651 57773 5676
rect 57707 5635 57773 5651
rect 57807 5753 57855 5797
rect 57841 5719 57855 5753
rect 57807 5685 57855 5719
rect 57841 5651 57855 5685
rect 57807 5635 57855 5651
rect 58693 5753 58747 5797
rect 58693 5719 58713 5753
rect 58693 5685 58747 5719
rect 58693 5651 58713 5685
rect 58693 5635 58747 5651
rect 58781 5753 58847 5763
rect 58781 5719 58797 5753
rect 58831 5719 58847 5753
rect 58781 5715 58847 5719
rect 58781 5681 58795 5715
rect 58829 5685 58847 5715
rect 58781 5651 58797 5681
rect 58831 5651 58847 5685
rect 58781 5635 58847 5651
rect 58881 5753 58929 5797
rect 58915 5719 58929 5753
rect 59278 5729 59294 5763
rect 59328 5729 59344 5763
rect 58881 5685 58929 5719
rect 58915 5651 58929 5685
rect 58881 5635 58929 5651
rect 59150 5667 59184 5686
rect 57617 5594 57637 5599
rect 57617 5560 57634 5594
rect 57671 5565 57687 5599
rect 57668 5560 57687 5565
rect 57617 5549 57687 5560
rect 57721 5515 57755 5635
rect 57789 5565 57805 5599
rect 57839 5590 57859 5599
rect 57789 5556 57807 5565
rect 57841 5556 57859 5590
rect 57789 5549 57859 5556
rect 58691 5592 58711 5599
rect 58691 5558 58709 5592
rect 58745 5565 58761 5599
rect 58743 5558 58761 5565
rect 58691 5549 58761 5558
rect 58795 5515 58829 5635
rect 59150 5599 59184 5601
rect 58863 5565 58879 5599
rect 58913 5592 58933 5599
rect 58863 5558 58883 5565
rect 58917 5558 58933 5592
rect 58863 5549 58933 5558
rect 59150 5563 59184 5565
rect 57294 5435 57560 5436
rect 57294 5401 57310 5435
rect 57344 5401 57560 5435
rect 57294 5400 57560 5401
rect 57619 5499 57685 5515
rect 57619 5465 57651 5499
rect 57721 5499 57857 5515
rect 57721 5481 57807 5499
rect 57619 5431 57685 5465
rect 56977 5363 57043 5397
rect 56977 5329 56993 5363
rect 57027 5329 57043 5363
rect 57619 5397 57651 5431
rect 57619 5363 57685 5397
rect 56977 5324 57043 5329
rect 57170 5329 57452 5362
rect 57170 5295 57260 5329
rect 57294 5327 57452 5329
rect 57294 5295 57379 5327
rect 57170 5293 57379 5295
rect 57413 5293 57452 5327
rect 57170 5287 57452 5293
rect 57619 5329 57651 5363
rect 57619 5287 57685 5329
rect 57791 5465 57807 5481
rect 57841 5465 57857 5499
rect 57791 5431 57857 5465
rect 57791 5397 57807 5431
rect 57841 5397 57857 5431
rect 57791 5363 57857 5397
rect 57791 5329 57807 5363
rect 57841 5329 57857 5363
rect 57791 5324 57857 5329
rect 58693 5499 58759 5515
rect 58693 5465 58725 5499
rect 58795 5499 58931 5515
rect 58795 5481 58881 5499
rect 58693 5431 58759 5465
rect 58693 5397 58725 5431
rect 58693 5363 58759 5397
rect 58693 5329 58725 5363
rect 58693 5287 58759 5329
rect 58865 5465 58881 5481
rect 58915 5465 58931 5499
rect 59150 5478 59184 5497
rect 59246 5667 59280 5686
rect 59246 5599 59280 5601
rect 59246 5563 59280 5565
rect 59246 5478 59280 5497
rect 59342 5667 59376 5686
rect 59342 5599 59376 5601
rect 59342 5563 59376 5565
rect 59342 5478 59376 5497
rect 58865 5431 58931 5465
rect 58865 5397 58881 5431
rect 58915 5397 58931 5431
rect 59182 5436 59248 5438
rect 59414 5436 59448 6050
rect 59499 5831 59533 6134
rect 59730 5831 59764 6042
rect 59488 5797 59517 5831
rect 59551 5797 59609 5831
rect 59643 5797 59701 5831
rect 59735 5797 59764 5831
rect 59507 5753 59561 5797
rect 59507 5719 59527 5753
rect 59507 5685 59561 5719
rect 59507 5651 59527 5685
rect 59507 5635 59561 5651
rect 59595 5753 59661 5763
rect 59595 5719 59611 5753
rect 59645 5719 59661 5753
rect 59595 5710 59661 5719
rect 59595 5685 59613 5710
rect 59595 5651 59611 5685
rect 59647 5676 59661 5710
rect 59645 5651 59661 5676
rect 59595 5635 59661 5651
rect 59695 5753 59743 5797
rect 59729 5719 59743 5753
rect 59695 5685 59743 5719
rect 59729 5651 59743 5685
rect 59695 5635 59743 5651
rect 59505 5594 59525 5599
rect 59505 5560 59522 5594
rect 59559 5565 59575 5599
rect 59556 5560 59575 5565
rect 59505 5549 59575 5560
rect 59609 5515 59643 5635
rect 59677 5565 59693 5599
rect 59727 5590 59747 5599
rect 59677 5556 59695 5565
rect 59729 5556 59747 5590
rect 59677 5549 59747 5556
rect 59182 5435 59448 5436
rect 59182 5401 59198 5435
rect 59232 5401 59448 5435
rect 59182 5400 59448 5401
rect 59507 5499 59573 5515
rect 59507 5465 59539 5499
rect 59609 5499 59745 5515
rect 59609 5481 59695 5499
rect 59507 5431 59573 5465
rect 58865 5363 58931 5397
rect 58865 5329 58881 5363
rect 58915 5329 58931 5363
rect 59507 5397 59539 5431
rect 59507 5363 59573 5397
rect 58865 5324 58931 5329
rect 59058 5329 59340 5362
rect 59058 5295 59148 5329
rect 59182 5327 59340 5329
rect 59182 5295 59267 5327
rect 59058 5293 59267 5295
rect 59301 5293 59340 5327
rect 59058 5287 59340 5293
rect 59507 5329 59539 5363
rect 59507 5287 59573 5329
rect 59679 5465 59695 5481
rect 59729 5465 59745 5499
rect 59679 5431 59745 5465
rect 59679 5397 59695 5431
rect 59729 5397 59745 5431
rect 59679 5363 59745 5397
rect 59679 5329 59695 5363
rect 59729 5329 59745 5363
rect 59679 5324 59745 5329
rect 158 5253 187 5287
rect 221 5253 279 5287
rect 313 5253 371 5287
rect 405 5253 1001 5287
rect 1035 5253 1093 5287
rect 1127 5253 1185 5287
rect 1219 5286 1248 5287
rect 1219 5253 1290 5286
rect 2046 5253 2075 5287
rect 2109 5253 2167 5287
rect 2201 5253 2259 5287
rect 2293 5253 2889 5287
rect 2923 5253 2981 5287
rect 3015 5253 3073 5287
rect 3107 5286 3136 5287
rect 3107 5253 3178 5286
rect 3934 5253 3963 5287
rect 3997 5253 4055 5287
rect 4089 5253 4147 5287
rect 4181 5253 4777 5287
rect 4811 5253 4869 5287
rect 4903 5253 4961 5287
rect 4995 5286 5024 5287
rect 4995 5253 5066 5286
rect 5822 5253 5851 5287
rect 5885 5253 5943 5287
rect 5977 5253 6035 5287
rect 6069 5253 6665 5287
rect 6699 5253 6757 5287
rect 6791 5253 6849 5287
rect 6883 5286 6912 5287
rect 6883 5253 6954 5286
rect 7710 5253 7739 5287
rect 7773 5253 7831 5287
rect 7865 5253 7923 5287
rect 7957 5253 8553 5287
rect 8587 5253 8645 5287
rect 8679 5253 8737 5287
rect 8771 5286 8800 5287
rect 8771 5253 8842 5286
rect 9598 5253 9627 5287
rect 9661 5253 9719 5287
rect 9753 5253 9811 5287
rect 9845 5253 10441 5287
rect 10475 5253 10533 5287
rect 10567 5253 10625 5287
rect 10659 5286 10688 5287
rect 10659 5253 10730 5286
rect 11486 5253 11515 5287
rect 11549 5253 11607 5287
rect 11641 5253 11699 5287
rect 11733 5253 12329 5287
rect 12363 5253 12421 5287
rect 12455 5253 12513 5287
rect 12547 5286 12576 5287
rect 12547 5253 12618 5286
rect 13374 5253 13403 5287
rect 13437 5253 13495 5287
rect 13529 5253 13587 5287
rect 13621 5253 14217 5287
rect 14251 5253 14309 5287
rect 14343 5253 14401 5287
rect 14435 5286 14464 5287
rect 14435 5253 14506 5286
rect 15256 5253 15285 5287
rect 15319 5253 15377 5287
rect 15411 5253 15469 5287
rect 15503 5253 16099 5287
rect 16133 5253 16191 5287
rect 16225 5253 16283 5287
rect 16317 5286 16346 5287
rect 16317 5253 16388 5286
rect 17144 5253 17173 5287
rect 17207 5253 17265 5287
rect 17299 5253 17357 5287
rect 17391 5253 17987 5287
rect 18021 5253 18079 5287
rect 18113 5253 18171 5287
rect 18205 5286 18234 5287
rect 18205 5253 18276 5286
rect 19032 5253 19061 5287
rect 19095 5253 19153 5287
rect 19187 5253 19245 5287
rect 19279 5253 19875 5287
rect 19909 5253 19967 5287
rect 20001 5253 20059 5287
rect 20093 5286 20122 5287
rect 20093 5253 20164 5286
rect 20920 5253 20949 5287
rect 20983 5253 21041 5287
rect 21075 5253 21133 5287
rect 21167 5253 21763 5287
rect 21797 5253 21855 5287
rect 21889 5253 21947 5287
rect 21981 5286 22010 5287
rect 21981 5253 22052 5286
rect 22808 5253 22837 5287
rect 22871 5253 22929 5287
rect 22963 5253 23021 5287
rect 23055 5253 23651 5287
rect 23685 5253 23743 5287
rect 23777 5253 23835 5287
rect 23869 5286 23898 5287
rect 23869 5253 23940 5286
rect 24696 5253 24725 5287
rect 24759 5253 24817 5287
rect 24851 5253 24909 5287
rect 24943 5253 25539 5287
rect 25573 5253 25631 5287
rect 25665 5253 25723 5287
rect 25757 5286 25786 5287
rect 25757 5253 25828 5286
rect 26584 5253 26613 5287
rect 26647 5253 26705 5287
rect 26739 5253 26797 5287
rect 26831 5253 27427 5287
rect 27461 5253 27519 5287
rect 27553 5253 27611 5287
rect 27645 5286 27674 5287
rect 27645 5253 27716 5286
rect 28472 5253 28501 5287
rect 28535 5253 28593 5287
rect 28627 5253 28685 5287
rect 28719 5253 29315 5287
rect 29349 5253 29407 5287
rect 29441 5253 29499 5287
rect 29533 5286 29562 5287
rect 29533 5253 29604 5286
rect 30360 5253 30389 5287
rect 30423 5253 30481 5287
rect 30515 5253 30573 5287
rect 30607 5253 31203 5287
rect 31237 5253 31295 5287
rect 31329 5253 31387 5287
rect 31421 5286 31450 5287
rect 31421 5253 31492 5286
rect 32248 5253 32277 5287
rect 32311 5253 32369 5287
rect 32403 5253 32461 5287
rect 32495 5253 33091 5287
rect 33125 5253 33183 5287
rect 33217 5253 33275 5287
rect 33309 5286 33338 5287
rect 33309 5253 33380 5286
rect 34136 5253 34165 5287
rect 34199 5253 34257 5287
rect 34291 5253 34349 5287
rect 34383 5253 34979 5287
rect 35013 5253 35071 5287
rect 35105 5253 35163 5287
rect 35197 5286 35226 5287
rect 35197 5253 35268 5286
rect 36024 5253 36053 5287
rect 36087 5253 36145 5287
rect 36179 5253 36237 5287
rect 36271 5253 36867 5287
rect 36901 5253 36959 5287
rect 36993 5253 37051 5287
rect 37085 5286 37114 5287
rect 37085 5253 37156 5286
rect 37912 5253 37941 5287
rect 37975 5253 38033 5287
rect 38067 5253 38125 5287
rect 38159 5253 38755 5287
rect 38789 5253 38847 5287
rect 38881 5253 38939 5287
rect 38973 5286 39002 5287
rect 38973 5253 39044 5286
rect 39800 5253 39829 5287
rect 39863 5253 39921 5287
rect 39955 5253 40013 5287
rect 40047 5253 40643 5287
rect 40677 5253 40735 5287
rect 40769 5253 40827 5287
rect 40861 5286 40890 5287
rect 40861 5253 40932 5286
rect 41688 5253 41717 5287
rect 41751 5253 41809 5287
rect 41843 5253 41901 5287
rect 41935 5253 42531 5287
rect 42565 5253 42623 5287
rect 42657 5253 42715 5287
rect 42749 5286 42778 5287
rect 42749 5253 42820 5286
rect 43576 5253 43605 5287
rect 43639 5253 43697 5287
rect 43731 5253 43789 5287
rect 43823 5253 44419 5287
rect 44453 5253 44511 5287
rect 44545 5253 44603 5287
rect 44637 5286 44666 5287
rect 44637 5253 44708 5286
rect 45458 5253 45487 5287
rect 45521 5253 45579 5287
rect 45613 5253 45671 5287
rect 45705 5253 46301 5287
rect 46335 5253 46393 5287
rect 46427 5253 46485 5287
rect 46519 5286 46548 5287
rect 46519 5253 46590 5286
rect 47346 5253 47375 5287
rect 47409 5253 47467 5287
rect 47501 5253 47559 5287
rect 47593 5253 48189 5287
rect 48223 5253 48281 5287
rect 48315 5253 48373 5287
rect 48407 5286 48436 5287
rect 48407 5253 48478 5286
rect 49234 5253 49263 5287
rect 49297 5253 49355 5287
rect 49389 5253 49447 5287
rect 49481 5253 50077 5287
rect 50111 5253 50169 5287
rect 50203 5253 50261 5287
rect 50295 5286 50324 5287
rect 50295 5253 50366 5286
rect 51122 5253 51151 5287
rect 51185 5253 51243 5287
rect 51277 5253 51335 5287
rect 51369 5253 51965 5287
rect 51999 5253 52057 5287
rect 52091 5253 52149 5287
rect 52183 5286 52212 5287
rect 52183 5253 52254 5286
rect 53010 5253 53039 5287
rect 53073 5253 53131 5287
rect 53165 5253 53223 5287
rect 53257 5253 53853 5287
rect 53887 5253 53945 5287
rect 53979 5253 54037 5287
rect 54071 5286 54100 5287
rect 54071 5253 54142 5286
rect 54898 5253 54927 5287
rect 54961 5253 55019 5287
rect 55053 5253 55111 5287
rect 55145 5253 55741 5287
rect 55775 5253 55833 5287
rect 55867 5253 55925 5287
rect 55959 5286 55988 5287
rect 55959 5253 56030 5286
rect 56786 5253 56815 5287
rect 56849 5253 56907 5287
rect 56941 5253 56999 5287
rect 57033 5253 57629 5287
rect 57663 5253 57721 5287
rect 57755 5253 57813 5287
rect 57847 5286 57876 5287
rect 57847 5253 57918 5286
rect 58674 5253 58703 5287
rect 58737 5253 58795 5287
rect 58829 5253 58887 5287
rect 58921 5253 59517 5287
rect 59551 5253 59609 5287
rect 59643 5253 59701 5287
rect 59735 5286 59764 5287
rect 59735 5253 59806 5286
rect 434 5252 824 5253
rect 1228 5252 1290 5253
rect 2322 5252 2712 5253
rect 3116 5252 3178 5253
rect 4210 5252 4600 5253
rect 5004 5252 5066 5253
rect 6098 5252 6488 5253
rect 6892 5252 6954 5253
rect 7986 5252 8376 5253
rect 8780 5252 8842 5253
rect 9874 5252 10264 5253
rect 10668 5252 10730 5253
rect 11762 5252 12152 5253
rect 12556 5252 12618 5253
rect 13650 5252 14040 5253
rect 14444 5252 14506 5253
rect 15532 5252 15922 5253
rect 16326 5252 16388 5253
rect 17420 5252 17810 5253
rect 18214 5252 18276 5253
rect 19308 5252 19698 5253
rect 20102 5252 20164 5253
rect 21196 5252 21586 5253
rect 21990 5252 22052 5253
rect 23084 5252 23474 5253
rect 23878 5252 23940 5253
rect 24972 5252 25362 5253
rect 25766 5252 25828 5253
rect 26860 5252 27250 5253
rect 27654 5252 27716 5253
rect 28748 5252 29138 5253
rect 29542 5252 29604 5253
rect 30636 5252 31026 5253
rect 31430 5252 31492 5253
rect 32524 5252 32914 5253
rect 33318 5252 33380 5253
rect 34412 5252 34802 5253
rect 35206 5252 35268 5253
rect 36300 5252 36690 5253
rect 37094 5252 37156 5253
rect 38188 5252 38578 5253
rect 38982 5252 39044 5253
rect 40076 5252 40466 5253
rect 40870 5252 40932 5253
rect 41964 5252 42354 5253
rect 42758 5252 42820 5253
rect 43852 5252 44242 5253
rect 44646 5252 44708 5253
rect 45734 5252 46124 5253
rect 46528 5252 46590 5253
rect 47622 5252 48012 5253
rect 48416 5252 48478 5253
rect 49510 5252 49900 5253
rect 50304 5252 50366 5253
rect 51398 5252 51788 5253
rect 52192 5252 52254 5253
rect 53286 5252 53676 5253
rect 54080 5252 54142 5253
rect 55174 5252 55564 5253
rect 55968 5252 56030 5253
rect 57062 5252 57452 5253
rect 57856 5252 57918 5253
rect 58950 5252 59340 5253
rect 59744 5252 59806 5253
rect 5664 5175 5693 5209
rect 5727 5175 5785 5209
rect 5819 5175 5877 5209
rect 5911 5175 5969 5209
rect 6003 5175 6061 5209
rect 6095 5175 6153 5209
rect 6187 5175 6245 5209
rect 6279 5175 6337 5209
rect 6371 5175 6429 5209
rect 6463 5175 6521 5209
rect 6555 5175 6613 5209
rect 6647 5175 6705 5209
rect 6739 5175 6797 5209
rect 6831 5175 6889 5209
rect 6923 5175 6981 5209
rect 7015 5175 7073 5209
rect 7107 5175 7136 5209
rect 5702 5133 5744 5175
rect 5702 5099 5710 5133
rect 5702 5065 5744 5099
rect 5702 5031 5710 5065
rect 5702 5015 5744 5031
rect 5778 5133 5844 5141
rect 5778 5099 5794 5133
rect 5828 5099 5844 5133
rect 5778 5065 5844 5099
rect 5778 5031 5794 5065
rect 5828 5031 5844 5065
rect 5778 5005 5844 5031
rect 5878 5133 5912 5175
rect 5878 5065 5912 5099
rect 5878 5015 5912 5031
rect 5946 5133 6012 5141
rect 5946 5099 5962 5133
rect 5996 5099 6012 5133
rect 5946 5065 6012 5099
rect 5946 5031 5962 5065
rect 5996 5031 6012 5065
rect 5778 4995 5799 5005
rect 5778 4961 5794 4995
rect 5833 4981 5844 5005
rect 5946 5009 6012 5031
rect 6046 5133 6080 5175
rect 6046 5065 6080 5099
rect 6046 5015 6080 5031
rect 6114 5133 6180 5141
rect 6114 5099 6130 5133
rect 6164 5099 6180 5133
rect 6114 5065 6180 5099
rect 6114 5031 6130 5065
rect 6164 5031 6180 5065
rect 5946 4981 5962 5009
rect 5833 4971 5962 4981
rect 5996 4981 6012 5009
rect 6114 5007 6180 5031
rect 6214 5133 6248 5175
rect 6214 5065 6248 5099
rect 6214 5015 6248 5031
rect 6282 5133 6348 5141
rect 6282 5099 6298 5133
rect 6332 5099 6348 5133
rect 6282 5065 6348 5099
rect 6282 5031 6298 5065
rect 6332 5031 6348 5065
rect 6114 4995 6132 5007
rect 6114 4981 6130 4995
rect 5828 4961 5962 4971
rect 5996 4961 6130 4981
rect 6166 4981 6180 5007
rect 6282 5007 6348 5031
rect 6382 5133 6416 5175
rect 6382 5065 6416 5099
rect 6382 5015 6416 5031
rect 6450 5133 6516 5141
rect 6450 5099 6466 5133
rect 6500 5099 6516 5133
rect 6450 5065 6516 5099
rect 6450 5031 6466 5065
rect 6500 5031 6516 5065
rect 6282 4981 6297 5007
rect 6331 4995 6348 5007
rect 6166 4973 6297 4981
rect 6332 4981 6348 4995
rect 6450 4995 6516 5031
rect 6550 5133 6584 5175
rect 6550 5065 6584 5099
rect 6550 5015 6584 5031
rect 6618 5133 6684 5141
rect 6618 5099 6634 5133
rect 6668 5099 6684 5133
rect 6618 5065 6684 5099
rect 6618 5031 6634 5065
rect 6668 5031 6684 5065
rect 6450 4981 6466 4995
rect 6164 4961 6298 4973
rect 6332 4961 6466 4981
rect 6500 4981 6516 4995
rect 6618 4996 6684 5031
rect 6718 5133 6752 5175
rect 6718 5065 6752 5099
rect 6718 5015 6752 5031
rect 6786 5133 6852 5141
rect 6786 5099 6802 5133
rect 6836 5099 6852 5133
rect 6786 5065 6852 5099
rect 6786 5031 6802 5065
rect 6836 5031 6852 5065
rect 6618 4995 6637 4996
rect 6618 4981 6634 4995
rect 6500 4961 6634 4981
rect 6671 4981 6684 4996
rect 6786 5001 6852 5031
rect 6886 5133 6920 5175
rect 6886 5065 6920 5099
rect 6886 5015 6920 5031
rect 6954 5133 7020 5141
rect 6954 5099 6970 5133
rect 7004 5099 7020 5133
rect 6954 5065 7020 5099
rect 6954 5031 6970 5065
rect 7004 5031 7020 5065
rect 6786 4981 6799 5001
rect 6833 4995 6852 5001
rect 6671 4967 6799 4981
rect 6836 4981 6852 4995
rect 6954 5002 7020 5031
rect 6954 4995 6972 5002
rect 6954 4981 6970 4995
rect 6671 4962 6802 4967
rect 6668 4961 6802 4962
rect 6836 4961 6970 4981
rect 7006 4968 7020 5002
rect 7004 4961 7020 4968
rect 5778 4959 6466 4961
rect 6500 4959 7020 4961
rect 5778 4947 7020 4959
rect 7054 5133 7096 5175
rect 7546 5173 7575 5207
rect 7609 5173 7667 5207
rect 7701 5173 7759 5207
rect 7793 5173 7851 5207
rect 7885 5173 7943 5207
rect 7977 5173 8035 5207
rect 8069 5173 8127 5207
rect 8161 5173 8219 5207
rect 8253 5173 8311 5207
rect 8345 5173 8403 5207
rect 8437 5173 8495 5207
rect 8529 5173 8587 5207
rect 8621 5173 8679 5207
rect 8713 5173 8771 5207
rect 8805 5173 8863 5207
rect 8897 5173 8955 5207
rect 8989 5173 9018 5207
rect 20762 5175 20791 5209
rect 20825 5175 20883 5209
rect 20917 5175 20975 5209
rect 21009 5175 21067 5209
rect 21101 5175 21159 5209
rect 21193 5175 21251 5209
rect 21285 5175 21343 5209
rect 21377 5175 21435 5209
rect 21469 5175 21527 5209
rect 21561 5175 21619 5209
rect 21653 5175 21711 5209
rect 21745 5175 21803 5209
rect 21837 5175 21895 5209
rect 21929 5175 21987 5209
rect 22021 5175 22079 5209
rect 22113 5175 22171 5209
rect 22205 5175 22234 5209
rect 7088 5099 7096 5133
rect 7054 5065 7096 5099
rect 7088 5031 7096 5065
rect 7054 4995 7096 5031
rect 7584 5131 7626 5173
rect 7584 5097 7592 5131
rect 7584 5063 7626 5097
rect 7584 5029 7592 5063
rect 7584 5013 7626 5029
rect 7660 5131 7726 5139
rect 7660 5097 7676 5131
rect 7710 5097 7726 5131
rect 7660 5063 7726 5097
rect 7660 5029 7676 5063
rect 7710 5029 7726 5063
rect 7088 4961 7096 4995
rect 5778 4829 5844 4947
rect 7054 4945 7096 4961
rect 7660 4993 7726 5029
rect 7760 5131 7794 5173
rect 7760 5063 7794 5097
rect 7760 5013 7794 5029
rect 7828 5131 7894 5139
rect 7828 5097 7844 5131
rect 7878 5097 7894 5131
rect 7828 5063 7894 5097
rect 7828 5029 7844 5063
rect 7878 5029 7894 5063
rect 7660 4959 7676 4993
rect 7710 4979 7726 4993
rect 7828 5003 7894 5029
rect 7928 5131 7962 5173
rect 7928 5063 7962 5097
rect 7928 5013 7962 5029
rect 7996 5131 8062 5139
rect 7996 5097 8012 5131
rect 8046 5097 8062 5131
rect 7996 5063 8062 5097
rect 7996 5029 8012 5063
rect 8046 5029 8062 5063
rect 7828 4993 7845 5003
rect 7828 4979 7844 4993
rect 7710 4959 7844 4979
rect 7879 4979 7894 5003
rect 7996 5012 8062 5029
rect 8096 5131 8130 5173
rect 8096 5063 8130 5097
rect 8096 5013 8130 5029
rect 8164 5131 8230 5139
rect 8164 5097 8180 5131
rect 8214 5097 8230 5131
rect 8164 5063 8230 5097
rect 8164 5029 8180 5063
rect 8214 5029 8230 5063
rect 7996 4993 8015 5012
rect 7996 4979 8012 4993
rect 7879 4969 8012 4979
rect 8049 4979 8062 5012
rect 8164 5010 8230 5029
rect 8264 5131 8298 5173
rect 8264 5063 8298 5097
rect 8264 5013 8298 5029
rect 8332 5131 8398 5139
rect 8332 5097 8348 5131
rect 8382 5097 8398 5131
rect 8332 5063 8398 5097
rect 8332 5029 8348 5063
rect 8382 5029 8398 5063
rect 8164 4993 8183 5010
rect 8164 4979 8180 4993
rect 8049 4978 8180 4979
rect 7878 4959 8012 4969
rect 8046 4959 8180 4978
rect 8217 4979 8230 5010
rect 8332 4997 8398 5029
rect 8432 5131 8466 5173
rect 8432 5063 8466 5097
rect 8432 5013 8466 5029
rect 8500 5131 8566 5139
rect 8500 5097 8516 5131
rect 8550 5097 8566 5131
rect 8500 5063 8566 5097
rect 8500 5029 8516 5063
rect 8550 5029 8566 5063
rect 8332 4993 8350 4997
rect 8332 4979 8348 4993
rect 8217 4976 8348 4979
rect 8214 4959 8348 4976
rect 8384 4979 8398 4997
rect 8500 5002 8566 5029
rect 8600 5131 8634 5173
rect 8600 5063 8634 5097
rect 8600 5013 8634 5029
rect 8668 5131 8734 5139
rect 8668 5097 8684 5131
rect 8718 5097 8734 5131
rect 8668 5063 8734 5097
rect 8668 5029 8684 5063
rect 8718 5029 8734 5063
rect 8500 4979 8515 5002
rect 8549 4993 8566 5002
rect 8384 4968 8515 4979
rect 8550 4979 8566 4993
rect 8668 5006 8734 5029
rect 8768 5131 8802 5173
rect 8768 5063 8802 5097
rect 8768 5013 8802 5029
rect 8836 5131 8902 5139
rect 8836 5097 8852 5131
rect 8886 5097 8902 5131
rect 8836 5063 8902 5097
rect 8836 5029 8852 5063
rect 8886 5029 8902 5063
rect 8668 4993 8688 5006
rect 8668 4979 8684 4993
rect 8384 4963 8516 4968
rect 8382 4959 8516 4963
rect 8550 4959 8684 4979
rect 8722 4979 8734 5006
rect 8836 5001 8902 5029
rect 8836 4979 8851 5001
rect 8885 4993 8902 5001
rect 8722 4972 8851 4979
rect 8718 4967 8851 4972
rect 8718 4959 8852 4967
rect 8886 4959 8902 4993
rect 7660 4945 8902 4959
rect 8936 5131 8978 5173
rect 8970 5097 8978 5131
rect 8936 5063 8978 5097
rect 8970 5029 8978 5063
rect 8936 4993 8978 5029
rect 20800 5133 20842 5175
rect 20800 5099 20808 5133
rect 20800 5065 20842 5099
rect 20800 5031 20808 5065
rect 20800 5015 20842 5031
rect 20876 5133 20942 5141
rect 20876 5099 20892 5133
rect 20926 5099 20942 5133
rect 20876 5065 20942 5099
rect 20876 5031 20892 5065
rect 20926 5031 20942 5065
rect 8970 4959 8978 4993
rect 6031 4900 7119 4911
rect 6031 4897 6318 4900
rect 6031 4863 6047 4897
rect 6081 4863 6214 4897
rect 6248 4866 6318 4897
rect 6352 4897 6426 4900
rect 6352 4866 6382 4897
rect 6248 4863 6382 4866
rect 6416 4866 6426 4897
rect 6460 4866 6534 4900
rect 6568 4897 6642 4900
rect 6583 4866 6642 4897
rect 6676 4897 6750 4900
rect 6676 4866 6718 4897
rect 6784 4866 6858 4900
rect 6892 4897 6966 4900
rect 6920 4866 6966 4897
rect 7000 4897 7074 4900
rect 7000 4866 7060 4897
rect 7108 4866 7119 4900
rect 6416 4863 6549 4866
rect 6583 4863 6718 4866
rect 6752 4863 6886 4866
rect 6920 4863 7060 4866
rect 7094 4863 7119 4866
rect 5702 4809 5744 4825
rect 5702 4775 5710 4809
rect 5702 4741 5744 4775
rect 5702 4707 5710 4741
rect 5702 4665 5744 4707
rect 5778 4809 7020 4829
rect 7660 4827 7726 4945
rect 8936 4943 8978 4959
rect 20876 4996 20942 5031
rect 20976 5133 21010 5175
rect 20976 5065 21010 5099
rect 20976 5015 21010 5031
rect 21044 5133 21110 5141
rect 21044 5099 21060 5133
rect 21094 5099 21110 5133
rect 21044 5065 21110 5099
rect 21044 5031 21060 5065
rect 21094 5031 21110 5065
rect 20876 4995 20901 4996
rect 20876 4961 20892 4995
rect 20935 4981 20942 4996
rect 21044 4998 21110 5031
rect 21144 5133 21178 5175
rect 21144 5065 21178 5099
rect 21144 5015 21178 5031
rect 21212 5133 21278 5141
rect 21212 5099 21228 5133
rect 21262 5099 21278 5133
rect 21212 5065 21278 5099
rect 21212 5031 21228 5065
rect 21262 5031 21278 5065
rect 21044 4981 21060 4998
rect 20935 4962 21060 4981
rect 21094 4981 21110 4998
rect 21212 5000 21278 5031
rect 21312 5133 21346 5175
rect 21312 5065 21346 5099
rect 21312 5015 21346 5031
rect 21380 5133 21446 5141
rect 21380 5099 21396 5133
rect 21430 5099 21446 5133
rect 21380 5065 21446 5099
rect 21380 5031 21396 5065
rect 21430 5031 21446 5065
rect 21212 4995 21230 5000
rect 21212 4981 21228 4995
rect 20926 4961 21060 4962
rect 21094 4961 21228 4981
rect 21264 4981 21278 5000
rect 21380 5006 21446 5031
rect 21480 5133 21514 5175
rect 21480 5065 21514 5099
rect 21480 5015 21514 5031
rect 21548 5133 21614 5141
rect 21548 5099 21564 5133
rect 21598 5099 21614 5133
rect 21548 5065 21614 5099
rect 21548 5031 21564 5065
rect 21598 5031 21614 5065
rect 21380 4995 21400 5006
rect 21380 4981 21396 4995
rect 21264 4966 21396 4981
rect 21434 4981 21446 5006
rect 21548 4995 21614 5031
rect 21648 5133 21682 5175
rect 21648 5065 21682 5099
rect 21648 5015 21682 5031
rect 21716 5133 21782 5141
rect 21716 5099 21732 5133
rect 21766 5099 21782 5133
rect 21716 5065 21782 5099
rect 21716 5031 21732 5065
rect 21766 5031 21782 5065
rect 21548 4981 21564 4995
rect 21434 4972 21564 4981
rect 21262 4961 21396 4966
rect 21430 4961 21564 4972
rect 21598 4981 21614 4995
rect 21716 5003 21782 5031
rect 21816 5133 21850 5175
rect 21816 5065 21850 5099
rect 21816 5015 21850 5031
rect 21884 5133 21950 5141
rect 21884 5099 21900 5133
rect 21934 5099 21950 5133
rect 21884 5065 21950 5099
rect 21884 5031 21900 5065
rect 21934 5031 21950 5065
rect 21716 4995 21733 5003
rect 21716 4981 21732 4995
rect 21598 4961 21732 4981
rect 21767 4981 21782 5003
rect 21884 4997 21950 5031
rect 21984 5133 22018 5175
rect 21984 5065 22018 5099
rect 21984 5015 22018 5031
rect 22052 5133 22118 5141
rect 22052 5099 22068 5133
rect 22102 5099 22118 5133
rect 22052 5065 22118 5099
rect 22052 5031 22068 5065
rect 22102 5031 22118 5065
rect 21884 4981 21900 4997
rect 21767 4969 21900 4981
rect 21766 4961 21900 4969
rect 21934 4981 21950 4997
rect 22052 4997 22118 5031
rect 22052 4981 22060 4997
rect 22094 4995 22118 4997
rect 21934 4963 22060 4981
rect 21934 4961 22068 4963
rect 22102 4961 22118 4995
rect 20876 4959 21564 4961
rect 21598 4959 22118 4961
rect 20876 4947 22118 4959
rect 22152 5133 22194 5175
rect 22644 5173 22673 5207
rect 22707 5173 22765 5207
rect 22799 5173 22857 5207
rect 22891 5173 22949 5207
rect 22983 5173 23041 5207
rect 23075 5173 23133 5207
rect 23167 5173 23225 5207
rect 23259 5173 23317 5207
rect 23351 5173 23409 5207
rect 23443 5173 23501 5207
rect 23535 5173 23593 5207
rect 23627 5173 23685 5207
rect 23719 5173 23777 5207
rect 23811 5173 23869 5207
rect 23903 5173 23961 5207
rect 23995 5173 24053 5207
rect 24087 5173 24116 5207
rect 35866 5175 35895 5209
rect 35929 5175 35987 5209
rect 36021 5175 36079 5209
rect 36113 5175 36171 5209
rect 36205 5175 36263 5209
rect 36297 5175 36355 5209
rect 36389 5175 36447 5209
rect 36481 5175 36539 5209
rect 36573 5175 36631 5209
rect 36665 5175 36723 5209
rect 36757 5175 36815 5209
rect 36849 5175 36907 5209
rect 36941 5175 36999 5209
rect 37033 5175 37091 5209
rect 37125 5175 37183 5209
rect 37217 5175 37275 5209
rect 37309 5175 37338 5209
rect 22186 5099 22194 5133
rect 22152 5065 22194 5099
rect 22186 5031 22194 5065
rect 22152 4995 22194 5031
rect 22682 5131 22724 5173
rect 22682 5097 22690 5131
rect 22682 5063 22724 5097
rect 22682 5029 22690 5063
rect 22682 5013 22724 5029
rect 22758 5131 22824 5139
rect 22758 5097 22774 5131
rect 22808 5097 22824 5131
rect 22758 5063 22824 5097
rect 22758 5029 22774 5063
rect 22808 5029 22824 5063
rect 22186 4961 22194 4995
rect 7913 4900 9001 4909
rect 7913 4895 7930 4900
rect 7913 4861 7929 4895
rect 7964 4866 8081 4900
rect 8115 4895 8178 4900
rect 8130 4866 8178 4895
rect 8212 4895 8275 4900
rect 8212 4866 8264 4895
rect 8309 4866 8372 4900
rect 8406 4895 8469 4900
rect 8406 4866 8431 4895
rect 7963 4861 8096 4866
rect 8130 4861 8264 4866
rect 8298 4861 8431 4866
rect 8465 4866 8469 4895
rect 8503 4866 8566 4900
rect 8600 4895 8663 4900
rect 8465 4861 8600 4866
rect 8634 4866 8663 4895
rect 8697 4866 8760 4900
rect 8794 4895 9001 4900
rect 8634 4861 8768 4866
rect 8802 4861 8942 4895
rect 8976 4861 9001 4895
rect 20876 4829 20942 4947
rect 22152 4945 22194 4961
rect 22758 4994 22824 5029
rect 22858 5131 22892 5173
rect 22858 5063 22892 5097
rect 22858 5013 22892 5029
rect 22926 5131 22992 5139
rect 22926 5097 22942 5131
rect 22976 5097 22992 5131
rect 22926 5063 22992 5097
rect 22926 5029 22942 5063
rect 22976 5029 22992 5063
rect 22758 4959 22774 4994
rect 22808 4979 22824 4994
rect 22926 4996 22992 5029
rect 23026 5131 23060 5173
rect 23026 5063 23060 5097
rect 23026 5013 23060 5029
rect 23094 5131 23160 5139
rect 23094 5097 23110 5131
rect 23144 5097 23160 5131
rect 23094 5063 23160 5097
rect 23094 5029 23110 5063
rect 23144 5029 23160 5063
rect 22926 4993 22944 4996
rect 22926 4979 22942 4993
rect 22808 4959 22942 4979
rect 22978 4979 22992 4996
rect 23094 5002 23160 5029
rect 23194 5131 23228 5173
rect 23194 5063 23228 5097
rect 23194 5013 23228 5029
rect 23262 5131 23328 5139
rect 23262 5097 23278 5131
rect 23312 5097 23328 5131
rect 23262 5063 23328 5097
rect 23262 5029 23278 5063
rect 23312 5029 23328 5063
rect 23094 4979 23110 5002
rect 22978 4962 23110 4979
rect 23144 4979 23160 5002
rect 23262 5001 23328 5029
rect 23362 5131 23396 5173
rect 23362 5063 23396 5097
rect 23362 5013 23396 5029
rect 23430 5131 23496 5139
rect 23430 5097 23446 5131
rect 23480 5097 23496 5131
rect 23430 5063 23496 5097
rect 23430 5029 23446 5063
rect 23480 5029 23496 5063
rect 23262 4993 23279 5001
rect 23262 4979 23278 4993
rect 22976 4959 23110 4962
rect 23144 4959 23278 4979
rect 23313 4979 23328 5001
rect 23430 4997 23496 5029
rect 23530 5131 23564 5173
rect 23530 5063 23564 5097
rect 23530 5013 23564 5029
rect 23598 5131 23664 5139
rect 23598 5097 23614 5131
rect 23648 5097 23664 5131
rect 23598 5063 23664 5097
rect 23598 5029 23614 5063
rect 23648 5029 23664 5063
rect 23430 4993 23448 4997
rect 23430 4979 23446 4993
rect 23313 4967 23446 4979
rect 23312 4959 23446 4967
rect 23482 4979 23496 4997
rect 23598 4999 23664 5029
rect 23698 5131 23732 5173
rect 23698 5063 23732 5097
rect 23698 5013 23732 5029
rect 23766 5131 23832 5139
rect 23766 5097 23782 5131
rect 23816 5097 23832 5131
rect 23766 5063 23832 5097
rect 23766 5029 23782 5063
rect 23816 5029 23832 5063
rect 23598 4993 23619 4999
rect 23598 4979 23614 4993
rect 23482 4963 23614 4979
rect 23653 4979 23664 4999
rect 23766 4997 23832 5029
rect 23866 5131 23900 5173
rect 23866 5063 23900 5097
rect 23866 5013 23900 5029
rect 23934 5131 24000 5139
rect 23934 5097 23950 5131
rect 23984 5097 24000 5131
rect 23934 5063 24000 5097
rect 23934 5029 23950 5063
rect 23984 5029 24000 5063
rect 23766 4993 23783 4997
rect 23766 4979 23782 4993
rect 23653 4965 23782 4979
rect 23480 4959 23614 4963
rect 23648 4959 23782 4965
rect 23817 4979 23832 4997
rect 23934 4995 24000 5029
rect 23934 4979 23949 4995
rect 23983 4993 24000 4995
rect 23817 4963 23949 4979
rect 23816 4961 23949 4963
rect 23816 4959 23950 4961
rect 23984 4959 24000 4993
rect 22758 4945 24000 4959
rect 24034 5131 24076 5173
rect 24068 5097 24076 5131
rect 24034 5063 24076 5097
rect 24068 5029 24076 5063
rect 24034 4993 24076 5029
rect 35904 5133 35946 5175
rect 35904 5099 35912 5133
rect 35904 5065 35946 5099
rect 35904 5031 35912 5065
rect 35904 5015 35946 5031
rect 35980 5133 36046 5141
rect 35980 5099 35996 5133
rect 36030 5099 36046 5133
rect 35980 5065 36046 5099
rect 35980 5031 35996 5065
rect 36030 5031 36046 5065
rect 24068 4959 24076 4993
rect 21129 4900 22217 4911
rect 21129 4897 21458 4900
rect 21492 4897 21577 4900
rect 21129 4863 21145 4897
rect 21179 4863 21312 4897
rect 21346 4866 21458 4897
rect 21514 4866 21577 4897
rect 21611 4897 21696 4900
rect 21611 4866 21647 4897
rect 21346 4863 21480 4866
rect 21514 4863 21647 4866
rect 21681 4866 21696 4897
rect 21730 4866 21815 4900
rect 21849 4897 21934 4900
rect 21850 4866 21934 4897
rect 21968 4897 22053 4900
rect 21968 4866 21984 4897
rect 21681 4863 21816 4866
rect 21850 4863 21984 4866
rect 22018 4866 22053 4897
rect 22087 4897 22172 4900
rect 22087 4866 22158 4897
rect 22206 4866 22217 4900
rect 22018 4863 22158 4866
rect 22192 4863 22217 4866
rect 5778 4775 5794 4809
rect 5828 4791 5962 4809
rect 5828 4775 5844 4791
rect 5778 4741 5844 4775
rect 5946 4775 5962 4791
rect 5996 4791 6130 4809
rect 5996 4775 6012 4791
rect 5778 4707 5794 4741
rect 5828 4707 5844 4741
rect 5778 4699 5844 4707
rect 5878 4741 5912 4757
rect 5878 4665 5912 4707
rect 5946 4741 6012 4775
rect 6114 4775 6130 4791
rect 6164 4791 6298 4809
rect 6164 4775 6180 4791
rect 5946 4707 5962 4741
rect 5996 4707 6012 4741
rect 5946 4699 6012 4707
rect 6046 4741 6080 4757
rect 6046 4665 6080 4707
rect 6114 4741 6180 4775
rect 6282 4775 6298 4791
rect 6332 4791 6466 4809
rect 6332 4775 6348 4791
rect 6114 4707 6130 4741
rect 6164 4707 6180 4741
rect 6114 4699 6180 4707
rect 6214 4741 6248 4757
rect 6214 4665 6248 4707
rect 6282 4741 6348 4775
rect 6450 4775 6466 4791
rect 6500 4791 6634 4809
rect 6500 4775 6516 4791
rect 6282 4707 6298 4741
rect 6332 4707 6348 4741
rect 6282 4699 6348 4707
rect 6382 4741 6416 4757
rect 6382 4665 6416 4707
rect 6450 4741 6516 4775
rect 6618 4775 6634 4791
rect 6668 4791 6802 4809
rect 6668 4775 6684 4791
rect 6450 4707 6466 4741
rect 6500 4707 6516 4741
rect 6450 4699 6516 4707
rect 6550 4741 6584 4757
rect 6550 4665 6584 4707
rect 6618 4741 6684 4775
rect 6786 4775 6802 4791
rect 6836 4791 6970 4809
rect 6836 4775 6852 4791
rect 6618 4707 6634 4741
rect 6668 4707 6684 4741
rect 6618 4699 6684 4707
rect 6718 4741 6752 4757
rect 6718 4665 6752 4707
rect 6786 4741 6852 4775
rect 6954 4775 6970 4791
rect 7004 4775 7020 4809
rect 6786 4707 6802 4741
rect 6836 4707 6852 4741
rect 6786 4699 6852 4707
rect 6886 4741 6920 4757
rect 6886 4665 6920 4707
rect 6954 4741 7020 4775
rect 6954 4707 6970 4741
rect 7004 4707 7020 4741
rect 6954 4699 7020 4707
rect 7054 4809 7100 4825
rect 7088 4775 7100 4809
rect 7054 4741 7100 4775
rect 7088 4707 7100 4741
rect 7054 4665 7100 4707
rect 7584 4807 7626 4823
rect 7584 4773 7592 4807
rect 7584 4739 7626 4773
rect 7584 4705 7592 4739
rect 5664 4631 5693 4665
rect 5727 4631 5785 4665
rect 5819 4631 5877 4665
rect 5911 4631 5969 4665
rect 6003 4631 6061 4665
rect 6095 4631 6153 4665
rect 6187 4631 6245 4665
rect 6279 4631 6337 4665
rect 6371 4631 6429 4665
rect 6463 4631 6521 4665
rect 6555 4631 6613 4665
rect 6647 4631 6705 4665
rect 6739 4631 6797 4665
rect 6831 4631 6889 4665
rect 6923 4631 6981 4665
rect 7015 4631 7073 4665
rect 7107 4631 7136 4665
rect 7584 4663 7626 4705
rect 7660 4807 8902 4827
rect 7660 4773 7676 4807
rect 7710 4789 7844 4807
rect 7710 4773 7726 4789
rect 7660 4739 7726 4773
rect 7828 4773 7844 4789
rect 7878 4789 8012 4807
rect 7878 4773 7894 4789
rect 7660 4705 7676 4739
rect 7710 4705 7726 4739
rect 7660 4697 7726 4705
rect 7760 4739 7794 4755
rect 7760 4663 7794 4705
rect 7828 4739 7894 4773
rect 7996 4773 8012 4789
rect 8046 4789 8180 4807
rect 8046 4773 8062 4789
rect 7828 4705 7844 4739
rect 7878 4705 7894 4739
rect 7828 4697 7894 4705
rect 7928 4739 7962 4755
rect 7928 4663 7962 4705
rect 7996 4739 8062 4773
rect 8164 4773 8180 4789
rect 8214 4789 8348 4807
rect 8214 4773 8230 4789
rect 7996 4705 8012 4739
rect 8046 4705 8062 4739
rect 7996 4697 8062 4705
rect 8096 4739 8130 4755
rect 8096 4663 8130 4705
rect 8164 4739 8230 4773
rect 8332 4773 8348 4789
rect 8382 4789 8516 4807
rect 8382 4773 8398 4789
rect 8164 4705 8180 4739
rect 8214 4705 8230 4739
rect 8164 4697 8230 4705
rect 8264 4739 8298 4755
rect 8264 4663 8298 4705
rect 8332 4739 8398 4773
rect 8500 4773 8516 4789
rect 8550 4789 8684 4807
rect 8550 4773 8566 4789
rect 8332 4705 8348 4739
rect 8382 4705 8398 4739
rect 8332 4697 8398 4705
rect 8432 4739 8466 4755
rect 8432 4663 8466 4705
rect 8500 4739 8566 4773
rect 8668 4773 8684 4789
rect 8718 4789 8852 4807
rect 8718 4773 8734 4789
rect 8500 4705 8516 4739
rect 8550 4705 8566 4739
rect 8500 4697 8566 4705
rect 8600 4739 8634 4755
rect 8600 4663 8634 4705
rect 8668 4739 8734 4773
rect 8836 4773 8852 4789
rect 8886 4773 8902 4807
rect 8668 4705 8684 4739
rect 8718 4705 8734 4739
rect 8668 4697 8734 4705
rect 8768 4739 8802 4755
rect 8768 4663 8802 4705
rect 8836 4739 8902 4773
rect 8836 4705 8852 4739
rect 8886 4705 8902 4739
rect 8836 4697 8902 4705
rect 8936 4807 8982 4823
rect 8970 4773 8982 4807
rect 8936 4739 8982 4773
rect 8970 4705 8982 4739
rect 8936 4663 8982 4705
rect 20800 4809 20842 4825
rect 20800 4775 20808 4809
rect 20800 4741 20842 4775
rect 20800 4707 20808 4741
rect 20800 4665 20842 4707
rect 20876 4809 22118 4829
rect 22758 4827 22824 4945
rect 24034 4943 24076 4959
rect 35980 5005 36046 5031
rect 36080 5133 36114 5175
rect 36080 5065 36114 5099
rect 36080 5015 36114 5031
rect 36148 5133 36214 5141
rect 36148 5099 36164 5133
rect 36198 5099 36214 5133
rect 36148 5065 36214 5099
rect 36148 5031 36164 5065
rect 36198 5031 36214 5065
rect 35980 4995 36001 5005
rect 35980 4961 35996 4995
rect 36035 4981 36046 5005
rect 36148 5009 36214 5031
rect 36248 5133 36282 5175
rect 36248 5065 36282 5099
rect 36248 5015 36282 5031
rect 36316 5133 36382 5141
rect 36316 5099 36332 5133
rect 36366 5099 36382 5133
rect 36316 5065 36382 5099
rect 36316 5031 36332 5065
rect 36366 5031 36382 5065
rect 36148 4981 36164 5009
rect 36035 4971 36164 4981
rect 36198 4981 36214 5009
rect 36316 5007 36382 5031
rect 36416 5133 36450 5175
rect 36416 5065 36450 5099
rect 36416 5015 36450 5031
rect 36484 5133 36550 5141
rect 36484 5099 36500 5133
rect 36534 5099 36550 5133
rect 36484 5065 36550 5099
rect 36484 5031 36500 5065
rect 36534 5031 36550 5065
rect 36316 4995 36334 5007
rect 36316 4981 36332 4995
rect 36030 4961 36164 4971
rect 36198 4961 36332 4981
rect 36368 4981 36382 5007
rect 36484 5007 36550 5031
rect 36584 5133 36618 5175
rect 36584 5065 36618 5099
rect 36584 5015 36618 5031
rect 36652 5133 36718 5141
rect 36652 5099 36668 5133
rect 36702 5099 36718 5133
rect 36652 5065 36718 5099
rect 36652 5031 36668 5065
rect 36702 5031 36718 5065
rect 36484 4981 36499 5007
rect 36533 4995 36550 5007
rect 36368 4973 36499 4981
rect 36534 4981 36550 4995
rect 36652 4995 36718 5031
rect 36752 5133 36786 5175
rect 36752 5065 36786 5099
rect 36752 5015 36786 5031
rect 36820 5133 36886 5141
rect 36820 5099 36836 5133
rect 36870 5099 36886 5133
rect 36820 5065 36886 5099
rect 36820 5031 36836 5065
rect 36870 5031 36886 5065
rect 36652 4981 36668 4995
rect 36366 4961 36500 4973
rect 36534 4961 36668 4981
rect 36702 4981 36718 4995
rect 36820 4996 36886 5031
rect 36920 5133 36954 5175
rect 36920 5065 36954 5099
rect 36920 5015 36954 5031
rect 36988 5133 37054 5141
rect 36988 5099 37004 5133
rect 37038 5099 37054 5133
rect 36988 5065 37054 5099
rect 36988 5031 37004 5065
rect 37038 5031 37054 5065
rect 36820 4995 36839 4996
rect 36820 4981 36836 4995
rect 36702 4961 36836 4981
rect 36873 4981 36886 4996
rect 36988 5001 37054 5031
rect 37088 5133 37122 5175
rect 37088 5065 37122 5099
rect 37088 5015 37122 5031
rect 37156 5133 37222 5141
rect 37156 5099 37172 5133
rect 37206 5099 37222 5133
rect 37156 5065 37222 5099
rect 37156 5031 37172 5065
rect 37206 5031 37222 5065
rect 36988 4981 37001 5001
rect 37035 4995 37054 5001
rect 36873 4967 37001 4981
rect 37038 4981 37054 4995
rect 37156 5002 37222 5031
rect 37156 4995 37174 5002
rect 37156 4981 37172 4995
rect 36873 4962 37004 4967
rect 36870 4961 37004 4962
rect 37038 4961 37172 4981
rect 37208 4968 37222 5002
rect 37206 4961 37222 4968
rect 35980 4959 36668 4961
rect 36702 4959 37222 4961
rect 35980 4947 37222 4959
rect 37256 5133 37298 5175
rect 37748 5173 37777 5207
rect 37811 5173 37869 5207
rect 37903 5173 37961 5207
rect 37995 5173 38053 5207
rect 38087 5173 38145 5207
rect 38179 5173 38237 5207
rect 38271 5173 38329 5207
rect 38363 5173 38421 5207
rect 38455 5173 38513 5207
rect 38547 5173 38605 5207
rect 38639 5173 38697 5207
rect 38731 5173 38789 5207
rect 38823 5173 38881 5207
rect 38915 5173 38973 5207
rect 39007 5173 39065 5207
rect 39099 5173 39157 5207
rect 39191 5173 39220 5207
rect 50964 5175 50993 5209
rect 51027 5175 51085 5209
rect 51119 5175 51177 5209
rect 51211 5175 51269 5209
rect 51303 5175 51361 5209
rect 51395 5175 51453 5209
rect 51487 5175 51545 5209
rect 51579 5175 51637 5209
rect 51671 5175 51729 5209
rect 51763 5175 51821 5209
rect 51855 5175 51913 5209
rect 51947 5175 52005 5209
rect 52039 5175 52097 5209
rect 52131 5175 52189 5209
rect 52223 5175 52281 5209
rect 52315 5175 52373 5209
rect 52407 5175 52436 5209
rect 37290 5099 37298 5133
rect 37256 5065 37298 5099
rect 37290 5031 37298 5065
rect 37256 4995 37298 5031
rect 37786 5131 37828 5173
rect 37786 5097 37794 5131
rect 37786 5063 37828 5097
rect 37786 5029 37794 5063
rect 37786 5013 37828 5029
rect 37862 5131 37928 5139
rect 37862 5097 37878 5131
rect 37912 5097 37928 5131
rect 37862 5063 37928 5097
rect 37862 5029 37878 5063
rect 37912 5029 37928 5063
rect 37290 4961 37298 4995
rect 23011 4900 24099 4909
rect 23011 4895 23028 4900
rect 23011 4861 23027 4895
rect 23062 4866 23132 4900
rect 23166 4895 23248 4900
rect 23166 4866 23194 4895
rect 23061 4861 23194 4866
rect 23228 4866 23248 4895
rect 23282 4866 23361 4900
rect 23395 4895 23474 4900
rect 23396 4866 23474 4895
rect 23508 4895 23587 4900
rect 23508 4866 23529 4895
rect 23228 4861 23362 4866
rect 23396 4861 23529 4866
rect 23563 4866 23587 4895
rect 23621 4895 23700 4900
rect 23621 4866 23698 4895
rect 23734 4866 23813 4900
rect 23847 4895 23926 4900
rect 23847 4866 23866 4895
rect 23563 4861 23698 4866
rect 23732 4861 23866 4866
rect 23900 4866 23926 4895
rect 23960 4895 24099 4900
rect 23960 4866 24040 4895
rect 23900 4861 24040 4866
rect 24074 4861 24099 4895
rect 35980 4829 36046 4947
rect 37256 4945 37298 4961
rect 37862 4993 37928 5029
rect 37962 5131 37996 5173
rect 37962 5063 37996 5097
rect 37962 5013 37996 5029
rect 38030 5131 38096 5139
rect 38030 5097 38046 5131
rect 38080 5097 38096 5131
rect 38030 5063 38096 5097
rect 38030 5029 38046 5063
rect 38080 5029 38096 5063
rect 37862 4959 37878 4993
rect 37912 4979 37928 4993
rect 38030 5003 38096 5029
rect 38130 5131 38164 5173
rect 38130 5063 38164 5097
rect 38130 5013 38164 5029
rect 38198 5131 38264 5139
rect 38198 5097 38214 5131
rect 38248 5097 38264 5131
rect 38198 5063 38264 5097
rect 38198 5029 38214 5063
rect 38248 5029 38264 5063
rect 38030 4993 38047 5003
rect 38030 4979 38046 4993
rect 37912 4959 38046 4979
rect 38081 4979 38096 5003
rect 38198 5012 38264 5029
rect 38298 5131 38332 5173
rect 38298 5063 38332 5097
rect 38298 5013 38332 5029
rect 38366 5131 38432 5139
rect 38366 5097 38382 5131
rect 38416 5097 38432 5131
rect 38366 5063 38432 5097
rect 38366 5029 38382 5063
rect 38416 5029 38432 5063
rect 38198 4993 38217 5012
rect 38198 4979 38214 4993
rect 38081 4969 38214 4979
rect 38251 4979 38264 5012
rect 38366 5010 38432 5029
rect 38466 5131 38500 5173
rect 38466 5063 38500 5097
rect 38466 5013 38500 5029
rect 38534 5131 38600 5139
rect 38534 5097 38550 5131
rect 38584 5097 38600 5131
rect 38534 5063 38600 5097
rect 38534 5029 38550 5063
rect 38584 5029 38600 5063
rect 38366 4993 38385 5010
rect 38366 4979 38382 4993
rect 38251 4978 38382 4979
rect 38080 4959 38214 4969
rect 38248 4959 38382 4978
rect 38419 4979 38432 5010
rect 38534 4997 38600 5029
rect 38634 5131 38668 5173
rect 38634 5063 38668 5097
rect 38634 5013 38668 5029
rect 38702 5131 38768 5139
rect 38702 5097 38718 5131
rect 38752 5097 38768 5131
rect 38702 5063 38768 5097
rect 38702 5029 38718 5063
rect 38752 5029 38768 5063
rect 38534 4993 38552 4997
rect 38534 4979 38550 4993
rect 38419 4976 38550 4979
rect 38416 4959 38550 4976
rect 38586 4979 38600 4997
rect 38702 5002 38768 5029
rect 38802 5131 38836 5173
rect 38802 5063 38836 5097
rect 38802 5013 38836 5029
rect 38870 5131 38936 5139
rect 38870 5097 38886 5131
rect 38920 5097 38936 5131
rect 38870 5063 38936 5097
rect 38870 5029 38886 5063
rect 38920 5029 38936 5063
rect 38702 4979 38717 5002
rect 38751 4993 38768 5002
rect 38586 4968 38717 4979
rect 38752 4979 38768 4993
rect 38870 5006 38936 5029
rect 38970 5131 39004 5173
rect 38970 5063 39004 5097
rect 38970 5013 39004 5029
rect 39038 5131 39104 5139
rect 39038 5097 39054 5131
rect 39088 5097 39104 5131
rect 39038 5063 39104 5097
rect 39038 5029 39054 5063
rect 39088 5029 39104 5063
rect 38870 4993 38890 5006
rect 38870 4979 38886 4993
rect 38586 4963 38718 4968
rect 38584 4959 38718 4963
rect 38752 4959 38886 4979
rect 38924 4979 38936 5006
rect 39038 5001 39104 5029
rect 39038 4979 39053 5001
rect 39087 4993 39104 5001
rect 38924 4972 39053 4979
rect 38920 4967 39053 4972
rect 38920 4959 39054 4967
rect 39088 4959 39104 4993
rect 37862 4945 39104 4959
rect 39138 5131 39180 5173
rect 39172 5097 39180 5131
rect 39138 5063 39180 5097
rect 39172 5029 39180 5063
rect 39138 4993 39180 5029
rect 51002 5133 51044 5175
rect 51002 5099 51010 5133
rect 51002 5065 51044 5099
rect 51002 5031 51010 5065
rect 51002 5015 51044 5031
rect 51078 5133 51144 5141
rect 51078 5099 51094 5133
rect 51128 5099 51144 5133
rect 51078 5065 51144 5099
rect 51078 5031 51094 5065
rect 51128 5031 51144 5065
rect 39172 4959 39180 4993
rect 36233 4900 37321 4911
rect 36233 4897 36520 4900
rect 36233 4863 36249 4897
rect 36283 4863 36416 4897
rect 36450 4866 36520 4897
rect 36554 4897 36628 4900
rect 36554 4866 36584 4897
rect 36450 4863 36584 4866
rect 36618 4866 36628 4897
rect 36662 4866 36736 4900
rect 36770 4897 36844 4900
rect 36785 4866 36844 4897
rect 36878 4897 36952 4900
rect 36878 4866 36920 4897
rect 36986 4866 37060 4900
rect 37094 4897 37168 4900
rect 37122 4866 37168 4897
rect 37202 4897 37276 4900
rect 37202 4866 37262 4897
rect 37310 4866 37321 4900
rect 36618 4863 36751 4866
rect 36785 4863 36920 4866
rect 36954 4863 37088 4866
rect 37122 4863 37262 4866
rect 37296 4863 37321 4866
rect 20876 4775 20892 4809
rect 20926 4791 21060 4809
rect 20926 4775 20942 4791
rect 20876 4741 20942 4775
rect 21044 4775 21060 4791
rect 21094 4791 21228 4809
rect 21094 4775 21110 4791
rect 20876 4707 20892 4741
rect 20926 4707 20942 4741
rect 20876 4699 20942 4707
rect 20976 4741 21010 4757
rect 20976 4665 21010 4707
rect 21044 4741 21110 4775
rect 21212 4775 21228 4791
rect 21262 4791 21396 4809
rect 21262 4775 21278 4791
rect 21044 4707 21060 4741
rect 21094 4707 21110 4741
rect 21044 4699 21110 4707
rect 21144 4741 21178 4757
rect 21144 4665 21178 4707
rect 21212 4741 21278 4775
rect 21380 4775 21396 4791
rect 21430 4791 21564 4809
rect 21430 4775 21446 4791
rect 21212 4707 21228 4741
rect 21262 4707 21278 4741
rect 21212 4699 21278 4707
rect 21312 4741 21346 4757
rect 21312 4665 21346 4707
rect 21380 4741 21446 4775
rect 21548 4775 21564 4791
rect 21598 4791 21732 4809
rect 21598 4775 21614 4791
rect 21380 4707 21396 4741
rect 21430 4707 21446 4741
rect 21380 4699 21446 4707
rect 21480 4741 21514 4757
rect 21480 4665 21514 4707
rect 21548 4741 21614 4775
rect 21716 4775 21732 4791
rect 21766 4791 21900 4809
rect 21766 4775 21782 4791
rect 21548 4707 21564 4741
rect 21598 4707 21614 4741
rect 21548 4699 21614 4707
rect 21648 4741 21682 4757
rect 21648 4665 21682 4707
rect 21716 4741 21782 4775
rect 21884 4775 21900 4791
rect 21934 4791 22068 4809
rect 21934 4775 21950 4791
rect 21716 4707 21732 4741
rect 21766 4707 21782 4741
rect 21716 4699 21782 4707
rect 21816 4741 21850 4757
rect 21816 4665 21850 4707
rect 21884 4741 21950 4775
rect 22052 4775 22068 4791
rect 22102 4775 22118 4809
rect 21884 4707 21900 4741
rect 21934 4707 21950 4741
rect 21884 4699 21950 4707
rect 21984 4741 22018 4757
rect 21984 4665 22018 4707
rect 22052 4741 22118 4775
rect 22052 4707 22068 4741
rect 22102 4707 22118 4741
rect 22052 4699 22118 4707
rect 22152 4809 22198 4825
rect 22186 4775 22198 4809
rect 22152 4741 22198 4775
rect 22186 4707 22198 4741
rect 22152 4665 22198 4707
rect 22682 4807 22724 4823
rect 22682 4773 22690 4807
rect 22682 4739 22724 4773
rect 22682 4705 22690 4739
rect 7546 4629 7575 4663
rect 7609 4629 7667 4663
rect 7701 4629 7759 4663
rect 7793 4629 7851 4663
rect 7885 4629 7943 4663
rect 7977 4629 8035 4663
rect 8069 4629 8127 4663
rect 8161 4629 8219 4663
rect 8253 4629 8311 4663
rect 8345 4629 8403 4663
rect 8437 4629 8495 4663
rect 8529 4629 8587 4663
rect 8621 4629 8679 4663
rect 8713 4629 8771 4663
rect 8805 4629 8863 4663
rect 8897 4629 8955 4663
rect 8989 4629 9018 4663
rect 20762 4631 20791 4665
rect 20825 4631 20883 4665
rect 20917 4631 20975 4665
rect 21009 4631 21067 4665
rect 21101 4631 21159 4665
rect 21193 4631 21251 4665
rect 21285 4631 21343 4665
rect 21377 4631 21435 4665
rect 21469 4631 21527 4665
rect 21561 4631 21619 4665
rect 21653 4631 21711 4665
rect 21745 4631 21803 4665
rect 21837 4631 21895 4665
rect 21929 4631 21987 4665
rect 22021 4631 22079 4665
rect 22113 4631 22171 4665
rect 22205 4631 22234 4665
rect 22682 4663 22724 4705
rect 22758 4807 24000 4827
rect 22758 4773 22774 4807
rect 22808 4789 22942 4807
rect 22808 4773 22824 4789
rect 22758 4739 22824 4773
rect 22926 4773 22942 4789
rect 22976 4789 23110 4807
rect 22976 4773 22992 4789
rect 22758 4705 22774 4739
rect 22808 4705 22824 4739
rect 22758 4697 22824 4705
rect 22858 4739 22892 4755
rect 22858 4663 22892 4705
rect 22926 4739 22992 4773
rect 23094 4773 23110 4789
rect 23144 4789 23278 4807
rect 23144 4773 23160 4789
rect 22926 4705 22942 4739
rect 22976 4705 22992 4739
rect 22926 4697 22992 4705
rect 23026 4739 23060 4755
rect 23026 4663 23060 4705
rect 23094 4739 23160 4773
rect 23262 4773 23278 4789
rect 23312 4789 23446 4807
rect 23312 4773 23328 4789
rect 23094 4705 23110 4739
rect 23144 4705 23160 4739
rect 23094 4697 23160 4705
rect 23194 4739 23228 4755
rect 23194 4663 23228 4705
rect 23262 4739 23328 4773
rect 23430 4773 23446 4789
rect 23480 4789 23614 4807
rect 23480 4773 23496 4789
rect 23262 4705 23278 4739
rect 23312 4705 23328 4739
rect 23262 4697 23328 4705
rect 23362 4739 23396 4755
rect 23362 4663 23396 4705
rect 23430 4739 23496 4773
rect 23598 4773 23614 4789
rect 23648 4789 23782 4807
rect 23648 4773 23664 4789
rect 23430 4705 23446 4739
rect 23480 4705 23496 4739
rect 23430 4697 23496 4705
rect 23530 4739 23564 4755
rect 23530 4663 23564 4705
rect 23598 4739 23664 4773
rect 23766 4773 23782 4789
rect 23816 4789 23950 4807
rect 23816 4773 23832 4789
rect 23598 4705 23614 4739
rect 23648 4705 23664 4739
rect 23598 4697 23664 4705
rect 23698 4739 23732 4755
rect 23698 4663 23732 4705
rect 23766 4739 23832 4773
rect 23934 4773 23950 4789
rect 23984 4773 24000 4807
rect 23766 4705 23782 4739
rect 23816 4705 23832 4739
rect 23766 4697 23832 4705
rect 23866 4739 23900 4755
rect 23866 4663 23900 4705
rect 23934 4739 24000 4773
rect 23934 4705 23950 4739
rect 23984 4705 24000 4739
rect 23934 4697 24000 4705
rect 24034 4807 24080 4823
rect 24068 4773 24080 4807
rect 24034 4739 24080 4773
rect 24068 4705 24080 4739
rect 24034 4663 24080 4705
rect 35904 4809 35946 4825
rect 35904 4775 35912 4809
rect 35904 4741 35946 4775
rect 35904 4707 35912 4741
rect 35904 4665 35946 4707
rect 35980 4809 37222 4829
rect 37862 4827 37928 4945
rect 39138 4943 39180 4959
rect 51078 4996 51144 5031
rect 51178 5133 51212 5175
rect 51178 5065 51212 5099
rect 51178 5015 51212 5031
rect 51246 5133 51312 5141
rect 51246 5099 51262 5133
rect 51296 5099 51312 5133
rect 51246 5065 51312 5099
rect 51246 5031 51262 5065
rect 51296 5031 51312 5065
rect 51078 4995 51103 4996
rect 51078 4961 51094 4995
rect 51137 4981 51144 4996
rect 51246 4998 51312 5031
rect 51346 5133 51380 5175
rect 51346 5065 51380 5099
rect 51346 5015 51380 5031
rect 51414 5133 51480 5141
rect 51414 5099 51430 5133
rect 51464 5099 51480 5133
rect 51414 5065 51480 5099
rect 51414 5031 51430 5065
rect 51464 5031 51480 5065
rect 51246 4981 51262 4998
rect 51137 4962 51262 4981
rect 51296 4981 51312 4998
rect 51414 5000 51480 5031
rect 51514 5133 51548 5175
rect 51514 5065 51548 5099
rect 51514 5015 51548 5031
rect 51582 5133 51648 5141
rect 51582 5099 51598 5133
rect 51632 5099 51648 5133
rect 51582 5065 51648 5099
rect 51582 5031 51598 5065
rect 51632 5031 51648 5065
rect 51414 4995 51432 5000
rect 51414 4981 51430 4995
rect 51128 4961 51262 4962
rect 51296 4961 51430 4981
rect 51466 4981 51480 5000
rect 51582 5006 51648 5031
rect 51682 5133 51716 5175
rect 51682 5065 51716 5099
rect 51682 5015 51716 5031
rect 51750 5133 51816 5141
rect 51750 5099 51766 5133
rect 51800 5099 51816 5133
rect 51750 5065 51816 5099
rect 51750 5031 51766 5065
rect 51800 5031 51816 5065
rect 51582 4995 51602 5006
rect 51582 4981 51598 4995
rect 51466 4966 51598 4981
rect 51636 4981 51648 5006
rect 51750 4995 51816 5031
rect 51850 5133 51884 5175
rect 51850 5065 51884 5099
rect 51850 5015 51884 5031
rect 51918 5133 51984 5141
rect 51918 5099 51934 5133
rect 51968 5099 51984 5133
rect 51918 5065 51984 5099
rect 51918 5031 51934 5065
rect 51968 5031 51984 5065
rect 51750 4981 51766 4995
rect 51636 4972 51766 4981
rect 51464 4961 51598 4966
rect 51632 4961 51766 4972
rect 51800 4981 51816 4995
rect 51918 5003 51984 5031
rect 52018 5133 52052 5175
rect 52018 5065 52052 5099
rect 52018 5015 52052 5031
rect 52086 5133 52152 5141
rect 52086 5099 52102 5133
rect 52136 5099 52152 5133
rect 52086 5065 52152 5099
rect 52086 5031 52102 5065
rect 52136 5031 52152 5065
rect 51918 4995 51935 5003
rect 51918 4981 51934 4995
rect 51800 4961 51934 4981
rect 51969 4981 51984 5003
rect 52086 4997 52152 5031
rect 52186 5133 52220 5175
rect 52186 5065 52220 5099
rect 52186 5015 52220 5031
rect 52254 5133 52320 5141
rect 52254 5099 52270 5133
rect 52304 5099 52320 5133
rect 52254 5065 52320 5099
rect 52254 5031 52270 5065
rect 52304 5031 52320 5065
rect 52086 4981 52102 4997
rect 51969 4969 52102 4981
rect 51968 4961 52102 4969
rect 52136 4981 52152 4997
rect 52254 4997 52320 5031
rect 52254 4981 52262 4997
rect 52296 4995 52320 4997
rect 52136 4963 52262 4981
rect 52136 4961 52270 4963
rect 52304 4961 52320 4995
rect 51078 4959 51766 4961
rect 51800 4959 52320 4961
rect 51078 4947 52320 4959
rect 52354 5133 52396 5175
rect 52846 5173 52875 5207
rect 52909 5173 52967 5207
rect 53001 5173 53059 5207
rect 53093 5173 53151 5207
rect 53185 5173 53243 5207
rect 53277 5173 53335 5207
rect 53369 5173 53427 5207
rect 53461 5173 53519 5207
rect 53553 5173 53611 5207
rect 53645 5173 53703 5207
rect 53737 5173 53795 5207
rect 53829 5173 53887 5207
rect 53921 5173 53979 5207
rect 54013 5173 54071 5207
rect 54105 5173 54163 5207
rect 54197 5173 54255 5207
rect 54289 5173 54318 5207
rect 52388 5099 52396 5133
rect 52354 5065 52396 5099
rect 52388 5031 52396 5065
rect 52354 4995 52396 5031
rect 52884 5131 52926 5173
rect 52884 5097 52892 5131
rect 52884 5063 52926 5097
rect 52884 5029 52892 5063
rect 52884 5013 52926 5029
rect 52960 5131 53026 5139
rect 52960 5097 52976 5131
rect 53010 5097 53026 5131
rect 52960 5063 53026 5097
rect 52960 5029 52976 5063
rect 53010 5029 53026 5063
rect 52388 4961 52396 4995
rect 38115 4900 39203 4909
rect 38115 4895 38132 4900
rect 38115 4861 38131 4895
rect 38166 4866 38283 4900
rect 38317 4895 38380 4900
rect 38332 4866 38380 4895
rect 38414 4895 38477 4900
rect 38414 4866 38466 4895
rect 38511 4866 38574 4900
rect 38608 4895 38671 4900
rect 38608 4866 38633 4895
rect 38165 4861 38298 4866
rect 38332 4861 38466 4866
rect 38500 4861 38633 4866
rect 38667 4866 38671 4895
rect 38705 4866 38768 4900
rect 38802 4895 38865 4900
rect 38667 4861 38802 4866
rect 38836 4866 38865 4895
rect 38899 4866 38962 4900
rect 38996 4895 39203 4900
rect 38836 4861 38970 4866
rect 39004 4861 39144 4895
rect 39178 4861 39203 4895
rect 51078 4829 51144 4947
rect 52354 4945 52396 4961
rect 52960 4994 53026 5029
rect 53060 5131 53094 5173
rect 53060 5063 53094 5097
rect 53060 5013 53094 5029
rect 53128 5131 53194 5139
rect 53128 5097 53144 5131
rect 53178 5097 53194 5131
rect 53128 5063 53194 5097
rect 53128 5029 53144 5063
rect 53178 5029 53194 5063
rect 52960 4959 52976 4994
rect 53010 4979 53026 4994
rect 53128 4996 53194 5029
rect 53228 5131 53262 5173
rect 53228 5063 53262 5097
rect 53228 5013 53262 5029
rect 53296 5131 53362 5139
rect 53296 5097 53312 5131
rect 53346 5097 53362 5131
rect 53296 5063 53362 5097
rect 53296 5029 53312 5063
rect 53346 5029 53362 5063
rect 53128 4993 53146 4996
rect 53128 4979 53144 4993
rect 53010 4959 53144 4979
rect 53180 4979 53194 4996
rect 53296 5002 53362 5029
rect 53396 5131 53430 5173
rect 53396 5063 53430 5097
rect 53396 5013 53430 5029
rect 53464 5131 53530 5139
rect 53464 5097 53480 5131
rect 53514 5097 53530 5131
rect 53464 5063 53530 5097
rect 53464 5029 53480 5063
rect 53514 5029 53530 5063
rect 53296 4979 53312 5002
rect 53180 4962 53312 4979
rect 53346 4979 53362 5002
rect 53464 5001 53530 5029
rect 53564 5131 53598 5173
rect 53564 5063 53598 5097
rect 53564 5013 53598 5029
rect 53632 5131 53698 5139
rect 53632 5097 53648 5131
rect 53682 5097 53698 5131
rect 53632 5063 53698 5097
rect 53632 5029 53648 5063
rect 53682 5029 53698 5063
rect 53464 4993 53481 5001
rect 53464 4979 53480 4993
rect 53178 4959 53312 4962
rect 53346 4959 53480 4979
rect 53515 4979 53530 5001
rect 53632 4997 53698 5029
rect 53732 5131 53766 5173
rect 53732 5063 53766 5097
rect 53732 5013 53766 5029
rect 53800 5131 53866 5139
rect 53800 5097 53816 5131
rect 53850 5097 53866 5131
rect 53800 5063 53866 5097
rect 53800 5029 53816 5063
rect 53850 5029 53866 5063
rect 53632 4993 53650 4997
rect 53632 4979 53648 4993
rect 53515 4967 53648 4979
rect 53514 4959 53648 4967
rect 53684 4979 53698 4997
rect 53800 4999 53866 5029
rect 53900 5131 53934 5173
rect 53900 5063 53934 5097
rect 53900 5013 53934 5029
rect 53968 5131 54034 5139
rect 53968 5097 53984 5131
rect 54018 5097 54034 5131
rect 53968 5063 54034 5097
rect 53968 5029 53984 5063
rect 54018 5029 54034 5063
rect 53800 4993 53821 4999
rect 53800 4979 53816 4993
rect 53684 4963 53816 4979
rect 53855 4979 53866 4999
rect 53968 4997 54034 5029
rect 54068 5131 54102 5173
rect 54068 5063 54102 5097
rect 54068 5013 54102 5029
rect 54136 5131 54202 5139
rect 54136 5097 54152 5131
rect 54186 5097 54202 5131
rect 54136 5063 54202 5097
rect 54136 5029 54152 5063
rect 54186 5029 54202 5063
rect 53968 4993 53985 4997
rect 53968 4979 53984 4993
rect 53855 4965 53984 4979
rect 53682 4959 53816 4963
rect 53850 4959 53984 4965
rect 54019 4979 54034 4997
rect 54136 4995 54202 5029
rect 54136 4979 54151 4995
rect 54185 4993 54202 4995
rect 54019 4963 54151 4979
rect 54018 4961 54151 4963
rect 54018 4959 54152 4961
rect 54186 4959 54202 4993
rect 52960 4945 54202 4959
rect 54236 5131 54278 5173
rect 54270 5097 54278 5131
rect 54236 5063 54278 5097
rect 54270 5029 54278 5063
rect 54236 4993 54278 5029
rect 54270 4959 54278 4993
rect 51331 4900 52419 4911
rect 51331 4897 51660 4900
rect 51694 4897 51779 4900
rect 51331 4863 51347 4897
rect 51381 4863 51514 4897
rect 51548 4866 51660 4897
rect 51716 4866 51779 4897
rect 51813 4897 51898 4900
rect 51813 4866 51849 4897
rect 51548 4863 51682 4866
rect 51716 4863 51849 4866
rect 51883 4866 51898 4897
rect 51932 4866 52017 4900
rect 52051 4897 52136 4900
rect 52052 4866 52136 4897
rect 52170 4897 52255 4900
rect 52170 4866 52186 4897
rect 51883 4863 52018 4866
rect 52052 4863 52186 4866
rect 52220 4866 52255 4897
rect 52289 4897 52374 4900
rect 52289 4866 52360 4897
rect 52408 4866 52419 4900
rect 52220 4863 52360 4866
rect 52394 4863 52419 4866
rect 35980 4775 35996 4809
rect 36030 4791 36164 4809
rect 36030 4775 36046 4791
rect 35980 4741 36046 4775
rect 36148 4775 36164 4791
rect 36198 4791 36332 4809
rect 36198 4775 36214 4791
rect 35980 4707 35996 4741
rect 36030 4707 36046 4741
rect 35980 4699 36046 4707
rect 36080 4741 36114 4757
rect 36080 4665 36114 4707
rect 36148 4741 36214 4775
rect 36316 4775 36332 4791
rect 36366 4791 36500 4809
rect 36366 4775 36382 4791
rect 36148 4707 36164 4741
rect 36198 4707 36214 4741
rect 36148 4699 36214 4707
rect 36248 4741 36282 4757
rect 36248 4665 36282 4707
rect 36316 4741 36382 4775
rect 36484 4775 36500 4791
rect 36534 4791 36668 4809
rect 36534 4775 36550 4791
rect 36316 4707 36332 4741
rect 36366 4707 36382 4741
rect 36316 4699 36382 4707
rect 36416 4741 36450 4757
rect 36416 4665 36450 4707
rect 36484 4741 36550 4775
rect 36652 4775 36668 4791
rect 36702 4791 36836 4809
rect 36702 4775 36718 4791
rect 36484 4707 36500 4741
rect 36534 4707 36550 4741
rect 36484 4699 36550 4707
rect 36584 4741 36618 4757
rect 36584 4665 36618 4707
rect 36652 4741 36718 4775
rect 36820 4775 36836 4791
rect 36870 4791 37004 4809
rect 36870 4775 36886 4791
rect 36652 4707 36668 4741
rect 36702 4707 36718 4741
rect 36652 4699 36718 4707
rect 36752 4741 36786 4757
rect 36752 4665 36786 4707
rect 36820 4741 36886 4775
rect 36988 4775 37004 4791
rect 37038 4791 37172 4809
rect 37038 4775 37054 4791
rect 36820 4707 36836 4741
rect 36870 4707 36886 4741
rect 36820 4699 36886 4707
rect 36920 4741 36954 4757
rect 36920 4665 36954 4707
rect 36988 4741 37054 4775
rect 37156 4775 37172 4791
rect 37206 4775 37222 4809
rect 36988 4707 37004 4741
rect 37038 4707 37054 4741
rect 36988 4699 37054 4707
rect 37088 4741 37122 4757
rect 37088 4665 37122 4707
rect 37156 4741 37222 4775
rect 37156 4707 37172 4741
rect 37206 4707 37222 4741
rect 37156 4699 37222 4707
rect 37256 4809 37302 4825
rect 37290 4775 37302 4809
rect 37256 4741 37302 4775
rect 37290 4707 37302 4741
rect 37256 4665 37302 4707
rect 37786 4807 37828 4823
rect 37786 4773 37794 4807
rect 37786 4739 37828 4773
rect 37786 4705 37794 4739
rect 22644 4629 22673 4663
rect 22707 4629 22765 4663
rect 22799 4629 22857 4663
rect 22891 4629 22949 4663
rect 22983 4629 23041 4663
rect 23075 4629 23133 4663
rect 23167 4629 23225 4663
rect 23259 4629 23317 4663
rect 23351 4629 23409 4663
rect 23443 4629 23501 4663
rect 23535 4629 23593 4663
rect 23627 4629 23685 4663
rect 23719 4629 23777 4663
rect 23811 4629 23869 4663
rect 23903 4629 23961 4663
rect 23995 4629 24053 4663
rect 24087 4629 24116 4663
rect 35866 4631 35895 4665
rect 35929 4631 35987 4665
rect 36021 4631 36079 4665
rect 36113 4631 36171 4665
rect 36205 4631 36263 4665
rect 36297 4631 36355 4665
rect 36389 4631 36447 4665
rect 36481 4631 36539 4665
rect 36573 4631 36631 4665
rect 36665 4631 36723 4665
rect 36757 4631 36815 4665
rect 36849 4631 36907 4665
rect 36941 4631 36999 4665
rect 37033 4631 37091 4665
rect 37125 4631 37183 4665
rect 37217 4631 37275 4665
rect 37309 4631 37338 4665
rect 37786 4663 37828 4705
rect 37862 4807 39104 4827
rect 37862 4773 37878 4807
rect 37912 4789 38046 4807
rect 37912 4773 37928 4789
rect 37862 4739 37928 4773
rect 38030 4773 38046 4789
rect 38080 4789 38214 4807
rect 38080 4773 38096 4789
rect 37862 4705 37878 4739
rect 37912 4705 37928 4739
rect 37862 4697 37928 4705
rect 37962 4739 37996 4755
rect 37962 4663 37996 4705
rect 38030 4739 38096 4773
rect 38198 4773 38214 4789
rect 38248 4789 38382 4807
rect 38248 4773 38264 4789
rect 38030 4705 38046 4739
rect 38080 4705 38096 4739
rect 38030 4697 38096 4705
rect 38130 4739 38164 4755
rect 38130 4663 38164 4705
rect 38198 4739 38264 4773
rect 38366 4773 38382 4789
rect 38416 4789 38550 4807
rect 38416 4773 38432 4789
rect 38198 4705 38214 4739
rect 38248 4705 38264 4739
rect 38198 4697 38264 4705
rect 38298 4739 38332 4755
rect 38298 4663 38332 4705
rect 38366 4739 38432 4773
rect 38534 4773 38550 4789
rect 38584 4789 38718 4807
rect 38584 4773 38600 4789
rect 38366 4705 38382 4739
rect 38416 4705 38432 4739
rect 38366 4697 38432 4705
rect 38466 4739 38500 4755
rect 38466 4663 38500 4705
rect 38534 4739 38600 4773
rect 38702 4773 38718 4789
rect 38752 4789 38886 4807
rect 38752 4773 38768 4789
rect 38534 4705 38550 4739
rect 38584 4705 38600 4739
rect 38534 4697 38600 4705
rect 38634 4739 38668 4755
rect 38634 4663 38668 4705
rect 38702 4739 38768 4773
rect 38870 4773 38886 4789
rect 38920 4789 39054 4807
rect 38920 4773 38936 4789
rect 38702 4705 38718 4739
rect 38752 4705 38768 4739
rect 38702 4697 38768 4705
rect 38802 4739 38836 4755
rect 38802 4663 38836 4705
rect 38870 4739 38936 4773
rect 39038 4773 39054 4789
rect 39088 4773 39104 4807
rect 38870 4705 38886 4739
rect 38920 4705 38936 4739
rect 38870 4697 38936 4705
rect 38970 4739 39004 4755
rect 38970 4663 39004 4705
rect 39038 4739 39104 4773
rect 39038 4705 39054 4739
rect 39088 4705 39104 4739
rect 39038 4697 39104 4705
rect 39138 4807 39184 4823
rect 39172 4773 39184 4807
rect 39138 4739 39184 4773
rect 39172 4705 39184 4739
rect 39138 4663 39184 4705
rect 51002 4809 51044 4825
rect 51002 4775 51010 4809
rect 51002 4741 51044 4775
rect 51002 4707 51010 4741
rect 51002 4665 51044 4707
rect 51078 4809 52320 4829
rect 52960 4827 53026 4945
rect 54236 4943 54278 4959
rect 53213 4900 54301 4909
rect 53213 4895 53230 4900
rect 53213 4861 53229 4895
rect 53264 4866 53334 4900
rect 53368 4895 53450 4900
rect 53368 4866 53396 4895
rect 53263 4861 53396 4866
rect 53430 4866 53450 4895
rect 53484 4866 53563 4900
rect 53597 4895 53676 4900
rect 53598 4866 53676 4895
rect 53710 4895 53789 4900
rect 53710 4866 53731 4895
rect 53430 4861 53564 4866
rect 53598 4861 53731 4866
rect 53765 4866 53789 4895
rect 53823 4895 53902 4900
rect 53823 4866 53900 4895
rect 53936 4866 54015 4900
rect 54049 4895 54128 4900
rect 54049 4866 54068 4895
rect 53765 4861 53900 4866
rect 53934 4861 54068 4866
rect 54102 4866 54128 4895
rect 54162 4895 54301 4900
rect 54162 4866 54242 4895
rect 54102 4861 54242 4866
rect 54276 4861 54301 4895
rect 51078 4775 51094 4809
rect 51128 4791 51262 4809
rect 51128 4775 51144 4791
rect 51078 4741 51144 4775
rect 51246 4775 51262 4791
rect 51296 4791 51430 4809
rect 51296 4775 51312 4791
rect 51078 4707 51094 4741
rect 51128 4707 51144 4741
rect 51078 4699 51144 4707
rect 51178 4741 51212 4757
rect 51178 4665 51212 4707
rect 51246 4741 51312 4775
rect 51414 4775 51430 4791
rect 51464 4791 51598 4809
rect 51464 4775 51480 4791
rect 51246 4707 51262 4741
rect 51296 4707 51312 4741
rect 51246 4699 51312 4707
rect 51346 4741 51380 4757
rect 51346 4665 51380 4707
rect 51414 4741 51480 4775
rect 51582 4775 51598 4791
rect 51632 4791 51766 4809
rect 51632 4775 51648 4791
rect 51414 4707 51430 4741
rect 51464 4707 51480 4741
rect 51414 4699 51480 4707
rect 51514 4741 51548 4757
rect 51514 4665 51548 4707
rect 51582 4741 51648 4775
rect 51750 4775 51766 4791
rect 51800 4791 51934 4809
rect 51800 4775 51816 4791
rect 51582 4707 51598 4741
rect 51632 4707 51648 4741
rect 51582 4699 51648 4707
rect 51682 4741 51716 4757
rect 51682 4665 51716 4707
rect 51750 4741 51816 4775
rect 51918 4775 51934 4791
rect 51968 4791 52102 4809
rect 51968 4775 51984 4791
rect 51750 4707 51766 4741
rect 51800 4707 51816 4741
rect 51750 4699 51816 4707
rect 51850 4741 51884 4757
rect 51850 4665 51884 4707
rect 51918 4741 51984 4775
rect 52086 4775 52102 4791
rect 52136 4791 52270 4809
rect 52136 4775 52152 4791
rect 51918 4707 51934 4741
rect 51968 4707 51984 4741
rect 51918 4699 51984 4707
rect 52018 4741 52052 4757
rect 52018 4665 52052 4707
rect 52086 4741 52152 4775
rect 52254 4775 52270 4791
rect 52304 4775 52320 4809
rect 52086 4707 52102 4741
rect 52136 4707 52152 4741
rect 52086 4699 52152 4707
rect 52186 4741 52220 4757
rect 52186 4665 52220 4707
rect 52254 4741 52320 4775
rect 52254 4707 52270 4741
rect 52304 4707 52320 4741
rect 52254 4699 52320 4707
rect 52354 4809 52400 4825
rect 52388 4775 52400 4809
rect 52354 4741 52400 4775
rect 52388 4707 52400 4741
rect 52354 4665 52400 4707
rect 52884 4807 52926 4823
rect 52884 4773 52892 4807
rect 52884 4739 52926 4773
rect 52884 4705 52892 4739
rect 37748 4629 37777 4663
rect 37811 4629 37869 4663
rect 37903 4629 37961 4663
rect 37995 4629 38053 4663
rect 38087 4629 38145 4663
rect 38179 4629 38237 4663
rect 38271 4629 38329 4663
rect 38363 4629 38421 4663
rect 38455 4629 38513 4663
rect 38547 4629 38605 4663
rect 38639 4629 38697 4663
rect 38731 4629 38789 4663
rect 38823 4629 38881 4663
rect 38915 4629 38973 4663
rect 39007 4629 39065 4663
rect 39099 4629 39157 4663
rect 39191 4629 39220 4663
rect 50964 4631 50993 4665
rect 51027 4631 51085 4665
rect 51119 4631 51177 4665
rect 51211 4631 51269 4665
rect 51303 4631 51361 4665
rect 51395 4631 51453 4665
rect 51487 4631 51545 4665
rect 51579 4631 51637 4665
rect 51671 4631 51729 4665
rect 51763 4631 51821 4665
rect 51855 4631 51913 4665
rect 51947 4631 52005 4665
rect 52039 4631 52097 4665
rect 52131 4631 52189 4665
rect 52223 4631 52281 4665
rect 52315 4631 52373 4665
rect 52407 4631 52436 4665
rect 52884 4663 52926 4705
rect 52960 4807 54202 4827
rect 52960 4773 52976 4807
rect 53010 4789 53144 4807
rect 53010 4773 53026 4789
rect 52960 4739 53026 4773
rect 53128 4773 53144 4789
rect 53178 4789 53312 4807
rect 53178 4773 53194 4789
rect 52960 4705 52976 4739
rect 53010 4705 53026 4739
rect 52960 4697 53026 4705
rect 53060 4739 53094 4755
rect 53060 4663 53094 4705
rect 53128 4739 53194 4773
rect 53296 4773 53312 4789
rect 53346 4789 53480 4807
rect 53346 4773 53362 4789
rect 53128 4705 53144 4739
rect 53178 4705 53194 4739
rect 53128 4697 53194 4705
rect 53228 4739 53262 4755
rect 53228 4663 53262 4705
rect 53296 4739 53362 4773
rect 53464 4773 53480 4789
rect 53514 4789 53648 4807
rect 53514 4773 53530 4789
rect 53296 4705 53312 4739
rect 53346 4705 53362 4739
rect 53296 4697 53362 4705
rect 53396 4739 53430 4755
rect 53396 4663 53430 4705
rect 53464 4739 53530 4773
rect 53632 4773 53648 4789
rect 53682 4789 53816 4807
rect 53682 4773 53698 4789
rect 53464 4705 53480 4739
rect 53514 4705 53530 4739
rect 53464 4697 53530 4705
rect 53564 4739 53598 4755
rect 53564 4663 53598 4705
rect 53632 4739 53698 4773
rect 53800 4773 53816 4789
rect 53850 4789 53984 4807
rect 53850 4773 53866 4789
rect 53632 4705 53648 4739
rect 53682 4705 53698 4739
rect 53632 4697 53698 4705
rect 53732 4739 53766 4755
rect 53732 4663 53766 4705
rect 53800 4739 53866 4773
rect 53968 4773 53984 4789
rect 54018 4789 54152 4807
rect 54018 4773 54034 4789
rect 53800 4705 53816 4739
rect 53850 4705 53866 4739
rect 53800 4697 53866 4705
rect 53900 4739 53934 4755
rect 53900 4663 53934 4705
rect 53968 4739 54034 4773
rect 54136 4773 54152 4789
rect 54186 4773 54202 4807
rect 53968 4705 53984 4739
rect 54018 4705 54034 4739
rect 53968 4697 54034 4705
rect 54068 4739 54102 4755
rect 54068 4663 54102 4705
rect 54136 4739 54202 4773
rect 54136 4705 54152 4739
rect 54186 4705 54202 4739
rect 54136 4697 54202 4705
rect 54236 4807 54282 4823
rect 54270 4773 54282 4807
rect 54236 4739 54282 4773
rect 54270 4705 54282 4739
rect 54236 4663 54282 4705
rect 52846 4629 52875 4663
rect 52909 4629 52967 4663
rect 53001 4629 53059 4663
rect 53093 4629 53151 4663
rect 53185 4629 53243 4663
rect 53277 4629 53335 4663
rect 53369 4629 53427 4663
rect 53461 4629 53519 4663
rect 53553 4629 53611 4663
rect 53645 4629 53703 4663
rect 53737 4629 53795 4663
rect 53829 4629 53887 4663
rect 53921 4629 53979 4663
rect 54013 4629 54071 4663
rect 54105 4629 54163 4663
rect 54197 4629 54255 4663
rect 54289 4629 54318 4663
rect 30027 4098 30056 4132
rect 30090 4098 30148 4132
rect 30182 4098 30240 4132
rect 30274 4098 30332 4132
rect 30366 4098 30424 4132
rect 30458 4098 30487 4132
rect 30555 4098 30584 4132
rect 30618 4098 30676 4132
rect 30710 4098 30768 4132
rect 30802 4098 30860 4132
rect 30894 4098 30952 4132
rect 30986 4098 31044 4132
rect 31078 4098 31136 4132
rect 31170 4098 31228 4132
rect 31262 4098 31320 4132
rect 31354 4098 31412 4132
rect 31446 4098 31504 4132
rect 31538 4098 31596 4132
rect 31630 4098 31688 4132
rect 31722 4098 31780 4132
rect 31814 4098 31872 4132
rect 31906 4098 31964 4132
rect 31998 4098 32027 4132
rect 30053 4056 30106 4098
rect 30053 4022 30072 4056
rect 30053 3988 30106 4022
rect 30053 3954 30072 3988
rect 30053 3920 30106 3954
rect 30053 3886 30072 3920
rect 30053 3870 30106 3886
rect 30140 4056 30206 4064
rect 30140 4022 30156 4056
rect 30190 4022 30206 4056
rect 30140 3988 30206 4022
rect 30140 3954 30156 3988
rect 30190 3954 30206 3988
rect 30140 3920 30206 3954
rect 30240 4056 30274 4098
rect 30240 3988 30274 4022
rect 30240 3938 30274 3954
rect 30308 4056 30374 4064
rect 30308 4022 30324 4056
rect 30358 4022 30374 4056
rect 30308 3988 30374 4022
rect 30408 4056 30450 4098
rect 30442 4022 30450 4056
rect 30408 4006 30450 4022
rect 30595 4056 30637 4098
rect 30595 4022 30603 4056
rect 30308 3954 30324 3988
rect 30358 3954 30374 3988
rect 30140 3886 30156 3920
rect 30190 3904 30206 3920
rect 30308 3920 30374 3954
rect 30308 3904 30324 3920
rect 30190 3886 30324 3904
rect 30358 3908 30374 3920
rect 30595 3988 30637 4022
rect 30595 3954 30603 3988
rect 30595 3918 30637 3954
rect 30358 3886 30461 3908
rect 30140 3870 30461 3886
rect 30408 3862 30461 3870
rect 30595 3884 30603 3918
rect 30595 3868 30637 3884
rect 30671 4056 30737 4064
rect 30671 4022 30687 4056
rect 30721 4022 30737 4056
rect 30671 3988 30737 4022
rect 30671 3954 30687 3988
rect 30721 3954 30737 3988
rect 30671 3918 30737 3954
rect 30771 4056 30805 4098
rect 30771 3988 30805 4022
rect 30771 3938 30805 3954
rect 30839 4056 30905 4064
rect 30839 4022 30855 4056
rect 30889 4022 30905 4056
rect 30839 3988 30905 4022
rect 30839 3954 30855 3988
rect 30889 3954 30905 3988
rect 30671 3884 30687 3918
rect 30721 3904 30737 3918
rect 30839 3918 30905 3954
rect 30939 4056 30973 4098
rect 30939 3988 30973 4022
rect 30939 3938 30973 3954
rect 31007 4056 31073 4064
rect 31007 4022 31023 4056
rect 31057 4022 31073 4056
rect 31007 3988 31073 4022
rect 31007 3954 31023 3988
rect 31057 3954 31073 3988
rect 30839 3904 30855 3918
rect 30721 3884 30855 3904
rect 30889 3904 30905 3918
rect 31007 3918 31073 3954
rect 31107 4056 31141 4098
rect 31107 3988 31141 4022
rect 31107 3938 31141 3954
rect 31175 4056 31241 4064
rect 31175 4022 31191 4056
rect 31225 4022 31241 4056
rect 31175 3988 31241 4022
rect 31175 3954 31191 3988
rect 31225 3954 31241 3988
rect 31007 3904 31023 3918
rect 30889 3884 31023 3904
rect 31057 3904 31073 3918
rect 31175 3918 31241 3954
rect 31275 4056 31309 4098
rect 31275 3988 31309 4022
rect 31275 3938 31309 3954
rect 31343 4056 31409 4064
rect 31343 4022 31359 4056
rect 31393 4022 31409 4056
rect 31343 3988 31409 4022
rect 31343 3954 31359 3988
rect 31393 3954 31409 3988
rect 31175 3904 31191 3918
rect 31057 3884 31191 3904
rect 31225 3904 31241 3918
rect 31343 3918 31409 3954
rect 31443 4056 31477 4098
rect 31443 3988 31477 4022
rect 31443 3938 31477 3954
rect 31511 4056 31577 4064
rect 31511 4022 31527 4056
rect 31561 4022 31577 4056
rect 31511 3988 31577 4022
rect 31511 3954 31527 3988
rect 31561 3954 31577 3988
rect 31343 3904 31359 3918
rect 31225 3884 31359 3904
rect 31393 3904 31409 3918
rect 31511 3918 31577 3954
rect 31611 4056 31645 4098
rect 31611 3988 31645 4022
rect 31611 3938 31645 3954
rect 31679 4056 31745 4064
rect 31679 4022 31695 4056
rect 31729 4022 31745 4056
rect 31679 3988 31745 4022
rect 31679 3954 31695 3988
rect 31729 3954 31745 3988
rect 31511 3904 31527 3918
rect 31393 3884 31527 3904
rect 31561 3904 31577 3918
rect 31679 3918 31745 3954
rect 31779 4056 31813 4098
rect 31779 3988 31813 4022
rect 31779 3938 31813 3954
rect 31847 4056 31913 4064
rect 31847 4022 31863 4056
rect 31897 4022 31913 4056
rect 31847 3988 31913 4022
rect 31847 3954 31863 3988
rect 31897 3954 31913 3988
rect 31679 3904 31695 3918
rect 31561 3884 31695 3904
rect 31729 3904 31745 3918
rect 31847 3918 31913 3954
rect 31947 4056 31989 4098
rect 31981 4038 31989 4056
rect 31981 4022 32102 4038
rect 31947 3988 32102 4022
rect 31981 3962 32102 3988
rect 31981 3954 31989 3962
rect 31947 3938 31989 3954
rect 31847 3904 31863 3918
rect 31729 3884 31863 3904
rect 31897 3884 31913 3918
rect 30671 3870 31913 3884
rect 43381 3882 43410 3916
rect 43444 3882 43502 3916
rect 43536 3882 43594 3916
rect 43628 3882 43686 3916
rect 43720 3882 43778 3916
rect 43812 3882 43870 3916
rect 43904 3882 43962 3916
rect 43996 3882 44054 3916
rect 44088 3882 44146 3916
rect 44180 3882 44238 3916
rect 44272 3882 44330 3916
rect 44364 3882 44422 3916
rect 44456 3882 44514 3916
rect 44548 3882 44606 3916
rect 44640 3882 44698 3916
rect 44732 3882 44790 3916
rect 44824 3882 44853 3916
rect 45311 3882 45340 3916
rect 45374 3882 45432 3916
rect 45466 3882 45524 3916
rect 45558 3882 45616 3916
rect 45650 3882 45708 3916
rect 45742 3882 45800 3916
rect 45834 3882 45892 3916
rect 45926 3882 45984 3916
rect 46018 3882 46076 3916
rect 46110 3882 46168 3916
rect 46202 3882 46260 3916
rect 46294 3882 46352 3916
rect 46386 3882 46444 3916
rect 46478 3882 46536 3916
rect 46570 3882 46628 3916
rect 46662 3882 46720 3916
rect 46754 3882 46783 3916
rect 29711 3820 30374 3836
rect 29711 3786 30064 3820
rect 30098 3786 30156 3820
rect 30190 3786 30240 3820
rect 30274 3786 30324 3820
rect 30358 3786 30374 3820
rect 30408 3828 30423 3862
rect 30457 3828 30461 3862
rect 30408 3782 30461 3828
rect 30572 3826 31660 3834
rect 30572 3820 30606 3826
rect 30572 3786 30597 3820
rect 30640 3792 30694 3826
rect 30728 3820 30782 3826
rect 30728 3792 30771 3820
rect 30816 3792 30870 3826
rect 30904 3820 30958 3826
rect 30904 3792 30939 3820
rect 30992 3792 31046 3826
rect 31080 3820 31134 3826
rect 31080 3792 31108 3820
rect 31168 3792 31222 3826
rect 31256 3820 31310 3826
rect 31256 3792 31275 3820
rect 30631 3786 30771 3792
rect 30805 3786 30939 3792
rect 30973 3786 31108 3792
rect 31142 3786 31275 3792
rect 31309 3792 31310 3820
rect 31344 3820 31660 3826
rect 31344 3792 31443 3820
rect 31309 3786 31443 3792
rect 31477 3786 31610 3820
rect 31644 3786 31660 3820
rect 13239 3722 13268 3756
rect 13302 3722 13360 3756
rect 13394 3722 13452 3756
rect 13486 3722 13544 3756
rect 13578 3722 13636 3756
rect 13670 3722 13728 3756
rect 13762 3722 13820 3756
rect 13854 3722 13912 3756
rect 13946 3722 14004 3756
rect 14038 3722 14096 3756
rect 14130 3722 14188 3756
rect 14222 3722 14280 3756
rect 14314 3722 14372 3756
rect 14406 3722 14464 3756
rect 14498 3722 14556 3756
rect 14590 3722 14648 3756
rect 14682 3722 14711 3756
rect 15169 3722 15198 3756
rect 15232 3722 15290 3756
rect 15324 3722 15382 3756
rect 15416 3722 15474 3756
rect 15508 3722 15566 3756
rect 15600 3722 15658 3756
rect 15692 3722 15750 3756
rect 15784 3722 15842 3756
rect 15876 3722 15934 3756
rect 15968 3722 16026 3756
rect 16060 3722 16118 3756
rect 16152 3722 16210 3756
rect 16244 3722 16302 3756
rect 16336 3722 16394 3756
rect 16428 3722 16486 3756
rect 16520 3722 16578 3756
rect 16612 3722 16641 3756
rect 30408 3752 30423 3782
rect 30140 3748 30423 3752
rect 30457 3748 30461 3782
rect 31847 3752 31913 3870
rect 13279 3680 13321 3722
rect 13279 3646 13287 3680
rect 13279 3612 13321 3646
rect 13279 3578 13287 3612
rect 13279 3542 13321 3578
rect 13279 3508 13287 3542
rect 13279 3492 13321 3508
rect 13355 3680 13421 3688
rect 13355 3646 13371 3680
rect 13405 3646 13421 3680
rect 13355 3612 13421 3646
rect 13355 3578 13371 3612
rect 13405 3578 13421 3612
rect 13355 3554 13421 3578
rect 13455 3680 13489 3722
rect 13455 3612 13489 3646
rect 13455 3562 13489 3578
rect 13523 3680 13589 3688
rect 13523 3646 13539 3680
rect 13573 3646 13589 3680
rect 13523 3612 13589 3646
rect 13523 3578 13539 3612
rect 13573 3578 13589 3612
rect 13355 3542 13372 3554
rect 13355 3508 13371 3542
rect 13406 3528 13421 3554
rect 13523 3561 13589 3578
rect 13623 3680 13657 3722
rect 13623 3612 13657 3646
rect 13623 3562 13657 3578
rect 13691 3680 13757 3688
rect 13691 3646 13707 3680
rect 13741 3646 13757 3680
rect 13691 3612 13757 3646
rect 13691 3578 13707 3612
rect 13741 3578 13757 3612
rect 13523 3542 13540 3561
rect 13523 3528 13539 3542
rect 13406 3509 13539 3528
rect 13574 3528 13589 3561
rect 13691 3551 13757 3578
rect 13791 3680 13825 3722
rect 13791 3612 13825 3646
rect 13791 3562 13825 3578
rect 13859 3680 13925 3688
rect 13859 3646 13875 3680
rect 13909 3646 13925 3680
rect 13859 3612 13925 3646
rect 13859 3578 13875 3612
rect 13909 3578 13925 3612
rect 13859 3563 13925 3578
rect 13691 3542 13708 3551
rect 13691 3528 13707 3542
rect 13574 3516 13707 3528
rect 13405 3508 13539 3509
rect 13573 3508 13707 3516
rect 13742 3528 13757 3551
rect 13859 3542 13876 3563
rect 13859 3528 13875 3542
rect 13742 3508 13875 3528
rect 13910 3528 13925 3563
rect 13959 3680 13993 3722
rect 13959 3612 13993 3646
rect 13959 3562 13993 3578
rect 14027 3680 14093 3688
rect 14027 3646 14043 3680
rect 14077 3646 14093 3680
rect 14027 3612 14093 3646
rect 14027 3578 14043 3612
rect 14077 3578 14093 3612
rect 14027 3561 14093 3578
rect 14127 3680 14161 3722
rect 14127 3612 14161 3646
rect 14127 3562 14161 3578
rect 14195 3680 14261 3688
rect 14195 3646 14211 3680
rect 14245 3646 14261 3680
rect 14195 3612 14261 3646
rect 14195 3578 14211 3612
rect 14245 3578 14261 3612
rect 14195 3563 14261 3578
rect 14027 3528 14042 3561
rect 14076 3542 14093 3561
rect 13910 3518 14042 3528
rect 13909 3516 14042 3518
rect 14077 3528 14093 3542
rect 14195 3528 14208 3563
rect 14242 3542 14261 3563
rect 14295 3680 14329 3722
rect 14295 3612 14329 3646
rect 14295 3562 14329 3578
rect 14363 3680 14429 3688
rect 14363 3646 14379 3680
rect 14413 3646 14429 3680
rect 14363 3612 14429 3646
rect 14363 3578 14379 3612
rect 14413 3578 14429 3612
rect 14363 3563 14429 3578
rect 14077 3518 14208 3528
rect 14245 3528 14261 3542
rect 14363 3528 14376 3563
rect 14410 3542 14429 3563
rect 14463 3680 14497 3722
rect 14463 3612 14497 3646
rect 14463 3562 14497 3578
rect 14531 3680 14597 3688
rect 14531 3646 14547 3680
rect 14581 3646 14597 3680
rect 14531 3612 14597 3646
rect 14531 3578 14547 3612
rect 14581 3578 14597 3612
rect 14245 3518 14376 3528
rect 14413 3528 14429 3542
rect 14531 3561 14597 3578
rect 14631 3680 14673 3722
rect 14665 3649 14673 3680
rect 15209 3680 15251 3722
rect 15209 3649 15217 3680
rect 14665 3646 15217 3649
rect 14631 3629 15251 3646
rect 14631 3612 14946 3629
rect 14665 3595 14946 3612
rect 14980 3612 15251 3629
rect 14980 3595 15217 3612
rect 14665 3578 15217 3595
rect 14631 3577 15251 3578
rect 14631 3562 14673 3577
rect 14531 3542 14550 3561
rect 14531 3528 14547 3542
rect 13909 3508 14043 3516
rect 14077 3508 14211 3518
rect 14245 3508 14379 3518
rect 14413 3508 14547 3528
rect 14584 3516 14597 3561
rect 14581 3508 14597 3516
rect 13355 3506 13708 3508
rect 13742 3506 14597 3508
rect 13355 3494 14597 3506
rect 13256 3452 14344 3458
rect 13256 3444 13572 3452
rect 13256 3410 13281 3444
rect 13315 3410 13455 3444
rect 13489 3418 13572 3444
rect 13606 3444 13672 3452
rect 13606 3418 13623 3444
rect 13489 3410 13623 3418
rect 13657 3418 13672 3444
rect 13706 3418 13772 3452
rect 13806 3444 13872 3452
rect 13826 3418 13872 3444
rect 13906 3444 13972 3452
rect 13906 3418 13959 3444
rect 14006 3418 14072 3452
rect 14106 3444 14172 3452
rect 14106 3418 14127 3444
rect 13657 3410 13792 3418
rect 13826 3410 13959 3418
rect 13993 3410 14127 3418
rect 14161 3418 14172 3444
rect 14206 3418 14272 3452
rect 14306 3444 14344 3452
rect 14161 3410 14294 3418
rect 14328 3410 14344 3444
rect 14531 3376 14597 3494
rect 15209 3542 15251 3577
rect 15209 3508 15217 3542
rect 15209 3492 15251 3508
rect 15285 3680 15351 3688
rect 15285 3646 15301 3680
rect 15335 3646 15351 3680
rect 15285 3612 15351 3646
rect 15285 3578 15301 3612
rect 15335 3578 15351 3612
rect 15285 3555 15351 3578
rect 15385 3680 15419 3722
rect 15385 3612 15419 3646
rect 15385 3562 15419 3578
rect 15453 3680 15519 3688
rect 15453 3646 15469 3680
rect 15503 3646 15519 3680
rect 15453 3612 15519 3646
rect 15453 3578 15469 3612
rect 15503 3578 15519 3612
rect 15285 3542 15306 3555
rect 15285 3508 15301 3542
rect 15340 3528 15351 3555
rect 15453 3559 15519 3578
rect 15553 3680 15587 3722
rect 15553 3612 15587 3646
rect 15553 3562 15587 3578
rect 15621 3680 15687 3688
rect 15621 3646 15637 3680
rect 15671 3646 15687 3680
rect 15621 3612 15687 3646
rect 15621 3578 15637 3612
rect 15671 3578 15687 3612
rect 15621 3563 15687 3578
rect 15453 3528 15468 3559
rect 15502 3542 15519 3559
rect 15340 3514 15468 3528
rect 15503 3528 15519 3542
rect 15621 3542 15638 3563
rect 15621 3528 15637 3542
rect 15340 3510 15469 3514
rect 15335 3508 15469 3510
rect 15503 3508 15637 3528
rect 15672 3528 15687 3563
rect 15721 3680 15755 3722
rect 15721 3612 15755 3646
rect 15721 3562 15755 3578
rect 15789 3680 15855 3688
rect 15789 3646 15805 3680
rect 15839 3646 15855 3680
rect 15789 3612 15855 3646
rect 15789 3578 15805 3612
rect 15839 3578 15855 3612
rect 15789 3559 15855 3578
rect 15889 3680 15923 3722
rect 15889 3612 15923 3646
rect 15889 3562 15923 3578
rect 15957 3680 16023 3688
rect 15957 3646 15973 3680
rect 16007 3646 16023 3680
rect 15957 3612 16023 3646
rect 15957 3578 15973 3612
rect 16007 3578 16023 3612
rect 15789 3528 15802 3559
rect 15836 3542 15855 3559
rect 15672 3518 15802 3528
rect 15671 3514 15802 3518
rect 15839 3528 15855 3542
rect 15957 3559 16023 3578
rect 16057 3680 16091 3722
rect 16057 3612 16091 3646
rect 16057 3562 16091 3578
rect 16125 3680 16191 3688
rect 16125 3646 16141 3680
rect 16175 3646 16191 3680
rect 16125 3612 16191 3646
rect 16125 3578 16141 3612
rect 16175 3578 16191 3612
rect 15957 3528 15972 3559
rect 16006 3542 16023 3559
rect 15839 3514 15972 3528
rect 16007 3528 16023 3542
rect 16125 3555 16191 3578
rect 16225 3680 16259 3722
rect 16225 3612 16259 3646
rect 16225 3562 16259 3578
rect 16293 3680 16359 3688
rect 16293 3646 16309 3680
rect 16343 3646 16359 3680
rect 16293 3612 16359 3646
rect 16293 3578 16309 3612
rect 16343 3578 16359 3612
rect 16125 3528 16140 3555
rect 16174 3542 16191 3555
rect 15671 3508 15805 3514
rect 15839 3508 15973 3514
rect 16007 3510 16140 3528
rect 16175 3528 16191 3542
rect 16293 3559 16359 3578
rect 16393 3680 16427 3722
rect 16393 3612 16427 3646
rect 16393 3562 16427 3578
rect 16461 3680 16527 3688
rect 16461 3646 16477 3680
rect 16511 3646 16527 3680
rect 16461 3612 16527 3646
rect 16461 3578 16477 3612
rect 16511 3578 16527 3612
rect 16293 3528 16308 3559
rect 16342 3542 16359 3559
rect 16175 3514 16308 3528
rect 16343 3528 16359 3542
rect 16461 3555 16527 3578
rect 16561 3680 16603 3722
rect 30140 3716 30461 3748
rect 30591 3732 30637 3748
rect 16595 3646 16603 3680
rect 16561 3612 16603 3646
rect 16595 3578 16603 3612
rect 30053 3664 30106 3680
rect 30053 3630 30072 3664
rect 30053 3588 30106 3630
rect 30140 3672 30206 3716
rect 30140 3638 30156 3672
rect 30190 3638 30206 3672
rect 30140 3622 30206 3638
rect 30240 3664 30274 3680
rect 30240 3588 30274 3630
rect 30308 3672 30374 3716
rect 30591 3698 30603 3732
rect 30308 3638 30324 3672
rect 30358 3638 30374 3672
rect 30308 3622 30374 3638
rect 30408 3665 30458 3681
rect 30442 3631 30458 3665
rect 30408 3588 30458 3631
rect 30591 3664 30637 3698
rect 30591 3630 30603 3664
rect 30591 3588 30637 3630
rect 30671 3732 31913 3752
rect 43421 3840 43463 3882
rect 43421 3806 43429 3840
rect 43421 3772 43463 3806
rect 30671 3698 30687 3732
rect 30721 3714 30855 3732
rect 30721 3698 30737 3714
rect 30671 3664 30737 3698
rect 30839 3698 30855 3714
rect 30889 3714 31023 3732
rect 31057 3724 31191 3732
rect 30889 3698 30905 3714
rect 30671 3630 30687 3664
rect 30721 3630 30737 3664
rect 30671 3622 30737 3630
rect 30771 3664 30805 3680
rect 30771 3588 30805 3630
rect 30839 3664 30905 3698
rect 31007 3698 31023 3714
rect 31063 3714 31191 3724
rect 31225 3720 31359 3732
rect 31393 3726 31527 3732
rect 31007 3690 31029 3698
rect 31063 3690 31073 3714
rect 30839 3630 30855 3664
rect 30889 3630 30905 3664
rect 30839 3622 30905 3630
rect 30939 3664 30973 3680
rect 30939 3588 30973 3630
rect 31007 3664 31073 3690
rect 31175 3698 31191 3714
rect 31229 3714 31359 3720
rect 31175 3686 31195 3698
rect 31229 3686 31241 3714
rect 31007 3630 31023 3664
rect 31057 3630 31073 3664
rect 31007 3622 31073 3630
rect 31107 3664 31141 3680
rect 31107 3588 31141 3630
rect 31175 3664 31241 3686
rect 31343 3698 31359 3714
rect 31397 3714 31527 3726
rect 31561 3724 31695 3732
rect 31729 3725 31863 3732
rect 31897 3726 31913 3732
rect 31343 3692 31363 3698
rect 31397 3692 31409 3714
rect 31175 3630 31191 3664
rect 31225 3630 31241 3664
rect 31175 3622 31241 3630
rect 31275 3664 31309 3680
rect 31275 3588 31309 3630
rect 31343 3664 31409 3692
rect 31511 3698 31527 3714
rect 31564 3714 31695 3724
rect 31511 3690 31530 3698
rect 31564 3690 31577 3714
rect 31343 3630 31359 3664
rect 31393 3630 31409 3664
rect 31343 3622 31409 3630
rect 31443 3664 31477 3680
rect 31443 3588 31477 3630
rect 31511 3664 31577 3690
rect 31679 3698 31695 3714
rect 31734 3714 31863 3725
rect 31679 3691 31700 3698
rect 31734 3691 31745 3714
rect 31511 3630 31527 3664
rect 31561 3630 31577 3664
rect 31511 3622 31577 3630
rect 31611 3664 31645 3680
rect 31611 3588 31645 3630
rect 31679 3664 31745 3691
rect 31847 3698 31863 3714
rect 31847 3692 31864 3698
rect 31898 3692 31913 3726
rect 31679 3630 31695 3664
rect 31729 3630 31745 3664
rect 31679 3622 31745 3630
rect 31779 3664 31813 3680
rect 31779 3588 31813 3630
rect 31847 3664 31913 3692
rect 31847 3630 31863 3664
rect 31897 3630 31913 3664
rect 31847 3622 31913 3630
rect 31947 3732 31989 3748
rect 31981 3698 31989 3732
rect 31947 3664 31989 3698
rect 31981 3630 31989 3664
rect 43421 3738 43429 3772
rect 43421 3702 43463 3738
rect 43421 3668 43429 3702
rect 43421 3652 43463 3668
rect 43497 3840 43563 3848
rect 43497 3806 43513 3840
rect 43547 3806 43563 3840
rect 43497 3772 43563 3806
rect 43497 3738 43513 3772
rect 43547 3738 43563 3772
rect 43497 3714 43563 3738
rect 43597 3840 43631 3882
rect 43597 3772 43631 3806
rect 43597 3722 43631 3738
rect 43665 3840 43731 3848
rect 43665 3806 43681 3840
rect 43715 3806 43731 3840
rect 43665 3772 43731 3806
rect 43665 3738 43681 3772
rect 43715 3738 43731 3772
rect 43497 3702 43514 3714
rect 43497 3668 43513 3702
rect 43548 3688 43563 3714
rect 43665 3721 43731 3738
rect 43765 3840 43799 3882
rect 43765 3772 43799 3806
rect 43765 3722 43799 3738
rect 43833 3840 43899 3848
rect 43833 3806 43849 3840
rect 43883 3806 43899 3840
rect 43833 3772 43899 3806
rect 43833 3738 43849 3772
rect 43883 3738 43899 3772
rect 43665 3702 43682 3721
rect 43665 3688 43681 3702
rect 43548 3669 43681 3688
rect 43716 3688 43731 3721
rect 43833 3711 43899 3738
rect 43933 3840 43967 3882
rect 43933 3772 43967 3806
rect 43933 3722 43967 3738
rect 44001 3840 44067 3848
rect 44001 3806 44017 3840
rect 44051 3806 44067 3840
rect 44001 3772 44067 3806
rect 44001 3738 44017 3772
rect 44051 3738 44067 3772
rect 44001 3723 44067 3738
rect 43833 3702 43850 3711
rect 43833 3688 43849 3702
rect 43716 3676 43849 3688
rect 43547 3668 43681 3669
rect 43715 3668 43849 3676
rect 43884 3688 43899 3711
rect 44001 3702 44018 3723
rect 44001 3688 44017 3702
rect 43884 3668 44017 3688
rect 44052 3688 44067 3723
rect 44101 3840 44135 3882
rect 44101 3772 44135 3806
rect 44101 3722 44135 3738
rect 44169 3840 44235 3848
rect 44169 3806 44185 3840
rect 44219 3806 44235 3840
rect 44169 3772 44235 3806
rect 44169 3738 44185 3772
rect 44219 3738 44235 3772
rect 44169 3721 44235 3738
rect 44269 3840 44303 3882
rect 44269 3772 44303 3806
rect 44269 3722 44303 3738
rect 44337 3840 44403 3848
rect 44337 3806 44353 3840
rect 44387 3806 44403 3840
rect 44337 3772 44403 3806
rect 44337 3738 44353 3772
rect 44387 3738 44403 3772
rect 44337 3723 44403 3738
rect 44169 3688 44184 3721
rect 44218 3702 44235 3721
rect 44052 3678 44184 3688
rect 44051 3676 44184 3678
rect 44219 3688 44235 3702
rect 44337 3688 44350 3723
rect 44384 3702 44403 3723
rect 44437 3840 44471 3882
rect 44437 3772 44471 3806
rect 44437 3722 44471 3738
rect 44505 3840 44571 3848
rect 44505 3806 44521 3840
rect 44555 3806 44571 3840
rect 44505 3772 44571 3806
rect 44505 3738 44521 3772
rect 44555 3738 44571 3772
rect 44505 3723 44571 3738
rect 44219 3678 44350 3688
rect 44387 3688 44403 3702
rect 44505 3688 44518 3723
rect 44552 3702 44571 3723
rect 44605 3840 44639 3882
rect 44605 3772 44639 3806
rect 44605 3722 44639 3738
rect 44673 3840 44739 3848
rect 44673 3806 44689 3840
rect 44723 3806 44739 3840
rect 44673 3772 44739 3806
rect 44673 3738 44689 3772
rect 44723 3738 44739 3772
rect 44387 3678 44518 3688
rect 44555 3688 44571 3702
rect 44673 3721 44739 3738
rect 44773 3840 44815 3882
rect 44807 3809 44815 3840
rect 45351 3840 45393 3882
rect 45351 3809 45359 3840
rect 44807 3806 45359 3809
rect 44773 3789 45393 3806
rect 44773 3772 45088 3789
rect 44807 3755 45088 3772
rect 45122 3772 45393 3789
rect 45122 3755 45359 3772
rect 44807 3738 45359 3755
rect 44773 3737 45393 3738
rect 44773 3722 44815 3737
rect 44673 3702 44692 3721
rect 44673 3688 44689 3702
rect 44051 3668 44185 3676
rect 44219 3668 44353 3678
rect 44387 3668 44521 3678
rect 44555 3668 44689 3688
rect 44726 3676 44739 3721
rect 44723 3668 44739 3676
rect 43497 3666 43850 3668
rect 43884 3666 44739 3668
rect 43497 3654 44739 3666
rect 31947 3588 31989 3630
rect 43398 3612 44486 3618
rect 43398 3604 43714 3612
rect 16561 3562 16603 3578
rect 16461 3542 16482 3555
rect 16461 3528 16477 3542
rect 16007 3508 16141 3510
rect 16175 3508 16309 3514
rect 16343 3508 16477 3528
rect 16516 3510 16527 3555
rect 30027 3554 30056 3588
rect 30090 3554 30148 3588
rect 30182 3554 30240 3588
rect 30274 3554 30332 3588
rect 30366 3554 30424 3588
rect 30458 3554 30487 3588
rect 30555 3554 30584 3588
rect 30618 3554 30676 3588
rect 30710 3554 30768 3588
rect 30802 3554 30860 3588
rect 30894 3554 30952 3588
rect 30986 3554 31044 3588
rect 31078 3554 31136 3588
rect 31170 3554 31228 3588
rect 31262 3554 31320 3588
rect 31354 3554 31412 3588
rect 31446 3554 31504 3588
rect 31538 3554 31596 3588
rect 31630 3554 31688 3588
rect 31722 3554 31780 3588
rect 31814 3554 31872 3588
rect 31906 3554 31964 3588
rect 31998 3554 32027 3588
rect 43398 3570 43423 3604
rect 43457 3570 43597 3604
rect 43631 3578 43714 3604
rect 43748 3604 43814 3612
rect 43748 3578 43765 3604
rect 43631 3570 43765 3578
rect 43799 3578 43814 3604
rect 43848 3578 43914 3612
rect 43948 3604 44014 3612
rect 43968 3578 44014 3604
rect 44048 3604 44114 3612
rect 44048 3578 44101 3604
rect 44148 3578 44214 3612
rect 44248 3604 44314 3612
rect 44248 3578 44269 3604
rect 43799 3570 43934 3578
rect 43968 3570 44101 3578
rect 44135 3570 44269 3578
rect 44303 3578 44314 3604
rect 44348 3578 44414 3612
rect 44448 3604 44486 3612
rect 44303 3570 44436 3578
rect 44470 3570 44486 3604
rect 44673 3536 44739 3654
rect 45351 3702 45393 3737
rect 45351 3668 45359 3702
rect 45351 3652 45393 3668
rect 45427 3840 45493 3848
rect 45427 3806 45443 3840
rect 45477 3806 45493 3840
rect 45427 3772 45493 3806
rect 45427 3738 45443 3772
rect 45477 3738 45493 3772
rect 45427 3715 45493 3738
rect 45527 3840 45561 3882
rect 45527 3772 45561 3806
rect 45527 3722 45561 3738
rect 45595 3840 45661 3848
rect 45595 3806 45611 3840
rect 45645 3806 45661 3840
rect 45595 3772 45661 3806
rect 45595 3738 45611 3772
rect 45645 3738 45661 3772
rect 45427 3702 45448 3715
rect 45427 3668 45443 3702
rect 45482 3688 45493 3715
rect 45595 3719 45661 3738
rect 45695 3840 45729 3882
rect 45695 3772 45729 3806
rect 45695 3722 45729 3738
rect 45763 3840 45829 3848
rect 45763 3806 45779 3840
rect 45813 3806 45829 3840
rect 45763 3772 45829 3806
rect 45763 3738 45779 3772
rect 45813 3738 45829 3772
rect 45763 3723 45829 3738
rect 45595 3688 45610 3719
rect 45644 3702 45661 3719
rect 45482 3674 45610 3688
rect 45645 3688 45661 3702
rect 45763 3702 45780 3723
rect 45763 3688 45779 3702
rect 45482 3670 45611 3674
rect 45477 3668 45611 3670
rect 45645 3668 45779 3688
rect 45814 3688 45829 3723
rect 45863 3840 45897 3882
rect 45863 3772 45897 3806
rect 45863 3722 45897 3738
rect 45931 3840 45997 3848
rect 45931 3806 45947 3840
rect 45981 3806 45997 3840
rect 45931 3772 45997 3806
rect 45931 3738 45947 3772
rect 45981 3738 45997 3772
rect 45931 3719 45997 3738
rect 46031 3840 46065 3882
rect 46031 3772 46065 3806
rect 46031 3722 46065 3738
rect 46099 3840 46165 3848
rect 46099 3806 46115 3840
rect 46149 3806 46165 3840
rect 46099 3772 46165 3806
rect 46099 3738 46115 3772
rect 46149 3738 46165 3772
rect 45931 3688 45944 3719
rect 45978 3702 45997 3719
rect 45814 3678 45944 3688
rect 45813 3674 45944 3678
rect 45981 3688 45997 3702
rect 46099 3719 46165 3738
rect 46199 3840 46233 3882
rect 46199 3772 46233 3806
rect 46199 3722 46233 3738
rect 46267 3840 46333 3848
rect 46267 3806 46283 3840
rect 46317 3806 46333 3840
rect 46267 3772 46333 3806
rect 46267 3738 46283 3772
rect 46317 3738 46333 3772
rect 46099 3688 46114 3719
rect 46148 3702 46165 3719
rect 45981 3674 46114 3688
rect 46149 3688 46165 3702
rect 46267 3715 46333 3738
rect 46367 3840 46401 3882
rect 46367 3772 46401 3806
rect 46367 3722 46401 3738
rect 46435 3840 46501 3848
rect 46435 3806 46451 3840
rect 46485 3806 46501 3840
rect 46435 3772 46501 3806
rect 46435 3738 46451 3772
rect 46485 3738 46501 3772
rect 46267 3688 46282 3715
rect 46316 3702 46333 3715
rect 45813 3668 45947 3674
rect 45981 3668 46115 3674
rect 46149 3670 46282 3688
rect 46317 3688 46333 3702
rect 46435 3719 46501 3738
rect 46535 3840 46569 3882
rect 46535 3772 46569 3806
rect 46535 3722 46569 3738
rect 46603 3840 46669 3848
rect 46603 3806 46619 3840
rect 46653 3806 46669 3840
rect 46603 3772 46669 3806
rect 46603 3738 46619 3772
rect 46653 3738 46669 3772
rect 46435 3688 46450 3719
rect 46484 3702 46501 3719
rect 46317 3674 46450 3688
rect 46485 3688 46501 3702
rect 46603 3715 46669 3738
rect 46703 3840 46745 3882
rect 46737 3806 46745 3840
rect 46703 3772 46745 3806
rect 46737 3738 46745 3772
rect 46703 3722 46745 3738
rect 46603 3702 46624 3715
rect 46603 3688 46619 3702
rect 46149 3668 46283 3670
rect 46317 3668 46451 3674
rect 46485 3668 46619 3688
rect 46658 3670 46669 3715
rect 46653 3668 46669 3670
rect 45427 3654 46669 3668
rect 45328 3612 46416 3618
rect 45328 3604 45374 3612
rect 45328 3570 45353 3604
rect 45408 3578 45474 3612
rect 45508 3604 45574 3612
rect 45508 3578 45527 3604
rect 45387 3570 45527 3578
rect 45561 3578 45574 3604
rect 45608 3578 45674 3612
rect 45708 3604 45774 3612
rect 45729 3578 45774 3604
rect 45808 3604 45874 3612
rect 45808 3578 45864 3604
rect 45908 3578 45974 3612
rect 46008 3604 46074 3612
rect 46008 3578 46031 3604
rect 45561 3570 45695 3578
rect 45729 3570 45864 3578
rect 45898 3570 46031 3578
rect 46065 3578 46074 3604
rect 46108 3604 46416 3612
rect 46108 3578 46199 3604
rect 46065 3570 46199 3578
rect 46233 3570 46366 3604
rect 46400 3570 46416 3604
rect 46603 3536 46669 3654
rect 16511 3508 16527 3510
rect 15285 3494 16527 3508
rect 15186 3452 16274 3458
rect 15186 3444 15232 3452
rect 15186 3410 15211 3444
rect 15266 3418 15332 3452
rect 15366 3444 15432 3452
rect 15366 3418 15385 3444
rect 15245 3410 15385 3418
rect 15419 3418 15432 3444
rect 15466 3418 15532 3452
rect 15566 3444 15632 3452
rect 15587 3418 15632 3444
rect 15666 3444 15732 3452
rect 15666 3418 15722 3444
rect 15766 3418 15832 3452
rect 15866 3444 15932 3452
rect 15866 3418 15889 3444
rect 15419 3410 15553 3418
rect 15587 3410 15722 3418
rect 15756 3410 15889 3418
rect 15923 3418 15932 3444
rect 15966 3444 16274 3452
rect 15966 3418 16057 3444
rect 15923 3410 16057 3418
rect 16091 3410 16224 3444
rect 16258 3410 16274 3444
rect 16461 3376 16527 3494
rect 13275 3356 13321 3372
rect 13275 3322 13287 3356
rect 13275 3288 13321 3322
rect 13275 3254 13287 3288
rect 13275 3212 13321 3254
rect 13355 3356 14597 3376
rect 13355 3322 13371 3356
rect 13405 3338 13539 3356
rect 13405 3322 13421 3338
rect 13355 3288 13421 3322
rect 13523 3322 13539 3338
rect 13573 3338 13707 3356
rect 13573 3322 13589 3338
rect 13355 3254 13371 3288
rect 13405 3254 13421 3288
rect 13355 3246 13421 3254
rect 13455 3288 13489 3304
rect 13455 3212 13489 3254
rect 13523 3288 13589 3322
rect 13691 3322 13707 3338
rect 13741 3338 13875 3356
rect 13741 3322 13757 3338
rect 13523 3254 13539 3288
rect 13573 3254 13589 3288
rect 13523 3246 13589 3254
rect 13623 3288 13657 3304
rect 13623 3212 13657 3254
rect 13691 3288 13757 3322
rect 13859 3322 13875 3338
rect 13909 3338 14043 3356
rect 13909 3322 13925 3338
rect 13691 3254 13707 3288
rect 13741 3254 13757 3288
rect 13691 3246 13757 3254
rect 13791 3288 13825 3304
rect 13791 3212 13825 3254
rect 13859 3288 13925 3322
rect 14027 3322 14043 3338
rect 14077 3338 14211 3356
rect 14077 3322 14093 3338
rect 13859 3254 13875 3288
rect 13909 3254 13925 3288
rect 13859 3246 13925 3254
rect 13959 3288 13993 3304
rect 13959 3212 13993 3254
rect 14027 3288 14093 3322
rect 14195 3322 14211 3338
rect 14245 3338 14379 3356
rect 14245 3322 14261 3338
rect 14027 3254 14043 3288
rect 14077 3254 14093 3288
rect 14027 3246 14093 3254
rect 14127 3288 14161 3304
rect 14127 3212 14161 3254
rect 14195 3288 14261 3322
rect 14363 3322 14379 3338
rect 14413 3338 14547 3356
rect 14413 3322 14429 3338
rect 14195 3254 14211 3288
rect 14245 3254 14261 3288
rect 14195 3246 14261 3254
rect 14295 3288 14329 3304
rect 14295 3212 14329 3254
rect 14363 3288 14429 3322
rect 14531 3322 14547 3338
rect 14581 3322 14597 3356
rect 14363 3254 14379 3288
rect 14413 3254 14429 3288
rect 14363 3246 14429 3254
rect 14463 3288 14497 3304
rect 14463 3212 14497 3254
rect 14531 3288 14597 3322
rect 14531 3254 14547 3288
rect 14581 3254 14597 3288
rect 14531 3246 14597 3254
rect 14631 3356 14673 3372
rect 14665 3322 14673 3356
rect 14631 3288 14673 3322
rect 14665 3254 14673 3288
rect 14631 3212 14673 3254
rect 15205 3356 15251 3372
rect 15205 3322 15217 3356
rect 15205 3288 15251 3322
rect 15205 3254 15217 3288
rect 15205 3212 15251 3254
rect 15285 3356 16527 3376
rect 43417 3516 43463 3532
rect 43417 3482 43429 3516
rect 43417 3448 43463 3482
rect 43417 3414 43429 3448
rect 43417 3372 43463 3414
rect 43497 3516 44739 3536
rect 43497 3482 43513 3516
rect 43547 3498 43681 3516
rect 43547 3482 43563 3498
rect 43497 3448 43563 3482
rect 43665 3482 43681 3498
rect 43715 3498 43849 3516
rect 43715 3482 43731 3498
rect 43497 3414 43513 3448
rect 43547 3414 43563 3448
rect 43497 3406 43563 3414
rect 43597 3448 43631 3464
rect 43597 3372 43631 3414
rect 43665 3448 43731 3482
rect 43833 3482 43849 3498
rect 43883 3498 44017 3516
rect 43883 3482 43899 3498
rect 43665 3414 43681 3448
rect 43715 3414 43731 3448
rect 43665 3406 43731 3414
rect 43765 3448 43799 3464
rect 43765 3372 43799 3414
rect 43833 3448 43899 3482
rect 44001 3482 44017 3498
rect 44051 3498 44185 3516
rect 44051 3482 44067 3498
rect 43833 3414 43849 3448
rect 43883 3414 43899 3448
rect 43833 3406 43899 3414
rect 43933 3448 43967 3464
rect 43933 3372 43967 3414
rect 44001 3448 44067 3482
rect 44169 3482 44185 3498
rect 44219 3498 44353 3516
rect 44219 3482 44235 3498
rect 44001 3414 44017 3448
rect 44051 3414 44067 3448
rect 44001 3406 44067 3414
rect 44101 3448 44135 3464
rect 44101 3372 44135 3414
rect 44169 3448 44235 3482
rect 44337 3482 44353 3498
rect 44387 3498 44521 3516
rect 44387 3482 44403 3498
rect 44169 3414 44185 3448
rect 44219 3414 44235 3448
rect 44169 3406 44235 3414
rect 44269 3448 44303 3464
rect 44269 3372 44303 3414
rect 44337 3448 44403 3482
rect 44505 3482 44521 3498
rect 44555 3498 44689 3516
rect 44555 3482 44571 3498
rect 44337 3414 44353 3448
rect 44387 3414 44403 3448
rect 44337 3406 44403 3414
rect 44437 3448 44471 3464
rect 44437 3372 44471 3414
rect 44505 3448 44571 3482
rect 44673 3482 44689 3498
rect 44723 3482 44739 3516
rect 44505 3414 44521 3448
rect 44555 3414 44571 3448
rect 44505 3406 44571 3414
rect 44605 3448 44639 3464
rect 44605 3372 44639 3414
rect 44673 3448 44739 3482
rect 44673 3414 44689 3448
rect 44723 3414 44739 3448
rect 44673 3406 44739 3414
rect 44773 3516 44815 3532
rect 44807 3482 44815 3516
rect 44773 3448 44815 3482
rect 44807 3414 44815 3448
rect 44773 3372 44815 3414
rect 45347 3516 45393 3532
rect 45347 3482 45359 3516
rect 45347 3448 45393 3482
rect 45347 3414 45359 3448
rect 45347 3372 45393 3414
rect 45427 3516 46669 3536
rect 45427 3482 45443 3516
rect 45477 3498 45611 3516
rect 45477 3482 45493 3498
rect 45427 3448 45493 3482
rect 45595 3482 45611 3498
rect 45645 3498 45779 3516
rect 45645 3482 45661 3498
rect 45427 3414 45443 3448
rect 45477 3414 45493 3448
rect 45427 3406 45493 3414
rect 45527 3448 45561 3464
rect 45527 3372 45561 3414
rect 45595 3448 45661 3482
rect 45763 3482 45779 3498
rect 45813 3498 45947 3516
rect 45813 3482 45829 3498
rect 45595 3414 45611 3448
rect 45645 3414 45661 3448
rect 45595 3406 45661 3414
rect 45695 3448 45729 3464
rect 45695 3372 45729 3414
rect 45763 3448 45829 3482
rect 45931 3482 45947 3498
rect 45981 3498 46115 3516
rect 45981 3482 45997 3498
rect 45763 3414 45779 3448
rect 45813 3414 45829 3448
rect 45763 3406 45829 3414
rect 45863 3448 45897 3464
rect 45863 3372 45897 3414
rect 45931 3448 45997 3482
rect 46099 3482 46115 3498
rect 46149 3498 46283 3516
rect 46149 3482 46165 3498
rect 45931 3414 45947 3448
rect 45981 3414 45997 3448
rect 45931 3406 45997 3414
rect 46031 3448 46065 3464
rect 46031 3372 46065 3414
rect 46099 3448 46165 3482
rect 46267 3482 46283 3498
rect 46317 3498 46451 3516
rect 46317 3482 46333 3498
rect 46099 3414 46115 3448
rect 46149 3414 46165 3448
rect 46099 3406 46165 3414
rect 46199 3448 46233 3464
rect 46199 3372 46233 3414
rect 46267 3448 46333 3482
rect 46435 3482 46451 3498
rect 46485 3498 46619 3516
rect 46485 3482 46501 3498
rect 46267 3414 46283 3448
rect 46317 3414 46333 3448
rect 46267 3406 46333 3414
rect 46367 3448 46401 3464
rect 46367 3372 46401 3414
rect 46435 3448 46501 3482
rect 46603 3482 46619 3498
rect 46653 3482 46669 3516
rect 46435 3414 46451 3448
rect 46485 3414 46501 3448
rect 46435 3406 46501 3414
rect 46535 3448 46569 3464
rect 46535 3372 46569 3414
rect 46603 3448 46669 3482
rect 46603 3414 46619 3448
rect 46653 3414 46669 3448
rect 46603 3406 46669 3414
rect 46703 3516 46745 3532
rect 46737 3482 46745 3516
rect 46703 3448 46745 3482
rect 46737 3414 46745 3448
rect 46703 3372 46745 3414
rect 15285 3322 15301 3356
rect 15335 3338 15469 3356
rect 15335 3322 15351 3338
rect 15285 3288 15351 3322
rect 15453 3322 15469 3338
rect 15503 3338 15637 3356
rect 15503 3322 15519 3338
rect 15285 3254 15301 3288
rect 15335 3254 15351 3288
rect 15285 3246 15351 3254
rect 15385 3288 15419 3304
rect 15385 3212 15419 3254
rect 15453 3288 15519 3322
rect 15621 3322 15637 3338
rect 15671 3338 15805 3356
rect 15671 3322 15687 3338
rect 15453 3254 15469 3288
rect 15503 3254 15519 3288
rect 15453 3246 15519 3254
rect 15553 3288 15587 3304
rect 15553 3212 15587 3254
rect 15621 3288 15687 3322
rect 15789 3322 15805 3338
rect 15839 3338 15973 3356
rect 15839 3322 15855 3338
rect 15621 3254 15637 3288
rect 15671 3254 15687 3288
rect 15621 3246 15687 3254
rect 15721 3288 15755 3304
rect 15721 3212 15755 3254
rect 15789 3288 15855 3322
rect 15957 3322 15973 3338
rect 16007 3338 16141 3356
rect 16007 3322 16023 3338
rect 15789 3254 15805 3288
rect 15839 3254 15855 3288
rect 15789 3246 15855 3254
rect 15889 3288 15923 3304
rect 15889 3212 15923 3254
rect 15957 3288 16023 3322
rect 16125 3322 16141 3338
rect 16175 3338 16309 3356
rect 16175 3322 16191 3338
rect 15957 3254 15973 3288
rect 16007 3254 16023 3288
rect 15957 3246 16023 3254
rect 16057 3288 16091 3304
rect 16057 3212 16091 3254
rect 16125 3288 16191 3322
rect 16293 3322 16309 3338
rect 16343 3338 16477 3356
rect 16343 3322 16359 3338
rect 16125 3254 16141 3288
rect 16175 3254 16191 3288
rect 16125 3246 16191 3254
rect 16225 3288 16259 3304
rect 16225 3212 16259 3254
rect 16293 3288 16359 3322
rect 16461 3322 16477 3338
rect 16511 3322 16527 3356
rect 16293 3254 16309 3288
rect 16343 3254 16359 3288
rect 16293 3246 16359 3254
rect 16393 3288 16427 3304
rect 16393 3212 16427 3254
rect 16461 3288 16527 3322
rect 16461 3254 16477 3288
rect 16511 3254 16527 3288
rect 16461 3246 16527 3254
rect 16561 3356 16603 3372
rect 16595 3322 16603 3356
rect 43381 3338 43410 3372
rect 43444 3338 43502 3372
rect 43536 3338 43594 3372
rect 43628 3338 43686 3372
rect 43720 3338 43778 3372
rect 43812 3338 43870 3372
rect 43904 3338 43962 3372
rect 43996 3338 44054 3372
rect 44088 3338 44146 3372
rect 44180 3338 44238 3372
rect 44272 3338 44330 3372
rect 44364 3338 44422 3372
rect 44456 3338 44514 3372
rect 44548 3338 44606 3372
rect 44640 3338 44698 3372
rect 44732 3338 44790 3372
rect 44824 3338 44853 3372
rect 45311 3338 45340 3372
rect 45374 3338 45432 3372
rect 45466 3338 45524 3372
rect 45558 3338 45616 3372
rect 45650 3338 45708 3372
rect 45742 3338 45800 3372
rect 45834 3338 45892 3372
rect 45926 3338 45984 3372
rect 46018 3338 46076 3372
rect 46110 3338 46168 3372
rect 46202 3338 46260 3372
rect 46294 3338 46352 3372
rect 46386 3338 46444 3372
rect 46478 3338 46536 3372
rect 46570 3338 46628 3372
rect 46662 3338 46720 3372
rect 46754 3338 46783 3372
rect 16561 3288 16603 3322
rect 16595 3254 16603 3288
rect 16561 3212 16603 3254
rect 13239 3178 13268 3212
rect 13302 3178 13360 3212
rect 13394 3178 13452 3212
rect 13486 3178 13544 3212
rect 13578 3178 13636 3212
rect 13670 3178 13728 3212
rect 13762 3178 13820 3212
rect 13854 3178 13912 3212
rect 13946 3178 14004 3212
rect 14038 3178 14096 3212
rect 14130 3178 14188 3212
rect 14222 3178 14280 3212
rect 14314 3178 14372 3212
rect 14406 3178 14464 3212
rect 14498 3178 14556 3212
rect 14590 3178 14648 3212
rect 14682 3178 14711 3212
rect 15169 3178 15198 3212
rect 15232 3178 15290 3212
rect 15324 3178 15382 3212
rect 15416 3178 15474 3212
rect 15508 3178 15566 3212
rect 15600 3178 15658 3212
rect 15692 3178 15750 3212
rect 15784 3178 15842 3212
rect 15876 3178 15934 3212
rect 15968 3178 16026 3212
rect 16060 3178 16118 3212
rect 16152 3178 16210 3212
rect 16244 3178 16302 3212
rect 16336 3178 16394 3212
rect 16428 3178 16486 3212
rect 16520 3178 16578 3212
rect 16612 3178 16641 3212
rect 5664 2777 5693 2811
rect 5727 2777 5785 2811
rect 5819 2777 5877 2811
rect 5911 2777 5969 2811
rect 6003 2777 6061 2811
rect 6095 2777 6153 2811
rect 6187 2777 6245 2811
rect 6279 2777 6337 2811
rect 6371 2777 6429 2811
rect 6463 2777 6521 2811
rect 6555 2777 6613 2811
rect 6647 2777 6705 2811
rect 6739 2777 6797 2811
rect 6831 2777 6889 2811
rect 6923 2777 6981 2811
rect 7015 2777 7073 2811
rect 7107 2777 7136 2811
rect 5700 2735 5746 2777
rect 5700 2701 5712 2735
rect 5700 2667 5746 2701
rect 5700 2633 5712 2667
rect 5700 2617 5746 2633
rect 5780 2735 5846 2743
rect 5780 2701 5796 2735
rect 5830 2701 5846 2735
rect 5780 2667 5846 2701
rect 5880 2735 5914 2777
rect 5880 2685 5914 2701
rect 5948 2735 6014 2743
rect 5948 2701 5964 2735
rect 5998 2701 6014 2735
rect 5780 2633 5796 2667
rect 5830 2651 5846 2667
rect 5948 2667 6014 2701
rect 6048 2735 6082 2777
rect 6048 2685 6082 2701
rect 6116 2735 6182 2743
rect 6116 2701 6132 2735
rect 6166 2701 6182 2735
rect 5948 2651 5964 2667
rect 5830 2633 5964 2651
rect 5998 2651 6014 2667
rect 6116 2667 6182 2701
rect 6216 2735 6250 2777
rect 6216 2685 6250 2701
rect 6284 2735 6350 2743
rect 6284 2701 6300 2735
rect 6334 2701 6350 2735
rect 6116 2651 6132 2667
rect 5998 2633 6132 2651
rect 6166 2651 6182 2667
rect 6284 2667 6350 2701
rect 6384 2735 6418 2777
rect 6384 2685 6418 2701
rect 6452 2735 6518 2743
rect 6452 2701 6468 2735
rect 6502 2701 6518 2735
rect 6284 2651 6300 2667
rect 6166 2633 6300 2651
rect 6334 2651 6350 2667
rect 6452 2667 6518 2701
rect 6552 2735 6586 2777
rect 6552 2685 6586 2701
rect 6620 2735 6686 2743
rect 6620 2701 6636 2735
rect 6670 2701 6686 2735
rect 6452 2651 6468 2667
rect 6334 2633 6468 2651
rect 6502 2651 6518 2667
rect 6620 2667 6686 2701
rect 6720 2735 6754 2777
rect 6720 2685 6754 2701
rect 6788 2735 6854 2743
rect 6788 2701 6804 2735
rect 6838 2701 6854 2735
rect 6620 2651 6636 2667
rect 6502 2633 6636 2651
rect 6670 2651 6686 2667
rect 6788 2667 6854 2701
rect 6888 2735 6922 2777
rect 6888 2685 6922 2701
rect 6956 2735 7022 2743
rect 6956 2701 6972 2735
rect 7006 2701 7022 2735
rect 6788 2651 6804 2667
rect 6670 2633 6804 2651
rect 6838 2651 6854 2667
rect 6956 2667 7022 2701
rect 6956 2651 6972 2667
rect 6838 2633 6972 2651
rect 7006 2633 7022 2667
rect 5780 2613 7022 2633
rect 7056 2735 7098 2777
rect 7546 2775 7575 2809
rect 7609 2775 7667 2809
rect 7701 2775 7759 2809
rect 7793 2775 7851 2809
rect 7885 2775 7943 2809
rect 7977 2775 8035 2809
rect 8069 2775 8127 2809
rect 8161 2775 8219 2809
rect 8253 2775 8311 2809
rect 8345 2775 8403 2809
rect 8437 2775 8495 2809
rect 8529 2775 8587 2809
rect 8621 2775 8679 2809
rect 8713 2775 8771 2809
rect 8805 2775 8863 2809
rect 8897 2775 8955 2809
rect 8989 2775 9018 2809
rect 20762 2777 20791 2811
rect 20825 2777 20883 2811
rect 20917 2777 20975 2811
rect 21009 2777 21067 2811
rect 21101 2777 21159 2811
rect 21193 2777 21251 2811
rect 21285 2777 21343 2811
rect 21377 2777 21435 2811
rect 21469 2777 21527 2811
rect 21561 2777 21619 2811
rect 21653 2777 21711 2811
rect 21745 2777 21803 2811
rect 21837 2777 21895 2811
rect 21929 2777 21987 2811
rect 22021 2777 22079 2811
rect 22113 2777 22171 2811
rect 22205 2777 22234 2811
rect 7090 2701 7098 2735
rect 7056 2667 7098 2701
rect 7090 2633 7098 2667
rect 7056 2617 7098 2633
rect 7582 2733 7628 2775
rect 7582 2699 7594 2733
rect 7582 2665 7628 2699
rect 7582 2631 7594 2665
rect 7582 2615 7628 2631
rect 7662 2733 7728 2741
rect 7662 2699 7678 2733
rect 7712 2699 7728 2733
rect 7662 2665 7728 2699
rect 7762 2733 7796 2775
rect 7762 2683 7796 2699
rect 7830 2733 7896 2741
rect 7830 2699 7846 2733
rect 7880 2699 7896 2733
rect 7662 2631 7678 2665
rect 7712 2649 7728 2665
rect 7830 2665 7896 2699
rect 7930 2733 7964 2775
rect 7930 2683 7964 2699
rect 7998 2733 8064 2741
rect 7998 2699 8014 2733
rect 8048 2699 8064 2733
rect 7830 2649 7846 2665
rect 7712 2631 7846 2649
rect 7880 2649 7896 2665
rect 7998 2665 8064 2699
rect 8098 2733 8132 2775
rect 8098 2683 8132 2699
rect 8166 2733 8232 2741
rect 8166 2699 8182 2733
rect 8216 2699 8232 2733
rect 7998 2649 8014 2665
rect 7880 2631 8014 2649
rect 8048 2649 8064 2665
rect 8166 2665 8232 2699
rect 8266 2733 8300 2775
rect 8266 2683 8300 2699
rect 8334 2733 8400 2741
rect 8334 2699 8350 2733
rect 8384 2699 8400 2733
rect 8166 2649 8182 2665
rect 8048 2631 8182 2649
rect 8216 2649 8232 2665
rect 8334 2665 8400 2699
rect 8434 2733 8468 2775
rect 8434 2683 8468 2699
rect 8502 2733 8568 2741
rect 8502 2699 8518 2733
rect 8552 2699 8568 2733
rect 8334 2649 8350 2665
rect 8216 2631 8350 2649
rect 8384 2649 8400 2665
rect 8502 2665 8568 2699
rect 8602 2733 8636 2775
rect 8602 2683 8636 2699
rect 8670 2733 8736 2741
rect 8670 2699 8686 2733
rect 8720 2699 8736 2733
rect 8502 2649 8518 2665
rect 8384 2631 8518 2649
rect 8552 2649 8568 2665
rect 8670 2665 8736 2699
rect 8770 2733 8804 2775
rect 8770 2683 8804 2699
rect 8838 2733 8904 2741
rect 8838 2699 8854 2733
rect 8888 2699 8904 2733
rect 8670 2649 8686 2665
rect 8552 2631 8686 2649
rect 8720 2649 8736 2665
rect 8838 2665 8904 2699
rect 8838 2649 8854 2665
rect 8720 2631 8854 2649
rect 8888 2631 8904 2665
rect 5681 2545 5706 2579
rect 5740 2574 5880 2579
rect 5740 2545 5820 2574
rect 5681 2540 5820 2545
rect 5854 2545 5880 2574
rect 5914 2574 6048 2579
rect 6082 2574 6217 2579
rect 5914 2545 5933 2574
rect 5854 2540 5933 2545
rect 5967 2540 6046 2574
rect 6082 2545 6159 2574
rect 6080 2540 6159 2545
rect 6193 2545 6217 2574
rect 6251 2574 6384 2579
rect 6418 2574 6552 2579
rect 6251 2545 6272 2574
rect 6193 2540 6272 2545
rect 6306 2545 6384 2574
rect 6306 2540 6385 2545
rect 6419 2540 6498 2574
rect 6532 2545 6552 2574
rect 6586 2574 6719 2579
rect 6586 2545 6614 2574
rect 6532 2540 6614 2545
rect 6648 2540 6718 2574
rect 6753 2545 6769 2579
rect 6752 2540 6769 2545
rect 5681 2531 6769 2540
rect 5704 2481 5746 2497
rect 6956 2495 7022 2613
rect 7662 2611 8904 2631
rect 8938 2733 8980 2775
rect 8972 2699 8980 2733
rect 8938 2665 8980 2699
rect 8972 2631 8980 2665
rect 8938 2615 8980 2631
rect 20798 2735 20844 2777
rect 20798 2701 20810 2735
rect 20798 2667 20844 2701
rect 20798 2633 20810 2667
rect 20798 2617 20844 2633
rect 20878 2735 20944 2743
rect 20878 2701 20894 2735
rect 20928 2701 20944 2735
rect 20878 2667 20944 2701
rect 20978 2735 21012 2777
rect 20978 2685 21012 2701
rect 21046 2735 21112 2743
rect 21046 2701 21062 2735
rect 21096 2701 21112 2735
rect 20878 2633 20894 2667
rect 20928 2651 20944 2667
rect 21046 2667 21112 2701
rect 21146 2735 21180 2777
rect 21146 2685 21180 2701
rect 21214 2735 21280 2743
rect 21214 2701 21230 2735
rect 21264 2701 21280 2735
rect 21046 2651 21062 2667
rect 20928 2633 21062 2651
rect 21096 2651 21112 2667
rect 21214 2667 21280 2701
rect 21314 2735 21348 2777
rect 21314 2685 21348 2701
rect 21382 2735 21448 2743
rect 21382 2701 21398 2735
rect 21432 2701 21448 2735
rect 21214 2651 21230 2667
rect 21096 2633 21230 2651
rect 21264 2651 21280 2667
rect 21382 2667 21448 2701
rect 21482 2735 21516 2777
rect 21482 2685 21516 2701
rect 21550 2735 21616 2743
rect 21550 2701 21566 2735
rect 21600 2701 21616 2735
rect 21382 2651 21398 2667
rect 21264 2633 21398 2651
rect 21432 2651 21448 2667
rect 21550 2667 21616 2701
rect 21650 2735 21684 2777
rect 21650 2685 21684 2701
rect 21718 2735 21784 2743
rect 21718 2701 21734 2735
rect 21768 2701 21784 2735
rect 21550 2651 21566 2667
rect 21432 2633 21566 2651
rect 21600 2651 21616 2667
rect 21718 2667 21784 2701
rect 21818 2735 21852 2777
rect 21818 2685 21852 2701
rect 21886 2735 21952 2743
rect 21886 2701 21902 2735
rect 21936 2701 21952 2735
rect 21718 2651 21734 2667
rect 21600 2633 21734 2651
rect 21768 2651 21784 2667
rect 21886 2667 21952 2701
rect 21986 2735 22020 2777
rect 21986 2685 22020 2701
rect 22054 2735 22120 2743
rect 22054 2701 22070 2735
rect 22104 2701 22120 2735
rect 21886 2651 21902 2667
rect 21768 2633 21902 2651
rect 21936 2651 21952 2667
rect 22054 2667 22120 2701
rect 22054 2651 22070 2667
rect 21936 2633 22070 2651
rect 22104 2633 22120 2667
rect 20878 2613 22120 2633
rect 22154 2735 22196 2777
rect 22644 2775 22673 2809
rect 22707 2775 22765 2809
rect 22799 2775 22857 2809
rect 22891 2775 22949 2809
rect 22983 2775 23041 2809
rect 23075 2775 23133 2809
rect 23167 2775 23225 2809
rect 23259 2775 23317 2809
rect 23351 2775 23409 2809
rect 23443 2775 23501 2809
rect 23535 2775 23593 2809
rect 23627 2775 23685 2809
rect 23719 2775 23777 2809
rect 23811 2775 23869 2809
rect 23903 2775 23961 2809
rect 23995 2775 24053 2809
rect 24087 2775 24116 2809
rect 35866 2777 35895 2811
rect 35929 2777 35987 2811
rect 36021 2777 36079 2811
rect 36113 2777 36171 2811
rect 36205 2777 36263 2811
rect 36297 2777 36355 2811
rect 36389 2777 36447 2811
rect 36481 2777 36539 2811
rect 36573 2777 36631 2811
rect 36665 2777 36723 2811
rect 36757 2777 36815 2811
rect 36849 2777 36907 2811
rect 36941 2777 36999 2811
rect 37033 2777 37091 2811
rect 37125 2777 37183 2811
rect 37217 2777 37275 2811
rect 37309 2777 37338 2811
rect 22188 2701 22196 2735
rect 22154 2667 22196 2701
rect 22188 2633 22196 2667
rect 22154 2617 22196 2633
rect 22680 2733 22726 2775
rect 22680 2699 22692 2733
rect 22680 2665 22726 2699
rect 22680 2631 22692 2665
rect 22680 2615 22726 2631
rect 22760 2733 22826 2741
rect 22760 2699 22776 2733
rect 22810 2699 22826 2733
rect 22760 2665 22826 2699
rect 22860 2733 22894 2775
rect 22860 2683 22894 2699
rect 22928 2733 22994 2741
rect 22928 2699 22944 2733
rect 22978 2699 22994 2733
rect 22760 2631 22776 2665
rect 22810 2649 22826 2665
rect 22928 2665 22994 2699
rect 23028 2733 23062 2775
rect 23028 2683 23062 2699
rect 23096 2733 23162 2741
rect 23096 2699 23112 2733
rect 23146 2699 23162 2733
rect 22928 2649 22944 2665
rect 22810 2631 22944 2649
rect 22978 2649 22994 2665
rect 23096 2665 23162 2699
rect 23196 2733 23230 2775
rect 23196 2683 23230 2699
rect 23264 2733 23330 2741
rect 23264 2699 23280 2733
rect 23314 2699 23330 2733
rect 23096 2649 23112 2665
rect 22978 2631 23112 2649
rect 23146 2649 23162 2665
rect 23264 2665 23330 2699
rect 23364 2733 23398 2775
rect 23364 2683 23398 2699
rect 23432 2733 23498 2741
rect 23432 2699 23448 2733
rect 23482 2699 23498 2733
rect 23264 2649 23280 2665
rect 23146 2631 23280 2649
rect 23314 2649 23330 2665
rect 23432 2665 23498 2699
rect 23532 2733 23566 2775
rect 23532 2683 23566 2699
rect 23600 2733 23666 2741
rect 23600 2699 23616 2733
rect 23650 2699 23666 2733
rect 23432 2649 23448 2665
rect 23314 2631 23448 2649
rect 23482 2649 23498 2665
rect 23600 2665 23666 2699
rect 23700 2733 23734 2775
rect 23700 2683 23734 2699
rect 23768 2733 23834 2741
rect 23768 2699 23784 2733
rect 23818 2699 23834 2733
rect 23600 2649 23616 2665
rect 23482 2631 23616 2649
rect 23650 2649 23666 2665
rect 23768 2665 23834 2699
rect 23868 2733 23902 2775
rect 23868 2683 23902 2699
rect 23936 2733 24002 2741
rect 23936 2699 23952 2733
rect 23986 2699 24002 2733
rect 23768 2649 23784 2665
rect 23650 2631 23784 2649
rect 23818 2649 23834 2665
rect 23936 2665 24002 2699
rect 23936 2649 23952 2665
rect 23818 2631 23952 2649
rect 23986 2631 24002 2665
rect 7563 2574 7588 2577
rect 7622 2574 7762 2577
rect 7563 2540 7574 2574
rect 7622 2543 7693 2574
rect 7608 2540 7693 2543
rect 7727 2543 7762 2574
rect 7796 2574 7930 2577
rect 7964 2574 8099 2577
rect 7796 2543 7812 2574
rect 7727 2540 7812 2543
rect 7846 2543 7930 2574
rect 7846 2540 7931 2543
rect 7965 2540 8050 2574
rect 8084 2543 8099 2574
rect 8133 2574 8266 2577
rect 8300 2574 8434 2577
rect 8133 2543 8169 2574
rect 8084 2540 8169 2543
rect 8203 2543 8266 2574
rect 8322 2543 8434 2574
rect 8468 2543 8601 2577
rect 8635 2543 8651 2577
rect 8203 2540 8288 2543
rect 8322 2540 8651 2543
rect 7563 2529 8651 2540
rect 5704 2447 5712 2481
rect 5704 2411 5746 2447
rect 5704 2377 5712 2411
rect 5704 2343 5746 2377
rect 5704 2309 5712 2343
rect 5704 2267 5746 2309
rect 5780 2481 7022 2495
rect 5780 2447 5796 2481
rect 5830 2479 5964 2481
rect 5831 2477 5964 2479
rect 5831 2461 5963 2477
rect 5780 2445 5797 2447
rect 5831 2445 5846 2461
rect 5780 2411 5846 2445
rect 5948 2443 5963 2461
rect 5998 2475 6132 2481
rect 6166 2477 6300 2481
rect 5998 2461 6127 2475
rect 5998 2447 6014 2461
rect 5997 2443 6014 2447
rect 5780 2377 5796 2411
rect 5830 2377 5846 2411
rect 5780 2343 5846 2377
rect 5780 2309 5796 2343
rect 5830 2309 5846 2343
rect 5780 2301 5846 2309
rect 5880 2411 5914 2427
rect 5880 2343 5914 2377
rect 5880 2267 5914 2309
rect 5948 2411 6014 2443
rect 6116 2441 6127 2461
rect 6166 2461 6298 2477
rect 6166 2447 6182 2461
rect 6161 2441 6182 2447
rect 5948 2377 5964 2411
rect 5998 2377 6014 2411
rect 5948 2343 6014 2377
rect 5948 2309 5964 2343
rect 5998 2309 6014 2343
rect 5948 2301 6014 2309
rect 6048 2411 6082 2427
rect 6048 2343 6082 2377
rect 6048 2267 6082 2309
rect 6116 2411 6182 2441
rect 6284 2443 6298 2461
rect 6334 2473 6468 2481
rect 6334 2461 6467 2473
rect 6334 2447 6350 2461
rect 6332 2443 6350 2447
rect 6116 2377 6132 2411
rect 6166 2377 6182 2411
rect 6116 2343 6182 2377
rect 6116 2309 6132 2343
rect 6166 2309 6182 2343
rect 6116 2301 6182 2309
rect 6216 2411 6250 2427
rect 6216 2343 6250 2377
rect 6216 2267 6250 2309
rect 6284 2411 6350 2443
rect 6452 2439 6467 2461
rect 6502 2461 6636 2481
rect 6670 2478 6804 2481
rect 6502 2447 6518 2461
rect 6501 2439 6518 2447
rect 6284 2377 6300 2411
rect 6334 2377 6350 2411
rect 6284 2343 6350 2377
rect 6284 2309 6300 2343
rect 6334 2309 6350 2343
rect 6284 2301 6350 2309
rect 6384 2411 6418 2427
rect 6384 2343 6418 2377
rect 6384 2267 6418 2309
rect 6452 2411 6518 2439
rect 6620 2438 6636 2461
rect 6670 2461 6802 2478
rect 6670 2438 6686 2461
rect 6452 2377 6468 2411
rect 6502 2377 6518 2411
rect 6452 2343 6518 2377
rect 6452 2309 6468 2343
rect 6502 2309 6518 2343
rect 6452 2301 6518 2309
rect 6552 2411 6586 2427
rect 6552 2343 6586 2377
rect 6552 2267 6586 2309
rect 6620 2411 6686 2438
rect 6788 2444 6802 2461
rect 6838 2461 6972 2481
rect 6838 2447 6854 2461
rect 6836 2444 6854 2447
rect 6620 2377 6636 2411
rect 6670 2377 6686 2411
rect 6620 2343 6686 2377
rect 6620 2309 6636 2343
rect 6670 2309 6686 2343
rect 6620 2301 6686 2309
rect 6720 2411 6754 2427
rect 6720 2343 6754 2377
rect 6720 2267 6754 2309
rect 6788 2411 6854 2444
rect 6956 2446 6972 2461
rect 7006 2446 7022 2481
rect 6788 2377 6804 2411
rect 6838 2377 6854 2411
rect 6788 2343 6854 2377
rect 6788 2309 6804 2343
rect 6838 2309 6854 2343
rect 6788 2301 6854 2309
rect 6888 2411 6922 2427
rect 6888 2343 6922 2377
rect 6888 2267 6922 2309
rect 6956 2411 7022 2446
rect 7586 2479 7628 2495
rect 8838 2493 8904 2611
rect 20779 2545 20804 2579
rect 20838 2545 20978 2579
rect 21012 2574 21146 2579
rect 20779 2540 20986 2545
rect 21020 2540 21083 2574
rect 21117 2545 21146 2574
rect 21180 2574 21315 2579
rect 21117 2540 21180 2545
rect 21214 2540 21277 2574
rect 21311 2545 21315 2574
rect 21349 2574 21482 2579
rect 21516 2574 21650 2579
rect 21684 2574 21817 2579
rect 21349 2545 21374 2574
rect 21311 2540 21374 2545
rect 21408 2540 21471 2574
rect 21516 2545 21568 2574
rect 21505 2540 21568 2545
rect 21602 2545 21650 2574
rect 21602 2540 21665 2545
rect 21699 2540 21816 2574
rect 21851 2545 21867 2579
rect 21850 2540 21867 2545
rect 20779 2531 21867 2540
rect 7586 2445 7594 2479
rect 6956 2377 6972 2411
rect 7006 2377 7022 2411
rect 6956 2343 7022 2377
rect 6956 2309 6972 2343
rect 7006 2309 7022 2343
rect 6956 2301 7022 2309
rect 7056 2411 7098 2427
rect 7090 2377 7098 2411
rect 7056 2343 7098 2377
rect 7090 2309 7098 2343
rect 7056 2267 7098 2309
rect 7586 2409 7628 2445
rect 7586 2375 7594 2409
rect 7586 2341 7628 2375
rect 7586 2307 7594 2341
rect 5664 2233 5693 2267
rect 5727 2233 5785 2267
rect 5819 2233 5877 2267
rect 5911 2233 5969 2267
rect 6003 2233 6061 2267
rect 6095 2233 6153 2267
rect 6187 2233 6245 2267
rect 6279 2233 6337 2267
rect 6371 2233 6429 2267
rect 6463 2233 6521 2267
rect 6555 2233 6613 2267
rect 6647 2233 6705 2267
rect 6739 2233 6797 2267
rect 6831 2233 6889 2267
rect 6923 2233 6981 2267
rect 7015 2233 7073 2267
rect 7107 2233 7136 2267
rect 7586 2265 7628 2307
rect 7662 2481 8904 2493
rect 7662 2479 8182 2481
rect 8216 2479 8904 2481
rect 7662 2445 7678 2479
rect 7712 2477 7846 2479
rect 7720 2459 7846 2477
rect 7662 2443 7686 2445
rect 7720 2443 7728 2459
rect 7662 2409 7728 2443
rect 7830 2443 7846 2459
rect 7880 2471 8014 2479
rect 7880 2459 8013 2471
rect 7880 2443 7896 2459
rect 7662 2375 7678 2409
rect 7712 2375 7728 2409
rect 7662 2341 7728 2375
rect 7662 2307 7678 2341
rect 7712 2307 7728 2341
rect 7662 2299 7728 2307
rect 7762 2409 7796 2425
rect 7762 2341 7796 2375
rect 7762 2265 7796 2307
rect 7830 2409 7896 2443
rect 7998 2437 8013 2459
rect 8048 2459 8182 2479
rect 8048 2445 8064 2459
rect 8047 2437 8064 2445
rect 7830 2375 7846 2409
rect 7880 2375 7896 2409
rect 7830 2341 7896 2375
rect 7830 2307 7846 2341
rect 7880 2307 7896 2341
rect 7830 2299 7896 2307
rect 7930 2409 7964 2425
rect 7930 2341 7964 2375
rect 7930 2265 7964 2307
rect 7998 2409 8064 2437
rect 8166 2445 8182 2459
rect 8216 2468 8350 2479
rect 8384 2474 8518 2479
rect 8216 2459 8346 2468
rect 8216 2445 8232 2459
rect 7998 2375 8014 2409
rect 8048 2375 8064 2409
rect 7998 2341 8064 2375
rect 7998 2307 8014 2341
rect 8048 2307 8064 2341
rect 7998 2299 8064 2307
rect 8098 2409 8132 2425
rect 8098 2341 8132 2375
rect 8098 2265 8132 2307
rect 8166 2409 8232 2445
rect 8334 2434 8346 2459
rect 8384 2459 8516 2474
rect 8384 2445 8400 2459
rect 8380 2434 8400 2445
rect 8166 2375 8182 2409
rect 8216 2375 8232 2409
rect 8166 2341 8232 2375
rect 8166 2307 8182 2341
rect 8216 2307 8232 2341
rect 8166 2299 8232 2307
rect 8266 2409 8300 2425
rect 8266 2341 8300 2375
rect 8266 2265 8300 2307
rect 8334 2409 8400 2434
rect 8502 2440 8516 2459
rect 8552 2459 8686 2479
rect 8720 2478 8854 2479
rect 8552 2445 8568 2459
rect 8550 2440 8568 2445
rect 8334 2375 8350 2409
rect 8384 2375 8400 2409
rect 8334 2341 8400 2375
rect 8334 2307 8350 2341
rect 8384 2307 8400 2341
rect 8334 2299 8400 2307
rect 8434 2409 8468 2425
rect 8434 2341 8468 2375
rect 8434 2265 8468 2307
rect 8502 2409 8568 2440
rect 8670 2442 8686 2459
rect 8720 2459 8845 2478
rect 8720 2442 8736 2459
rect 8502 2375 8518 2409
rect 8552 2375 8568 2409
rect 8502 2341 8568 2375
rect 8502 2307 8518 2341
rect 8552 2307 8568 2341
rect 8502 2299 8568 2307
rect 8602 2409 8636 2425
rect 8602 2341 8636 2375
rect 8602 2265 8636 2307
rect 8670 2409 8736 2442
rect 8838 2444 8845 2459
rect 8888 2445 8904 2479
rect 8879 2444 8904 2445
rect 8670 2375 8686 2409
rect 8720 2375 8736 2409
rect 8670 2341 8736 2375
rect 8670 2307 8686 2341
rect 8720 2307 8736 2341
rect 8670 2299 8736 2307
rect 8770 2409 8804 2425
rect 8770 2341 8804 2375
rect 8770 2265 8804 2307
rect 8838 2409 8904 2444
rect 20802 2481 20844 2497
rect 22054 2495 22120 2613
rect 22760 2611 24002 2631
rect 24036 2733 24078 2775
rect 24070 2699 24078 2733
rect 24036 2665 24078 2699
rect 24070 2631 24078 2665
rect 24036 2615 24078 2631
rect 35902 2735 35948 2777
rect 35902 2701 35914 2735
rect 35902 2667 35948 2701
rect 35902 2633 35914 2667
rect 35902 2617 35948 2633
rect 35982 2735 36048 2743
rect 35982 2701 35998 2735
rect 36032 2701 36048 2735
rect 35982 2667 36048 2701
rect 36082 2735 36116 2777
rect 36082 2685 36116 2701
rect 36150 2735 36216 2743
rect 36150 2701 36166 2735
rect 36200 2701 36216 2735
rect 35982 2633 35998 2667
rect 36032 2651 36048 2667
rect 36150 2667 36216 2701
rect 36250 2735 36284 2777
rect 36250 2685 36284 2701
rect 36318 2735 36384 2743
rect 36318 2701 36334 2735
rect 36368 2701 36384 2735
rect 36150 2651 36166 2667
rect 36032 2633 36166 2651
rect 36200 2651 36216 2667
rect 36318 2667 36384 2701
rect 36418 2735 36452 2777
rect 36418 2685 36452 2701
rect 36486 2735 36552 2743
rect 36486 2701 36502 2735
rect 36536 2701 36552 2735
rect 36318 2651 36334 2667
rect 36200 2633 36334 2651
rect 36368 2651 36384 2667
rect 36486 2667 36552 2701
rect 36586 2735 36620 2777
rect 36586 2685 36620 2701
rect 36654 2735 36720 2743
rect 36654 2701 36670 2735
rect 36704 2701 36720 2735
rect 36486 2651 36502 2667
rect 36368 2633 36502 2651
rect 36536 2651 36552 2667
rect 36654 2667 36720 2701
rect 36754 2735 36788 2777
rect 36754 2685 36788 2701
rect 36822 2735 36888 2743
rect 36822 2701 36838 2735
rect 36872 2701 36888 2735
rect 36654 2651 36670 2667
rect 36536 2633 36670 2651
rect 36704 2651 36720 2667
rect 36822 2667 36888 2701
rect 36922 2735 36956 2777
rect 36922 2685 36956 2701
rect 36990 2735 37056 2743
rect 36990 2701 37006 2735
rect 37040 2701 37056 2735
rect 36822 2651 36838 2667
rect 36704 2633 36838 2651
rect 36872 2651 36888 2667
rect 36990 2667 37056 2701
rect 37090 2735 37124 2777
rect 37090 2685 37124 2701
rect 37158 2735 37224 2743
rect 37158 2701 37174 2735
rect 37208 2701 37224 2735
rect 36990 2651 37006 2667
rect 36872 2633 37006 2651
rect 37040 2651 37056 2667
rect 37158 2667 37224 2701
rect 37158 2651 37174 2667
rect 37040 2633 37174 2651
rect 37208 2633 37224 2667
rect 35982 2613 37224 2633
rect 37258 2735 37300 2777
rect 37748 2775 37777 2809
rect 37811 2775 37869 2809
rect 37903 2775 37961 2809
rect 37995 2775 38053 2809
rect 38087 2775 38145 2809
rect 38179 2775 38237 2809
rect 38271 2775 38329 2809
rect 38363 2775 38421 2809
rect 38455 2775 38513 2809
rect 38547 2775 38605 2809
rect 38639 2775 38697 2809
rect 38731 2775 38789 2809
rect 38823 2775 38881 2809
rect 38915 2775 38973 2809
rect 39007 2775 39065 2809
rect 39099 2775 39157 2809
rect 39191 2775 39220 2809
rect 50964 2777 50993 2811
rect 51027 2777 51085 2811
rect 51119 2777 51177 2811
rect 51211 2777 51269 2811
rect 51303 2777 51361 2811
rect 51395 2777 51453 2811
rect 51487 2777 51545 2811
rect 51579 2777 51637 2811
rect 51671 2777 51729 2811
rect 51763 2777 51821 2811
rect 51855 2777 51913 2811
rect 51947 2777 52005 2811
rect 52039 2777 52097 2811
rect 52131 2777 52189 2811
rect 52223 2777 52281 2811
rect 52315 2777 52373 2811
rect 52407 2777 52436 2811
rect 37292 2701 37300 2735
rect 37258 2667 37300 2701
rect 37292 2633 37300 2667
rect 37258 2617 37300 2633
rect 37784 2733 37830 2775
rect 37784 2699 37796 2733
rect 37784 2665 37830 2699
rect 37784 2631 37796 2665
rect 37784 2615 37830 2631
rect 37864 2733 37930 2741
rect 37864 2699 37880 2733
rect 37914 2699 37930 2733
rect 37864 2665 37930 2699
rect 37964 2733 37998 2775
rect 37964 2683 37998 2699
rect 38032 2733 38098 2741
rect 38032 2699 38048 2733
rect 38082 2699 38098 2733
rect 37864 2631 37880 2665
rect 37914 2649 37930 2665
rect 38032 2665 38098 2699
rect 38132 2733 38166 2775
rect 38132 2683 38166 2699
rect 38200 2733 38266 2741
rect 38200 2699 38216 2733
rect 38250 2699 38266 2733
rect 38032 2649 38048 2665
rect 37914 2631 38048 2649
rect 38082 2649 38098 2665
rect 38200 2665 38266 2699
rect 38300 2733 38334 2775
rect 38300 2683 38334 2699
rect 38368 2733 38434 2741
rect 38368 2699 38384 2733
rect 38418 2699 38434 2733
rect 38200 2649 38216 2665
rect 38082 2631 38216 2649
rect 38250 2649 38266 2665
rect 38368 2665 38434 2699
rect 38468 2733 38502 2775
rect 38468 2683 38502 2699
rect 38536 2733 38602 2741
rect 38536 2699 38552 2733
rect 38586 2699 38602 2733
rect 38368 2649 38384 2665
rect 38250 2631 38384 2649
rect 38418 2649 38434 2665
rect 38536 2665 38602 2699
rect 38636 2733 38670 2775
rect 38636 2683 38670 2699
rect 38704 2733 38770 2741
rect 38704 2699 38720 2733
rect 38754 2699 38770 2733
rect 38536 2649 38552 2665
rect 38418 2631 38552 2649
rect 38586 2649 38602 2665
rect 38704 2665 38770 2699
rect 38804 2733 38838 2775
rect 38804 2683 38838 2699
rect 38872 2733 38938 2741
rect 38872 2699 38888 2733
rect 38922 2699 38938 2733
rect 38704 2649 38720 2665
rect 38586 2631 38720 2649
rect 38754 2649 38770 2665
rect 38872 2665 38938 2699
rect 38972 2733 39006 2775
rect 38972 2683 39006 2699
rect 39040 2733 39106 2741
rect 39040 2699 39056 2733
rect 39090 2699 39106 2733
rect 38872 2649 38888 2665
rect 38754 2631 38888 2649
rect 38922 2649 38938 2665
rect 39040 2665 39106 2699
rect 39040 2649 39056 2665
rect 38922 2631 39056 2649
rect 39090 2631 39106 2665
rect 22661 2574 22686 2577
rect 22720 2574 22860 2577
rect 22894 2574 23028 2577
rect 23062 2574 23197 2577
rect 23231 2574 23364 2577
rect 22661 2540 22672 2574
rect 22720 2543 22780 2574
rect 22706 2540 22780 2543
rect 22814 2543 22860 2574
rect 22814 2540 22888 2543
rect 22922 2540 22996 2574
rect 23062 2543 23104 2574
rect 23030 2540 23104 2543
rect 23138 2543 23197 2574
rect 23138 2540 23212 2543
rect 23246 2540 23320 2574
rect 23354 2543 23364 2574
rect 23398 2574 23532 2577
rect 23398 2543 23428 2574
rect 23354 2540 23428 2543
rect 23462 2543 23532 2574
rect 23566 2543 23699 2577
rect 23733 2543 23749 2577
rect 23462 2540 23749 2543
rect 22661 2529 23749 2540
rect 20802 2447 20810 2481
rect 8838 2375 8854 2409
rect 8888 2375 8904 2409
rect 8838 2341 8904 2375
rect 8838 2307 8854 2341
rect 8888 2307 8904 2341
rect 8838 2299 8904 2307
rect 8938 2409 8980 2425
rect 8972 2375 8980 2409
rect 8938 2341 8980 2375
rect 8972 2307 8980 2341
rect 8938 2265 8980 2307
rect 20802 2411 20844 2447
rect 20802 2377 20810 2411
rect 20802 2343 20844 2377
rect 20802 2309 20810 2343
rect 20802 2267 20844 2309
rect 20878 2481 22120 2495
rect 20878 2447 20894 2481
rect 20928 2473 21062 2481
rect 20929 2468 21062 2473
rect 20929 2461 21058 2468
rect 20878 2439 20895 2447
rect 20929 2439 20944 2461
rect 20878 2411 20944 2439
rect 21046 2434 21058 2461
rect 21096 2461 21230 2481
rect 21264 2477 21398 2481
rect 21264 2472 21396 2477
rect 21096 2447 21112 2461
rect 21092 2434 21112 2447
rect 20878 2377 20894 2411
rect 20928 2377 20944 2411
rect 20878 2343 20944 2377
rect 20878 2309 20894 2343
rect 20928 2309 20944 2343
rect 20878 2301 20944 2309
rect 20978 2411 21012 2427
rect 20978 2343 21012 2377
rect 20978 2267 21012 2309
rect 21046 2411 21112 2434
rect 21214 2447 21230 2461
rect 21265 2461 21396 2472
rect 21214 2438 21231 2447
rect 21265 2438 21280 2461
rect 21046 2377 21062 2411
rect 21096 2377 21112 2411
rect 21046 2343 21112 2377
rect 21046 2309 21062 2343
rect 21096 2309 21112 2343
rect 21046 2301 21112 2309
rect 21146 2411 21180 2427
rect 21146 2343 21180 2377
rect 21146 2267 21180 2309
rect 21214 2411 21280 2438
rect 21382 2443 21396 2461
rect 21432 2464 21566 2481
rect 21432 2461 21563 2464
rect 21432 2447 21448 2461
rect 21430 2443 21448 2447
rect 21214 2377 21230 2411
rect 21264 2377 21280 2411
rect 21214 2343 21280 2377
rect 21214 2309 21230 2343
rect 21264 2309 21280 2343
rect 21214 2301 21280 2309
rect 21314 2411 21348 2427
rect 21314 2343 21348 2377
rect 21314 2267 21348 2309
rect 21382 2411 21448 2443
rect 21550 2430 21563 2461
rect 21600 2462 21734 2481
rect 21768 2471 21902 2481
rect 21600 2461 21731 2462
rect 21600 2447 21616 2461
rect 21597 2430 21616 2447
rect 21382 2377 21398 2411
rect 21432 2377 21448 2411
rect 21382 2343 21448 2377
rect 21382 2309 21398 2343
rect 21432 2309 21448 2343
rect 21382 2301 21448 2309
rect 21482 2411 21516 2427
rect 21482 2343 21516 2377
rect 21482 2267 21516 2309
rect 21550 2411 21616 2430
rect 21718 2428 21731 2461
rect 21768 2461 21901 2471
rect 21768 2447 21784 2461
rect 21765 2428 21784 2447
rect 21550 2377 21566 2411
rect 21600 2377 21616 2411
rect 21550 2343 21616 2377
rect 21550 2309 21566 2343
rect 21600 2309 21616 2343
rect 21550 2301 21616 2309
rect 21650 2411 21684 2427
rect 21650 2343 21684 2377
rect 21650 2267 21684 2309
rect 21718 2411 21784 2428
rect 21886 2437 21901 2461
rect 21936 2461 22070 2481
rect 21936 2447 21952 2461
rect 21935 2437 21952 2447
rect 21718 2377 21734 2411
rect 21768 2377 21784 2411
rect 21718 2343 21784 2377
rect 21718 2309 21734 2343
rect 21768 2309 21784 2343
rect 21718 2301 21784 2309
rect 21818 2411 21852 2427
rect 21818 2343 21852 2377
rect 21818 2267 21852 2309
rect 21886 2411 21952 2437
rect 22054 2447 22070 2461
rect 22104 2447 22120 2481
rect 21886 2377 21902 2411
rect 21936 2377 21952 2411
rect 21886 2343 21952 2377
rect 21886 2309 21902 2343
rect 21936 2309 21952 2343
rect 21886 2301 21952 2309
rect 21986 2411 22020 2427
rect 21986 2343 22020 2377
rect 21986 2267 22020 2309
rect 22054 2411 22120 2447
rect 22684 2479 22726 2495
rect 23936 2493 24002 2611
rect 35883 2545 35908 2579
rect 35942 2574 36082 2579
rect 35942 2545 36022 2574
rect 35883 2540 36022 2545
rect 36056 2545 36082 2574
rect 36116 2574 36250 2579
rect 36284 2574 36419 2579
rect 36116 2545 36135 2574
rect 36056 2540 36135 2545
rect 36169 2540 36248 2574
rect 36284 2545 36361 2574
rect 36282 2540 36361 2545
rect 36395 2545 36419 2574
rect 36453 2574 36586 2579
rect 36620 2574 36754 2579
rect 36453 2545 36474 2574
rect 36395 2540 36474 2545
rect 36508 2545 36586 2574
rect 36508 2540 36587 2545
rect 36621 2540 36700 2574
rect 36734 2545 36754 2574
rect 36788 2574 36921 2579
rect 36788 2545 36816 2574
rect 36734 2540 36816 2545
rect 36850 2540 36920 2574
rect 36955 2545 36971 2579
rect 36954 2540 36971 2545
rect 35883 2531 36971 2540
rect 22684 2445 22692 2479
rect 22054 2377 22070 2411
rect 22104 2377 22120 2411
rect 22054 2343 22120 2377
rect 22054 2309 22070 2343
rect 22104 2309 22120 2343
rect 22054 2301 22120 2309
rect 22154 2411 22196 2427
rect 22188 2377 22196 2411
rect 22154 2343 22196 2377
rect 22188 2309 22196 2343
rect 22154 2267 22196 2309
rect 22684 2409 22726 2445
rect 22684 2375 22692 2409
rect 22684 2341 22726 2375
rect 22684 2307 22692 2341
rect 7546 2231 7575 2265
rect 7609 2231 7667 2265
rect 7701 2231 7759 2265
rect 7793 2231 7851 2265
rect 7885 2231 7943 2265
rect 7977 2231 8035 2265
rect 8069 2231 8127 2265
rect 8161 2231 8219 2265
rect 8253 2231 8311 2265
rect 8345 2231 8403 2265
rect 8437 2231 8495 2265
rect 8529 2231 8587 2265
rect 8621 2231 8679 2265
rect 8713 2231 8771 2265
rect 8805 2231 8863 2265
rect 8897 2231 8955 2265
rect 8989 2231 9018 2265
rect 20762 2233 20791 2267
rect 20825 2233 20883 2267
rect 20917 2233 20975 2267
rect 21009 2233 21067 2267
rect 21101 2233 21159 2267
rect 21193 2233 21251 2267
rect 21285 2233 21343 2267
rect 21377 2233 21435 2267
rect 21469 2233 21527 2267
rect 21561 2233 21619 2267
rect 21653 2233 21711 2267
rect 21745 2233 21803 2267
rect 21837 2233 21895 2267
rect 21929 2233 21987 2267
rect 22021 2233 22079 2267
rect 22113 2233 22171 2267
rect 22205 2233 22234 2267
rect 22684 2265 22726 2307
rect 22760 2481 24002 2493
rect 22760 2479 23280 2481
rect 23314 2479 24002 2481
rect 22760 2472 22776 2479
rect 22760 2438 22774 2472
rect 22810 2459 22944 2479
rect 22978 2478 23112 2479
rect 22978 2473 23109 2478
rect 22810 2445 22826 2459
rect 22808 2438 22826 2445
rect 22760 2409 22826 2438
rect 22928 2445 22944 2459
rect 22981 2459 23109 2473
rect 22928 2439 22947 2445
rect 22981 2439 22994 2459
rect 22760 2375 22776 2409
rect 22810 2375 22826 2409
rect 22760 2341 22826 2375
rect 22760 2307 22776 2341
rect 22810 2307 22826 2341
rect 22760 2299 22826 2307
rect 22860 2409 22894 2425
rect 22860 2341 22894 2375
rect 22860 2265 22894 2307
rect 22928 2409 22994 2439
rect 23096 2444 23109 2459
rect 23146 2459 23280 2479
rect 23146 2445 23162 2459
rect 23143 2444 23162 2445
rect 22928 2375 22944 2409
rect 22978 2375 22994 2409
rect 22928 2341 22994 2375
rect 22928 2307 22944 2341
rect 22978 2307 22994 2341
rect 22928 2299 22994 2307
rect 23028 2409 23062 2425
rect 23028 2341 23062 2375
rect 23028 2265 23062 2307
rect 23096 2409 23162 2444
rect 23264 2445 23280 2459
rect 23314 2459 23448 2479
rect 23482 2467 23616 2479
rect 23314 2445 23330 2459
rect 23096 2375 23112 2409
rect 23146 2375 23162 2409
rect 23096 2341 23162 2375
rect 23096 2307 23112 2341
rect 23146 2307 23162 2341
rect 23096 2299 23162 2307
rect 23196 2409 23230 2425
rect 23196 2341 23230 2375
rect 23196 2265 23230 2307
rect 23264 2409 23330 2445
rect 23432 2445 23448 2459
rect 23483 2459 23614 2467
rect 23432 2433 23449 2445
rect 23483 2433 23498 2459
rect 23264 2375 23280 2409
rect 23314 2375 23330 2409
rect 23264 2341 23330 2375
rect 23264 2307 23280 2341
rect 23314 2307 23330 2341
rect 23264 2299 23330 2307
rect 23364 2409 23398 2425
rect 23364 2341 23398 2375
rect 23364 2265 23398 2307
rect 23432 2409 23498 2433
rect 23600 2433 23614 2459
rect 23650 2459 23784 2479
rect 23818 2469 23952 2479
rect 23650 2445 23666 2459
rect 23648 2433 23666 2445
rect 23432 2375 23448 2409
rect 23482 2375 23498 2409
rect 23432 2341 23498 2375
rect 23432 2307 23448 2341
rect 23482 2307 23498 2341
rect 23432 2299 23498 2307
rect 23532 2409 23566 2425
rect 23532 2341 23566 2375
rect 23532 2265 23566 2307
rect 23600 2409 23666 2433
rect 23768 2431 23784 2459
rect 23818 2459 23947 2469
rect 23818 2431 23834 2459
rect 23600 2375 23616 2409
rect 23650 2375 23666 2409
rect 23600 2341 23666 2375
rect 23600 2307 23616 2341
rect 23650 2307 23666 2341
rect 23600 2299 23666 2307
rect 23700 2409 23734 2425
rect 23700 2341 23734 2375
rect 23700 2265 23734 2307
rect 23768 2409 23834 2431
rect 23936 2435 23947 2459
rect 23986 2445 24002 2479
rect 23981 2435 24002 2445
rect 23768 2375 23784 2409
rect 23818 2375 23834 2409
rect 23768 2341 23834 2375
rect 23768 2307 23784 2341
rect 23818 2307 23834 2341
rect 23768 2299 23834 2307
rect 23868 2409 23902 2425
rect 23868 2341 23902 2375
rect 23868 2265 23902 2307
rect 23936 2409 24002 2435
rect 35906 2481 35948 2497
rect 37158 2495 37224 2613
rect 37864 2611 39106 2631
rect 39140 2733 39182 2775
rect 39174 2699 39182 2733
rect 39140 2665 39182 2699
rect 39174 2631 39182 2665
rect 39140 2615 39182 2631
rect 51000 2735 51046 2777
rect 51000 2701 51012 2735
rect 51000 2667 51046 2701
rect 51000 2633 51012 2667
rect 51000 2617 51046 2633
rect 51080 2735 51146 2743
rect 51080 2701 51096 2735
rect 51130 2701 51146 2735
rect 51080 2667 51146 2701
rect 51180 2735 51214 2777
rect 51180 2685 51214 2701
rect 51248 2735 51314 2743
rect 51248 2701 51264 2735
rect 51298 2701 51314 2735
rect 51080 2633 51096 2667
rect 51130 2651 51146 2667
rect 51248 2667 51314 2701
rect 51348 2735 51382 2777
rect 51348 2685 51382 2701
rect 51416 2735 51482 2743
rect 51416 2701 51432 2735
rect 51466 2701 51482 2735
rect 51248 2651 51264 2667
rect 51130 2633 51264 2651
rect 51298 2651 51314 2667
rect 51416 2667 51482 2701
rect 51516 2735 51550 2777
rect 51516 2685 51550 2701
rect 51584 2735 51650 2743
rect 51584 2701 51600 2735
rect 51634 2701 51650 2735
rect 51416 2651 51432 2667
rect 51298 2633 51432 2651
rect 51466 2651 51482 2667
rect 51584 2667 51650 2701
rect 51684 2735 51718 2777
rect 51684 2685 51718 2701
rect 51752 2735 51818 2743
rect 51752 2701 51768 2735
rect 51802 2701 51818 2735
rect 51584 2651 51600 2667
rect 51466 2633 51600 2651
rect 51634 2651 51650 2667
rect 51752 2667 51818 2701
rect 51852 2735 51886 2777
rect 51852 2685 51886 2701
rect 51920 2735 51986 2743
rect 51920 2701 51936 2735
rect 51970 2701 51986 2735
rect 51752 2651 51768 2667
rect 51634 2633 51768 2651
rect 51802 2651 51818 2667
rect 51920 2667 51986 2701
rect 52020 2735 52054 2777
rect 52020 2685 52054 2701
rect 52088 2735 52154 2743
rect 52088 2701 52104 2735
rect 52138 2701 52154 2735
rect 51920 2651 51936 2667
rect 51802 2633 51936 2651
rect 51970 2651 51986 2667
rect 52088 2667 52154 2701
rect 52188 2735 52222 2777
rect 52188 2685 52222 2701
rect 52256 2735 52322 2743
rect 52256 2701 52272 2735
rect 52306 2701 52322 2735
rect 52088 2651 52104 2667
rect 51970 2633 52104 2651
rect 52138 2651 52154 2667
rect 52256 2667 52322 2701
rect 52256 2651 52272 2667
rect 52138 2633 52272 2651
rect 52306 2633 52322 2667
rect 51080 2613 52322 2633
rect 52356 2735 52398 2777
rect 52846 2775 52875 2809
rect 52909 2775 52967 2809
rect 53001 2775 53059 2809
rect 53093 2775 53151 2809
rect 53185 2775 53243 2809
rect 53277 2775 53335 2809
rect 53369 2775 53427 2809
rect 53461 2775 53519 2809
rect 53553 2775 53611 2809
rect 53645 2775 53703 2809
rect 53737 2775 53795 2809
rect 53829 2775 53887 2809
rect 53921 2775 53979 2809
rect 54013 2775 54071 2809
rect 54105 2775 54163 2809
rect 54197 2775 54255 2809
rect 54289 2775 54318 2809
rect 52390 2701 52398 2735
rect 52356 2667 52398 2701
rect 52390 2633 52398 2667
rect 52356 2617 52398 2633
rect 52882 2733 52928 2775
rect 52882 2699 52894 2733
rect 52882 2665 52928 2699
rect 52882 2631 52894 2665
rect 52882 2615 52928 2631
rect 52962 2733 53028 2741
rect 52962 2699 52978 2733
rect 53012 2699 53028 2733
rect 52962 2665 53028 2699
rect 53062 2733 53096 2775
rect 53062 2683 53096 2699
rect 53130 2733 53196 2741
rect 53130 2699 53146 2733
rect 53180 2699 53196 2733
rect 52962 2631 52978 2665
rect 53012 2649 53028 2665
rect 53130 2665 53196 2699
rect 53230 2733 53264 2775
rect 53230 2683 53264 2699
rect 53298 2733 53364 2741
rect 53298 2699 53314 2733
rect 53348 2699 53364 2733
rect 53130 2649 53146 2665
rect 53012 2631 53146 2649
rect 53180 2649 53196 2665
rect 53298 2665 53364 2699
rect 53398 2733 53432 2775
rect 53398 2683 53432 2699
rect 53466 2733 53532 2741
rect 53466 2699 53482 2733
rect 53516 2699 53532 2733
rect 53298 2649 53314 2665
rect 53180 2631 53314 2649
rect 53348 2649 53364 2665
rect 53466 2665 53532 2699
rect 53566 2733 53600 2775
rect 53566 2683 53600 2699
rect 53634 2733 53700 2741
rect 53634 2699 53650 2733
rect 53684 2699 53700 2733
rect 53466 2649 53482 2665
rect 53348 2631 53482 2649
rect 53516 2649 53532 2665
rect 53634 2665 53700 2699
rect 53734 2733 53768 2775
rect 53734 2683 53768 2699
rect 53802 2733 53868 2741
rect 53802 2699 53818 2733
rect 53852 2699 53868 2733
rect 53634 2649 53650 2665
rect 53516 2631 53650 2649
rect 53684 2649 53700 2665
rect 53802 2665 53868 2699
rect 53902 2733 53936 2775
rect 53902 2683 53936 2699
rect 53970 2733 54036 2741
rect 53970 2699 53986 2733
rect 54020 2699 54036 2733
rect 53802 2649 53818 2665
rect 53684 2631 53818 2649
rect 53852 2649 53868 2665
rect 53970 2665 54036 2699
rect 54070 2733 54104 2775
rect 54070 2683 54104 2699
rect 54138 2733 54204 2741
rect 54138 2699 54154 2733
rect 54188 2699 54204 2733
rect 53970 2649 53986 2665
rect 53852 2631 53986 2649
rect 54020 2649 54036 2665
rect 54138 2665 54204 2699
rect 54138 2649 54154 2665
rect 54020 2631 54154 2649
rect 54188 2631 54204 2665
rect 37765 2574 37790 2577
rect 37824 2574 37964 2577
rect 37765 2540 37776 2574
rect 37824 2543 37895 2574
rect 37810 2540 37895 2543
rect 37929 2543 37964 2574
rect 37998 2574 38132 2577
rect 38166 2574 38301 2577
rect 37998 2543 38014 2574
rect 37929 2540 38014 2543
rect 38048 2543 38132 2574
rect 38048 2540 38133 2543
rect 38167 2540 38252 2574
rect 38286 2543 38301 2574
rect 38335 2574 38468 2577
rect 38502 2574 38636 2577
rect 38335 2543 38371 2574
rect 38286 2540 38371 2543
rect 38405 2543 38468 2574
rect 38524 2543 38636 2574
rect 38670 2543 38803 2577
rect 38837 2543 38853 2577
rect 38405 2540 38490 2543
rect 38524 2540 38853 2543
rect 37765 2529 38853 2540
rect 35906 2447 35914 2481
rect 23936 2375 23952 2409
rect 23986 2375 24002 2409
rect 23936 2341 24002 2375
rect 23936 2307 23952 2341
rect 23986 2307 24002 2341
rect 23936 2299 24002 2307
rect 24036 2409 24078 2425
rect 24070 2375 24078 2409
rect 24036 2341 24078 2375
rect 24070 2307 24078 2341
rect 24036 2265 24078 2307
rect 35906 2411 35948 2447
rect 35906 2377 35914 2411
rect 35906 2343 35948 2377
rect 35906 2309 35914 2343
rect 35906 2267 35948 2309
rect 35982 2481 37224 2495
rect 35982 2447 35998 2481
rect 36032 2479 36166 2481
rect 36033 2477 36166 2479
rect 36033 2461 36165 2477
rect 35982 2445 35999 2447
rect 36033 2445 36048 2461
rect 35982 2411 36048 2445
rect 36150 2443 36165 2461
rect 36200 2475 36334 2481
rect 36368 2477 36502 2481
rect 36200 2461 36329 2475
rect 36200 2447 36216 2461
rect 36199 2443 36216 2447
rect 35982 2377 35998 2411
rect 36032 2377 36048 2411
rect 35982 2343 36048 2377
rect 35982 2309 35998 2343
rect 36032 2309 36048 2343
rect 35982 2301 36048 2309
rect 36082 2411 36116 2427
rect 36082 2343 36116 2377
rect 36082 2267 36116 2309
rect 36150 2411 36216 2443
rect 36318 2441 36329 2461
rect 36368 2461 36500 2477
rect 36368 2447 36384 2461
rect 36363 2441 36384 2447
rect 36150 2377 36166 2411
rect 36200 2377 36216 2411
rect 36150 2343 36216 2377
rect 36150 2309 36166 2343
rect 36200 2309 36216 2343
rect 36150 2301 36216 2309
rect 36250 2411 36284 2427
rect 36250 2343 36284 2377
rect 36250 2267 36284 2309
rect 36318 2411 36384 2441
rect 36486 2443 36500 2461
rect 36536 2473 36670 2481
rect 36536 2461 36669 2473
rect 36536 2447 36552 2461
rect 36534 2443 36552 2447
rect 36318 2377 36334 2411
rect 36368 2377 36384 2411
rect 36318 2343 36384 2377
rect 36318 2309 36334 2343
rect 36368 2309 36384 2343
rect 36318 2301 36384 2309
rect 36418 2411 36452 2427
rect 36418 2343 36452 2377
rect 36418 2267 36452 2309
rect 36486 2411 36552 2443
rect 36654 2439 36669 2461
rect 36704 2461 36838 2481
rect 36872 2478 37006 2481
rect 36704 2447 36720 2461
rect 36703 2439 36720 2447
rect 36486 2377 36502 2411
rect 36536 2377 36552 2411
rect 36486 2343 36552 2377
rect 36486 2309 36502 2343
rect 36536 2309 36552 2343
rect 36486 2301 36552 2309
rect 36586 2411 36620 2427
rect 36586 2343 36620 2377
rect 36586 2267 36620 2309
rect 36654 2411 36720 2439
rect 36822 2438 36838 2461
rect 36872 2461 37004 2478
rect 36872 2438 36888 2461
rect 36654 2377 36670 2411
rect 36704 2377 36720 2411
rect 36654 2343 36720 2377
rect 36654 2309 36670 2343
rect 36704 2309 36720 2343
rect 36654 2301 36720 2309
rect 36754 2411 36788 2427
rect 36754 2343 36788 2377
rect 36754 2267 36788 2309
rect 36822 2411 36888 2438
rect 36990 2444 37004 2461
rect 37040 2461 37174 2481
rect 37040 2447 37056 2461
rect 37038 2444 37056 2447
rect 36822 2377 36838 2411
rect 36872 2377 36888 2411
rect 36822 2343 36888 2377
rect 36822 2309 36838 2343
rect 36872 2309 36888 2343
rect 36822 2301 36888 2309
rect 36922 2411 36956 2427
rect 36922 2343 36956 2377
rect 36922 2267 36956 2309
rect 36990 2411 37056 2444
rect 37158 2446 37174 2461
rect 37208 2446 37224 2481
rect 36990 2377 37006 2411
rect 37040 2377 37056 2411
rect 36990 2343 37056 2377
rect 36990 2309 37006 2343
rect 37040 2309 37056 2343
rect 36990 2301 37056 2309
rect 37090 2411 37124 2427
rect 37090 2343 37124 2377
rect 37090 2267 37124 2309
rect 37158 2411 37224 2446
rect 37788 2479 37830 2495
rect 39040 2493 39106 2611
rect 50981 2545 51006 2579
rect 51040 2545 51180 2579
rect 51214 2574 51348 2579
rect 50981 2540 51188 2545
rect 51222 2540 51285 2574
rect 51319 2545 51348 2574
rect 51382 2574 51517 2579
rect 51319 2540 51382 2545
rect 51416 2540 51479 2574
rect 51513 2545 51517 2574
rect 51551 2574 51684 2579
rect 51718 2574 51852 2579
rect 51886 2574 52019 2579
rect 51551 2545 51576 2574
rect 51513 2540 51576 2545
rect 51610 2540 51673 2574
rect 51718 2545 51770 2574
rect 51707 2540 51770 2545
rect 51804 2545 51852 2574
rect 51804 2540 51867 2545
rect 51901 2540 52018 2574
rect 52053 2545 52069 2579
rect 52052 2540 52069 2545
rect 50981 2531 52069 2540
rect 37788 2445 37796 2479
rect 37158 2377 37174 2411
rect 37208 2377 37224 2411
rect 37158 2343 37224 2377
rect 37158 2309 37174 2343
rect 37208 2309 37224 2343
rect 37158 2301 37224 2309
rect 37258 2411 37300 2427
rect 37292 2377 37300 2411
rect 37258 2343 37300 2377
rect 37292 2309 37300 2343
rect 37258 2267 37300 2309
rect 37788 2409 37830 2445
rect 37788 2375 37796 2409
rect 37788 2341 37830 2375
rect 37788 2307 37796 2341
rect 22644 2231 22673 2265
rect 22707 2231 22765 2265
rect 22799 2231 22857 2265
rect 22891 2231 22949 2265
rect 22983 2231 23041 2265
rect 23075 2231 23133 2265
rect 23167 2231 23225 2265
rect 23259 2231 23317 2265
rect 23351 2231 23409 2265
rect 23443 2231 23501 2265
rect 23535 2231 23593 2265
rect 23627 2231 23685 2265
rect 23719 2231 23777 2265
rect 23811 2231 23869 2265
rect 23903 2231 23961 2265
rect 23995 2231 24053 2265
rect 24087 2231 24116 2265
rect 35866 2233 35895 2267
rect 35929 2233 35987 2267
rect 36021 2233 36079 2267
rect 36113 2233 36171 2267
rect 36205 2233 36263 2267
rect 36297 2233 36355 2267
rect 36389 2233 36447 2267
rect 36481 2233 36539 2267
rect 36573 2233 36631 2267
rect 36665 2233 36723 2267
rect 36757 2233 36815 2267
rect 36849 2233 36907 2267
rect 36941 2233 36999 2267
rect 37033 2233 37091 2267
rect 37125 2233 37183 2267
rect 37217 2233 37275 2267
rect 37309 2233 37338 2267
rect 37788 2265 37830 2307
rect 37864 2481 39106 2493
rect 37864 2479 38384 2481
rect 38418 2479 39106 2481
rect 37864 2445 37880 2479
rect 37914 2477 38048 2479
rect 37922 2459 38048 2477
rect 37864 2443 37888 2445
rect 37922 2443 37930 2459
rect 37864 2409 37930 2443
rect 38032 2443 38048 2459
rect 38082 2471 38216 2479
rect 38082 2459 38215 2471
rect 38082 2443 38098 2459
rect 37864 2375 37880 2409
rect 37914 2375 37930 2409
rect 37864 2341 37930 2375
rect 37864 2307 37880 2341
rect 37914 2307 37930 2341
rect 37864 2299 37930 2307
rect 37964 2409 37998 2425
rect 37964 2341 37998 2375
rect 37964 2265 37998 2307
rect 38032 2409 38098 2443
rect 38200 2437 38215 2459
rect 38250 2459 38384 2479
rect 38250 2445 38266 2459
rect 38249 2437 38266 2445
rect 38032 2375 38048 2409
rect 38082 2375 38098 2409
rect 38032 2341 38098 2375
rect 38032 2307 38048 2341
rect 38082 2307 38098 2341
rect 38032 2299 38098 2307
rect 38132 2409 38166 2425
rect 38132 2341 38166 2375
rect 38132 2265 38166 2307
rect 38200 2409 38266 2437
rect 38368 2445 38384 2459
rect 38418 2468 38552 2479
rect 38586 2474 38720 2479
rect 38418 2459 38548 2468
rect 38418 2445 38434 2459
rect 38200 2375 38216 2409
rect 38250 2375 38266 2409
rect 38200 2341 38266 2375
rect 38200 2307 38216 2341
rect 38250 2307 38266 2341
rect 38200 2299 38266 2307
rect 38300 2409 38334 2425
rect 38300 2341 38334 2375
rect 38300 2265 38334 2307
rect 38368 2409 38434 2445
rect 38536 2434 38548 2459
rect 38586 2459 38718 2474
rect 38586 2445 38602 2459
rect 38582 2434 38602 2445
rect 38368 2375 38384 2409
rect 38418 2375 38434 2409
rect 38368 2341 38434 2375
rect 38368 2307 38384 2341
rect 38418 2307 38434 2341
rect 38368 2299 38434 2307
rect 38468 2409 38502 2425
rect 38468 2341 38502 2375
rect 38468 2265 38502 2307
rect 38536 2409 38602 2434
rect 38704 2440 38718 2459
rect 38754 2459 38888 2479
rect 38922 2478 39056 2479
rect 38754 2445 38770 2459
rect 38752 2440 38770 2445
rect 38536 2375 38552 2409
rect 38586 2375 38602 2409
rect 38536 2341 38602 2375
rect 38536 2307 38552 2341
rect 38586 2307 38602 2341
rect 38536 2299 38602 2307
rect 38636 2409 38670 2425
rect 38636 2341 38670 2375
rect 38636 2265 38670 2307
rect 38704 2409 38770 2440
rect 38872 2442 38888 2459
rect 38922 2459 39047 2478
rect 38922 2442 38938 2459
rect 38704 2375 38720 2409
rect 38754 2375 38770 2409
rect 38704 2341 38770 2375
rect 38704 2307 38720 2341
rect 38754 2307 38770 2341
rect 38704 2299 38770 2307
rect 38804 2409 38838 2425
rect 38804 2341 38838 2375
rect 38804 2265 38838 2307
rect 38872 2409 38938 2442
rect 39040 2444 39047 2459
rect 39090 2445 39106 2479
rect 39081 2444 39106 2445
rect 38872 2375 38888 2409
rect 38922 2375 38938 2409
rect 38872 2341 38938 2375
rect 38872 2307 38888 2341
rect 38922 2307 38938 2341
rect 38872 2299 38938 2307
rect 38972 2409 39006 2425
rect 38972 2341 39006 2375
rect 38972 2265 39006 2307
rect 39040 2409 39106 2444
rect 51004 2481 51046 2497
rect 52256 2495 52322 2613
rect 52962 2611 54204 2631
rect 54238 2733 54280 2775
rect 54272 2699 54280 2733
rect 54238 2665 54280 2699
rect 54272 2631 54280 2665
rect 54238 2615 54280 2631
rect 52863 2574 52888 2577
rect 52922 2574 53062 2577
rect 53096 2574 53230 2577
rect 53264 2574 53399 2577
rect 53433 2574 53566 2577
rect 52863 2540 52874 2574
rect 52922 2543 52982 2574
rect 52908 2540 52982 2543
rect 53016 2543 53062 2574
rect 53016 2540 53090 2543
rect 53124 2540 53198 2574
rect 53264 2543 53306 2574
rect 53232 2540 53306 2543
rect 53340 2543 53399 2574
rect 53340 2540 53414 2543
rect 53448 2540 53522 2574
rect 53556 2543 53566 2574
rect 53600 2574 53734 2577
rect 53600 2543 53630 2574
rect 53556 2540 53630 2543
rect 53664 2543 53734 2574
rect 53768 2543 53901 2577
rect 53935 2543 53951 2577
rect 53664 2540 53951 2543
rect 52863 2529 53951 2540
rect 51004 2447 51012 2481
rect 39040 2375 39056 2409
rect 39090 2375 39106 2409
rect 39040 2341 39106 2375
rect 39040 2307 39056 2341
rect 39090 2307 39106 2341
rect 39040 2299 39106 2307
rect 39140 2409 39182 2425
rect 39174 2375 39182 2409
rect 39140 2341 39182 2375
rect 39174 2307 39182 2341
rect 39140 2265 39182 2307
rect 51004 2411 51046 2447
rect 51004 2377 51012 2411
rect 51004 2343 51046 2377
rect 51004 2309 51012 2343
rect 51004 2267 51046 2309
rect 51080 2481 52322 2495
rect 51080 2447 51096 2481
rect 51130 2473 51264 2481
rect 51131 2468 51264 2473
rect 51131 2461 51260 2468
rect 51080 2439 51097 2447
rect 51131 2439 51146 2461
rect 51080 2411 51146 2439
rect 51248 2434 51260 2461
rect 51298 2461 51432 2481
rect 51466 2477 51600 2481
rect 51466 2472 51598 2477
rect 51298 2447 51314 2461
rect 51294 2434 51314 2447
rect 51080 2377 51096 2411
rect 51130 2377 51146 2411
rect 51080 2343 51146 2377
rect 51080 2309 51096 2343
rect 51130 2309 51146 2343
rect 51080 2301 51146 2309
rect 51180 2411 51214 2427
rect 51180 2343 51214 2377
rect 51180 2267 51214 2309
rect 51248 2411 51314 2434
rect 51416 2447 51432 2461
rect 51467 2461 51598 2472
rect 51416 2438 51433 2447
rect 51467 2438 51482 2461
rect 51248 2377 51264 2411
rect 51298 2377 51314 2411
rect 51248 2343 51314 2377
rect 51248 2309 51264 2343
rect 51298 2309 51314 2343
rect 51248 2301 51314 2309
rect 51348 2411 51382 2427
rect 51348 2343 51382 2377
rect 51348 2267 51382 2309
rect 51416 2411 51482 2438
rect 51584 2443 51598 2461
rect 51634 2464 51768 2481
rect 51634 2461 51765 2464
rect 51634 2447 51650 2461
rect 51632 2443 51650 2447
rect 51416 2377 51432 2411
rect 51466 2377 51482 2411
rect 51416 2343 51482 2377
rect 51416 2309 51432 2343
rect 51466 2309 51482 2343
rect 51416 2301 51482 2309
rect 51516 2411 51550 2427
rect 51516 2343 51550 2377
rect 51516 2267 51550 2309
rect 51584 2411 51650 2443
rect 51752 2430 51765 2461
rect 51802 2462 51936 2481
rect 51970 2471 52104 2481
rect 51802 2461 51933 2462
rect 51802 2447 51818 2461
rect 51799 2430 51818 2447
rect 51584 2377 51600 2411
rect 51634 2377 51650 2411
rect 51584 2343 51650 2377
rect 51584 2309 51600 2343
rect 51634 2309 51650 2343
rect 51584 2301 51650 2309
rect 51684 2411 51718 2427
rect 51684 2343 51718 2377
rect 51684 2267 51718 2309
rect 51752 2411 51818 2430
rect 51920 2428 51933 2461
rect 51970 2461 52103 2471
rect 51970 2447 51986 2461
rect 51967 2428 51986 2447
rect 51752 2377 51768 2411
rect 51802 2377 51818 2411
rect 51752 2343 51818 2377
rect 51752 2309 51768 2343
rect 51802 2309 51818 2343
rect 51752 2301 51818 2309
rect 51852 2411 51886 2427
rect 51852 2343 51886 2377
rect 51852 2267 51886 2309
rect 51920 2411 51986 2428
rect 52088 2437 52103 2461
rect 52138 2461 52272 2481
rect 52138 2447 52154 2461
rect 52137 2437 52154 2447
rect 51920 2377 51936 2411
rect 51970 2377 51986 2411
rect 51920 2343 51986 2377
rect 51920 2309 51936 2343
rect 51970 2309 51986 2343
rect 51920 2301 51986 2309
rect 52020 2411 52054 2427
rect 52020 2343 52054 2377
rect 52020 2267 52054 2309
rect 52088 2411 52154 2437
rect 52256 2447 52272 2461
rect 52306 2447 52322 2481
rect 52088 2377 52104 2411
rect 52138 2377 52154 2411
rect 52088 2343 52154 2377
rect 52088 2309 52104 2343
rect 52138 2309 52154 2343
rect 52088 2301 52154 2309
rect 52188 2411 52222 2427
rect 52188 2343 52222 2377
rect 52188 2267 52222 2309
rect 52256 2411 52322 2447
rect 52886 2479 52928 2495
rect 54138 2493 54204 2611
rect 52886 2445 52894 2479
rect 52256 2377 52272 2411
rect 52306 2377 52322 2411
rect 52256 2343 52322 2377
rect 52256 2309 52272 2343
rect 52306 2309 52322 2343
rect 52256 2301 52322 2309
rect 52356 2411 52398 2427
rect 52390 2377 52398 2411
rect 52356 2343 52398 2377
rect 52390 2309 52398 2343
rect 52356 2267 52398 2309
rect 52886 2409 52928 2445
rect 52886 2375 52894 2409
rect 52886 2341 52928 2375
rect 52886 2307 52894 2341
rect 37748 2231 37777 2265
rect 37811 2231 37869 2265
rect 37903 2231 37961 2265
rect 37995 2231 38053 2265
rect 38087 2231 38145 2265
rect 38179 2231 38237 2265
rect 38271 2231 38329 2265
rect 38363 2231 38421 2265
rect 38455 2231 38513 2265
rect 38547 2231 38605 2265
rect 38639 2231 38697 2265
rect 38731 2231 38789 2265
rect 38823 2231 38881 2265
rect 38915 2231 38973 2265
rect 39007 2231 39065 2265
rect 39099 2231 39157 2265
rect 39191 2231 39220 2265
rect 50964 2233 50993 2267
rect 51027 2233 51085 2267
rect 51119 2233 51177 2267
rect 51211 2233 51269 2267
rect 51303 2233 51361 2267
rect 51395 2233 51453 2267
rect 51487 2233 51545 2267
rect 51579 2233 51637 2267
rect 51671 2233 51729 2267
rect 51763 2233 51821 2267
rect 51855 2233 51913 2267
rect 51947 2233 52005 2267
rect 52039 2233 52097 2267
rect 52131 2233 52189 2267
rect 52223 2233 52281 2267
rect 52315 2233 52373 2267
rect 52407 2233 52436 2267
rect 52886 2265 52928 2307
rect 52962 2481 54204 2493
rect 52962 2479 53482 2481
rect 53516 2479 54204 2481
rect 52962 2472 52978 2479
rect 52962 2438 52976 2472
rect 53012 2459 53146 2479
rect 53180 2478 53314 2479
rect 53180 2473 53311 2478
rect 53012 2445 53028 2459
rect 53010 2438 53028 2445
rect 52962 2409 53028 2438
rect 53130 2445 53146 2459
rect 53183 2459 53311 2473
rect 53130 2439 53149 2445
rect 53183 2439 53196 2459
rect 52962 2375 52978 2409
rect 53012 2375 53028 2409
rect 52962 2341 53028 2375
rect 52962 2307 52978 2341
rect 53012 2307 53028 2341
rect 52962 2299 53028 2307
rect 53062 2409 53096 2425
rect 53062 2341 53096 2375
rect 53062 2265 53096 2307
rect 53130 2409 53196 2439
rect 53298 2444 53311 2459
rect 53348 2459 53482 2479
rect 53348 2445 53364 2459
rect 53345 2444 53364 2445
rect 53130 2375 53146 2409
rect 53180 2375 53196 2409
rect 53130 2341 53196 2375
rect 53130 2307 53146 2341
rect 53180 2307 53196 2341
rect 53130 2299 53196 2307
rect 53230 2409 53264 2425
rect 53230 2341 53264 2375
rect 53230 2265 53264 2307
rect 53298 2409 53364 2444
rect 53466 2445 53482 2459
rect 53516 2459 53650 2479
rect 53684 2467 53818 2479
rect 53516 2445 53532 2459
rect 53298 2375 53314 2409
rect 53348 2375 53364 2409
rect 53298 2341 53364 2375
rect 53298 2307 53314 2341
rect 53348 2307 53364 2341
rect 53298 2299 53364 2307
rect 53398 2409 53432 2425
rect 53398 2341 53432 2375
rect 53398 2265 53432 2307
rect 53466 2409 53532 2445
rect 53634 2445 53650 2459
rect 53685 2459 53816 2467
rect 53634 2433 53651 2445
rect 53685 2433 53700 2459
rect 53466 2375 53482 2409
rect 53516 2375 53532 2409
rect 53466 2341 53532 2375
rect 53466 2307 53482 2341
rect 53516 2307 53532 2341
rect 53466 2299 53532 2307
rect 53566 2409 53600 2425
rect 53566 2341 53600 2375
rect 53566 2265 53600 2307
rect 53634 2409 53700 2433
rect 53802 2433 53816 2459
rect 53852 2459 53986 2479
rect 54020 2469 54154 2479
rect 53852 2445 53868 2459
rect 53850 2433 53868 2445
rect 53634 2375 53650 2409
rect 53684 2375 53700 2409
rect 53634 2341 53700 2375
rect 53634 2307 53650 2341
rect 53684 2307 53700 2341
rect 53634 2299 53700 2307
rect 53734 2409 53768 2425
rect 53734 2341 53768 2375
rect 53734 2265 53768 2307
rect 53802 2409 53868 2433
rect 53970 2431 53986 2459
rect 54020 2459 54149 2469
rect 54020 2431 54036 2459
rect 53802 2375 53818 2409
rect 53852 2375 53868 2409
rect 53802 2341 53868 2375
rect 53802 2307 53818 2341
rect 53852 2307 53868 2341
rect 53802 2299 53868 2307
rect 53902 2409 53936 2425
rect 53902 2341 53936 2375
rect 53902 2265 53936 2307
rect 53970 2409 54036 2431
rect 54138 2435 54149 2459
rect 54188 2445 54204 2479
rect 54183 2435 54204 2445
rect 53970 2375 53986 2409
rect 54020 2375 54036 2409
rect 53970 2341 54036 2375
rect 53970 2307 53986 2341
rect 54020 2307 54036 2341
rect 53970 2299 54036 2307
rect 54070 2409 54104 2425
rect 54070 2341 54104 2375
rect 54070 2265 54104 2307
rect 54138 2409 54204 2435
rect 54138 2375 54154 2409
rect 54188 2375 54204 2409
rect 54138 2341 54204 2375
rect 54138 2307 54154 2341
rect 54188 2307 54204 2341
rect 54138 2299 54204 2307
rect 54238 2409 54280 2425
rect 54272 2375 54280 2409
rect 54238 2341 54280 2375
rect 54272 2307 54280 2341
rect 54238 2265 54280 2307
rect 52846 2231 52875 2265
rect 52909 2231 52967 2265
rect 53001 2231 53059 2265
rect 53093 2231 53151 2265
rect 53185 2231 53243 2265
rect 53277 2231 53335 2265
rect 53369 2231 53427 2265
rect 53461 2231 53519 2265
rect 53553 2231 53611 2265
rect 53645 2231 53703 2265
rect 53737 2231 53795 2265
rect 53829 2231 53887 2265
rect 53921 2231 53979 2265
rect 54013 2231 54071 2265
rect 54105 2231 54163 2265
rect 54197 2231 54255 2265
rect 54289 2231 54318 2265
rect 176 2187 238 2188
rect 642 2187 1032 2188
rect 2064 2187 2126 2188
rect 2530 2187 2920 2188
rect 3952 2187 4014 2188
rect 4418 2187 4808 2188
rect 5840 2187 5902 2188
rect 6306 2187 6696 2188
rect 7728 2187 7790 2188
rect 8194 2187 8584 2188
rect 9616 2187 9678 2188
rect 10082 2187 10472 2188
rect 11504 2187 11566 2188
rect 11970 2187 12360 2188
rect 13392 2187 13454 2188
rect 13858 2187 14248 2188
rect 15274 2187 15336 2188
rect 15740 2187 16130 2188
rect 17162 2187 17224 2188
rect 17628 2187 18018 2188
rect 19050 2187 19112 2188
rect 19516 2187 19906 2188
rect 20938 2187 21000 2188
rect 21404 2187 21794 2188
rect 22826 2187 22888 2188
rect 23292 2187 23682 2188
rect 24714 2187 24776 2188
rect 25180 2187 25570 2188
rect 26602 2187 26664 2188
rect 27068 2187 27458 2188
rect 28490 2187 28552 2188
rect 28956 2187 29346 2188
rect 30378 2187 30440 2188
rect 30844 2187 31234 2188
rect 32266 2187 32328 2188
rect 32732 2187 33122 2188
rect 34154 2187 34216 2188
rect 34620 2187 35010 2188
rect 36042 2187 36104 2188
rect 36508 2187 36898 2188
rect 37930 2187 37992 2188
rect 38396 2187 38786 2188
rect 39818 2187 39880 2188
rect 40284 2187 40674 2188
rect 41706 2187 41768 2188
rect 42172 2187 42562 2188
rect 43594 2187 43656 2188
rect 44060 2187 44450 2188
rect 45476 2187 45538 2188
rect 45942 2187 46332 2188
rect 47364 2187 47426 2188
rect 47830 2187 48220 2188
rect 49252 2187 49314 2188
rect 49718 2187 50108 2188
rect 51140 2187 51202 2188
rect 51606 2187 51996 2188
rect 53028 2187 53090 2188
rect 53494 2187 53884 2188
rect 54916 2187 54978 2188
rect 55382 2187 55772 2188
rect 56804 2187 56866 2188
rect 57270 2187 57660 2188
rect 58692 2187 58754 2188
rect 59158 2187 59548 2188
rect 176 2154 247 2187
rect 218 2153 247 2154
rect 281 2153 339 2187
rect 373 2153 431 2187
rect 465 2153 1061 2187
rect 1095 2153 1153 2187
rect 1187 2153 1245 2187
rect 1279 2153 1308 2187
rect 2064 2154 2135 2187
rect 2106 2153 2135 2154
rect 2169 2153 2227 2187
rect 2261 2153 2319 2187
rect 2353 2153 2949 2187
rect 2983 2153 3041 2187
rect 3075 2153 3133 2187
rect 3167 2153 3196 2187
rect 3952 2154 4023 2187
rect 3994 2153 4023 2154
rect 4057 2153 4115 2187
rect 4149 2153 4207 2187
rect 4241 2153 4837 2187
rect 4871 2153 4929 2187
rect 4963 2153 5021 2187
rect 5055 2153 5084 2187
rect 5840 2154 5911 2187
rect 5882 2153 5911 2154
rect 5945 2153 6003 2187
rect 6037 2153 6095 2187
rect 6129 2153 6725 2187
rect 6759 2153 6817 2187
rect 6851 2153 6909 2187
rect 6943 2153 6972 2187
rect 7728 2154 7799 2187
rect 7770 2153 7799 2154
rect 7833 2153 7891 2187
rect 7925 2153 7983 2187
rect 8017 2153 8613 2187
rect 8647 2153 8705 2187
rect 8739 2153 8797 2187
rect 8831 2153 8860 2187
rect 9616 2154 9687 2187
rect 9658 2153 9687 2154
rect 9721 2153 9779 2187
rect 9813 2153 9871 2187
rect 9905 2153 10501 2187
rect 10535 2153 10593 2187
rect 10627 2153 10685 2187
rect 10719 2153 10748 2187
rect 11504 2154 11575 2187
rect 11546 2153 11575 2154
rect 11609 2153 11667 2187
rect 11701 2153 11759 2187
rect 11793 2153 12389 2187
rect 12423 2153 12481 2187
rect 12515 2153 12573 2187
rect 12607 2153 12636 2187
rect 13392 2154 13463 2187
rect 13434 2153 13463 2154
rect 13497 2153 13555 2187
rect 13589 2153 13647 2187
rect 13681 2153 14277 2187
rect 14311 2153 14369 2187
rect 14403 2153 14461 2187
rect 14495 2153 14524 2187
rect 15274 2154 15345 2187
rect 15316 2153 15345 2154
rect 15379 2153 15437 2187
rect 15471 2153 15529 2187
rect 15563 2153 16159 2187
rect 16193 2153 16251 2187
rect 16285 2153 16343 2187
rect 16377 2153 16406 2187
rect 17162 2154 17233 2187
rect 17204 2153 17233 2154
rect 17267 2153 17325 2187
rect 17359 2153 17417 2187
rect 17451 2153 18047 2187
rect 18081 2153 18139 2187
rect 18173 2153 18231 2187
rect 18265 2153 18294 2187
rect 19050 2154 19121 2187
rect 19092 2153 19121 2154
rect 19155 2153 19213 2187
rect 19247 2153 19305 2187
rect 19339 2153 19935 2187
rect 19969 2153 20027 2187
rect 20061 2153 20119 2187
rect 20153 2153 20182 2187
rect 20938 2154 21009 2187
rect 20980 2153 21009 2154
rect 21043 2153 21101 2187
rect 21135 2153 21193 2187
rect 21227 2153 21823 2187
rect 21857 2153 21915 2187
rect 21949 2153 22007 2187
rect 22041 2153 22070 2187
rect 22826 2154 22897 2187
rect 22868 2153 22897 2154
rect 22931 2153 22989 2187
rect 23023 2153 23081 2187
rect 23115 2153 23711 2187
rect 23745 2153 23803 2187
rect 23837 2153 23895 2187
rect 23929 2153 23958 2187
rect 24714 2154 24785 2187
rect 24756 2153 24785 2154
rect 24819 2153 24877 2187
rect 24911 2153 24969 2187
rect 25003 2153 25599 2187
rect 25633 2153 25691 2187
rect 25725 2153 25783 2187
rect 25817 2153 25846 2187
rect 26602 2154 26673 2187
rect 26644 2153 26673 2154
rect 26707 2153 26765 2187
rect 26799 2153 26857 2187
rect 26891 2153 27487 2187
rect 27521 2153 27579 2187
rect 27613 2153 27671 2187
rect 27705 2153 27734 2187
rect 28490 2154 28561 2187
rect 28532 2153 28561 2154
rect 28595 2153 28653 2187
rect 28687 2153 28745 2187
rect 28779 2153 29375 2187
rect 29409 2153 29467 2187
rect 29501 2153 29559 2187
rect 29593 2153 29622 2187
rect 30378 2154 30449 2187
rect 30420 2153 30449 2154
rect 30483 2153 30541 2187
rect 30575 2153 30633 2187
rect 30667 2153 31263 2187
rect 31297 2153 31355 2187
rect 31389 2153 31447 2187
rect 31481 2153 31510 2187
rect 32266 2154 32337 2187
rect 32308 2153 32337 2154
rect 32371 2153 32429 2187
rect 32463 2153 32521 2187
rect 32555 2153 33151 2187
rect 33185 2153 33243 2187
rect 33277 2153 33335 2187
rect 33369 2153 33398 2187
rect 34154 2154 34225 2187
rect 34196 2153 34225 2154
rect 34259 2153 34317 2187
rect 34351 2153 34409 2187
rect 34443 2153 35039 2187
rect 35073 2153 35131 2187
rect 35165 2153 35223 2187
rect 35257 2153 35286 2187
rect 36042 2154 36113 2187
rect 36084 2153 36113 2154
rect 36147 2153 36205 2187
rect 36239 2153 36297 2187
rect 36331 2153 36927 2187
rect 36961 2153 37019 2187
rect 37053 2153 37111 2187
rect 37145 2153 37174 2187
rect 37930 2154 38001 2187
rect 37972 2153 38001 2154
rect 38035 2153 38093 2187
rect 38127 2153 38185 2187
rect 38219 2153 38815 2187
rect 38849 2153 38907 2187
rect 38941 2153 38999 2187
rect 39033 2153 39062 2187
rect 39818 2154 39889 2187
rect 39860 2153 39889 2154
rect 39923 2153 39981 2187
rect 40015 2153 40073 2187
rect 40107 2153 40703 2187
rect 40737 2153 40795 2187
rect 40829 2153 40887 2187
rect 40921 2153 40950 2187
rect 41706 2154 41777 2187
rect 41748 2153 41777 2154
rect 41811 2153 41869 2187
rect 41903 2153 41961 2187
rect 41995 2153 42591 2187
rect 42625 2153 42683 2187
rect 42717 2153 42775 2187
rect 42809 2153 42838 2187
rect 43594 2154 43665 2187
rect 43636 2153 43665 2154
rect 43699 2153 43757 2187
rect 43791 2153 43849 2187
rect 43883 2153 44479 2187
rect 44513 2153 44571 2187
rect 44605 2153 44663 2187
rect 44697 2153 44726 2187
rect 45476 2154 45547 2187
rect 45518 2153 45547 2154
rect 45581 2153 45639 2187
rect 45673 2153 45731 2187
rect 45765 2153 46361 2187
rect 46395 2153 46453 2187
rect 46487 2153 46545 2187
rect 46579 2153 46608 2187
rect 47364 2154 47435 2187
rect 47406 2153 47435 2154
rect 47469 2153 47527 2187
rect 47561 2153 47619 2187
rect 47653 2153 48249 2187
rect 48283 2153 48341 2187
rect 48375 2153 48433 2187
rect 48467 2153 48496 2187
rect 49252 2154 49323 2187
rect 49294 2153 49323 2154
rect 49357 2153 49415 2187
rect 49449 2153 49507 2187
rect 49541 2153 50137 2187
rect 50171 2153 50229 2187
rect 50263 2153 50321 2187
rect 50355 2153 50384 2187
rect 51140 2154 51211 2187
rect 51182 2153 51211 2154
rect 51245 2153 51303 2187
rect 51337 2153 51395 2187
rect 51429 2153 52025 2187
rect 52059 2153 52117 2187
rect 52151 2153 52209 2187
rect 52243 2153 52272 2187
rect 53028 2154 53099 2187
rect 53070 2153 53099 2154
rect 53133 2153 53191 2187
rect 53225 2153 53283 2187
rect 53317 2153 53913 2187
rect 53947 2153 54005 2187
rect 54039 2153 54097 2187
rect 54131 2153 54160 2187
rect 54916 2154 54987 2187
rect 54958 2153 54987 2154
rect 55021 2153 55079 2187
rect 55113 2153 55171 2187
rect 55205 2153 55801 2187
rect 55835 2153 55893 2187
rect 55927 2153 55985 2187
rect 56019 2153 56048 2187
rect 56804 2154 56875 2187
rect 56846 2153 56875 2154
rect 56909 2153 56967 2187
rect 57001 2153 57059 2187
rect 57093 2153 57689 2187
rect 57723 2153 57781 2187
rect 57815 2153 57873 2187
rect 57907 2153 57936 2187
rect 58692 2154 58763 2187
rect 58734 2153 58763 2154
rect 58797 2153 58855 2187
rect 58889 2153 58947 2187
rect 58981 2153 59577 2187
rect 59611 2153 59669 2187
rect 59703 2153 59761 2187
rect 59795 2153 59824 2187
rect 237 2111 303 2116
rect 237 2077 253 2111
rect 287 2077 303 2111
rect 237 2043 303 2077
rect 237 2009 253 2043
rect 287 2009 303 2043
rect 237 1975 303 2009
rect 237 1941 253 1975
rect 287 1959 303 1975
rect 409 2111 475 2153
rect 443 2077 475 2111
rect 642 2147 924 2153
rect 642 2113 681 2147
rect 715 2145 924 2147
rect 715 2113 800 2145
rect 642 2111 800 2113
rect 834 2111 924 2145
rect 642 2078 924 2111
rect 1051 2111 1117 2116
rect 409 2043 475 2077
rect 443 2009 475 2043
rect 1051 2077 1067 2111
rect 1101 2077 1117 2111
rect 1051 2043 1117 2077
rect 409 1975 475 2009
rect 287 1941 373 1959
rect 237 1925 373 1941
rect 443 1941 475 1975
rect 409 1925 475 1941
rect 534 2039 800 2040
rect 534 2005 750 2039
rect 784 2005 800 2039
rect 534 2004 800 2005
rect 235 1884 305 1891
rect 235 1850 253 1884
rect 287 1875 305 1884
rect 235 1841 255 1850
rect 289 1841 305 1875
rect 339 1805 373 1925
rect 407 1880 477 1891
rect 407 1875 426 1880
rect 407 1841 423 1875
rect 460 1846 477 1880
rect 457 1841 477 1846
rect 239 1789 287 1805
rect 239 1755 253 1789
rect 239 1721 287 1755
rect 239 1687 253 1721
rect 239 1643 287 1687
rect 321 1789 387 1805
rect 321 1764 337 1789
rect 321 1730 335 1764
rect 371 1755 387 1789
rect 369 1730 387 1755
rect 321 1721 387 1730
rect 321 1687 337 1721
rect 371 1687 387 1721
rect 321 1677 387 1687
rect 421 1789 475 1805
rect 455 1755 475 1789
rect 421 1721 475 1755
rect 455 1687 475 1721
rect 421 1643 475 1687
rect 218 1609 247 1643
rect 281 1609 339 1643
rect 373 1609 431 1643
rect 465 1609 494 1643
rect 218 1398 252 1609
rect 449 1306 483 1609
rect 534 1390 568 2004
rect 734 2002 800 2004
rect 1051 2009 1067 2043
rect 1101 2009 1117 2043
rect 1051 1975 1117 2009
rect 606 1943 640 1962
rect 606 1875 640 1877
rect 606 1839 640 1841
rect 606 1754 640 1773
rect 702 1943 736 1962
rect 702 1875 736 1877
rect 702 1839 736 1841
rect 702 1754 736 1773
rect 798 1943 832 1962
rect 1051 1941 1067 1975
rect 1101 1959 1117 1975
rect 1223 2111 1289 2153
rect 1257 2077 1289 2111
rect 1223 2043 1289 2077
rect 1257 2009 1289 2043
rect 1223 1975 1289 2009
rect 1101 1941 1187 1959
rect 1051 1925 1187 1941
rect 1257 1941 1289 1975
rect 1223 1925 1289 1941
rect 2125 2111 2191 2116
rect 2125 2077 2141 2111
rect 2175 2077 2191 2111
rect 2125 2043 2191 2077
rect 2125 2009 2141 2043
rect 2175 2009 2191 2043
rect 2125 1975 2191 2009
rect 2125 1941 2141 1975
rect 2175 1959 2191 1975
rect 2297 2111 2363 2153
rect 2331 2077 2363 2111
rect 2530 2147 2812 2153
rect 2530 2113 2569 2147
rect 2603 2145 2812 2147
rect 2603 2113 2688 2145
rect 2530 2111 2688 2113
rect 2722 2111 2812 2145
rect 2530 2078 2812 2111
rect 2939 2111 3005 2116
rect 2297 2043 2363 2077
rect 2331 2009 2363 2043
rect 2939 2077 2955 2111
rect 2989 2077 3005 2111
rect 2939 2043 3005 2077
rect 2297 1975 2363 2009
rect 2175 1941 2261 1959
rect 2125 1925 2261 1941
rect 2331 1941 2363 1975
rect 2297 1925 2363 1941
rect 2422 2039 2688 2040
rect 2422 2005 2638 2039
rect 2672 2005 2688 2039
rect 2422 2004 2688 2005
rect 798 1875 832 1877
rect 1049 1882 1119 1891
rect 1049 1848 1065 1882
rect 1099 1875 1119 1882
rect 1049 1841 1069 1848
rect 1103 1841 1119 1875
rect 798 1839 832 1841
rect 1153 1805 1187 1925
rect 1221 1882 1291 1891
rect 1221 1875 1239 1882
rect 1221 1841 1237 1875
rect 1273 1848 1291 1882
rect 1271 1841 1291 1848
rect 2123 1884 2193 1891
rect 2123 1850 2141 1884
rect 2175 1875 2193 1884
rect 2123 1841 2143 1850
rect 2177 1841 2193 1875
rect 2227 1805 2261 1925
rect 2295 1880 2365 1891
rect 2295 1875 2314 1880
rect 2295 1841 2311 1875
rect 2348 1846 2365 1880
rect 2345 1841 2365 1846
rect 798 1754 832 1773
rect 1053 1789 1101 1805
rect 1053 1755 1067 1789
rect 1053 1721 1101 1755
rect 638 1677 654 1711
rect 688 1677 704 1711
rect 1053 1687 1067 1721
rect 1053 1643 1101 1687
rect 1135 1789 1201 1805
rect 1135 1755 1151 1789
rect 1185 1759 1201 1789
rect 1135 1725 1153 1755
rect 1187 1725 1201 1759
rect 1135 1721 1201 1725
rect 1135 1687 1151 1721
rect 1185 1687 1201 1721
rect 1135 1677 1201 1687
rect 1235 1789 1289 1805
rect 1269 1755 1289 1789
rect 1235 1721 1289 1755
rect 1269 1687 1289 1721
rect 1235 1643 1289 1687
rect 2127 1789 2175 1805
rect 2127 1755 2141 1789
rect 2127 1721 2175 1755
rect 2127 1687 2141 1721
rect 2127 1643 2175 1687
rect 2209 1789 2275 1805
rect 2209 1764 2225 1789
rect 2209 1730 2223 1764
rect 2259 1755 2275 1789
rect 2257 1730 2275 1755
rect 2209 1721 2275 1730
rect 2209 1687 2225 1721
rect 2259 1687 2275 1721
rect 2209 1677 2275 1687
rect 2309 1789 2363 1805
rect 2343 1755 2363 1789
rect 2309 1721 2363 1755
rect 2343 1687 2363 1721
rect 2309 1643 2363 1687
rect 750 1596 766 1630
rect 800 1596 816 1630
rect 1032 1609 1061 1643
rect 1095 1609 1153 1643
rect 1187 1609 1245 1643
rect 1279 1609 1308 1643
rect 2106 1609 2135 1643
rect 2169 1609 2227 1643
rect 2261 1609 2319 1643
rect 2353 1609 2382 1643
rect 622 1546 656 1562
rect 622 1476 656 1510
rect 622 1424 656 1440
rect 718 1546 752 1562
rect 718 1476 752 1510
rect 718 1424 752 1440
rect 814 1546 848 1562
rect 814 1476 848 1510
rect 848 1440 1196 1464
rect 814 1424 1196 1440
rect 534 1356 670 1390
rect 704 1356 720 1390
rect 449 1286 844 1306
rect 449 1281 711 1286
rect 449 1272 590 1281
rect 574 1247 590 1272
rect 624 1252 711 1281
rect 745 1262 844 1286
rect 1016 1264 1062 1266
rect 1016 1262 1020 1264
rect 745 1252 1020 1262
rect 624 1247 1020 1252
rect 574 1230 1020 1247
rect 1054 1230 1062 1264
rect 574 1228 1062 1230
rect 1016 1222 1062 1228
rect 115 1133 149 1140
rect 40 1099 69 1133
rect 103 1099 161 1133
rect 195 1099 253 1133
rect 287 1099 316 1133
rect 416 1109 432 1143
rect 466 1109 482 1143
rect 640 1130 754 1132
rect 108 1057 150 1099
rect 640 1091 922 1130
rect 1062 1109 1078 1143
rect 1112 1109 1128 1143
rect 640 1066 679 1091
rect 108 1023 116 1057
rect 108 989 150 1023
rect 108 955 116 989
rect 108 921 150 955
rect 108 887 116 921
rect 108 871 150 887
rect 184 1057 250 1065
rect 184 1023 200 1057
rect 234 1023 250 1057
rect 184 989 250 1023
rect 184 955 200 989
rect 234 955 250 989
rect 184 921 250 955
rect 184 887 200 921
rect 234 887 250 921
rect 184 869 250 887
rect 104 832 170 835
rect 104 798 118 832
rect 152 821 170 832
rect 104 787 120 798
rect 154 787 170 821
rect 104 737 150 753
rect 204 749 250 869
rect 388 1047 422 1066
rect 474 1057 679 1066
rect 713 1089 922 1091
rect 713 1057 798 1089
rect 474 1055 798 1057
rect 832 1066 922 1089
rect 1162 1066 1196 1424
rect 2106 1398 2140 1609
rect 2337 1306 2371 1609
rect 2422 1390 2456 2004
rect 2622 2002 2688 2004
rect 2939 2009 2955 2043
rect 2989 2009 3005 2043
rect 2939 1975 3005 2009
rect 2494 1943 2528 1962
rect 2494 1875 2528 1877
rect 2494 1839 2528 1841
rect 2494 1754 2528 1773
rect 2590 1943 2624 1962
rect 2590 1875 2624 1877
rect 2590 1839 2624 1841
rect 2590 1754 2624 1773
rect 2686 1943 2720 1962
rect 2939 1941 2955 1975
rect 2989 1959 3005 1975
rect 3111 2111 3177 2153
rect 3145 2077 3177 2111
rect 3111 2043 3177 2077
rect 3145 2009 3177 2043
rect 3111 1975 3177 2009
rect 2989 1941 3075 1959
rect 2939 1925 3075 1941
rect 3145 1941 3177 1975
rect 3111 1925 3177 1941
rect 4013 2111 4079 2116
rect 4013 2077 4029 2111
rect 4063 2077 4079 2111
rect 4013 2043 4079 2077
rect 4013 2009 4029 2043
rect 4063 2009 4079 2043
rect 4013 1975 4079 2009
rect 4013 1941 4029 1975
rect 4063 1959 4079 1975
rect 4185 2111 4251 2153
rect 4219 2077 4251 2111
rect 4418 2147 4700 2153
rect 4418 2113 4457 2147
rect 4491 2145 4700 2147
rect 4491 2113 4576 2145
rect 4418 2111 4576 2113
rect 4610 2111 4700 2145
rect 4418 2078 4700 2111
rect 4827 2111 4893 2116
rect 4185 2043 4251 2077
rect 4219 2009 4251 2043
rect 4827 2077 4843 2111
rect 4877 2077 4893 2111
rect 4827 2043 4893 2077
rect 4185 1975 4251 2009
rect 4063 1941 4149 1959
rect 4013 1925 4149 1941
rect 4219 1941 4251 1975
rect 4185 1925 4251 1941
rect 4310 2039 4576 2040
rect 4310 2005 4526 2039
rect 4560 2005 4576 2039
rect 4310 2004 4576 2005
rect 2686 1875 2720 1877
rect 2937 1882 3007 1891
rect 2937 1848 2953 1882
rect 2987 1875 3007 1882
rect 2937 1841 2957 1848
rect 2991 1841 3007 1875
rect 2686 1839 2720 1841
rect 3041 1805 3075 1925
rect 3109 1882 3179 1891
rect 3109 1875 3127 1882
rect 3109 1841 3125 1875
rect 3161 1848 3179 1882
rect 3159 1841 3179 1848
rect 4011 1884 4081 1891
rect 4011 1850 4029 1884
rect 4063 1875 4081 1884
rect 4011 1841 4031 1850
rect 4065 1841 4081 1875
rect 4115 1805 4149 1925
rect 4183 1880 4253 1891
rect 4183 1875 4202 1880
rect 4183 1841 4199 1875
rect 4236 1846 4253 1880
rect 4233 1841 4253 1846
rect 2686 1754 2720 1773
rect 2941 1789 2989 1805
rect 2941 1755 2955 1789
rect 2941 1721 2989 1755
rect 2526 1677 2542 1711
rect 2576 1677 2592 1711
rect 2941 1687 2955 1721
rect 2941 1643 2989 1687
rect 3023 1789 3089 1805
rect 3023 1755 3039 1789
rect 3073 1759 3089 1789
rect 3023 1725 3041 1755
rect 3075 1725 3089 1759
rect 3023 1721 3089 1725
rect 3023 1687 3039 1721
rect 3073 1687 3089 1721
rect 3023 1677 3089 1687
rect 3123 1789 3177 1805
rect 3157 1755 3177 1789
rect 3123 1721 3177 1755
rect 3157 1687 3177 1721
rect 3123 1643 3177 1687
rect 4015 1789 4063 1805
rect 4015 1755 4029 1789
rect 4015 1721 4063 1755
rect 4015 1687 4029 1721
rect 4015 1643 4063 1687
rect 4097 1789 4163 1805
rect 4097 1764 4113 1789
rect 4097 1730 4111 1764
rect 4147 1755 4163 1789
rect 4145 1730 4163 1755
rect 4097 1721 4163 1730
rect 4097 1687 4113 1721
rect 4147 1687 4163 1721
rect 4097 1677 4163 1687
rect 4197 1789 4251 1805
rect 4231 1755 4251 1789
rect 4197 1721 4251 1755
rect 4231 1687 4251 1721
rect 4197 1643 4251 1687
rect 2638 1596 2654 1630
rect 2688 1596 2704 1630
rect 2920 1609 2949 1643
rect 2983 1609 3041 1643
rect 3075 1609 3133 1643
rect 3167 1609 3196 1643
rect 3994 1609 4023 1643
rect 4057 1609 4115 1643
rect 4149 1609 4207 1643
rect 4241 1609 4270 1643
rect 2510 1546 2544 1562
rect 2510 1476 2544 1510
rect 2510 1424 2544 1440
rect 2606 1546 2640 1562
rect 2606 1476 2640 1510
rect 2606 1424 2640 1440
rect 2702 1546 2736 1562
rect 2702 1476 2736 1510
rect 2736 1440 3084 1464
rect 2702 1424 3084 1440
rect 2422 1356 2558 1390
rect 2592 1356 2608 1390
rect 2337 1286 2732 1306
rect 2337 1281 2599 1286
rect 2337 1272 2478 1281
rect 2462 1247 2478 1272
rect 2512 1252 2599 1281
rect 2633 1262 2732 1286
rect 2904 1264 2950 1266
rect 2904 1262 2908 1264
rect 2633 1252 2908 1262
rect 2512 1247 2908 1252
rect 2462 1230 2908 1247
rect 2942 1230 2950 1264
rect 2462 1228 2950 1230
rect 2904 1222 2950 1228
rect 1236 1107 1265 1141
rect 1299 1107 1357 1141
rect 1391 1107 1449 1141
rect 1483 1107 1512 1141
rect 832 1055 1068 1066
rect 474 1047 1068 1055
rect 474 1022 476 1047
rect 388 979 422 981
rect 388 943 422 945
rect 388 858 422 877
rect 510 1022 1034 1047
rect 1120 1047 1196 1066
rect 1120 1026 1122 1047
rect 476 979 510 981
rect 732 949 748 983
rect 782 949 798 983
rect 1034 979 1068 981
rect 476 943 510 945
rect 1034 943 1068 945
rect 476 858 510 877
rect 604 887 638 906
rect 604 819 638 821
rect 416 781 432 815
rect 466 781 482 815
rect 604 783 638 785
rect 104 703 116 737
rect 104 669 150 703
rect 104 635 116 669
rect 104 589 150 635
rect 184 737 250 749
rect 184 703 200 737
rect 234 703 250 737
rect 184 690 250 703
rect 604 698 638 717
rect 700 887 734 906
rect 700 819 734 821
rect 700 783 734 785
rect 700 698 734 717
rect 796 887 830 906
rect 1034 858 1068 877
rect 1156 1026 1196 1047
rect 1304 1065 1346 1107
rect 1582 1105 1611 1139
rect 1645 1105 1703 1139
rect 1737 1105 1795 1139
rect 1829 1105 1858 1139
rect 2003 1133 2037 1140
rect 1304 1031 1312 1065
rect 1122 979 1156 981
rect 1122 943 1156 945
rect 1304 997 1346 1031
rect 1304 963 1312 997
rect 1304 929 1346 963
rect 1304 895 1312 929
rect 1304 879 1346 895
rect 1380 1065 1446 1073
rect 1380 1031 1396 1065
rect 1430 1031 1446 1065
rect 1380 997 1446 1031
rect 1380 963 1396 997
rect 1430 963 1446 997
rect 1380 929 1446 963
rect 1380 895 1396 929
rect 1430 895 1446 929
rect 1380 877 1446 895
rect 1615 1055 1651 1071
rect 1615 1021 1617 1055
rect 1615 987 1651 1021
rect 1615 953 1617 987
rect 1687 1055 1753 1105
rect 1928 1099 1957 1133
rect 1991 1099 2049 1133
rect 2083 1099 2141 1133
rect 2175 1099 2204 1133
rect 2304 1109 2320 1143
rect 2354 1109 2370 1143
rect 2528 1130 2642 1132
rect 1687 1021 1703 1055
rect 1737 1021 1753 1055
rect 1687 987 1753 1021
rect 1687 953 1703 987
rect 1737 953 1753 987
rect 1787 1055 1841 1071
rect 1787 1021 1789 1055
rect 1823 1021 1841 1055
rect 1787 974 1841 1021
rect 1615 919 1651 953
rect 1787 940 1789 974
rect 1823 940 1841 974
rect 1615 885 1750 919
rect 1787 890 1841 940
rect 1122 858 1156 877
rect 796 819 830 821
rect 1208 843 1352 844
rect 1208 829 1366 843
rect 796 783 830 785
rect 1062 816 1128 818
rect 1208 816 1316 829
rect 1062 815 1316 816
rect 1062 781 1078 815
rect 1112 802 1316 815
rect 1112 782 1248 802
rect 1300 795 1316 802
rect 1350 795 1366 829
rect 1112 781 1128 782
rect 1300 745 1346 761
rect 1400 757 1446 877
rect 1716 856 1750 885
rect 1603 827 1671 849
rect 1603 826 1619 827
rect 1603 792 1617 826
rect 1653 793 1671 827
rect 1651 792 1671 793
rect 1603 775 1671 792
rect 1716 840 1771 856
rect 1716 806 1737 840
rect 1716 790 1771 806
rect 1805 840 1841 890
rect 1996 1057 2038 1099
rect 2528 1091 2810 1130
rect 2950 1109 2966 1143
rect 3000 1109 3016 1143
rect 2528 1066 2567 1091
rect 1996 1023 2004 1057
rect 1996 989 2038 1023
rect 1996 955 2004 989
rect 1996 921 2038 955
rect 1996 887 2004 921
rect 1996 871 2038 887
rect 2072 1057 2138 1065
rect 2072 1023 2088 1057
rect 2122 1023 2138 1057
rect 2072 989 2138 1023
rect 2072 955 2088 989
rect 2122 955 2138 989
rect 2072 921 2138 955
rect 2072 887 2088 921
rect 2122 887 2138 921
rect 2072 869 2138 887
rect 1805 838 1846 840
rect 1805 804 1810 838
rect 1844 804 1846 838
rect 1805 802 1846 804
rect 1992 832 2058 835
rect 830 717 1076 734
rect 796 700 1076 717
rect 796 698 830 700
rect 184 669 526 690
rect 184 635 200 669
rect 234 658 526 669
rect 234 655 702 658
rect 234 654 652 655
rect 234 635 256 654
rect 184 630 256 635
rect 184 623 250 630
rect 490 622 652 654
rect 636 621 652 622
rect 686 621 702 655
rect 1028 612 1076 700
rect 40 555 69 589
rect 103 555 161 589
rect 195 555 253 589
rect 287 555 316 589
rect 398 584 444 594
rect 398 550 404 584
rect 438 564 444 584
rect 1028 578 1036 612
rect 1070 578 1076 612
rect 1300 711 1312 745
rect 1300 677 1346 711
rect 1300 643 1312 677
rect 1300 597 1346 643
rect 1380 745 1446 757
rect 1380 694 1396 745
rect 1430 694 1446 745
rect 1716 739 1750 790
rect 1380 677 1446 694
rect 1380 643 1396 677
rect 1430 643 1446 677
rect 1380 631 1446 643
rect 1617 705 1750 739
rect 1805 730 1841 802
rect 1992 798 2006 832
rect 2040 821 2058 832
rect 1992 787 2008 798
rect 2042 787 2058 821
rect 1617 684 1651 705
rect 1789 701 1841 730
rect 1617 629 1651 650
rect 1687 637 1703 671
rect 1737 637 1753 671
rect 438 550 448 564
rect 398 480 448 550
rect 748 540 764 574
rect 798 540 814 574
rect 1028 566 1076 578
rect 1236 563 1265 597
rect 1299 563 1357 597
rect 1391 563 1449 597
rect 1483 563 1512 597
rect 1687 595 1753 637
rect 1823 667 1841 701
rect 1789 629 1841 667
rect 1992 737 2038 753
rect 2092 749 2138 869
rect 2276 1047 2310 1066
rect 2362 1057 2567 1066
rect 2601 1089 2810 1091
rect 2601 1057 2686 1089
rect 2362 1055 2686 1057
rect 2720 1066 2810 1089
rect 3050 1066 3084 1424
rect 3994 1398 4028 1609
rect 4225 1306 4259 1609
rect 4310 1390 4344 2004
rect 4510 2002 4576 2004
rect 4827 2009 4843 2043
rect 4877 2009 4893 2043
rect 4827 1975 4893 2009
rect 4382 1943 4416 1962
rect 4382 1875 4416 1877
rect 4382 1839 4416 1841
rect 4382 1754 4416 1773
rect 4478 1943 4512 1962
rect 4478 1875 4512 1877
rect 4478 1839 4512 1841
rect 4478 1754 4512 1773
rect 4574 1943 4608 1962
rect 4827 1941 4843 1975
rect 4877 1959 4893 1975
rect 4999 2111 5065 2153
rect 5033 2077 5065 2111
rect 4999 2043 5065 2077
rect 5033 2009 5065 2043
rect 4999 1975 5065 2009
rect 4877 1941 4963 1959
rect 4827 1925 4963 1941
rect 5033 1941 5065 1975
rect 4999 1925 5065 1941
rect 5901 2111 5967 2116
rect 5901 2077 5917 2111
rect 5951 2077 5967 2111
rect 5901 2043 5967 2077
rect 5901 2009 5917 2043
rect 5951 2009 5967 2043
rect 5901 1975 5967 2009
rect 5901 1941 5917 1975
rect 5951 1959 5967 1975
rect 6073 2111 6139 2153
rect 6107 2077 6139 2111
rect 6306 2147 6588 2153
rect 6306 2113 6345 2147
rect 6379 2145 6588 2147
rect 6379 2113 6464 2145
rect 6306 2111 6464 2113
rect 6498 2111 6588 2145
rect 6306 2078 6588 2111
rect 6715 2111 6781 2116
rect 6073 2043 6139 2077
rect 6107 2009 6139 2043
rect 6715 2077 6731 2111
rect 6765 2077 6781 2111
rect 6715 2043 6781 2077
rect 6073 1975 6139 2009
rect 5951 1941 6037 1959
rect 5901 1925 6037 1941
rect 6107 1941 6139 1975
rect 6073 1925 6139 1941
rect 6198 2039 6464 2040
rect 6198 2005 6414 2039
rect 6448 2005 6464 2039
rect 6198 2004 6464 2005
rect 4574 1875 4608 1877
rect 4825 1882 4895 1891
rect 4825 1848 4841 1882
rect 4875 1875 4895 1882
rect 4825 1841 4845 1848
rect 4879 1841 4895 1875
rect 4574 1839 4608 1841
rect 4929 1805 4963 1925
rect 4997 1882 5067 1891
rect 4997 1875 5015 1882
rect 4997 1841 5013 1875
rect 5049 1848 5067 1882
rect 5047 1841 5067 1848
rect 5899 1884 5969 1891
rect 5899 1850 5917 1884
rect 5951 1875 5969 1884
rect 5899 1841 5919 1850
rect 5953 1841 5969 1875
rect 6003 1805 6037 1925
rect 6071 1880 6141 1891
rect 6071 1875 6090 1880
rect 6071 1841 6087 1875
rect 6124 1846 6141 1880
rect 6121 1841 6141 1846
rect 4574 1754 4608 1773
rect 4829 1789 4877 1805
rect 4829 1755 4843 1789
rect 4829 1721 4877 1755
rect 4414 1677 4430 1711
rect 4464 1677 4480 1711
rect 4829 1687 4843 1721
rect 4829 1643 4877 1687
rect 4911 1789 4977 1805
rect 4911 1755 4927 1789
rect 4961 1759 4977 1789
rect 4911 1725 4929 1755
rect 4963 1725 4977 1759
rect 4911 1721 4977 1725
rect 4911 1687 4927 1721
rect 4961 1687 4977 1721
rect 4911 1677 4977 1687
rect 5011 1789 5065 1805
rect 5045 1755 5065 1789
rect 5011 1721 5065 1755
rect 5045 1687 5065 1721
rect 5011 1643 5065 1687
rect 5903 1789 5951 1805
rect 5903 1755 5917 1789
rect 5903 1721 5951 1755
rect 5903 1687 5917 1721
rect 5903 1643 5951 1687
rect 5985 1789 6051 1805
rect 5985 1764 6001 1789
rect 5985 1730 5999 1764
rect 6035 1755 6051 1789
rect 6033 1730 6051 1755
rect 5985 1721 6051 1730
rect 5985 1687 6001 1721
rect 6035 1687 6051 1721
rect 5985 1677 6051 1687
rect 6085 1789 6139 1805
rect 6119 1755 6139 1789
rect 6085 1721 6139 1755
rect 6119 1687 6139 1721
rect 6085 1643 6139 1687
rect 4526 1596 4542 1630
rect 4576 1596 4592 1630
rect 4808 1609 4837 1643
rect 4871 1609 4929 1643
rect 4963 1609 5021 1643
rect 5055 1609 5084 1643
rect 5882 1609 5911 1643
rect 5945 1609 6003 1643
rect 6037 1609 6095 1643
rect 6129 1609 6158 1643
rect 4398 1546 4432 1562
rect 4398 1476 4432 1510
rect 4398 1424 4432 1440
rect 4494 1546 4528 1562
rect 4494 1476 4528 1510
rect 4494 1424 4528 1440
rect 4590 1546 4624 1562
rect 4590 1476 4624 1510
rect 4624 1440 4972 1464
rect 4590 1424 4972 1440
rect 4310 1356 4446 1390
rect 4480 1356 4496 1390
rect 4225 1286 4620 1306
rect 4225 1281 4487 1286
rect 4225 1272 4366 1281
rect 4350 1247 4366 1272
rect 4400 1252 4487 1281
rect 4521 1262 4620 1286
rect 4792 1264 4838 1266
rect 4792 1262 4796 1264
rect 4521 1252 4796 1262
rect 4400 1247 4796 1252
rect 4350 1230 4796 1247
rect 4830 1230 4838 1264
rect 4350 1228 4838 1230
rect 4792 1222 4838 1228
rect 3124 1107 3153 1141
rect 3187 1107 3245 1141
rect 3279 1107 3337 1141
rect 3371 1107 3400 1141
rect 2720 1055 2956 1066
rect 2362 1047 2956 1055
rect 2362 1022 2364 1047
rect 2276 979 2310 981
rect 2276 943 2310 945
rect 2276 858 2310 877
rect 2398 1022 2922 1047
rect 3008 1047 3084 1066
rect 3008 1026 3010 1047
rect 2364 979 2398 981
rect 2620 949 2636 983
rect 2670 949 2686 983
rect 2922 979 2956 981
rect 2364 943 2398 945
rect 2922 943 2956 945
rect 2364 858 2398 877
rect 2492 887 2526 906
rect 2492 819 2526 821
rect 2304 781 2320 815
rect 2354 781 2370 815
rect 2492 783 2526 785
rect 1992 703 2004 737
rect 1992 669 2038 703
rect 1992 635 2004 669
rect 1582 561 1611 595
rect 1645 561 1703 595
rect 1737 561 1795 595
rect 1829 561 1858 595
rect 1992 589 2038 635
rect 2072 737 2138 749
rect 2072 703 2088 737
rect 2122 703 2138 737
rect 2072 690 2138 703
rect 2492 698 2526 717
rect 2588 887 2622 906
rect 2588 819 2622 821
rect 2588 783 2622 785
rect 2588 698 2622 717
rect 2684 887 2718 906
rect 2922 858 2956 877
rect 3044 1026 3084 1047
rect 3192 1065 3234 1107
rect 3470 1105 3499 1139
rect 3533 1105 3591 1139
rect 3625 1105 3683 1139
rect 3717 1105 3746 1139
rect 3891 1133 3925 1140
rect 3192 1031 3200 1065
rect 3010 979 3044 981
rect 3010 943 3044 945
rect 3192 997 3234 1031
rect 3192 963 3200 997
rect 3192 929 3234 963
rect 3192 895 3200 929
rect 3192 879 3234 895
rect 3268 1065 3334 1073
rect 3268 1031 3284 1065
rect 3318 1031 3334 1065
rect 3268 997 3334 1031
rect 3268 963 3284 997
rect 3318 963 3334 997
rect 3268 929 3334 963
rect 3268 895 3284 929
rect 3318 895 3334 929
rect 3268 877 3334 895
rect 3503 1055 3539 1071
rect 3503 1021 3505 1055
rect 3503 987 3539 1021
rect 3503 953 3505 987
rect 3575 1055 3641 1105
rect 3816 1099 3845 1133
rect 3879 1099 3937 1133
rect 3971 1099 4029 1133
rect 4063 1099 4092 1133
rect 4192 1109 4208 1143
rect 4242 1109 4258 1143
rect 4416 1130 4530 1132
rect 3575 1021 3591 1055
rect 3625 1021 3641 1055
rect 3575 987 3641 1021
rect 3575 953 3591 987
rect 3625 953 3641 987
rect 3675 1055 3729 1071
rect 3675 1021 3677 1055
rect 3711 1021 3729 1055
rect 3675 974 3729 1021
rect 3503 919 3539 953
rect 3675 940 3677 974
rect 3711 940 3729 974
rect 3503 885 3638 919
rect 3675 890 3729 940
rect 3010 858 3044 877
rect 2684 819 2718 821
rect 3096 843 3240 844
rect 3096 829 3254 843
rect 2684 783 2718 785
rect 2950 816 3016 818
rect 3096 816 3204 829
rect 2950 815 3204 816
rect 2950 781 2966 815
rect 3000 802 3204 815
rect 3000 782 3136 802
rect 3188 795 3204 802
rect 3238 795 3254 829
rect 3000 781 3016 782
rect 3188 745 3234 761
rect 3288 757 3334 877
rect 3604 856 3638 885
rect 3491 827 3559 849
rect 3491 826 3507 827
rect 3491 792 3505 826
rect 3541 793 3559 827
rect 3539 792 3559 793
rect 3491 775 3559 792
rect 3604 840 3659 856
rect 3604 806 3625 840
rect 3604 790 3659 806
rect 3693 840 3729 890
rect 3884 1057 3926 1099
rect 4416 1091 4698 1130
rect 4838 1109 4854 1143
rect 4888 1109 4904 1143
rect 4416 1066 4455 1091
rect 3884 1023 3892 1057
rect 3884 989 3926 1023
rect 3884 955 3892 989
rect 3884 921 3926 955
rect 3884 887 3892 921
rect 3884 871 3926 887
rect 3960 1057 4026 1065
rect 3960 1023 3976 1057
rect 4010 1023 4026 1057
rect 3960 989 4026 1023
rect 3960 955 3976 989
rect 4010 955 4026 989
rect 3960 921 4026 955
rect 3960 887 3976 921
rect 4010 887 4026 921
rect 3960 869 4026 887
rect 3693 838 3734 840
rect 3693 804 3698 838
rect 3732 804 3734 838
rect 3693 802 3734 804
rect 3880 832 3946 835
rect 2718 717 2964 734
rect 2684 700 2964 717
rect 2684 698 2718 700
rect 2072 669 2414 690
rect 2072 635 2088 669
rect 2122 658 2414 669
rect 2122 655 2590 658
rect 2122 654 2540 655
rect 2122 635 2144 654
rect 2072 630 2144 635
rect 2072 623 2138 630
rect 2378 622 2540 654
rect 2524 621 2540 622
rect 2574 621 2590 655
rect 2916 612 2964 700
rect 1928 555 1957 589
rect 1991 555 2049 589
rect 2083 555 2141 589
rect 2175 555 2204 589
rect 2286 584 2332 594
rect 2286 550 2292 584
rect 2326 564 2332 584
rect 2916 578 2924 612
rect 2958 578 2964 612
rect 3188 711 3200 745
rect 3188 677 3234 711
rect 3188 643 3200 677
rect 3188 597 3234 643
rect 3268 745 3334 757
rect 3268 694 3284 745
rect 3318 694 3334 745
rect 3604 739 3638 790
rect 3268 677 3334 694
rect 3268 643 3284 677
rect 3318 643 3334 677
rect 3268 631 3334 643
rect 3505 705 3638 739
rect 3693 730 3729 802
rect 3880 798 3894 832
rect 3928 821 3946 832
rect 3880 787 3896 798
rect 3930 787 3946 821
rect 3505 684 3539 705
rect 3677 701 3729 730
rect 3505 629 3539 650
rect 3575 637 3591 671
rect 3625 637 3641 671
rect 2326 550 2336 564
rect 316 444 448 480
rect 620 490 654 506
rect 716 490 750 506
rect 654 454 655 455
rect 316 396 352 444
rect 620 420 655 454
rect 654 418 655 420
rect 716 420 750 454
rect 500 396 620 418
rect 316 384 620 396
rect 654 384 656 418
rect 316 382 656 384
rect 316 360 536 382
rect 620 368 654 382
rect 716 368 750 384
rect 812 490 846 506
rect 2286 480 2336 550
rect 2636 540 2652 574
rect 2686 540 2702 574
rect 2916 566 2964 578
rect 3124 563 3153 597
rect 3187 563 3245 597
rect 3279 563 3337 597
rect 3371 563 3400 597
rect 3575 595 3641 637
rect 3711 667 3729 701
rect 3677 629 3729 667
rect 3880 737 3926 753
rect 3980 749 4026 869
rect 4164 1047 4198 1066
rect 4250 1057 4455 1066
rect 4489 1089 4698 1091
rect 4489 1057 4574 1089
rect 4250 1055 4574 1057
rect 4608 1066 4698 1089
rect 4938 1066 4972 1424
rect 5882 1398 5916 1609
rect 6113 1306 6147 1609
rect 6198 1390 6232 2004
rect 6398 2002 6464 2004
rect 6715 2009 6731 2043
rect 6765 2009 6781 2043
rect 6715 1975 6781 2009
rect 6270 1943 6304 1962
rect 6270 1875 6304 1877
rect 6270 1839 6304 1841
rect 6270 1754 6304 1773
rect 6366 1943 6400 1962
rect 6366 1875 6400 1877
rect 6366 1839 6400 1841
rect 6366 1754 6400 1773
rect 6462 1943 6496 1962
rect 6715 1941 6731 1975
rect 6765 1959 6781 1975
rect 6887 2111 6953 2153
rect 6921 2077 6953 2111
rect 6887 2043 6953 2077
rect 6921 2009 6953 2043
rect 6887 1975 6953 2009
rect 6765 1941 6851 1959
rect 6715 1925 6851 1941
rect 6921 1941 6953 1975
rect 6887 1925 6953 1941
rect 7789 2111 7855 2116
rect 7789 2077 7805 2111
rect 7839 2077 7855 2111
rect 7789 2043 7855 2077
rect 7789 2009 7805 2043
rect 7839 2009 7855 2043
rect 7789 1975 7855 2009
rect 7789 1941 7805 1975
rect 7839 1959 7855 1975
rect 7961 2111 8027 2153
rect 7995 2077 8027 2111
rect 8194 2147 8476 2153
rect 8194 2113 8233 2147
rect 8267 2145 8476 2147
rect 8267 2113 8352 2145
rect 8194 2111 8352 2113
rect 8386 2111 8476 2145
rect 8194 2078 8476 2111
rect 8603 2111 8669 2116
rect 7961 2043 8027 2077
rect 7995 2009 8027 2043
rect 8603 2077 8619 2111
rect 8653 2077 8669 2111
rect 8603 2043 8669 2077
rect 7961 1975 8027 2009
rect 7839 1941 7925 1959
rect 7789 1925 7925 1941
rect 7995 1941 8027 1975
rect 7961 1925 8027 1941
rect 8086 2039 8352 2040
rect 8086 2005 8302 2039
rect 8336 2005 8352 2039
rect 8086 2004 8352 2005
rect 6462 1875 6496 1877
rect 6713 1882 6783 1891
rect 6713 1848 6729 1882
rect 6763 1875 6783 1882
rect 6713 1841 6733 1848
rect 6767 1841 6783 1875
rect 6462 1839 6496 1841
rect 6817 1805 6851 1925
rect 6885 1882 6955 1891
rect 6885 1875 6903 1882
rect 6885 1841 6901 1875
rect 6937 1848 6955 1882
rect 6935 1841 6955 1848
rect 7787 1884 7857 1891
rect 7787 1850 7805 1884
rect 7839 1875 7857 1884
rect 7787 1841 7807 1850
rect 7841 1841 7857 1875
rect 7891 1805 7925 1925
rect 7959 1880 8029 1891
rect 7959 1875 7978 1880
rect 7959 1841 7975 1875
rect 8012 1846 8029 1880
rect 8009 1841 8029 1846
rect 6462 1754 6496 1773
rect 6717 1789 6765 1805
rect 6717 1755 6731 1789
rect 6717 1721 6765 1755
rect 6302 1677 6318 1711
rect 6352 1677 6368 1711
rect 6717 1687 6731 1721
rect 6717 1643 6765 1687
rect 6799 1789 6865 1805
rect 6799 1755 6815 1789
rect 6849 1759 6865 1789
rect 6799 1725 6817 1755
rect 6851 1725 6865 1759
rect 6799 1721 6865 1725
rect 6799 1687 6815 1721
rect 6849 1687 6865 1721
rect 6799 1677 6865 1687
rect 6899 1789 6953 1805
rect 6933 1755 6953 1789
rect 6899 1721 6953 1755
rect 6933 1687 6953 1721
rect 6899 1643 6953 1687
rect 7791 1789 7839 1805
rect 7791 1755 7805 1789
rect 7791 1721 7839 1755
rect 7791 1687 7805 1721
rect 7791 1643 7839 1687
rect 7873 1789 7939 1805
rect 7873 1764 7889 1789
rect 7873 1730 7887 1764
rect 7923 1755 7939 1789
rect 7921 1730 7939 1755
rect 7873 1721 7939 1730
rect 7873 1687 7889 1721
rect 7923 1687 7939 1721
rect 7873 1677 7939 1687
rect 7973 1789 8027 1805
rect 8007 1755 8027 1789
rect 7973 1721 8027 1755
rect 8007 1687 8027 1721
rect 7973 1643 8027 1687
rect 6414 1596 6430 1630
rect 6464 1596 6480 1630
rect 6696 1609 6725 1643
rect 6759 1609 6817 1643
rect 6851 1609 6909 1643
rect 6943 1609 6972 1643
rect 7770 1609 7799 1643
rect 7833 1609 7891 1643
rect 7925 1609 7983 1643
rect 8017 1609 8046 1643
rect 6286 1546 6320 1562
rect 6286 1476 6320 1510
rect 6286 1424 6320 1440
rect 6382 1546 6416 1562
rect 6382 1476 6416 1510
rect 6382 1424 6416 1440
rect 6478 1546 6512 1562
rect 6478 1476 6512 1510
rect 6512 1440 6860 1464
rect 6478 1424 6860 1440
rect 6198 1356 6334 1390
rect 6368 1356 6384 1390
rect 6113 1286 6508 1306
rect 6113 1281 6375 1286
rect 6113 1272 6254 1281
rect 6238 1247 6254 1272
rect 6288 1252 6375 1281
rect 6409 1262 6508 1286
rect 6680 1264 6726 1266
rect 6680 1262 6684 1264
rect 6409 1252 6684 1262
rect 6288 1247 6684 1252
rect 6238 1230 6684 1247
rect 6718 1230 6726 1264
rect 6238 1228 6726 1230
rect 6680 1222 6726 1228
rect 5012 1107 5041 1141
rect 5075 1107 5133 1141
rect 5167 1107 5225 1141
rect 5259 1107 5288 1141
rect 4608 1055 4844 1066
rect 4250 1047 4844 1055
rect 4250 1022 4252 1047
rect 4164 979 4198 981
rect 4164 943 4198 945
rect 4164 858 4198 877
rect 4286 1022 4810 1047
rect 4896 1047 4972 1066
rect 4896 1026 4898 1047
rect 4252 979 4286 981
rect 4508 949 4524 983
rect 4558 949 4574 983
rect 4810 979 4844 981
rect 4252 943 4286 945
rect 4810 943 4844 945
rect 4252 858 4286 877
rect 4380 887 4414 906
rect 4380 819 4414 821
rect 4192 781 4208 815
rect 4242 781 4258 815
rect 4380 783 4414 785
rect 3880 703 3892 737
rect 3880 669 3926 703
rect 3880 635 3892 669
rect 3470 561 3499 595
rect 3533 561 3591 595
rect 3625 561 3683 595
rect 3717 561 3746 595
rect 3880 589 3926 635
rect 3960 737 4026 749
rect 3960 703 3976 737
rect 4010 703 4026 737
rect 3960 690 4026 703
rect 4380 698 4414 717
rect 4476 887 4510 906
rect 4476 819 4510 821
rect 4476 783 4510 785
rect 4476 698 4510 717
rect 4572 887 4606 906
rect 4810 858 4844 877
rect 4932 1026 4972 1047
rect 5080 1065 5122 1107
rect 5358 1105 5387 1139
rect 5421 1105 5479 1139
rect 5513 1105 5571 1139
rect 5605 1105 5634 1139
rect 5779 1133 5813 1140
rect 5080 1031 5088 1065
rect 4898 979 4932 981
rect 4898 943 4932 945
rect 5080 997 5122 1031
rect 5080 963 5088 997
rect 5080 929 5122 963
rect 5080 895 5088 929
rect 5080 879 5122 895
rect 5156 1065 5222 1073
rect 5156 1031 5172 1065
rect 5206 1031 5222 1065
rect 5156 997 5222 1031
rect 5156 963 5172 997
rect 5206 963 5222 997
rect 5156 929 5222 963
rect 5156 895 5172 929
rect 5206 895 5222 929
rect 5156 877 5222 895
rect 5391 1055 5427 1071
rect 5391 1021 5393 1055
rect 5391 987 5427 1021
rect 5391 953 5393 987
rect 5463 1055 5529 1105
rect 5704 1099 5733 1133
rect 5767 1099 5825 1133
rect 5859 1099 5917 1133
rect 5951 1099 5980 1133
rect 6080 1109 6096 1143
rect 6130 1109 6146 1143
rect 6304 1130 6418 1132
rect 5463 1021 5479 1055
rect 5513 1021 5529 1055
rect 5463 987 5529 1021
rect 5463 953 5479 987
rect 5513 953 5529 987
rect 5563 1055 5617 1071
rect 5563 1021 5565 1055
rect 5599 1021 5617 1055
rect 5563 974 5617 1021
rect 5391 919 5427 953
rect 5563 940 5565 974
rect 5599 940 5617 974
rect 5391 885 5526 919
rect 5563 890 5617 940
rect 4898 858 4932 877
rect 4572 819 4606 821
rect 4984 843 5128 844
rect 4984 829 5142 843
rect 4572 783 4606 785
rect 4838 816 4904 818
rect 4984 816 5092 829
rect 4838 815 5092 816
rect 4838 781 4854 815
rect 4888 802 5092 815
rect 4888 782 5024 802
rect 5076 795 5092 802
rect 5126 795 5142 829
rect 4888 781 4904 782
rect 5076 745 5122 761
rect 5176 757 5222 877
rect 5492 856 5526 885
rect 5379 827 5447 849
rect 5379 826 5395 827
rect 5379 792 5393 826
rect 5429 793 5447 827
rect 5427 792 5447 793
rect 5379 775 5447 792
rect 5492 840 5547 856
rect 5492 806 5513 840
rect 5492 790 5547 806
rect 5581 840 5617 890
rect 5772 1057 5814 1099
rect 6304 1091 6586 1130
rect 6726 1109 6742 1143
rect 6776 1109 6792 1143
rect 6304 1066 6343 1091
rect 5772 1023 5780 1057
rect 5772 989 5814 1023
rect 5772 955 5780 989
rect 5772 921 5814 955
rect 5772 887 5780 921
rect 5772 871 5814 887
rect 5848 1057 5914 1065
rect 5848 1023 5864 1057
rect 5898 1023 5914 1057
rect 5848 989 5914 1023
rect 5848 955 5864 989
rect 5898 955 5914 989
rect 5848 921 5914 955
rect 5848 887 5864 921
rect 5898 887 5914 921
rect 5848 869 5914 887
rect 5581 838 5622 840
rect 5581 804 5586 838
rect 5620 804 5622 838
rect 5581 802 5622 804
rect 5768 832 5834 835
rect 4606 717 4852 734
rect 4572 700 4852 717
rect 4572 698 4606 700
rect 3960 669 4302 690
rect 3960 635 3976 669
rect 4010 658 4302 669
rect 4010 655 4478 658
rect 4010 654 4428 655
rect 4010 635 4032 654
rect 3960 630 4032 635
rect 3960 623 4026 630
rect 4266 622 4428 654
rect 4412 621 4428 622
rect 4462 621 4478 655
rect 4804 612 4852 700
rect 3816 555 3845 589
rect 3879 555 3937 589
rect 3971 555 4029 589
rect 4063 555 4092 589
rect 4174 584 4220 594
rect 4174 550 4180 584
rect 4214 564 4220 584
rect 4804 578 4812 612
rect 4846 578 4852 612
rect 5076 711 5088 745
rect 5076 677 5122 711
rect 5076 643 5088 677
rect 5076 597 5122 643
rect 5156 745 5222 757
rect 5156 694 5172 745
rect 5206 694 5222 745
rect 5492 739 5526 790
rect 5156 677 5222 694
rect 5156 643 5172 677
rect 5206 643 5222 677
rect 5156 631 5222 643
rect 5393 705 5526 739
rect 5581 730 5617 802
rect 5768 798 5782 832
rect 5816 821 5834 832
rect 5768 787 5784 798
rect 5818 787 5834 821
rect 5393 684 5427 705
rect 5565 701 5617 730
rect 5393 629 5427 650
rect 5463 637 5479 671
rect 5513 637 5529 671
rect 4214 550 4224 564
rect 812 420 846 454
rect 812 368 846 384
rect 2204 444 2336 480
rect 2508 490 2542 506
rect 2604 490 2638 506
rect 2542 454 2543 455
rect 2204 396 2240 444
rect 2508 420 2543 454
rect 2542 418 2543 420
rect 2604 420 2638 454
rect 2388 396 2508 418
rect 2204 384 2508 396
rect 2542 384 2544 418
rect 2204 382 2544 384
rect 2204 360 2424 382
rect 2508 368 2542 382
rect 2604 368 2638 384
rect 2700 490 2734 506
rect 4174 480 4224 550
rect 4524 540 4540 574
rect 4574 540 4590 574
rect 4804 566 4852 578
rect 5012 563 5041 597
rect 5075 563 5133 597
rect 5167 563 5225 597
rect 5259 563 5288 597
rect 5463 595 5529 637
rect 5599 667 5617 701
rect 5565 629 5617 667
rect 5768 737 5814 753
rect 5868 749 5914 869
rect 6052 1047 6086 1066
rect 6138 1057 6343 1066
rect 6377 1089 6586 1091
rect 6377 1057 6462 1089
rect 6138 1055 6462 1057
rect 6496 1066 6586 1089
rect 6826 1066 6860 1424
rect 7770 1398 7804 1609
rect 8001 1306 8035 1609
rect 8086 1390 8120 2004
rect 8286 2002 8352 2004
rect 8603 2009 8619 2043
rect 8653 2009 8669 2043
rect 8603 1975 8669 2009
rect 8158 1943 8192 1962
rect 8158 1875 8192 1877
rect 8158 1839 8192 1841
rect 8158 1754 8192 1773
rect 8254 1943 8288 1962
rect 8254 1875 8288 1877
rect 8254 1839 8288 1841
rect 8254 1754 8288 1773
rect 8350 1943 8384 1962
rect 8603 1941 8619 1975
rect 8653 1959 8669 1975
rect 8775 2111 8841 2153
rect 8809 2077 8841 2111
rect 8775 2043 8841 2077
rect 8809 2009 8841 2043
rect 8775 1975 8841 2009
rect 8653 1941 8739 1959
rect 8603 1925 8739 1941
rect 8809 1941 8841 1975
rect 8775 1925 8841 1941
rect 9677 2111 9743 2116
rect 9677 2077 9693 2111
rect 9727 2077 9743 2111
rect 9677 2043 9743 2077
rect 9677 2009 9693 2043
rect 9727 2009 9743 2043
rect 9677 1975 9743 2009
rect 9677 1941 9693 1975
rect 9727 1959 9743 1975
rect 9849 2111 9915 2153
rect 9883 2077 9915 2111
rect 10082 2147 10364 2153
rect 10082 2113 10121 2147
rect 10155 2145 10364 2147
rect 10155 2113 10240 2145
rect 10082 2111 10240 2113
rect 10274 2111 10364 2145
rect 10082 2078 10364 2111
rect 10491 2111 10557 2116
rect 9849 2043 9915 2077
rect 9883 2009 9915 2043
rect 10491 2077 10507 2111
rect 10541 2077 10557 2111
rect 10491 2043 10557 2077
rect 9849 1975 9915 2009
rect 9727 1941 9813 1959
rect 9677 1925 9813 1941
rect 9883 1941 9915 1975
rect 9849 1925 9915 1941
rect 9974 2039 10240 2040
rect 9974 2005 10190 2039
rect 10224 2005 10240 2039
rect 9974 2004 10240 2005
rect 8350 1875 8384 1877
rect 8601 1882 8671 1891
rect 8601 1848 8617 1882
rect 8651 1875 8671 1882
rect 8601 1841 8621 1848
rect 8655 1841 8671 1875
rect 8350 1839 8384 1841
rect 8705 1805 8739 1925
rect 8773 1882 8843 1891
rect 8773 1875 8791 1882
rect 8773 1841 8789 1875
rect 8825 1848 8843 1882
rect 8823 1841 8843 1848
rect 9675 1884 9745 1891
rect 9675 1850 9693 1884
rect 9727 1875 9745 1884
rect 9675 1841 9695 1850
rect 9729 1841 9745 1875
rect 9779 1805 9813 1925
rect 9847 1880 9917 1891
rect 9847 1875 9866 1880
rect 9847 1841 9863 1875
rect 9900 1846 9917 1880
rect 9897 1841 9917 1846
rect 8350 1754 8384 1773
rect 8605 1789 8653 1805
rect 8605 1755 8619 1789
rect 8605 1721 8653 1755
rect 8190 1677 8206 1711
rect 8240 1677 8256 1711
rect 8605 1687 8619 1721
rect 8605 1643 8653 1687
rect 8687 1789 8753 1805
rect 8687 1755 8703 1789
rect 8737 1759 8753 1789
rect 8687 1725 8705 1755
rect 8739 1725 8753 1759
rect 8687 1721 8753 1725
rect 8687 1687 8703 1721
rect 8737 1687 8753 1721
rect 8687 1677 8753 1687
rect 8787 1789 8841 1805
rect 8821 1755 8841 1789
rect 8787 1721 8841 1755
rect 8821 1687 8841 1721
rect 8787 1643 8841 1687
rect 9679 1789 9727 1805
rect 9679 1755 9693 1789
rect 9679 1721 9727 1755
rect 9679 1687 9693 1721
rect 9679 1643 9727 1687
rect 9761 1789 9827 1805
rect 9761 1764 9777 1789
rect 9761 1730 9775 1764
rect 9811 1755 9827 1789
rect 9809 1730 9827 1755
rect 9761 1721 9827 1730
rect 9761 1687 9777 1721
rect 9811 1687 9827 1721
rect 9761 1677 9827 1687
rect 9861 1789 9915 1805
rect 9895 1755 9915 1789
rect 9861 1721 9915 1755
rect 9895 1687 9915 1721
rect 9861 1643 9915 1687
rect 8302 1596 8318 1630
rect 8352 1596 8368 1630
rect 8584 1609 8613 1643
rect 8647 1609 8705 1643
rect 8739 1609 8797 1643
rect 8831 1609 8860 1643
rect 9658 1609 9687 1643
rect 9721 1609 9779 1643
rect 9813 1609 9871 1643
rect 9905 1609 9934 1643
rect 8174 1546 8208 1562
rect 8174 1476 8208 1510
rect 8174 1424 8208 1440
rect 8270 1546 8304 1562
rect 8270 1476 8304 1510
rect 8270 1424 8304 1440
rect 8366 1546 8400 1562
rect 8366 1476 8400 1510
rect 8400 1440 8748 1464
rect 8366 1424 8748 1440
rect 8086 1356 8222 1390
rect 8256 1356 8272 1390
rect 8001 1286 8396 1306
rect 8001 1281 8263 1286
rect 8001 1272 8142 1281
rect 8126 1247 8142 1272
rect 8176 1252 8263 1281
rect 8297 1262 8396 1286
rect 8568 1264 8614 1266
rect 8568 1262 8572 1264
rect 8297 1252 8572 1262
rect 8176 1247 8572 1252
rect 8126 1230 8572 1247
rect 8606 1230 8614 1264
rect 8126 1228 8614 1230
rect 8568 1222 8614 1228
rect 6900 1107 6929 1141
rect 6963 1107 7021 1141
rect 7055 1107 7113 1141
rect 7147 1107 7176 1141
rect 6496 1055 6732 1066
rect 6138 1047 6732 1055
rect 6138 1022 6140 1047
rect 6052 979 6086 981
rect 6052 943 6086 945
rect 6052 858 6086 877
rect 6174 1022 6698 1047
rect 6784 1047 6860 1066
rect 6784 1026 6786 1047
rect 6140 979 6174 981
rect 6396 949 6412 983
rect 6446 949 6462 983
rect 6698 979 6732 981
rect 6140 943 6174 945
rect 6698 943 6732 945
rect 6140 858 6174 877
rect 6268 887 6302 906
rect 6268 819 6302 821
rect 6080 781 6096 815
rect 6130 781 6146 815
rect 6268 783 6302 785
rect 5768 703 5780 737
rect 5768 669 5814 703
rect 5768 635 5780 669
rect 5358 561 5387 595
rect 5421 561 5479 595
rect 5513 561 5571 595
rect 5605 561 5634 595
rect 5768 589 5814 635
rect 5848 737 5914 749
rect 5848 703 5864 737
rect 5898 703 5914 737
rect 5848 690 5914 703
rect 6268 698 6302 717
rect 6364 887 6398 906
rect 6364 819 6398 821
rect 6364 783 6398 785
rect 6364 698 6398 717
rect 6460 887 6494 906
rect 6698 858 6732 877
rect 6820 1026 6860 1047
rect 6968 1065 7010 1107
rect 7246 1105 7275 1139
rect 7309 1105 7367 1139
rect 7401 1105 7459 1139
rect 7493 1105 7522 1139
rect 7667 1133 7701 1140
rect 6968 1031 6976 1065
rect 6786 979 6820 981
rect 6786 943 6820 945
rect 6968 997 7010 1031
rect 6968 963 6976 997
rect 6968 929 7010 963
rect 6968 895 6976 929
rect 6968 879 7010 895
rect 7044 1065 7110 1073
rect 7044 1031 7060 1065
rect 7094 1031 7110 1065
rect 7044 997 7110 1031
rect 7044 963 7060 997
rect 7094 963 7110 997
rect 7044 929 7110 963
rect 7044 895 7060 929
rect 7094 895 7110 929
rect 7044 877 7110 895
rect 7279 1055 7315 1071
rect 7279 1021 7281 1055
rect 7279 987 7315 1021
rect 7279 953 7281 987
rect 7351 1055 7417 1105
rect 7592 1099 7621 1133
rect 7655 1099 7713 1133
rect 7747 1099 7805 1133
rect 7839 1099 7868 1133
rect 7968 1109 7984 1143
rect 8018 1109 8034 1143
rect 8192 1130 8306 1132
rect 7351 1021 7367 1055
rect 7401 1021 7417 1055
rect 7351 987 7417 1021
rect 7351 953 7367 987
rect 7401 953 7417 987
rect 7451 1055 7505 1071
rect 7451 1021 7453 1055
rect 7487 1021 7505 1055
rect 7451 974 7505 1021
rect 7279 919 7315 953
rect 7451 940 7453 974
rect 7487 940 7505 974
rect 7279 885 7414 919
rect 7451 890 7505 940
rect 6786 858 6820 877
rect 6460 819 6494 821
rect 6872 843 7016 844
rect 6872 829 7030 843
rect 6460 783 6494 785
rect 6726 816 6792 818
rect 6872 816 6980 829
rect 6726 815 6980 816
rect 6726 781 6742 815
rect 6776 802 6980 815
rect 6776 782 6912 802
rect 6964 795 6980 802
rect 7014 795 7030 829
rect 6776 781 6792 782
rect 6964 745 7010 761
rect 7064 757 7110 877
rect 7380 856 7414 885
rect 7267 827 7335 849
rect 7267 826 7283 827
rect 7267 792 7281 826
rect 7317 793 7335 827
rect 7315 792 7335 793
rect 7267 775 7335 792
rect 7380 840 7435 856
rect 7380 806 7401 840
rect 7380 790 7435 806
rect 7469 840 7505 890
rect 7660 1057 7702 1099
rect 8192 1091 8474 1130
rect 8614 1109 8630 1143
rect 8664 1109 8680 1143
rect 8192 1066 8231 1091
rect 7660 1023 7668 1057
rect 7660 989 7702 1023
rect 7660 955 7668 989
rect 7660 921 7702 955
rect 7660 887 7668 921
rect 7660 871 7702 887
rect 7736 1057 7802 1065
rect 7736 1023 7752 1057
rect 7786 1023 7802 1057
rect 7736 989 7802 1023
rect 7736 955 7752 989
rect 7786 955 7802 989
rect 7736 921 7802 955
rect 7736 887 7752 921
rect 7786 887 7802 921
rect 7736 869 7802 887
rect 7469 838 7510 840
rect 7469 804 7474 838
rect 7508 804 7510 838
rect 7469 802 7510 804
rect 7656 832 7722 835
rect 6494 717 6740 734
rect 6460 700 6740 717
rect 6460 698 6494 700
rect 5848 669 6190 690
rect 5848 635 5864 669
rect 5898 658 6190 669
rect 5898 655 6366 658
rect 5898 654 6316 655
rect 5898 635 5920 654
rect 5848 630 5920 635
rect 5848 623 5914 630
rect 6154 622 6316 654
rect 6300 621 6316 622
rect 6350 621 6366 655
rect 6692 612 6740 700
rect 5704 555 5733 589
rect 5767 555 5825 589
rect 5859 555 5917 589
rect 5951 555 5980 589
rect 6062 584 6108 594
rect 6062 550 6068 584
rect 6102 564 6108 584
rect 6692 578 6700 612
rect 6734 578 6740 612
rect 6964 711 6976 745
rect 6964 677 7010 711
rect 6964 643 6976 677
rect 6964 597 7010 643
rect 7044 745 7110 757
rect 7044 694 7060 745
rect 7094 694 7110 745
rect 7380 739 7414 790
rect 7044 677 7110 694
rect 7044 643 7060 677
rect 7094 643 7110 677
rect 7044 631 7110 643
rect 7281 705 7414 739
rect 7469 730 7505 802
rect 7656 798 7670 832
rect 7704 821 7722 832
rect 7656 787 7672 798
rect 7706 787 7722 821
rect 7281 684 7315 705
rect 7453 701 7505 730
rect 7281 629 7315 650
rect 7351 637 7367 671
rect 7401 637 7417 671
rect 6102 550 6112 564
rect 2700 420 2734 454
rect 2700 368 2734 384
rect 4092 444 4224 480
rect 4396 490 4430 506
rect 4492 490 4526 506
rect 4430 454 4431 455
rect 4092 396 4128 444
rect 4396 420 4431 454
rect 4430 418 4431 420
rect 4492 420 4526 454
rect 4276 396 4396 418
rect 4092 384 4396 396
rect 4430 384 4432 418
rect 4092 382 4432 384
rect 4092 360 4312 382
rect 4396 368 4430 382
rect 4492 368 4526 384
rect 4588 490 4622 506
rect 6062 480 6112 550
rect 6412 540 6428 574
rect 6462 540 6478 574
rect 6692 566 6740 578
rect 6900 563 6929 597
rect 6963 563 7021 597
rect 7055 563 7113 597
rect 7147 563 7176 597
rect 7351 595 7417 637
rect 7487 667 7505 701
rect 7453 629 7505 667
rect 7656 737 7702 753
rect 7756 749 7802 869
rect 7940 1047 7974 1066
rect 8026 1057 8231 1066
rect 8265 1089 8474 1091
rect 8265 1057 8350 1089
rect 8026 1055 8350 1057
rect 8384 1066 8474 1089
rect 8714 1066 8748 1424
rect 9658 1398 9692 1609
rect 9889 1306 9923 1609
rect 9974 1390 10008 2004
rect 10174 2002 10240 2004
rect 10491 2009 10507 2043
rect 10541 2009 10557 2043
rect 10491 1975 10557 2009
rect 10046 1943 10080 1962
rect 10046 1875 10080 1877
rect 10046 1839 10080 1841
rect 10046 1754 10080 1773
rect 10142 1943 10176 1962
rect 10142 1875 10176 1877
rect 10142 1839 10176 1841
rect 10142 1754 10176 1773
rect 10238 1943 10272 1962
rect 10491 1941 10507 1975
rect 10541 1959 10557 1975
rect 10663 2111 10729 2153
rect 10697 2077 10729 2111
rect 10663 2043 10729 2077
rect 10697 2009 10729 2043
rect 10663 1975 10729 2009
rect 10541 1941 10627 1959
rect 10491 1925 10627 1941
rect 10697 1941 10729 1975
rect 10663 1925 10729 1941
rect 11565 2111 11631 2116
rect 11565 2077 11581 2111
rect 11615 2077 11631 2111
rect 11565 2043 11631 2077
rect 11565 2009 11581 2043
rect 11615 2009 11631 2043
rect 11565 1975 11631 2009
rect 11565 1941 11581 1975
rect 11615 1959 11631 1975
rect 11737 2111 11803 2153
rect 11771 2077 11803 2111
rect 11970 2147 12252 2153
rect 11970 2113 12009 2147
rect 12043 2145 12252 2147
rect 12043 2113 12128 2145
rect 11970 2111 12128 2113
rect 12162 2111 12252 2145
rect 11970 2078 12252 2111
rect 12379 2111 12445 2116
rect 11737 2043 11803 2077
rect 11771 2009 11803 2043
rect 12379 2077 12395 2111
rect 12429 2077 12445 2111
rect 12379 2043 12445 2077
rect 11737 1975 11803 2009
rect 11615 1941 11701 1959
rect 11565 1925 11701 1941
rect 11771 1941 11803 1975
rect 11737 1925 11803 1941
rect 11862 2039 12128 2040
rect 11862 2005 12078 2039
rect 12112 2005 12128 2039
rect 11862 2004 12128 2005
rect 10238 1875 10272 1877
rect 10489 1882 10559 1891
rect 10489 1848 10505 1882
rect 10539 1875 10559 1882
rect 10489 1841 10509 1848
rect 10543 1841 10559 1875
rect 10238 1839 10272 1841
rect 10593 1805 10627 1925
rect 10661 1882 10731 1891
rect 10661 1875 10679 1882
rect 10661 1841 10677 1875
rect 10713 1848 10731 1882
rect 10711 1841 10731 1848
rect 11563 1884 11633 1891
rect 11563 1850 11581 1884
rect 11615 1875 11633 1884
rect 11563 1841 11583 1850
rect 11617 1841 11633 1875
rect 11667 1805 11701 1925
rect 11735 1880 11805 1891
rect 11735 1875 11754 1880
rect 11735 1841 11751 1875
rect 11788 1846 11805 1880
rect 11785 1841 11805 1846
rect 10238 1754 10272 1773
rect 10493 1789 10541 1805
rect 10493 1755 10507 1789
rect 10493 1721 10541 1755
rect 10078 1677 10094 1711
rect 10128 1677 10144 1711
rect 10493 1687 10507 1721
rect 10493 1643 10541 1687
rect 10575 1789 10641 1805
rect 10575 1755 10591 1789
rect 10625 1759 10641 1789
rect 10575 1725 10593 1755
rect 10627 1725 10641 1759
rect 10575 1721 10641 1725
rect 10575 1687 10591 1721
rect 10625 1687 10641 1721
rect 10575 1677 10641 1687
rect 10675 1789 10729 1805
rect 10709 1755 10729 1789
rect 10675 1721 10729 1755
rect 10709 1687 10729 1721
rect 10675 1643 10729 1687
rect 11567 1789 11615 1805
rect 11567 1755 11581 1789
rect 11567 1721 11615 1755
rect 11567 1687 11581 1721
rect 11567 1643 11615 1687
rect 11649 1789 11715 1805
rect 11649 1764 11665 1789
rect 11649 1730 11663 1764
rect 11699 1755 11715 1789
rect 11697 1730 11715 1755
rect 11649 1721 11715 1730
rect 11649 1687 11665 1721
rect 11699 1687 11715 1721
rect 11649 1677 11715 1687
rect 11749 1789 11803 1805
rect 11783 1755 11803 1789
rect 11749 1721 11803 1755
rect 11783 1687 11803 1721
rect 11749 1643 11803 1687
rect 10190 1596 10206 1630
rect 10240 1596 10256 1630
rect 10472 1609 10501 1643
rect 10535 1609 10593 1643
rect 10627 1609 10685 1643
rect 10719 1609 10748 1643
rect 11546 1609 11575 1643
rect 11609 1609 11667 1643
rect 11701 1609 11759 1643
rect 11793 1609 11822 1643
rect 10062 1546 10096 1562
rect 10062 1476 10096 1510
rect 10062 1424 10096 1440
rect 10158 1546 10192 1562
rect 10158 1476 10192 1510
rect 10158 1424 10192 1440
rect 10254 1546 10288 1562
rect 10254 1476 10288 1510
rect 10288 1440 10636 1464
rect 10254 1424 10636 1440
rect 9974 1356 10110 1390
rect 10144 1356 10160 1390
rect 9889 1286 10284 1306
rect 9889 1281 10151 1286
rect 9889 1272 10030 1281
rect 10014 1247 10030 1272
rect 10064 1252 10151 1281
rect 10185 1262 10284 1286
rect 10456 1264 10502 1266
rect 10456 1262 10460 1264
rect 10185 1252 10460 1262
rect 10064 1247 10460 1252
rect 10014 1230 10460 1247
rect 10494 1230 10502 1264
rect 10014 1228 10502 1230
rect 10456 1222 10502 1228
rect 8788 1107 8817 1141
rect 8851 1107 8909 1141
rect 8943 1107 9001 1141
rect 9035 1107 9064 1141
rect 8384 1055 8620 1066
rect 8026 1047 8620 1055
rect 8026 1022 8028 1047
rect 7940 979 7974 981
rect 7940 943 7974 945
rect 7940 858 7974 877
rect 8062 1022 8586 1047
rect 8672 1047 8748 1066
rect 8672 1026 8674 1047
rect 8028 979 8062 981
rect 8284 949 8300 983
rect 8334 949 8350 983
rect 8586 979 8620 981
rect 8028 943 8062 945
rect 8586 943 8620 945
rect 8028 858 8062 877
rect 8156 887 8190 906
rect 8156 819 8190 821
rect 7968 781 7984 815
rect 8018 781 8034 815
rect 8156 783 8190 785
rect 7656 703 7668 737
rect 7656 669 7702 703
rect 7656 635 7668 669
rect 7246 561 7275 595
rect 7309 561 7367 595
rect 7401 561 7459 595
rect 7493 561 7522 595
rect 7656 589 7702 635
rect 7736 737 7802 749
rect 7736 703 7752 737
rect 7786 703 7802 737
rect 7736 690 7802 703
rect 8156 698 8190 717
rect 8252 887 8286 906
rect 8252 819 8286 821
rect 8252 783 8286 785
rect 8252 698 8286 717
rect 8348 887 8382 906
rect 8586 858 8620 877
rect 8708 1026 8748 1047
rect 8856 1065 8898 1107
rect 9134 1105 9163 1139
rect 9197 1105 9255 1139
rect 9289 1105 9347 1139
rect 9381 1105 9410 1139
rect 9555 1133 9589 1140
rect 8856 1031 8864 1065
rect 8674 979 8708 981
rect 8674 943 8708 945
rect 8856 997 8898 1031
rect 8856 963 8864 997
rect 8856 929 8898 963
rect 8856 895 8864 929
rect 8856 879 8898 895
rect 8932 1065 8998 1073
rect 8932 1031 8948 1065
rect 8982 1031 8998 1065
rect 8932 997 8998 1031
rect 8932 963 8948 997
rect 8982 963 8998 997
rect 8932 929 8998 963
rect 8932 895 8948 929
rect 8982 895 8998 929
rect 8932 877 8998 895
rect 9167 1055 9203 1071
rect 9167 1021 9169 1055
rect 9167 987 9203 1021
rect 9167 953 9169 987
rect 9239 1055 9305 1105
rect 9480 1099 9509 1133
rect 9543 1099 9601 1133
rect 9635 1099 9693 1133
rect 9727 1099 9756 1133
rect 9856 1109 9872 1143
rect 9906 1109 9922 1143
rect 10080 1130 10194 1132
rect 9239 1021 9255 1055
rect 9289 1021 9305 1055
rect 9239 987 9305 1021
rect 9239 953 9255 987
rect 9289 953 9305 987
rect 9339 1055 9393 1071
rect 9339 1021 9341 1055
rect 9375 1021 9393 1055
rect 9339 974 9393 1021
rect 9167 919 9203 953
rect 9339 940 9341 974
rect 9375 940 9393 974
rect 9167 885 9302 919
rect 9339 890 9393 940
rect 8674 858 8708 877
rect 8348 819 8382 821
rect 8760 843 8904 844
rect 8760 829 8918 843
rect 8348 783 8382 785
rect 8614 816 8680 818
rect 8760 816 8868 829
rect 8614 815 8868 816
rect 8614 781 8630 815
rect 8664 802 8868 815
rect 8664 782 8800 802
rect 8852 795 8868 802
rect 8902 795 8918 829
rect 8664 781 8680 782
rect 8852 745 8898 761
rect 8952 757 8998 877
rect 9268 856 9302 885
rect 9155 827 9223 849
rect 9155 826 9171 827
rect 9155 792 9169 826
rect 9205 793 9223 827
rect 9203 792 9223 793
rect 9155 775 9223 792
rect 9268 840 9323 856
rect 9268 806 9289 840
rect 9268 790 9323 806
rect 9357 840 9393 890
rect 9548 1057 9590 1099
rect 10080 1091 10362 1130
rect 10502 1109 10518 1143
rect 10552 1109 10568 1143
rect 10080 1066 10119 1091
rect 9548 1023 9556 1057
rect 9548 989 9590 1023
rect 9548 955 9556 989
rect 9548 921 9590 955
rect 9548 887 9556 921
rect 9548 871 9590 887
rect 9624 1057 9690 1065
rect 9624 1023 9640 1057
rect 9674 1023 9690 1057
rect 9624 989 9690 1023
rect 9624 955 9640 989
rect 9674 955 9690 989
rect 9624 921 9690 955
rect 9624 887 9640 921
rect 9674 887 9690 921
rect 9624 869 9690 887
rect 9357 838 9398 840
rect 9357 804 9362 838
rect 9396 804 9398 838
rect 9357 802 9398 804
rect 9544 832 9610 835
rect 8382 717 8628 734
rect 8348 700 8628 717
rect 8348 698 8382 700
rect 7736 669 8078 690
rect 7736 635 7752 669
rect 7786 658 8078 669
rect 7786 655 8254 658
rect 7786 654 8204 655
rect 7786 635 7808 654
rect 7736 630 7808 635
rect 7736 623 7802 630
rect 8042 622 8204 654
rect 8188 621 8204 622
rect 8238 621 8254 655
rect 8580 612 8628 700
rect 7592 555 7621 589
rect 7655 555 7713 589
rect 7747 555 7805 589
rect 7839 555 7868 589
rect 7950 584 7996 594
rect 7950 550 7956 584
rect 7990 564 7996 584
rect 8580 578 8588 612
rect 8622 578 8628 612
rect 8852 711 8864 745
rect 8852 677 8898 711
rect 8852 643 8864 677
rect 8852 597 8898 643
rect 8932 745 8998 757
rect 8932 694 8948 745
rect 8982 694 8998 745
rect 9268 739 9302 790
rect 8932 677 8998 694
rect 8932 643 8948 677
rect 8982 643 8998 677
rect 8932 631 8998 643
rect 9169 705 9302 739
rect 9357 730 9393 802
rect 9544 798 9558 832
rect 9592 821 9610 832
rect 9544 787 9560 798
rect 9594 787 9610 821
rect 9169 684 9203 705
rect 9341 701 9393 730
rect 9169 629 9203 650
rect 9239 637 9255 671
rect 9289 637 9305 671
rect 7990 550 8000 564
rect 4588 420 4622 454
rect 4588 368 4622 384
rect 5980 444 6112 480
rect 6284 490 6318 506
rect 6380 490 6414 506
rect 6318 454 6319 455
rect 5980 396 6016 444
rect 6284 420 6319 454
rect 6318 418 6319 420
rect 6380 420 6414 454
rect 6164 396 6284 418
rect 5980 384 6284 396
rect 6318 384 6320 418
rect 5980 382 6320 384
rect 5980 360 6200 382
rect 6284 368 6318 382
rect 6380 368 6414 384
rect 6476 490 6510 506
rect 7950 480 8000 550
rect 8300 540 8316 574
rect 8350 540 8366 574
rect 8580 566 8628 578
rect 8788 563 8817 597
rect 8851 563 8909 597
rect 8943 563 9001 597
rect 9035 563 9064 597
rect 9239 595 9305 637
rect 9375 667 9393 701
rect 9341 629 9393 667
rect 9544 737 9590 753
rect 9644 749 9690 869
rect 9828 1047 9862 1066
rect 9914 1057 10119 1066
rect 10153 1089 10362 1091
rect 10153 1057 10238 1089
rect 9914 1055 10238 1057
rect 10272 1066 10362 1089
rect 10602 1066 10636 1424
rect 11546 1398 11580 1609
rect 11777 1306 11811 1609
rect 11862 1390 11896 2004
rect 12062 2002 12128 2004
rect 12379 2009 12395 2043
rect 12429 2009 12445 2043
rect 12379 1975 12445 2009
rect 11934 1943 11968 1962
rect 11934 1875 11968 1877
rect 11934 1839 11968 1841
rect 11934 1754 11968 1773
rect 12030 1943 12064 1962
rect 12030 1875 12064 1877
rect 12030 1839 12064 1841
rect 12030 1754 12064 1773
rect 12126 1943 12160 1962
rect 12379 1941 12395 1975
rect 12429 1959 12445 1975
rect 12551 2111 12617 2153
rect 12585 2077 12617 2111
rect 12551 2043 12617 2077
rect 12585 2009 12617 2043
rect 12551 1975 12617 2009
rect 12429 1941 12515 1959
rect 12379 1925 12515 1941
rect 12585 1941 12617 1975
rect 12551 1925 12617 1941
rect 13453 2111 13519 2116
rect 13453 2077 13469 2111
rect 13503 2077 13519 2111
rect 13453 2043 13519 2077
rect 13453 2009 13469 2043
rect 13503 2009 13519 2043
rect 13453 1975 13519 2009
rect 13453 1941 13469 1975
rect 13503 1959 13519 1975
rect 13625 2111 13691 2153
rect 13659 2077 13691 2111
rect 13858 2147 14140 2153
rect 13858 2113 13897 2147
rect 13931 2145 14140 2147
rect 13931 2113 14016 2145
rect 13858 2111 14016 2113
rect 14050 2111 14140 2145
rect 13858 2078 14140 2111
rect 14267 2111 14333 2116
rect 13625 2043 13691 2077
rect 13659 2009 13691 2043
rect 14267 2077 14283 2111
rect 14317 2077 14333 2111
rect 14267 2043 14333 2077
rect 13625 1975 13691 2009
rect 13503 1941 13589 1959
rect 13453 1925 13589 1941
rect 13659 1941 13691 1975
rect 13625 1925 13691 1941
rect 13750 2039 14016 2040
rect 13750 2005 13966 2039
rect 14000 2005 14016 2039
rect 13750 2004 14016 2005
rect 12126 1875 12160 1877
rect 12377 1882 12447 1891
rect 12377 1848 12393 1882
rect 12427 1875 12447 1882
rect 12377 1841 12397 1848
rect 12431 1841 12447 1875
rect 12126 1839 12160 1841
rect 12481 1805 12515 1925
rect 12549 1882 12619 1891
rect 12549 1875 12567 1882
rect 12549 1841 12565 1875
rect 12601 1848 12619 1882
rect 12599 1841 12619 1848
rect 13451 1884 13521 1891
rect 13451 1850 13469 1884
rect 13503 1875 13521 1884
rect 13451 1841 13471 1850
rect 13505 1841 13521 1875
rect 13555 1805 13589 1925
rect 13623 1880 13693 1891
rect 13623 1875 13642 1880
rect 13623 1841 13639 1875
rect 13676 1846 13693 1880
rect 13673 1841 13693 1846
rect 12126 1754 12160 1773
rect 12381 1789 12429 1805
rect 12381 1755 12395 1789
rect 12381 1721 12429 1755
rect 11966 1677 11982 1711
rect 12016 1677 12032 1711
rect 12381 1687 12395 1721
rect 12381 1643 12429 1687
rect 12463 1789 12529 1805
rect 12463 1755 12479 1789
rect 12513 1759 12529 1789
rect 12463 1725 12481 1755
rect 12515 1725 12529 1759
rect 12463 1721 12529 1725
rect 12463 1687 12479 1721
rect 12513 1687 12529 1721
rect 12463 1677 12529 1687
rect 12563 1789 12617 1805
rect 12597 1755 12617 1789
rect 12563 1721 12617 1755
rect 12597 1687 12617 1721
rect 12563 1643 12617 1687
rect 13455 1789 13503 1805
rect 13455 1755 13469 1789
rect 13455 1721 13503 1755
rect 13455 1687 13469 1721
rect 13455 1643 13503 1687
rect 13537 1789 13603 1805
rect 13537 1764 13553 1789
rect 13537 1730 13551 1764
rect 13587 1755 13603 1789
rect 13585 1730 13603 1755
rect 13537 1721 13603 1730
rect 13537 1687 13553 1721
rect 13587 1687 13603 1721
rect 13537 1677 13603 1687
rect 13637 1789 13691 1805
rect 13671 1755 13691 1789
rect 13637 1721 13691 1755
rect 13671 1687 13691 1721
rect 13637 1643 13691 1687
rect 12078 1596 12094 1630
rect 12128 1596 12144 1630
rect 12360 1609 12389 1643
rect 12423 1609 12481 1643
rect 12515 1609 12573 1643
rect 12607 1609 12636 1643
rect 13434 1609 13463 1643
rect 13497 1609 13555 1643
rect 13589 1609 13647 1643
rect 13681 1609 13710 1643
rect 11950 1546 11984 1562
rect 11950 1476 11984 1510
rect 11950 1424 11984 1440
rect 12046 1546 12080 1562
rect 12046 1476 12080 1510
rect 12046 1424 12080 1440
rect 12142 1546 12176 1562
rect 12142 1476 12176 1510
rect 12176 1440 12524 1464
rect 12142 1424 12524 1440
rect 11862 1356 11998 1390
rect 12032 1356 12048 1390
rect 11777 1286 12172 1306
rect 11777 1281 12039 1286
rect 11777 1272 11918 1281
rect 11902 1247 11918 1272
rect 11952 1252 12039 1281
rect 12073 1262 12172 1286
rect 12344 1264 12390 1266
rect 12344 1262 12348 1264
rect 12073 1252 12348 1262
rect 11952 1247 12348 1252
rect 11902 1230 12348 1247
rect 12382 1230 12390 1264
rect 11902 1228 12390 1230
rect 12344 1222 12390 1228
rect 10676 1107 10705 1141
rect 10739 1107 10797 1141
rect 10831 1107 10889 1141
rect 10923 1107 10952 1141
rect 10272 1055 10508 1066
rect 9914 1047 10508 1055
rect 9914 1022 9916 1047
rect 9828 979 9862 981
rect 9828 943 9862 945
rect 9828 858 9862 877
rect 9950 1022 10474 1047
rect 10560 1047 10636 1066
rect 10560 1026 10562 1047
rect 9916 979 9950 981
rect 10172 949 10188 983
rect 10222 949 10238 983
rect 10474 979 10508 981
rect 9916 943 9950 945
rect 10474 943 10508 945
rect 9916 858 9950 877
rect 10044 887 10078 906
rect 10044 819 10078 821
rect 9856 781 9872 815
rect 9906 781 9922 815
rect 10044 783 10078 785
rect 9544 703 9556 737
rect 9544 669 9590 703
rect 9544 635 9556 669
rect 9134 561 9163 595
rect 9197 561 9255 595
rect 9289 561 9347 595
rect 9381 561 9410 595
rect 9544 589 9590 635
rect 9624 737 9690 749
rect 9624 703 9640 737
rect 9674 703 9690 737
rect 9624 690 9690 703
rect 10044 698 10078 717
rect 10140 887 10174 906
rect 10140 819 10174 821
rect 10140 783 10174 785
rect 10140 698 10174 717
rect 10236 887 10270 906
rect 10474 858 10508 877
rect 10596 1026 10636 1047
rect 10744 1065 10786 1107
rect 11022 1105 11051 1139
rect 11085 1105 11143 1139
rect 11177 1105 11235 1139
rect 11269 1105 11298 1139
rect 11443 1133 11477 1140
rect 10744 1031 10752 1065
rect 10562 979 10596 981
rect 10562 943 10596 945
rect 10744 997 10786 1031
rect 10744 963 10752 997
rect 10744 929 10786 963
rect 10744 895 10752 929
rect 10744 879 10786 895
rect 10820 1065 10886 1073
rect 10820 1031 10836 1065
rect 10870 1031 10886 1065
rect 10820 997 10886 1031
rect 10820 963 10836 997
rect 10870 963 10886 997
rect 10820 929 10886 963
rect 10820 895 10836 929
rect 10870 895 10886 929
rect 10820 877 10886 895
rect 11055 1055 11091 1071
rect 11055 1021 11057 1055
rect 11055 987 11091 1021
rect 11055 953 11057 987
rect 11127 1055 11193 1105
rect 11368 1099 11397 1133
rect 11431 1099 11489 1133
rect 11523 1099 11581 1133
rect 11615 1099 11644 1133
rect 11744 1109 11760 1143
rect 11794 1109 11810 1143
rect 11968 1130 12082 1132
rect 11127 1021 11143 1055
rect 11177 1021 11193 1055
rect 11127 987 11193 1021
rect 11127 953 11143 987
rect 11177 953 11193 987
rect 11227 1055 11281 1071
rect 11227 1021 11229 1055
rect 11263 1021 11281 1055
rect 11227 974 11281 1021
rect 11055 919 11091 953
rect 11227 940 11229 974
rect 11263 940 11281 974
rect 11055 885 11190 919
rect 11227 890 11281 940
rect 10562 858 10596 877
rect 10236 819 10270 821
rect 10648 843 10792 844
rect 10648 829 10806 843
rect 10236 783 10270 785
rect 10502 816 10568 818
rect 10648 816 10756 829
rect 10502 815 10756 816
rect 10502 781 10518 815
rect 10552 802 10756 815
rect 10552 782 10688 802
rect 10740 795 10756 802
rect 10790 795 10806 829
rect 10552 781 10568 782
rect 10740 745 10786 761
rect 10840 757 10886 877
rect 11156 856 11190 885
rect 11043 827 11111 849
rect 11043 826 11059 827
rect 11043 792 11057 826
rect 11093 793 11111 827
rect 11091 792 11111 793
rect 11043 775 11111 792
rect 11156 840 11211 856
rect 11156 806 11177 840
rect 11156 790 11211 806
rect 11245 840 11281 890
rect 11436 1057 11478 1099
rect 11968 1091 12250 1130
rect 12390 1109 12406 1143
rect 12440 1109 12456 1143
rect 11968 1066 12007 1091
rect 11436 1023 11444 1057
rect 11436 989 11478 1023
rect 11436 955 11444 989
rect 11436 921 11478 955
rect 11436 887 11444 921
rect 11436 871 11478 887
rect 11512 1057 11578 1065
rect 11512 1023 11528 1057
rect 11562 1023 11578 1057
rect 11512 989 11578 1023
rect 11512 955 11528 989
rect 11562 955 11578 989
rect 11512 921 11578 955
rect 11512 887 11528 921
rect 11562 887 11578 921
rect 11512 869 11578 887
rect 11245 838 11286 840
rect 11245 804 11250 838
rect 11284 804 11286 838
rect 11245 802 11286 804
rect 11432 832 11498 835
rect 10270 717 10516 734
rect 10236 700 10516 717
rect 10236 698 10270 700
rect 9624 669 9966 690
rect 9624 635 9640 669
rect 9674 658 9966 669
rect 9674 655 10142 658
rect 9674 654 10092 655
rect 9674 635 9696 654
rect 9624 630 9696 635
rect 9624 623 9690 630
rect 9930 622 10092 654
rect 10076 621 10092 622
rect 10126 621 10142 655
rect 10468 612 10516 700
rect 9480 555 9509 589
rect 9543 555 9601 589
rect 9635 555 9693 589
rect 9727 555 9756 589
rect 9838 584 9884 594
rect 9838 550 9844 584
rect 9878 564 9884 584
rect 10468 578 10476 612
rect 10510 578 10516 612
rect 10740 711 10752 745
rect 10740 677 10786 711
rect 10740 643 10752 677
rect 10740 597 10786 643
rect 10820 745 10886 757
rect 10820 694 10836 745
rect 10870 694 10886 745
rect 11156 739 11190 790
rect 10820 677 10886 694
rect 10820 643 10836 677
rect 10870 643 10886 677
rect 10820 631 10886 643
rect 11057 705 11190 739
rect 11245 730 11281 802
rect 11432 798 11446 832
rect 11480 821 11498 832
rect 11432 787 11448 798
rect 11482 787 11498 821
rect 11057 684 11091 705
rect 11229 701 11281 730
rect 11057 629 11091 650
rect 11127 637 11143 671
rect 11177 637 11193 671
rect 9878 550 9888 564
rect 6476 420 6510 454
rect 6476 368 6510 384
rect 7868 444 8000 480
rect 8172 490 8206 506
rect 8268 490 8302 506
rect 8206 454 8207 455
rect 7868 396 7904 444
rect 8172 420 8207 454
rect 8206 418 8207 420
rect 8268 420 8302 454
rect 8052 396 8172 418
rect 7868 384 8172 396
rect 8206 384 8208 418
rect 7868 382 8208 384
rect 7868 360 8088 382
rect 8172 368 8206 382
rect 8268 368 8302 384
rect 8364 490 8398 506
rect 9838 480 9888 550
rect 10188 540 10204 574
rect 10238 540 10254 574
rect 10468 566 10516 578
rect 10676 563 10705 597
rect 10739 563 10797 597
rect 10831 563 10889 597
rect 10923 563 10952 597
rect 11127 595 11193 637
rect 11263 667 11281 701
rect 11229 629 11281 667
rect 11432 737 11478 753
rect 11532 749 11578 869
rect 11716 1047 11750 1066
rect 11802 1057 12007 1066
rect 12041 1089 12250 1091
rect 12041 1057 12126 1089
rect 11802 1055 12126 1057
rect 12160 1066 12250 1089
rect 12490 1066 12524 1424
rect 13434 1398 13468 1609
rect 13665 1306 13699 1609
rect 13750 1390 13784 2004
rect 13950 2002 14016 2004
rect 14267 2009 14283 2043
rect 14317 2009 14333 2043
rect 14267 1975 14333 2009
rect 13822 1943 13856 1962
rect 13822 1875 13856 1877
rect 13822 1839 13856 1841
rect 13822 1754 13856 1773
rect 13918 1943 13952 1962
rect 13918 1875 13952 1877
rect 13918 1839 13952 1841
rect 13918 1754 13952 1773
rect 14014 1943 14048 1962
rect 14267 1941 14283 1975
rect 14317 1959 14333 1975
rect 14439 2111 14505 2153
rect 14473 2077 14505 2111
rect 14439 2043 14505 2077
rect 14473 2009 14505 2043
rect 14439 1975 14505 2009
rect 14317 1941 14403 1959
rect 14267 1925 14403 1941
rect 14473 1941 14505 1975
rect 14439 1925 14505 1941
rect 15335 2111 15401 2116
rect 15335 2077 15351 2111
rect 15385 2077 15401 2111
rect 15335 2043 15401 2077
rect 15335 2009 15351 2043
rect 15385 2009 15401 2043
rect 15335 1975 15401 2009
rect 15335 1941 15351 1975
rect 15385 1959 15401 1975
rect 15507 2111 15573 2153
rect 15541 2077 15573 2111
rect 15740 2147 16022 2153
rect 15740 2113 15779 2147
rect 15813 2145 16022 2147
rect 15813 2113 15898 2145
rect 15740 2111 15898 2113
rect 15932 2111 16022 2145
rect 15740 2078 16022 2111
rect 16149 2111 16215 2116
rect 15507 2043 15573 2077
rect 15541 2009 15573 2043
rect 16149 2077 16165 2111
rect 16199 2077 16215 2111
rect 16149 2043 16215 2077
rect 15507 1975 15573 2009
rect 15385 1941 15471 1959
rect 15335 1925 15471 1941
rect 15541 1941 15573 1975
rect 15507 1925 15573 1941
rect 15632 2039 15898 2040
rect 15632 2005 15848 2039
rect 15882 2005 15898 2039
rect 15632 2004 15898 2005
rect 14014 1875 14048 1877
rect 14265 1882 14335 1891
rect 14265 1848 14281 1882
rect 14315 1875 14335 1882
rect 14265 1841 14285 1848
rect 14319 1841 14335 1875
rect 14014 1839 14048 1841
rect 14369 1805 14403 1925
rect 14437 1882 14507 1891
rect 14437 1875 14455 1882
rect 14437 1841 14453 1875
rect 14489 1848 14507 1882
rect 14487 1841 14507 1848
rect 15333 1884 15403 1891
rect 15333 1850 15351 1884
rect 15385 1875 15403 1884
rect 15333 1841 15353 1850
rect 15387 1841 15403 1875
rect 15437 1805 15471 1925
rect 15505 1880 15575 1891
rect 15505 1875 15524 1880
rect 15505 1841 15521 1875
rect 15558 1846 15575 1880
rect 15555 1841 15575 1846
rect 14014 1754 14048 1773
rect 14269 1789 14317 1805
rect 14269 1755 14283 1789
rect 14269 1721 14317 1755
rect 13854 1677 13870 1711
rect 13904 1677 13920 1711
rect 14269 1687 14283 1721
rect 14269 1643 14317 1687
rect 14351 1789 14417 1805
rect 14351 1755 14367 1789
rect 14401 1759 14417 1789
rect 14351 1725 14369 1755
rect 14403 1725 14417 1759
rect 14351 1721 14417 1725
rect 14351 1687 14367 1721
rect 14401 1687 14417 1721
rect 14351 1677 14417 1687
rect 14451 1789 14505 1805
rect 14485 1755 14505 1789
rect 14451 1721 14505 1755
rect 14485 1687 14505 1721
rect 14451 1643 14505 1687
rect 15337 1789 15385 1805
rect 15337 1755 15351 1789
rect 15337 1721 15385 1755
rect 15337 1687 15351 1721
rect 15337 1643 15385 1687
rect 15419 1789 15485 1805
rect 15419 1764 15435 1789
rect 15419 1730 15433 1764
rect 15469 1755 15485 1789
rect 15467 1730 15485 1755
rect 15419 1721 15485 1730
rect 15419 1687 15435 1721
rect 15469 1687 15485 1721
rect 15419 1677 15485 1687
rect 15519 1789 15573 1805
rect 15553 1755 15573 1789
rect 15519 1721 15573 1755
rect 15553 1687 15573 1721
rect 15519 1643 15573 1687
rect 13966 1596 13982 1630
rect 14016 1596 14032 1630
rect 14248 1609 14277 1643
rect 14311 1609 14369 1643
rect 14403 1609 14461 1643
rect 14495 1609 14524 1643
rect 15316 1609 15345 1643
rect 15379 1609 15437 1643
rect 15471 1609 15529 1643
rect 15563 1609 15592 1643
rect 13838 1546 13872 1562
rect 13838 1476 13872 1510
rect 13838 1424 13872 1440
rect 13934 1546 13968 1562
rect 13934 1476 13968 1510
rect 13934 1424 13968 1440
rect 14030 1546 14064 1562
rect 14030 1476 14064 1510
rect 14064 1440 14412 1464
rect 14030 1424 14412 1440
rect 13750 1356 13886 1390
rect 13920 1356 13936 1390
rect 13665 1286 14060 1306
rect 13665 1281 13927 1286
rect 13665 1272 13806 1281
rect 13790 1247 13806 1272
rect 13840 1252 13927 1281
rect 13961 1262 14060 1286
rect 14232 1264 14278 1266
rect 14232 1262 14236 1264
rect 13961 1252 14236 1262
rect 13840 1247 14236 1252
rect 13790 1230 14236 1247
rect 14270 1230 14278 1264
rect 13790 1228 14278 1230
rect 14232 1222 14278 1228
rect 12564 1107 12593 1141
rect 12627 1107 12685 1141
rect 12719 1107 12777 1141
rect 12811 1107 12840 1141
rect 12160 1055 12396 1066
rect 11802 1047 12396 1055
rect 11802 1022 11804 1047
rect 11716 979 11750 981
rect 11716 943 11750 945
rect 11716 858 11750 877
rect 11838 1022 12362 1047
rect 12448 1047 12524 1066
rect 12448 1026 12450 1047
rect 11804 979 11838 981
rect 12060 949 12076 983
rect 12110 949 12126 983
rect 12362 979 12396 981
rect 11804 943 11838 945
rect 12362 943 12396 945
rect 11804 858 11838 877
rect 11932 887 11966 906
rect 11932 819 11966 821
rect 11744 781 11760 815
rect 11794 781 11810 815
rect 11932 783 11966 785
rect 11432 703 11444 737
rect 11432 669 11478 703
rect 11432 635 11444 669
rect 11022 561 11051 595
rect 11085 561 11143 595
rect 11177 561 11235 595
rect 11269 561 11298 595
rect 11432 589 11478 635
rect 11512 737 11578 749
rect 11512 703 11528 737
rect 11562 703 11578 737
rect 11512 690 11578 703
rect 11932 698 11966 717
rect 12028 887 12062 906
rect 12028 819 12062 821
rect 12028 783 12062 785
rect 12028 698 12062 717
rect 12124 887 12158 906
rect 12362 858 12396 877
rect 12484 1026 12524 1047
rect 12632 1065 12674 1107
rect 12910 1105 12939 1139
rect 12973 1105 13031 1139
rect 13065 1105 13123 1139
rect 13157 1105 13186 1139
rect 13331 1133 13365 1140
rect 12632 1031 12640 1065
rect 12450 979 12484 981
rect 12450 943 12484 945
rect 12632 997 12674 1031
rect 12632 963 12640 997
rect 12632 929 12674 963
rect 12632 895 12640 929
rect 12632 879 12674 895
rect 12708 1065 12774 1073
rect 12708 1031 12724 1065
rect 12758 1031 12774 1065
rect 12708 997 12774 1031
rect 12708 963 12724 997
rect 12758 963 12774 997
rect 12708 929 12774 963
rect 12708 895 12724 929
rect 12758 895 12774 929
rect 12708 877 12774 895
rect 12943 1055 12979 1071
rect 12943 1021 12945 1055
rect 12943 987 12979 1021
rect 12943 953 12945 987
rect 13015 1055 13081 1105
rect 13256 1099 13285 1133
rect 13319 1099 13377 1133
rect 13411 1099 13469 1133
rect 13503 1099 13532 1133
rect 13632 1109 13648 1143
rect 13682 1109 13698 1143
rect 13856 1130 13970 1132
rect 13015 1021 13031 1055
rect 13065 1021 13081 1055
rect 13015 987 13081 1021
rect 13015 953 13031 987
rect 13065 953 13081 987
rect 13115 1055 13169 1071
rect 13115 1021 13117 1055
rect 13151 1021 13169 1055
rect 13115 974 13169 1021
rect 12943 919 12979 953
rect 13115 940 13117 974
rect 13151 940 13169 974
rect 12943 885 13078 919
rect 13115 890 13169 940
rect 12450 858 12484 877
rect 12124 819 12158 821
rect 12536 843 12680 844
rect 12536 829 12694 843
rect 12124 783 12158 785
rect 12390 816 12456 818
rect 12536 816 12644 829
rect 12390 815 12644 816
rect 12390 781 12406 815
rect 12440 802 12644 815
rect 12440 782 12576 802
rect 12628 795 12644 802
rect 12678 795 12694 829
rect 12440 781 12456 782
rect 12628 745 12674 761
rect 12728 757 12774 877
rect 13044 856 13078 885
rect 12931 827 12999 849
rect 12931 826 12947 827
rect 12931 792 12945 826
rect 12981 793 12999 827
rect 12979 792 12999 793
rect 12931 775 12999 792
rect 13044 840 13099 856
rect 13044 806 13065 840
rect 13044 790 13099 806
rect 13133 840 13169 890
rect 13324 1057 13366 1099
rect 13856 1091 14138 1130
rect 14278 1109 14294 1143
rect 14328 1109 14344 1143
rect 13856 1066 13895 1091
rect 13324 1023 13332 1057
rect 13324 989 13366 1023
rect 13324 955 13332 989
rect 13324 921 13366 955
rect 13324 887 13332 921
rect 13324 871 13366 887
rect 13400 1057 13466 1065
rect 13400 1023 13416 1057
rect 13450 1023 13466 1057
rect 13400 989 13466 1023
rect 13400 955 13416 989
rect 13450 955 13466 989
rect 13400 921 13466 955
rect 13400 887 13416 921
rect 13450 887 13466 921
rect 13400 869 13466 887
rect 13133 838 13174 840
rect 13133 804 13138 838
rect 13172 804 13174 838
rect 13133 802 13174 804
rect 13320 832 13386 835
rect 12158 717 12404 734
rect 12124 700 12404 717
rect 12124 698 12158 700
rect 11512 669 11854 690
rect 11512 635 11528 669
rect 11562 658 11854 669
rect 11562 655 12030 658
rect 11562 654 11980 655
rect 11562 635 11584 654
rect 11512 630 11584 635
rect 11512 623 11578 630
rect 11818 622 11980 654
rect 11964 621 11980 622
rect 12014 621 12030 655
rect 12356 612 12404 700
rect 11368 555 11397 589
rect 11431 555 11489 589
rect 11523 555 11581 589
rect 11615 555 11644 589
rect 11726 584 11772 594
rect 11726 550 11732 584
rect 11766 564 11772 584
rect 12356 578 12364 612
rect 12398 578 12404 612
rect 12628 711 12640 745
rect 12628 677 12674 711
rect 12628 643 12640 677
rect 12628 597 12674 643
rect 12708 745 12774 757
rect 12708 694 12724 745
rect 12758 694 12774 745
rect 13044 739 13078 790
rect 12708 677 12774 694
rect 12708 643 12724 677
rect 12758 643 12774 677
rect 12708 631 12774 643
rect 12945 705 13078 739
rect 13133 730 13169 802
rect 13320 798 13334 832
rect 13368 821 13386 832
rect 13320 787 13336 798
rect 13370 787 13386 821
rect 12945 684 12979 705
rect 13117 701 13169 730
rect 12945 629 12979 650
rect 13015 637 13031 671
rect 13065 637 13081 671
rect 11766 550 11776 564
rect 8364 420 8398 454
rect 8364 368 8398 384
rect 9756 444 9888 480
rect 10060 490 10094 506
rect 10156 490 10190 506
rect 10094 454 10095 455
rect 9756 396 9792 444
rect 10060 420 10095 454
rect 10094 418 10095 420
rect 10156 420 10190 454
rect 9940 396 10060 418
rect 9756 384 10060 396
rect 10094 384 10096 418
rect 9756 382 10096 384
rect 9756 360 9976 382
rect 10060 368 10094 382
rect 10156 368 10190 384
rect 10252 490 10286 506
rect 11726 480 11776 550
rect 12076 540 12092 574
rect 12126 540 12142 574
rect 12356 566 12404 578
rect 12564 563 12593 597
rect 12627 563 12685 597
rect 12719 563 12777 597
rect 12811 563 12840 597
rect 13015 595 13081 637
rect 13151 667 13169 701
rect 13117 629 13169 667
rect 13320 737 13366 753
rect 13420 749 13466 869
rect 13604 1047 13638 1066
rect 13690 1057 13895 1066
rect 13929 1089 14138 1091
rect 13929 1057 14014 1089
rect 13690 1055 14014 1057
rect 14048 1066 14138 1089
rect 14378 1066 14412 1424
rect 15316 1398 15350 1609
rect 15547 1306 15581 1609
rect 15632 1390 15666 2004
rect 15832 2002 15898 2004
rect 16149 2009 16165 2043
rect 16199 2009 16215 2043
rect 16149 1975 16215 2009
rect 15704 1943 15738 1962
rect 15704 1875 15738 1877
rect 15704 1839 15738 1841
rect 15704 1754 15738 1773
rect 15800 1943 15834 1962
rect 15800 1875 15834 1877
rect 15800 1839 15834 1841
rect 15800 1754 15834 1773
rect 15896 1943 15930 1962
rect 16149 1941 16165 1975
rect 16199 1959 16215 1975
rect 16321 2111 16387 2153
rect 16355 2077 16387 2111
rect 16321 2043 16387 2077
rect 16355 2009 16387 2043
rect 16321 1975 16387 2009
rect 16199 1941 16285 1959
rect 16149 1925 16285 1941
rect 16355 1941 16387 1975
rect 16321 1925 16387 1941
rect 17223 2111 17289 2116
rect 17223 2077 17239 2111
rect 17273 2077 17289 2111
rect 17223 2043 17289 2077
rect 17223 2009 17239 2043
rect 17273 2009 17289 2043
rect 17223 1975 17289 2009
rect 17223 1941 17239 1975
rect 17273 1959 17289 1975
rect 17395 2111 17461 2153
rect 17429 2077 17461 2111
rect 17628 2147 17910 2153
rect 17628 2113 17667 2147
rect 17701 2145 17910 2147
rect 17701 2113 17786 2145
rect 17628 2111 17786 2113
rect 17820 2111 17910 2145
rect 17628 2078 17910 2111
rect 18037 2111 18103 2116
rect 17395 2043 17461 2077
rect 17429 2009 17461 2043
rect 18037 2077 18053 2111
rect 18087 2077 18103 2111
rect 18037 2043 18103 2077
rect 17395 1975 17461 2009
rect 17273 1941 17359 1959
rect 17223 1925 17359 1941
rect 17429 1941 17461 1975
rect 17395 1925 17461 1941
rect 17520 2039 17786 2040
rect 17520 2005 17736 2039
rect 17770 2005 17786 2039
rect 17520 2004 17786 2005
rect 15896 1875 15930 1877
rect 16147 1882 16217 1891
rect 16147 1848 16163 1882
rect 16197 1875 16217 1882
rect 16147 1841 16167 1848
rect 16201 1841 16217 1875
rect 15896 1839 15930 1841
rect 16251 1805 16285 1925
rect 16319 1882 16389 1891
rect 16319 1875 16337 1882
rect 16319 1841 16335 1875
rect 16371 1848 16389 1882
rect 16369 1841 16389 1848
rect 17221 1884 17291 1891
rect 17221 1850 17239 1884
rect 17273 1875 17291 1884
rect 17221 1841 17241 1850
rect 17275 1841 17291 1875
rect 17325 1805 17359 1925
rect 17393 1880 17463 1891
rect 17393 1875 17412 1880
rect 17393 1841 17409 1875
rect 17446 1846 17463 1880
rect 17443 1841 17463 1846
rect 15896 1754 15930 1773
rect 16151 1789 16199 1805
rect 16151 1755 16165 1789
rect 16151 1721 16199 1755
rect 15736 1677 15752 1711
rect 15786 1677 15802 1711
rect 16151 1687 16165 1721
rect 16151 1643 16199 1687
rect 16233 1789 16299 1805
rect 16233 1755 16249 1789
rect 16283 1759 16299 1789
rect 16233 1725 16251 1755
rect 16285 1725 16299 1759
rect 16233 1721 16299 1725
rect 16233 1687 16249 1721
rect 16283 1687 16299 1721
rect 16233 1677 16299 1687
rect 16333 1789 16387 1805
rect 16367 1755 16387 1789
rect 16333 1721 16387 1755
rect 16367 1687 16387 1721
rect 16333 1643 16387 1687
rect 17225 1789 17273 1805
rect 17225 1755 17239 1789
rect 17225 1721 17273 1755
rect 17225 1687 17239 1721
rect 17225 1643 17273 1687
rect 17307 1789 17373 1805
rect 17307 1764 17323 1789
rect 17307 1730 17321 1764
rect 17357 1755 17373 1789
rect 17355 1730 17373 1755
rect 17307 1721 17373 1730
rect 17307 1687 17323 1721
rect 17357 1687 17373 1721
rect 17307 1677 17373 1687
rect 17407 1789 17461 1805
rect 17441 1755 17461 1789
rect 17407 1721 17461 1755
rect 17441 1687 17461 1721
rect 17407 1643 17461 1687
rect 15848 1596 15864 1630
rect 15898 1596 15914 1630
rect 16130 1609 16159 1643
rect 16193 1609 16251 1643
rect 16285 1609 16343 1643
rect 16377 1609 16406 1643
rect 17204 1609 17233 1643
rect 17267 1609 17325 1643
rect 17359 1609 17417 1643
rect 17451 1609 17480 1643
rect 15720 1546 15754 1562
rect 15720 1476 15754 1510
rect 15720 1424 15754 1440
rect 15816 1546 15850 1562
rect 15816 1476 15850 1510
rect 15816 1424 15850 1440
rect 15912 1546 15946 1562
rect 15912 1476 15946 1510
rect 15946 1440 16294 1464
rect 15912 1424 16294 1440
rect 15632 1356 15768 1390
rect 15802 1356 15818 1390
rect 15547 1286 15942 1306
rect 15547 1281 15809 1286
rect 15547 1272 15688 1281
rect 15672 1247 15688 1272
rect 15722 1252 15809 1281
rect 15843 1262 15942 1286
rect 16114 1264 16160 1266
rect 16114 1262 16118 1264
rect 15843 1252 16118 1262
rect 15722 1247 16118 1252
rect 15672 1230 16118 1247
rect 16152 1230 16160 1264
rect 15672 1228 16160 1230
rect 16114 1222 16160 1228
rect 14452 1107 14481 1141
rect 14515 1107 14573 1141
rect 14607 1107 14665 1141
rect 14699 1107 14728 1141
rect 14048 1055 14284 1066
rect 13690 1047 14284 1055
rect 13690 1022 13692 1047
rect 13604 979 13638 981
rect 13604 943 13638 945
rect 13604 858 13638 877
rect 13726 1022 14250 1047
rect 14336 1047 14412 1066
rect 14336 1026 14338 1047
rect 13692 979 13726 981
rect 13948 949 13964 983
rect 13998 949 14014 983
rect 14250 979 14284 981
rect 13692 943 13726 945
rect 14250 943 14284 945
rect 13692 858 13726 877
rect 13820 887 13854 906
rect 13820 819 13854 821
rect 13632 781 13648 815
rect 13682 781 13698 815
rect 13820 783 13854 785
rect 13320 703 13332 737
rect 13320 669 13366 703
rect 13320 635 13332 669
rect 12910 561 12939 595
rect 12973 561 13031 595
rect 13065 561 13123 595
rect 13157 561 13186 595
rect 13320 589 13366 635
rect 13400 737 13466 749
rect 13400 703 13416 737
rect 13450 703 13466 737
rect 13400 690 13466 703
rect 13820 698 13854 717
rect 13916 887 13950 906
rect 13916 819 13950 821
rect 13916 783 13950 785
rect 13916 698 13950 717
rect 14012 887 14046 906
rect 14250 858 14284 877
rect 14372 1026 14412 1047
rect 14520 1065 14562 1107
rect 14798 1105 14827 1139
rect 14861 1105 14919 1139
rect 14953 1105 15011 1139
rect 15045 1105 15074 1139
rect 15213 1133 15247 1140
rect 14520 1031 14528 1065
rect 14338 979 14372 981
rect 14338 943 14372 945
rect 14520 997 14562 1031
rect 14520 963 14528 997
rect 14520 929 14562 963
rect 14520 895 14528 929
rect 14520 879 14562 895
rect 14596 1065 14662 1073
rect 14596 1031 14612 1065
rect 14646 1031 14662 1065
rect 14596 997 14662 1031
rect 14596 963 14612 997
rect 14646 963 14662 997
rect 14596 929 14662 963
rect 14596 895 14612 929
rect 14646 895 14662 929
rect 14596 877 14662 895
rect 14831 1055 14867 1071
rect 14831 1021 14833 1055
rect 14831 987 14867 1021
rect 14831 953 14833 987
rect 14903 1055 14969 1105
rect 15138 1099 15167 1133
rect 15201 1099 15259 1133
rect 15293 1099 15351 1133
rect 15385 1099 15414 1133
rect 15514 1109 15530 1143
rect 15564 1109 15580 1143
rect 15738 1130 15852 1132
rect 14903 1021 14919 1055
rect 14953 1021 14969 1055
rect 14903 987 14969 1021
rect 14903 953 14919 987
rect 14953 953 14969 987
rect 15003 1055 15057 1071
rect 15003 1021 15005 1055
rect 15039 1021 15057 1055
rect 15003 974 15057 1021
rect 14831 919 14867 953
rect 15003 940 15005 974
rect 15039 940 15057 974
rect 14831 885 14966 919
rect 15003 890 15057 940
rect 14338 858 14372 877
rect 14012 819 14046 821
rect 14424 843 14568 844
rect 14424 829 14582 843
rect 14012 783 14046 785
rect 14278 816 14344 818
rect 14424 816 14532 829
rect 14278 815 14532 816
rect 14278 781 14294 815
rect 14328 802 14532 815
rect 14328 782 14464 802
rect 14516 795 14532 802
rect 14566 795 14582 829
rect 14328 781 14344 782
rect 14516 745 14562 761
rect 14616 757 14662 877
rect 14932 856 14966 885
rect 14819 827 14887 849
rect 14819 826 14835 827
rect 14819 792 14833 826
rect 14869 793 14887 827
rect 14867 792 14887 793
rect 14819 775 14887 792
rect 14932 840 14987 856
rect 14932 806 14953 840
rect 14932 790 14987 806
rect 15021 840 15057 890
rect 15206 1057 15248 1099
rect 15738 1091 16020 1130
rect 16160 1109 16176 1143
rect 16210 1109 16226 1143
rect 15738 1066 15777 1091
rect 15206 1023 15214 1057
rect 15206 989 15248 1023
rect 15206 955 15214 989
rect 15206 921 15248 955
rect 15206 887 15214 921
rect 15206 871 15248 887
rect 15282 1057 15348 1065
rect 15282 1023 15298 1057
rect 15332 1023 15348 1057
rect 15282 989 15348 1023
rect 15282 955 15298 989
rect 15332 955 15348 989
rect 15282 921 15348 955
rect 15282 887 15298 921
rect 15332 887 15348 921
rect 15282 869 15348 887
rect 15021 838 15062 840
rect 15021 804 15026 838
rect 15060 804 15062 838
rect 15021 802 15062 804
rect 15202 832 15268 835
rect 14046 717 14292 734
rect 14012 700 14292 717
rect 14012 698 14046 700
rect 13400 669 13742 690
rect 13400 635 13416 669
rect 13450 658 13742 669
rect 13450 655 13918 658
rect 13450 654 13868 655
rect 13450 635 13472 654
rect 13400 630 13472 635
rect 13400 623 13466 630
rect 13706 622 13868 654
rect 13852 621 13868 622
rect 13902 621 13918 655
rect 14244 612 14292 700
rect 13256 555 13285 589
rect 13319 555 13377 589
rect 13411 555 13469 589
rect 13503 555 13532 589
rect 13614 584 13660 594
rect 13614 550 13620 584
rect 13654 564 13660 584
rect 14244 578 14252 612
rect 14286 578 14292 612
rect 14516 711 14528 745
rect 14516 677 14562 711
rect 14516 643 14528 677
rect 14516 597 14562 643
rect 14596 745 14662 757
rect 14596 694 14612 745
rect 14646 694 14662 745
rect 14932 739 14966 790
rect 14596 677 14662 694
rect 14596 643 14612 677
rect 14646 643 14662 677
rect 14596 631 14662 643
rect 14833 705 14966 739
rect 15021 730 15057 802
rect 15202 798 15216 832
rect 15250 821 15268 832
rect 15202 787 15218 798
rect 15252 787 15268 821
rect 14833 684 14867 705
rect 15005 701 15057 730
rect 14833 629 14867 650
rect 14903 637 14919 671
rect 14953 637 14969 671
rect 13654 550 13664 564
rect 10252 420 10286 454
rect 10252 368 10286 384
rect 11644 444 11776 480
rect 11948 490 11982 506
rect 12044 490 12078 506
rect 11982 454 11983 455
rect 11644 396 11680 444
rect 11948 420 11983 454
rect 11982 418 11983 420
rect 12044 420 12078 454
rect 11828 396 11948 418
rect 11644 384 11948 396
rect 11982 384 11984 418
rect 11644 382 11984 384
rect 11644 360 11864 382
rect 11948 368 11982 382
rect 12044 368 12078 384
rect 12140 490 12174 506
rect 13614 480 13664 550
rect 13964 540 13980 574
rect 14014 540 14030 574
rect 14244 566 14292 578
rect 14452 563 14481 597
rect 14515 563 14573 597
rect 14607 563 14665 597
rect 14699 563 14728 597
rect 14903 595 14969 637
rect 15039 667 15057 701
rect 15005 629 15057 667
rect 15202 737 15248 753
rect 15302 749 15348 869
rect 15486 1047 15520 1066
rect 15572 1057 15777 1066
rect 15811 1089 16020 1091
rect 15811 1057 15896 1089
rect 15572 1055 15896 1057
rect 15930 1066 16020 1089
rect 16260 1066 16294 1424
rect 17204 1398 17238 1609
rect 17435 1306 17469 1609
rect 17520 1390 17554 2004
rect 17720 2002 17786 2004
rect 18037 2009 18053 2043
rect 18087 2009 18103 2043
rect 18037 1975 18103 2009
rect 17592 1943 17626 1962
rect 17592 1875 17626 1877
rect 17592 1839 17626 1841
rect 17592 1754 17626 1773
rect 17688 1943 17722 1962
rect 17688 1875 17722 1877
rect 17688 1839 17722 1841
rect 17688 1754 17722 1773
rect 17784 1943 17818 1962
rect 18037 1941 18053 1975
rect 18087 1959 18103 1975
rect 18209 2111 18275 2153
rect 18243 2077 18275 2111
rect 18209 2043 18275 2077
rect 18243 2009 18275 2043
rect 18209 1975 18275 2009
rect 18087 1941 18173 1959
rect 18037 1925 18173 1941
rect 18243 1941 18275 1975
rect 18209 1925 18275 1941
rect 19111 2111 19177 2116
rect 19111 2077 19127 2111
rect 19161 2077 19177 2111
rect 19111 2043 19177 2077
rect 19111 2009 19127 2043
rect 19161 2009 19177 2043
rect 19111 1975 19177 2009
rect 19111 1941 19127 1975
rect 19161 1959 19177 1975
rect 19283 2111 19349 2153
rect 19317 2077 19349 2111
rect 19516 2147 19798 2153
rect 19516 2113 19555 2147
rect 19589 2145 19798 2147
rect 19589 2113 19674 2145
rect 19516 2111 19674 2113
rect 19708 2111 19798 2145
rect 19516 2078 19798 2111
rect 19925 2111 19991 2116
rect 19283 2043 19349 2077
rect 19317 2009 19349 2043
rect 19925 2077 19941 2111
rect 19975 2077 19991 2111
rect 19925 2043 19991 2077
rect 19283 1975 19349 2009
rect 19161 1941 19247 1959
rect 19111 1925 19247 1941
rect 19317 1941 19349 1975
rect 19283 1925 19349 1941
rect 19408 2039 19674 2040
rect 19408 2005 19624 2039
rect 19658 2005 19674 2039
rect 19408 2004 19674 2005
rect 17784 1875 17818 1877
rect 18035 1882 18105 1891
rect 18035 1848 18051 1882
rect 18085 1875 18105 1882
rect 18035 1841 18055 1848
rect 18089 1841 18105 1875
rect 17784 1839 17818 1841
rect 18139 1805 18173 1925
rect 18207 1882 18277 1891
rect 18207 1875 18225 1882
rect 18207 1841 18223 1875
rect 18259 1848 18277 1882
rect 18257 1841 18277 1848
rect 19109 1884 19179 1891
rect 19109 1850 19127 1884
rect 19161 1875 19179 1884
rect 19109 1841 19129 1850
rect 19163 1841 19179 1875
rect 19213 1805 19247 1925
rect 19281 1880 19351 1891
rect 19281 1875 19300 1880
rect 19281 1841 19297 1875
rect 19334 1846 19351 1880
rect 19331 1841 19351 1846
rect 17784 1754 17818 1773
rect 18039 1789 18087 1805
rect 18039 1755 18053 1789
rect 18039 1721 18087 1755
rect 17624 1677 17640 1711
rect 17674 1677 17690 1711
rect 18039 1687 18053 1721
rect 18039 1643 18087 1687
rect 18121 1789 18187 1805
rect 18121 1755 18137 1789
rect 18171 1759 18187 1789
rect 18121 1725 18139 1755
rect 18173 1725 18187 1759
rect 18121 1721 18187 1725
rect 18121 1687 18137 1721
rect 18171 1687 18187 1721
rect 18121 1677 18187 1687
rect 18221 1789 18275 1805
rect 18255 1755 18275 1789
rect 18221 1721 18275 1755
rect 18255 1687 18275 1721
rect 18221 1643 18275 1687
rect 19113 1789 19161 1805
rect 19113 1755 19127 1789
rect 19113 1721 19161 1755
rect 19113 1687 19127 1721
rect 19113 1643 19161 1687
rect 19195 1789 19261 1805
rect 19195 1764 19211 1789
rect 19195 1730 19209 1764
rect 19245 1755 19261 1789
rect 19243 1730 19261 1755
rect 19195 1721 19261 1730
rect 19195 1687 19211 1721
rect 19245 1687 19261 1721
rect 19195 1677 19261 1687
rect 19295 1789 19349 1805
rect 19329 1755 19349 1789
rect 19295 1721 19349 1755
rect 19329 1687 19349 1721
rect 19295 1643 19349 1687
rect 17736 1596 17752 1630
rect 17786 1596 17802 1630
rect 18018 1609 18047 1643
rect 18081 1609 18139 1643
rect 18173 1609 18231 1643
rect 18265 1609 18294 1643
rect 19092 1609 19121 1643
rect 19155 1609 19213 1643
rect 19247 1609 19305 1643
rect 19339 1609 19368 1643
rect 17608 1546 17642 1562
rect 17608 1476 17642 1510
rect 17608 1424 17642 1440
rect 17704 1546 17738 1562
rect 17704 1476 17738 1510
rect 17704 1424 17738 1440
rect 17800 1546 17834 1562
rect 17800 1476 17834 1510
rect 17834 1440 18182 1464
rect 17800 1424 18182 1440
rect 17520 1356 17656 1390
rect 17690 1356 17706 1390
rect 17435 1286 17830 1306
rect 17435 1281 17697 1286
rect 17435 1272 17576 1281
rect 17560 1247 17576 1272
rect 17610 1252 17697 1281
rect 17731 1262 17830 1286
rect 18002 1264 18048 1266
rect 18002 1262 18006 1264
rect 17731 1252 18006 1262
rect 17610 1247 18006 1252
rect 17560 1230 18006 1247
rect 18040 1230 18048 1264
rect 17560 1228 18048 1230
rect 18002 1222 18048 1228
rect 16334 1107 16363 1141
rect 16397 1107 16455 1141
rect 16489 1107 16547 1141
rect 16581 1107 16610 1141
rect 15930 1055 16166 1066
rect 15572 1047 16166 1055
rect 15572 1022 15574 1047
rect 15486 979 15520 981
rect 15486 943 15520 945
rect 15486 858 15520 877
rect 15608 1022 16132 1047
rect 16218 1047 16294 1066
rect 16218 1026 16220 1047
rect 15574 979 15608 981
rect 15830 949 15846 983
rect 15880 949 15896 983
rect 16132 979 16166 981
rect 15574 943 15608 945
rect 16132 943 16166 945
rect 15574 858 15608 877
rect 15702 887 15736 906
rect 15702 819 15736 821
rect 15514 781 15530 815
rect 15564 781 15580 815
rect 15702 783 15736 785
rect 15202 703 15214 737
rect 15202 669 15248 703
rect 15202 635 15214 669
rect 14798 561 14827 595
rect 14861 561 14919 595
rect 14953 561 15011 595
rect 15045 561 15074 595
rect 15202 589 15248 635
rect 15282 737 15348 749
rect 15282 703 15298 737
rect 15332 703 15348 737
rect 15282 690 15348 703
rect 15702 698 15736 717
rect 15798 887 15832 906
rect 15798 819 15832 821
rect 15798 783 15832 785
rect 15798 698 15832 717
rect 15894 887 15928 906
rect 16132 858 16166 877
rect 16254 1026 16294 1047
rect 16402 1065 16444 1107
rect 16680 1105 16709 1139
rect 16743 1105 16801 1139
rect 16835 1105 16893 1139
rect 16927 1105 16956 1139
rect 17101 1133 17135 1140
rect 16402 1031 16410 1065
rect 16220 979 16254 981
rect 16220 943 16254 945
rect 16402 997 16444 1031
rect 16402 963 16410 997
rect 16402 929 16444 963
rect 16402 895 16410 929
rect 16402 879 16444 895
rect 16478 1065 16544 1073
rect 16478 1031 16494 1065
rect 16528 1031 16544 1065
rect 16478 997 16544 1031
rect 16478 963 16494 997
rect 16528 963 16544 997
rect 16478 929 16544 963
rect 16478 895 16494 929
rect 16528 895 16544 929
rect 16478 877 16544 895
rect 16713 1055 16749 1071
rect 16713 1021 16715 1055
rect 16713 987 16749 1021
rect 16713 953 16715 987
rect 16785 1055 16851 1105
rect 17026 1099 17055 1133
rect 17089 1099 17147 1133
rect 17181 1099 17239 1133
rect 17273 1099 17302 1133
rect 17402 1109 17418 1143
rect 17452 1109 17468 1143
rect 17626 1130 17740 1132
rect 16785 1021 16801 1055
rect 16835 1021 16851 1055
rect 16785 987 16851 1021
rect 16785 953 16801 987
rect 16835 953 16851 987
rect 16885 1055 16939 1071
rect 16885 1021 16887 1055
rect 16921 1021 16939 1055
rect 16885 974 16939 1021
rect 16713 919 16749 953
rect 16885 940 16887 974
rect 16921 940 16939 974
rect 16713 885 16848 919
rect 16885 890 16939 940
rect 16220 858 16254 877
rect 15894 819 15928 821
rect 16306 843 16450 844
rect 16306 829 16464 843
rect 15894 783 15928 785
rect 16160 816 16226 818
rect 16306 816 16414 829
rect 16160 815 16414 816
rect 16160 781 16176 815
rect 16210 802 16414 815
rect 16210 782 16346 802
rect 16398 795 16414 802
rect 16448 795 16464 829
rect 16210 781 16226 782
rect 16398 745 16444 761
rect 16498 757 16544 877
rect 16814 856 16848 885
rect 16701 827 16769 849
rect 16701 826 16717 827
rect 16701 792 16715 826
rect 16751 793 16769 827
rect 16749 792 16769 793
rect 16701 775 16769 792
rect 16814 840 16869 856
rect 16814 806 16835 840
rect 16814 790 16869 806
rect 16903 840 16939 890
rect 17094 1057 17136 1099
rect 17626 1091 17908 1130
rect 18048 1109 18064 1143
rect 18098 1109 18114 1143
rect 17626 1066 17665 1091
rect 17094 1023 17102 1057
rect 17094 989 17136 1023
rect 17094 955 17102 989
rect 17094 921 17136 955
rect 17094 887 17102 921
rect 17094 871 17136 887
rect 17170 1057 17236 1065
rect 17170 1023 17186 1057
rect 17220 1023 17236 1057
rect 17170 989 17236 1023
rect 17170 955 17186 989
rect 17220 955 17236 989
rect 17170 921 17236 955
rect 17170 887 17186 921
rect 17220 887 17236 921
rect 17170 869 17236 887
rect 16903 838 16944 840
rect 16903 804 16908 838
rect 16942 804 16944 838
rect 16903 802 16944 804
rect 17090 832 17156 835
rect 15928 717 16174 734
rect 15894 700 16174 717
rect 15894 698 15928 700
rect 15282 669 15624 690
rect 15282 635 15298 669
rect 15332 658 15624 669
rect 15332 655 15800 658
rect 15332 654 15750 655
rect 15332 635 15354 654
rect 15282 630 15354 635
rect 15282 623 15348 630
rect 15588 622 15750 654
rect 15734 621 15750 622
rect 15784 621 15800 655
rect 16126 612 16174 700
rect 15138 555 15167 589
rect 15201 555 15259 589
rect 15293 555 15351 589
rect 15385 555 15414 589
rect 15496 584 15542 594
rect 15496 550 15502 584
rect 15536 564 15542 584
rect 16126 578 16134 612
rect 16168 578 16174 612
rect 16398 711 16410 745
rect 16398 677 16444 711
rect 16398 643 16410 677
rect 16398 597 16444 643
rect 16478 745 16544 757
rect 16478 694 16494 745
rect 16528 694 16544 745
rect 16814 739 16848 790
rect 16478 677 16544 694
rect 16478 643 16494 677
rect 16528 643 16544 677
rect 16478 631 16544 643
rect 16715 705 16848 739
rect 16903 730 16939 802
rect 17090 798 17104 832
rect 17138 821 17156 832
rect 17090 787 17106 798
rect 17140 787 17156 821
rect 16715 684 16749 705
rect 16887 701 16939 730
rect 16715 629 16749 650
rect 16785 637 16801 671
rect 16835 637 16851 671
rect 15536 550 15546 564
rect 12140 420 12174 454
rect 12140 368 12174 384
rect 13532 444 13664 480
rect 13836 490 13870 506
rect 13932 490 13966 506
rect 13870 454 13871 455
rect 13532 396 13568 444
rect 13836 420 13871 454
rect 13870 418 13871 420
rect 13932 420 13966 454
rect 13716 396 13836 418
rect 13532 384 13836 396
rect 13870 384 13872 418
rect 13532 382 13872 384
rect 13532 360 13752 382
rect 13836 368 13870 382
rect 13932 368 13966 384
rect 14028 490 14062 506
rect 15496 480 15546 550
rect 15846 540 15862 574
rect 15896 540 15912 574
rect 16126 566 16174 578
rect 16334 563 16363 597
rect 16397 563 16455 597
rect 16489 563 16547 597
rect 16581 563 16610 597
rect 16785 595 16851 637
rect 16921 667 16939 701
rect 16887 629 16939 667
rect 17090 737 17136 753
rect 17190 749 17236 869
rect 17374 1047 17408 1066
rect 17460 1057 17665 1066
rect 17699 1089 17908 1091
rect 17699 1057 17784 1089
rect 17460 1055 17784 1057
rect 17818 1066 17908 1089
rect 18148 1066 18182 1424
rect 19092 1398 19126 1609
rect 19323 1306 19357 1609
rect 19408 1390 19442 2004
rect 19608 2002 19674 2004
rect 19925 2009 19941 2043
rect 19975 2009 19991 2043
rect 19925 1975 19991 2009
rect 19480 1943 19514 1962
rect 19480 1875 19514 1877
rect 19480 1839 19514 1841
rect 19480 1754 19514 1773
rect 19576 1943 19610 1962
rect 19576 1875 19610 1877
rect 19576 1839 19610 1841
rect 19576 1754 19610 1773
rect 19672 1943 19706 1962
rect 19925 1941 19941 1975
rect 19975 1959 19991 1975
rect 20097 2111 20163 2153
rect 20131 2077 20163 2111
rect 20097 2043 20163 2077
rect 20131 2009 20163 2043
rect 20097 1975 20163 2009
rect 19975 1941 20061 1959
rect 19925 1925 20061 1941
rect 20131 1941 20163 1975
rect 20097 1925 20163 1941
rect 20999 2111 21065 2116
rect 20999 2077 21015 2111
rect 21049 2077 21065 2111
rect 20999 2043 21065 2077
rect 20999 2009 21015 2043
rect 21049 2009 21065 2043
rect 20999 1975 21065 2009
rect 20999 1941 21015 1975
rect 21049 1959 21065 1975
rect 21171 2111 21237 2153
rect 21205 2077 21237 2111
rect 21404 2147 21686 2153
rect 21404 2113 21443 2147
rect 21477 2145 21686 2147
rect 21477 2113 21562 2145
rect 21404 2111 21562 2113
rect 21596 2111 21686 2145
rect 21404 2078 21686 2111
rect 21813 2111 21879 2116
rect 21171 2043 21237 2077
rect 21205 2009 21237 2043
rect 21813 2077 21829 2111
rect 21863 2077 21879 2111
rect 21813 2043 21879 2077
rect 21171 1975 21237 2009
rect 21049 1941 21135 1959
rect 20999 1925 21135 1941
rect 21205 1941 21237 1975
rect 21171 1925 21237 1941
rect 21296 2039 21562 2040
rect 21296 2005 21512 2039
rect 21546 2005 21562 2039
rect 21296 2004 21562 2005
rect 19672 1875 19706 1877
rect 19923 1882 19993 1891
rect 19923 1848 19939 1882
rect 19973 1875 19993 1882
rect 19923 1841 19943 1848
rect 19977 1841 19993 1875
rect 19672 1839 19706 1841
rect 20027 1805 20061 1925
rect 20095 1882 20165 1891
rect 20095 1875 20113 1882
rect 20095 1841 20111 1875
rect 20147 1848 20165 1882
rect 20145 1841 20165 1848
rect 20997 1884 21067 1891
rect 20997 1850 21015 1884
rect 21049 1875 21067 1884
rect 20997 1841 21017 1850
rect 21051 1841 21067 1875
rect 21101 1805 21135 1925
rect 21169 1880 21239 1891
rect 21169 1875 21188 1880
rect 21169 1841 21185 1875
rect 21222 1846 21239 1880
rect 21219 1841 21239 1846
rect 19672 1754 19706 1773
rect 19927 1789 19975 1805
rect 19927 1755 19941 1789
rect 19927 1721 19975 1755
rect 19512 1677 19528 1711
rect 19562 1677 19578 1711
rect 19927 1687 19941 1721
rect 19927 1643 19975 1687
rect 20009 1789 20075 1805
rect 20009 1755 20025 1789
rect 20059 1759 20075 1789
rect 20009 1725 20027 1755
rect 20061 1725 20075 1759
rect 20009 1721 20075 1725
rect 20009 1687 20025 1721
rect 20059 1687 20075 1721
rect 20009 1677 20075 1687
rect 20109 1789 20163 1805
rect 20143 1755 20163 1789
rect 20109 1721 20163 1755
rect 20143 1687 20163 1721
rect 20109 1643 20163 1687
rect 21001 1789 21049 1805
rect 21001 1755 21015 1789
rect 21001 1721 21049 1755
rect 21001 1687 21015 1721
rect 21001 1643 21049 1687
rect 21083 1789 21149 1805
rect 21083 1764 21099 1789
rect 21083 1730 21097 1764
rect 21133 1755 21149 1789
rect 21131 1730 21149 1755
rect 21083 1721 21149 1730
rect 21083 1687 21099 1721
rect 21133 1687 21149 1721
rect 21083 1677 21149 1687
rect 21183 1789 21237 1805
rect 21217 1755 21237 1789
rect 21183 1721 21237 1755
rect 21217 1687 21237 1721
rect 21183 1643 21237 1687
rect 19624 1596 19640 1630
rect 19674 1596 19690 1630
rect 19906 1609 19935 1643
rect 19969 1609 20027 1643
rect 20061 1609 20119 1643
rect 20153 1609 20182 1643
rect 20980 1609 21009 1643
rect 21043 1609 21101 1643
rect 21135 1609 21193 1643
rect 21227 1609 21256 1643
rect 19496 1546 19530 1562
rect 19496 1476 19530 1510
rect 19496 1424 19530 1440
rect 19592 1546 19626 1562
rect 19592 1476 19626 1510
rect 19592 1424 19626 1440
rect 19688 1546 19722 1562
rect 19688 1476 19722 1510
rect 19722 1440 20070 1464
rect 19688 1424 20070 1440
rect 19408 1356 19544 1390
rect 19578 1356 19594 1390
rect 19323 1286 19718 1306
rect 19323 1281 19585 1286
rect 19323 1272 19464 1281
rect 19448 1247 19464 1272
rect 19498 1252 19585 1281
rect 19619 1262 19718 1286
rect 19890 1264 19936 1266
rect 19890 1262 19894 1264
rect 19619 1252 19894 1262
rect 19498 1247 19894 1252
rect 19448 1230 19894 1247
rect 19928 1230 19936 1264
rect 19448 1228 19936 1230
rect 19890 1222 19936 1228
rect 18222 1107 18251 1141
rect 18285 1107 18343 1141
rect 18377 1107 18435 1141
rect 18469 1107 18498 1141
rect 17818 1055 18054 1066
rect 17460 1047 18054 1055
rect 17460 1022 17462 1047
rect 17374 979 17408 981
rect 17374 943 17408 945
rect 17374 858 17408 877
rect 17496 1022 18020 1047
rect 18106 1047 18182 1066
rect 18106 1026 18108 1047
rect 17462 979 17496 981
rect 17718 949 17734 983
rect 17768 949 17784 983
rect 18020 979 18054 981
rect 17462 943 17496 945
rect 18020 943 18054 945
rect 17462 858 17496 877
rect 17590 887 17624 906
rect 17590 819 17624 821
rect 17402 781 17418 815
rect 17452 781 17468 815
rect 17590 783 17624 785
rect 17090 703 17102 737
rect 17090 669 17136 703
rect 17090 635 17102 669
rect 16680 561 16709 595
rect 16743 561 16801 595
rect 16835 561 16893 595
rect 16927 561 16956 595
rect 17090 589 17136 635
rect 17170 737 17236 749
rect 17170 703 17186 737
rect 17220 703 17236 737
rect 17170 690 17236 703
rect 17590 698 17624 717
rect 17686 887 17720 906
rect 17686 819 17720 821
rect 17686 783 17720 785
rect 17686 698 17720 717
rect 17782 887 17816 906
rect 18020 858 18054 877
rect 18142 1026 18182 1047
rect 18290 1065 18332 1107
rect 18568 1105 18597 1139
rect 18631 1105 18689 1139
rect 18723 1105 18781 1139
rect 18815 1105 18844 1139
rect 18989 1133 19023 1140
rect 18290 1031 18298 1065
rect 18108 979 18142 981
rect 18108 943 18142 945
rect 18290 997 18332 1031
rect 18290 963 18298 997
rect 18290 929 18332 963
rect 18290 895 18298 929
rect 18290 879 18332 895
rect 18366 1065 18432 1073
rect 18366 1031 18382 1065
rect 18416 1031 18432 1065
rect 18366 997 18432 1031
rect 18366 963 18382 997
rect 18416 963 18432 997
rect 18366 929 18432 963
rect 18366 895 18382 929
rect 18416 895 18432 929
rect 18366 877 18432 895
rect 18601 1055 18637 1071
rect 18601 1021 18603 1055
rect 18601 987 18637 1021
rect 18601 953 18603 987
rect 18673 1055 18739 1105
rect 18914 1099 18943 1133
rect 18977 1099 19035 1133
rect 19069 1099 19127 1133
rect 19161 1099 19190 1133
rect 19290 1109 19306 1143
rect 19340 1109 19356 1143
rect 19514 1130 19628 1132
rect 18673 1021 18689 1055
rect 18723 1021 18739 1055
rect 18673 987 18739 1021
rect 18673 953 18689 987
rect 18723 953 18739 987
rect 18773 1055 18827 1071
rect 18773 1021 18775 1055
rect 18809 1021 18827 1055
rect 18773 974 18827 1021
rect 18601 919 18637 953
rect 18773 940 18775 974
rect 18809 940 18827 974
rect 18601 885 18736 919
rect 18773 890 18827 940
rect 18108 858 18142 877
rect 17782 819 17816 821
rect 18194 843 18338 844
rect 18194 829 18352 843
rect 17782 783 17816 785
rect 18048 816 18114 818
rect 18194 816 18302 829
rect 18048 815 18302 816
rect 18048 781 18064 815
rect 18098 802 18302 815
rect 18098 782 18234 802
rect 18286 795 18302 802
rect 18336 795 18352 829
rect 18098 781 18114 782
rect 18286 745 18332 761
rect 18386 757 18432 877
rect 18702 856 18736 885
rect 18589 827 18657 849
rect 18589 826 18605 827
rect 18589 792 18603 826
rect 18639 793 18657 827
rect 18637 792 18657 793
rect 18589 775 18657 792
rect 18702 840 18757 856
rect 18702 806 18723 840
rect 18702 790 18757 806
rect 18791 840 18827 890
rect 18982 1057 19024 1099
rect 19514 1091 19796 1130
rect 19936 1109 19952 1143
rect 19986 1109 20002 1143
rect 19514 1066 19553 1091
rect 18982 1023 18990 1057
rect 18982 989 19024 1023
rect 18982 955 18990 989
rect 18982 921 19024 955
rect 18982 887 18990 921
rect 18982 871 19024 887
rect 19058 1057 19124 1065
rect 19058 1023 19074 1057
rect 19108 1023 19124 1057
rect 19058 989 19124 1023
rect 19058 955 19074 989
rect 19108 955 19124 989
rect 19058 921 19124 955
rect 19058 887 19074 921
rect 19108 887 19124 921
rect 19058 869 19124 887
rect 18791 838 18832 840
rect 18791 804 18796 838
rect 18830 804 18832 838
rect 18791 802 18832 804
rect 18978 832 19044 835
rect 17816 717 18062 734
rect 17782 700 18062 717
rect 17782 698 17816 700
rect 17170 669 17512 690
rect 17170 635 17186 669
rect 17220 658 17512 669
rect 17220 655 17688 658
rect 17220 654 17638 655
rect 17220 635 17242 654
rect 17170 630 17242 635
rect 17170 623 17236 630
rect 17476 622 17638 654
rect 17622 621 17638 622
rect 17672 621 17688 655
rect 18014 612 18062 700
rect 17026 555 17055 589
rect 17089 555 17147 589
rect 17181 555 17239 589
rect 17273 555 17302 589
rect 17384 584 17430 594
rect 17384 550 17390 584
rect 17424 564 17430 584
rect 18014 578 18022 612
rect 18056 578 18062 612
rect 18286 711 18298 745
rect 18286 677 18332 711
rect 18286 643 18298 677
rect 18286 597 18332 643
rect 18366 745 18432 757
rect 18366 694 18382 745
rect 18416 694 18432 745
rect 18702 739 18736 790
rect 18366 677 18432 694
rect 18366 643 18382 677
rect 18416 643 18432 677
rect 18366 631 18432 643
rect 18603 705 18736 739
rect 18791 730 18827 802
rect 18978 798 18992 832
rect 19026 821 19044 832
rect 18978 787 18994 798
rect 19028 787 19044 821
rect 18603 684 18637 705
rect 18775 701 18827 730
rect 18603 629 18637 650
rect 18673 637 18689 671
rect 18723 637 18739 671
rect 17424 550 17434 564
rect 14028 420 14062 454
rect 14028 368 14062 384
rect 15414 444 15546 480
rect 15718 490 15752 506
rect 15814 490 15848 506
rect 15752 454 15753 455
rect 15414 396 15450 444
rect 15718 420 15753 454
rect 15752 418 15753 420
rect 15814 420 15848 454
rect 15598 396 15718 418
rect 15414 384 15718 396
rect 15752 384 15754 418
rect 15414 382 15754 384
rect 15414 360 15634 382
rect 15718 368 15752 382
rect 15814 368 15848 384
rect 15910 490 15944 506
rect 17384 480 17434 550
rect 17734 540 17750 574
rect 17784 540 17800 574
rect 18014 566 18062 578
rect 18222 563 18251 597
rect 18285 563 18343 597
rect 18377 563 18435 597
rect 18469 563 18498 597
rect 18673 595 18739 637
rect 18809 667 18827 701
rect 18775 629 18827 667
rect 18978 737 19024 753
rect 19078 749 19124 869
rect 19262 1047 19296 1066
rect 19348 1057 19553 1066
rect 19587 1089 19796 1091
rect 19587 1057 19672 1089
rect 19348 1055 19672 1057
rect 19706 1066 19796 1089
rect 20036 1066 20070 1424
rect 20980 1398 21014 1609
rect 21211 1306 21245 1609
rect 21296 1390 21330 2004
rect 21496 2002 21562 2004
rect 21813 2009 21829 2043
rect 21863 2009 21879 2043
rect 21813 1975 21879 2009
rect 21368 1943 21402 1962
rect 21368 1875 21402 1877
rect 21368 1839 21402 1841
rect 21368 1754 21402 1773
rect 21464 1943 21498 1962
rect 21464 1875 21498 1877
rect 21464 1839 21498 1841
rect 21464 1754 21498 1773
rect 21560 1943 21594 1962
rect 21813 1941 21829 1975
rect 21863 1959 21879 1975
rect 21985 2111 22051 2153
rect 22019 2077 22051 2111
rect 21985 2043 22051 2077
rect 22019 2009 22051 2043
rect 21985 1975 22051 2009
rect 21863 1941 21949 1959
rect 21813 1925 21949 1941
rect 22019 1941 22051 1975
rect 21985 1925 22051 1941
rect 22887 2111 22953 2116
rect 22887 2077 22903 2111
rect 22937 2077 22953 2111
rect 22887 2043 22953 2077
rect 22887 2009 22903 2043
rect 22937 2009 22953 2043
rect 22887 1975 22953 2009
rect 22887 1941 22903 1975
rect 22937 1959 22953 1975
rect 23059 2111 23125 2153
rect 23093 2077 23125 2111
rect 23292 2147 23574 2153
rect 23292 2113 23331 2147
rect 23365 2145 23574 2147
rect 23365 2113 23450 2145
rect 23292 2111 23450 2113
rect 23484 2111 23574 2145
rect 23292 2078 23574 2111
rect 23701 2111 23767 2116
rect 23059 2043 23125 2077
rect 23093 2009 23125 2043
rect 23701 2077 23717 2111
rect 23751 2077 23767 2111
rect 23701 2043 23767 2077
rect 23059 1975 23125 2009
rect 22937 1941 23023 1959
rect 22887 1925 23023 1941
rect 23093 1941 23125 1975
rect 23059 1925 23125 1941
rect 23184 2039 23450 2040
rect 23184 2005 23400 2039
rect 23434 2005 23450 2039
rect 23184 2004 23450 2005
rect 21560 1875 21594 1877
rect 21811 1882 21881 1891
rect 21811 1848 21827 1882
rect 21861 1875 21881 1882
rect 21811 1841 21831 1848
rect 21865 1841 21881 1875
rect 21560 1839 21594 1841
rect 21915 1805 21949 1925
rect 21983 1882 22053 1891
rect 21983 1875 22001 1882
rect 21983 1841 21999 1875
rect 22035 1848 22053 1882
rect 22033 1841 22053 1848
rect 22885 1884 22955 1891
rect 22885 1850 22903 1884
rect 22937 1875 22955 1884
rect 22885 1841 22905 1850
rect 22939 1841 22955 1875
rect 22989 1805 23023 1925
rect 23057 1880 23127 1891
rect 23057 1875 23076 1880
rect 23057 1841 23073 1875
rect 23110 1846 23127 1880
rect 23107 1841 23127 1846
rect 21560 1754 21594 1773
rect 21815 1789 21863 1805
rect 21815 1755 21829 1789
rect 21815 1721 21863 1755
rect 21400 1677 21416 1711
rect 21450 1677 21466 1711
rect 21815 1687 21829 1721
rect 21815 1643 21863 1687
rect 21897 1789 21963 1805
rect 21897 1755 21913 1789
rect 21947 1759 21963 1789
rect 21897 1725 21915 1755
rect 21949 1725 21963 1759
rect 21897 1721 21963 1725
rect 21897 1687 21913 1721
rect 21947 1687 21963 1721
rect 21897 1677 21963 1687
rect 21997 1789 22051 1805
rect 22031 1755 22051 1789
rect 21997 1721 22051 1755
rect 22031 1687 22051 1721
rect 21997 1643 22051 1687
rect 22889 1789 22937 1805
rect 22889 1755 22903 1789
rect 22889 1721 22937 1755
rect 22889 1687 22903 1721
rect 22889 1643 22937 1687
rect 22971 1789 23037 1805
rect 22971 1764 22987 1789
rect 22971 1730 22985 1764
rect 23021 1755 23037 1789
rect 23019 1730 23037 1755
rect 22971 1721 23037 1730
rect 22971 1687 22987 1721
rect 23021 1687 23037 1721
rect 22971 1677 23037 1687
rect 23071 1789 23125 1805
rect 23105 1755 23125 1789
rect 23071 1721 23125 1755
rect 23105 1687 23125 1721
rect 23071 1643 23125 1687
rect 21512 1596 21528 1630
rect 21562 1596 21578 1630
rect 21794 1609 21823 1643
rect 21857 1609 21915 1643
rect 21949 1609 22007 1643
rect 22041 1609 22070 1643
rect 22868 1609 22897 1643
rect 22931 1609 22989 1643
rect 23023 1609 23081 1643
rect 23115 1609 23144 1643
rect 21384 1546 21418 1562
rect 21384 1476 21418 1510
rect 21384 1424 21418 1440
rect 21480 1546 21514 1562
rect 21480 1476 21514 1510
rect 21480 1424 21514 1440
rect 21576 1546 21610 1562
rect 21576 1476 21610 1510
rect 21610 1440 21958 1464
rect 21576 1424 21958 1440
rect 21296 1356 21432 1390
rect 21466 1356 21482 1390
rect 21211 1286 21606 1306
rect 21211 1281 21473 1286
rect 21211 1272 21352 1281
rect 21336 1247 21352 1272
rect 21386 1252 21473 1281
rect 21507 1262 21606 1286
rect 21778 1264 21824 1266
rect 21778 1262 21782 1264
rect 21507 1252 21782 1262
rect 21386 1247 21782 1252
rect 21336 1230 21782 1247
rect 21816 1230 21824 1264
rect 21336 1228 21824 1230
rect 21778 1222 21824 1228
rect 20110 1107 20139 1141
rect 20173 1107 20231 1141
rect 20265 1107 20323 1141
rect 20357 1107 20386 1141
rect 19706 1055 19942 1066
rect 19348 1047 19942 1055
rect 19348 1022 19350 1047
rect 19262 979 19296 981
rect 19262 943 19296 945
rect 19262 858 19296 877
rect 19384 1022 19908 1047
rect 19994 1047 20070 1066
rect 19994 1026 19996 1047
rect 19350 979 19384 981
rect 19606 949 19622 983
rect 19656 949 19672 983
rect 19908 979 19942 981
rect 19350 943 19384 945
rect 19908 943 19942 945
rect 19350 858 19384 877
rect 19478 887 19512 906
rect 19478 819 19512 821
rect 19290 781 19306 815
rect 19340 781 19356 815
rect 19478 783 19512 785
rect 18978 703 18990 737
rect 18978 669 19024 703
rect 18978 635 18990 669
rect 18568 561 18597 595
rect 18631 561 18689 595
rect 18723 561 18781 595
rect 18815 561 18844 595
rect 18978 589 19024 635
rect 19058 737 19124 749
rect 19058 703 19074 737
rect 19108 703 19124 737
rect 19058 690 19124 703
rect 19478 698 19512 717
rect 19574 887 19608 906
rect 19574 819 19608 821
rect 19574 783 19608 785
rect 19574 698 19608 717
rect 19670 887 19704 906
rect 19908 858 19942 877
rect 20030 1026 20070 1047
rect 20178 1065 20220 1107
rect 20456 1105 20485 1139
rect 20519 1105 20577 1139
rect 20611 1105 20669 1139
rect 20703 1105 20732 1139
rect 20877 1133 20911 1140
rect 20178 1031 20186 1065
rect 19996 979 20030 981
rect 19996 943 20030 945
rect 20178 997 20220 1031
rect 20178 963 20186 997
rect 20178 929 20220 963
rect 20178 895 20186 929
rect 20178 879 20220 895
rect 20254 1065 20320 1073
rect 20254 1031 20270 1065
rect 20304 1031 20320 1065
rect 20254 997 20320 1031
rect 20254 963 20270 997
rect 20304 963 20320 997
rect 20254 929 20320 963
rect 20254 895 20270 929
rect 20304 895 20320 929
rect 20254 877 20320 895
rect 20489 1055 20525 1071
rect 20489 1021 20491 1055
rect 20489 987 20525 1021
rect 20489 953 20491 987
rect 20561 1055 20627 1105
rect 20802 1099 20831 1133
rect 20865 1099 20923 1133
rect 20957 1099 21015 1133
rect 21049 1099 21078 1133
rect 21178 1109 21194 1143
rect 21228 1109 21244 1143
rect 21402 1130 21516 1132
rect 20561 1021 20577 1055
rect 20611 1021 20627 1055
rect 20561 987 20627 1021
rect 20561 953 20577 987
rect 20611 953 20627 987
rect 20661 1055 20715 1071
rect 20661 1021 20663 1055
rect 20697 1021 20715 1055
rect 20661 974 20715 1021
rect 20489 919 20525 953
rect 20661 940 20663 974
rect 20697 940 20715 974
rect 20489 885 20624 919
rect 20661 890 20715 940
rect 19996 858 20030 877
rect 19670 819 19704 821
rect 20082 843 20226 844
rect 20082 829 20240 843
rect 19670 783 19704 785
rect 19936 816 20002 818
rect 20082 816 20190 829
rect 19936 815 20190 816
rect 19936 781 19952 815
rect 19986 802 20190 815
rect 19986 782 20122 802
rect 20174 795 20190 802
rect 20224 795 20240 829
rect 19986 781 20002 782
rect 20174 745 20220 761
rect 20274 757 20320 877
rect 20590 856 20624 885
rect 20477 827 20545 849
rect 20477 826 20493 827
rect 20477 792 20491 826
rect 20527 793 20545 827
rect 20525 792 20545 793
rect 20477 775 20545 792
rect 20590 840 20645 856
rect 20590 806 20611 840
rect 20590 790 20645 806
rect 20679 840 20715 890
rect 20870 1057 20912 1099
rect 21402 1091 21684 1130
rect 21824 1109 21840 1143
rect 21874 1109 21890 1143
rect 21402 1066 21441 1091
rect 20870 1023 20878 1057
rect 20870 989 20912 1023
rect 20870 955 20878 989
rect 20870 921 20912 955
rect 20870 887 20878 921
rect 20870 871 20912 887
rect 20946 1057 21012 1065
rect 20946 1023 20962 1057
rect 20996 1023 21012 1057
rect 20946 989 21012 1023
rect 20946 955 20962 989
rect 20996 955 21012 989
rect 20946 921 21012 955
rect 20946 887 20962 921
rect 20996 887 21012 921
rect 20946 869 21012 887
rect 20679 838 20720 840
rect 20679 804 20684 838
rect 20718 804 20720 838
rect 20679 802 20720 804
rect 20866 832 20932 835
rect 19704 717 19950 734
rect 19670 700 19950 717
rect 19670 698 19704 700
rect 19058 669 19400 690
rect 19058 635 19074 669
rect 19108 658 19400 669
rect 19108 655 19576 658
rect 19108 654 19526 655
rect 19108 635 19130 654
rect 19058 630 19130 635
rect 19058 623 19124 630
rect 19364 622 19526 654
rect 19510 621 19526 622
rect 19560 621 19576 655
rect 19902 612 19950 700
rect 18914 555 18943 589
rect 18977 555 19035 589
rect 19069 555 19127 589
rect 19161 555 19190 589
rect 19272 584 19318 594
rect 19272 550 19278 584
rect 19312 564 19318 584
rect 19902 578 19910 612
rect 19944 578 19950 612
rect 20174 711 20186 745
rect 20174 677 20220 711
rect 20174 643 20186 677
rect 20174 597 20220 643
rect 20254 745 20320 757
rect 20254 694 20270 745
rect 20304 694 20320 745
rect 20590 739 20624 790
rect 20254 677 20320 694
rect 20254 643 20270 677
rect 20304 643 20320 677
rect 20254 631 20320 643
rect 20491 705 20624 739
rect 20679 730 20715 802
rect 20866 798 20880 832
rect 20914 821 20932 832
rect 20866 787 20882 798
rect 20916 787 20932 821
rect 20491 684 20525 705
rect 20663 701 20715 730
rect 20491 629 20525 650
rect 20561 637 20577 671
rect 20611 637 20627 671
rect 19312 550 19322 564
rect 15910 420 15944 454
rect 15910 368 15944 384
rect 17302 444 17434 480
rect 17606 490 17640 506
rect 17702 490 17736 506
rect 17640 454 17641 455
rect 17302 396 17338 444
rect 17606 420 17641 454
rect 17640 418 17641 420
rect 17702 420 17736 454
rect 17486 396 17606 418
rect 17302 384 17606 396
rect 17640 384 17642 418
rect 17302 382 17642 384
rect 17302 360 17522 382
rect 17606 368 17640 382
rect 17702 368 17736 384
rect 17798 490 17832 506
rect 19272 480 19322 550
rect 19622 540 19638 574
rect 19672 540 19688 574
rect 19902 566 19950 578
rect 20110 563 20139 597
rect 20173 563 20231 597
rect 20265 563 20323 597
rect 20357 563 20386 597
rect 20561 595 20627 637
rect 20697 667 20715 701
rect 20663 629 20715 667
rect 20866 737 20912 753
rect 20966 749 21012 869
rect 21150 1047 21184 1066
rect 21236 1057 21441 1066
rect 21475 1089 21684 1091
rect 21475 1057 21560 1089
rect 21236 1055 21560 1057
rect 21594 1066 21684 1089
rect 21924 1066 21958 1424
rect 22868 1398 22902 1609
rect 23099 1306 23133 1609
rect 23184 1390 23218 2004
rect 23384 2002 23450 2004
rect 23701 2009 23717 2043
rect 23751 2009 23767 2043
rect 23701 1975 23767 2009
rect 23256 1943 23290 1962
rect 23256 1875 23290 1877
rect 23256 1839 23290 1841
rect 23256 1754 23290 1773
rect 23352 1943 23386 1962
rect 23352 1875 23386 1877
rect 23352 1839 23386 1841
rect 23352 1754 23386 1773
rect 23448 1943 23482 1962
rect 23701 1941 23717 1975
rect 23751 1959 23767 1975
rect 23873 2111 23939 2153
rect 23907 2077 23939 2111
rect 23873 2043 23939 2077
rect 23907 2009 23939 2043
rect 23873 1975 23939 2009
rect 23751 1941 23837 1959
rect 23701 1925 23837 1941
rect 23907 1941 23939 1975
rect 23873 1925 23939 1941
rect 24775 2111 24841 2116
rect 24775 2077 24791 2111
rect 24825 2077 24841 2111
rect 24775 2043 24841 2077
rect 24775 2009 24791 2043
rect 24825 2009 24841 2043
rect 24775 1975 24841 2009
rect 24775 1941 24791 1975
rect 24825 1959 24841 1975
rect 24947 2111 25013 2153
rect 24981 2077 25013 2111
rect 25180 2147 25462 2153
rect 25180 2113 25219 2147
rect 25253 2145 25462 2147
rect 25253 2113 25338 2145
rect 25180 2111 25338 2113
rect 25372 2111 25462 2145
rect 25180 2078 25462 2111
rect 25589 2111 25655 2116
rect 24947 2043 25013 2077
rect 24981 2009 25013 2043
rect 25589 2077 25605 2111
rect 25639 2077 25655 2111
rect 25589 2043 25655 2077
rect 24947 1975 25013 2009
rect 24825 1941 24911 1959
rect 24775 1925 24911 1941
rect 24981 1941 25013 1975
rect 24947 1925 25013 1941
rect 25072 2039 25338 2040
rect 25072 2005 25288 2039
rect 25322 2005 25338 2039
rect 25072 2004 25338 2005
rect 23448 1875 23482 1877
rect 23699 1882 23769 1891
rect 23699 1848 23715 1882
rect 23749 1875 23769 1882
rect 23699 1841 23719 1848
rect 23753 1841 23769 1875
rect 23448 1839 23482 1841
rect 23803 1805 23837 1925
rect 23871 1882 23941 1891
rect 23871 1875 23889 1882
rect 23871 1841 23887 1875
rect 23923 1848 23941 1882
rect 23921 1841 23941 1848
rect 24773 1884 24843 1891
rect 24773 1850 24791 1884
rect 24825 1875 24843 1884
rect 24773 1841 24793 1850
rect 24827 1841 24843 1875
rect 24877 1805 24911 1925
rect 24945 1880 25015 1891
rect 24945 1875 24964 1880
rect 24945 1841 24961 1875
rect 24998 1846 25015 1880
rect 24995 1841 25015 1846
rect 23448 1754 23482 1773
rect 23703 1789 23751 1805
rect 23703 1755 23717 1789
rect 23703 1721 23751 1755
rect 23288 1677 23304 1711
rect 23338 1677 23354 1711
rect 23703 1687 23717 1721
rect 23703 1643 23751 1687
rect 23785 1789 23851 1805
rect 23785 1755 23801 1789
rect 23835 1759 23851 1789
rect 23785 1725 23803 1755
rect 23837 1725 23851 1759
rect 23785 1721 23851 1725
rect 23785 1687 23801 1721
rect 23835 1687 23851 1721
rect 23785 1677 23851 1687
rect 23885 1789 23939 1805
rect 23919 1755 23939 1789
rect 23885 1721 23939 1755
rect 23919 1687 23939 1721
rect 23885 1643 23939 1687
rect 24777 1789 24825 1805
rect 24777 1755 24791 1789
rect 24777 1721 24825 1755
rect 24777 1687 24791 1721
rect 24777 1643 24825 1687
rect 24859 1789 24925 1805
rect 24859 1764 24875 1789
rect 24859 1730 24873 1764
rect 24909 1755 24925 1789
rect 24907 1730 24925 1755
rect 24859 1721 24925 1730
rect 24859 1687 24875 1721
rect 24909 1687 24925 1721
rect 24859 1677 24925 1687
rect 24959 1789 25013 1805
rect 24993 1755 25013 1789
rect 24959 1721 25013 1755
rect 24993 1687 25013 1721
rect 24959 1643 25013 1687
rect 23400 1596 23416 1630
rect 23450 1596 23466 1630
rect 23682 1609 23711 1643
rect 23745 1609 23803 1643
rect 23837 1609 23895 1643
rect 23929 1609 23958 1643
rect 24756 1609 24785 1643
rect 24819 1609 24877 1643
rect 24911 1609 24969 1643
rect 25003 1609 25032 1643
rect 23272 1546 23306 1562
rect 23272 1476 23306 1510
rect 23272 1424 23306 1440
rect 23368 1546 23402 1562
rect 23368 1476 23402 1510
rect 23368 1424 23402 1440
rect 23464 1546 23498 1562
rect 23464 1476 23498 1510
rect 23498 1440 23846 1464
rect 23464 1424 23846 1440
rect 23184 1356 23320 1390
rect 23354 1356 23370 1390
rect 23099 1286 23494 1306
rect 23099 1281 23361 1286
rect 23099 1272 23240 1281
rect 23224 1247 23240 1272
rect 23274 1252 23361 1281
rect 23395 1262 23494 1286
rect 23666 1264 23712 1266
rect 23666 1262 23670 1264
rect 23395 1252 23670 1262
rect 23274 1247 23670 1252
rect 23224 1230 23670 1247
rect 23704 1230 23712 1264
rect 23224 1228 23712 1230
rect 23666 1222 23712 1228
rect 21998 1107 22027 1141
rect 22061 1107 22119 1141
rect 22153 1107 22211 1141
rect 22245 1107 22274 1141
rect 21594 1055 21830 1066
rect 21236 1047 21830 1055
rect 21236 1022 21238 1047
rect 21150 979 21184 981
rect 21150 943 21184 945
rect 21150 858 21184 877
rect 21272 1022 21796 1047
rect 21882 1047 21958 1066
rect 21882 1026 21884 1047
rect 21238 979 21272 981
rect 21494 949 21510 983
rect 21544 949 21560 983
rect 21796 979 21830 981
rect 21238 943 21272 945
rect 21796 943 21830 945
rect 21238 858 21272 877
rect 21366 887 21400 906
rect 21366 819 21400 821
rect 21178 781 21194 815
rect 21228 781 21244 815
rect 21366 783 21400 785
rect 20866 703 20878 737
rect 20866 669 20912 703
rect 20866 635 20878 669
rect 20456 561 20485 595
rect 20519 561 20577 595
rect 20611 561 20669 595
rect 20703 561 20732 595
rect 20866 589 20912 635
rect 20946 737 21012 749
rect 20946 703 20962 737
rect 20996 703 21012 737
rect 20946 690 21012 703
rect 21366 698 21400 717
rect 21462 887 21496 906
rect 21462 819 21496 821
rect 21462 783 21496 785
rect 21462 698 21496 717
rect 21558 887 21592 906
rect 21796 858 21830 877
rect 21918 1026 21958 1047
rect 22066 1065 22108 1107
rect 22344 1105 22373 1139
rect 22407 1105 22465 1139
rect 22499 1105 22557 1139
rect 22591 1105 22620 1139
rect 22765 1133 22799 1140
rect 22066 1031 22074 1065
rect 21884 979 21918 981
rect 21884 943 21918 945
rect 22066 997 22108 1031
rect 22066 963 22074 997
rect 22066 929 22108 963
rect 22066 895 22074 929
rect 22066 879 22108 895
rect 22142 1065 22208 1073
rect 22142 1031 22158 1065
rect 22192 1031 22208 1065
rect 22142 997 22208 1031
rect 22142 963 22158 997
rect 22192 963 22208 997
rect 22142 929 22208 963
rect 22142 895 22158 929
rect 22192 895 22208 929
rect 22142 877 22208 895
rect 22377 1055 22413 1071
rect 22377 1021 22379 1055
rect 22377 987 22413 1021
rect 22377 953 22379 987
rect 22449 1055 22515 1105
rect 22690 1099 22719 1133
rect 22753 1099 22811 1133
rect 22845 1099 22903 1133
rect 22937 1099 22966 1133
rect 23066 1109 23082 1143
rect 23116 1109 23132 1143
rect 23290 1130 23404 1132
rect 22449 1021 22465 1055
rect 22499 1021 22515 1055
rect 22449 987 22515 1021
rect 22449 953 22465 987
rect 22499 953 22515 987
rect 22549 1055 22603 1071
rect 22549 1021 22551 1055
rect 22585 1021 22603 1055
rect 22549 974 22603 1021
rect 22377 919 22413 953
rect 22549 940 22551 974
rect 22585 940 22603 974
rect 22377 885 22512 919
rect 22549 890 22603 940
rect 21884 858 21918 877
rect 21558 819 21592 821
rect 21970 843 22114 844
rect 21970 829 22128 843
rect 21558 783 21592 785
rect 21824 816 21890 818
rect 21970 816 22078 829
rect 21824 815 22078 816
rect 21824 781 21840 815
rect 21874 802 22078 815
rect 21874 782 22010 802
rect 22062 795 22078 802
rect 22112 795 22128 829
rect 21874 781 21890 782
rect 22062 745 22108 761
rect 22162 757 22208 877
rect 22478 856 22512 885
rect 22365 827 22433 849
rect 22365 826 22381 827
rect 22365 792 22379 826
rect 22415 793 22433 827
rect 22413 792 22433 793
rect 22365 775 22433 792
rect 22478 840 22533 856
rect 22478 806 22499 840
rect 22478 790 22533 806
rect 22567 840 22603 890
rect 22758 1057 22800 1099
rect 23290 1091 23572 1130
rect 23712 1109 23728 1143
rect 23762 1109 23778 1143
rect 23290 1066 23329 1091
rect 22758 1023 22766 1057
rect 22758 989 22800 1023
rect 22758 955 22766 989
rect 22758 921 22800 955
rect 22758 887 22766 921
rect 22758 871 22800 887
rect 22834 1057 22900 1065
rect 22834 1023 22850 1057
rect 22884 1023 22900 1057
rect 22834 989 22900 1023
rect 22834 955 22850 989
rect 22884 955 22900 989
rect 22834 921 22900 955
rect 22834 887 22850 921
rect 22884 887 22900 921
rect 22834 869 22900 887
rect 22567 838 22608 840
rect 22567 804 22572 838
rect 22606 804 22608 838
rect 22567 802 22608 804
rect 22754 832 22820 835
rect 21592 717 21838 734
rect 21558 700 21838 717
rect 21558 698 21592 700
rect 20946 669 21288 690
rect 20946 635 20962 669
rect 20996 658 21288 669
rect 20996 655 21464 658
rect 20996 654 21414 655
rect 20996 635 21018 654
rect 20946 630 21018 635
rect 20946 623 21012 630
rect 21252 622 21414 654
rect 21398 621 21414 622
rect 21448 621 21464 655
rect 21790 612 21838 700
rect 20802 555 20831 589
rect 20865 555 20923 589
rect 20957 555 21015 589
rect 21049 555 21078 589
rect 21160 584 21206 594
rect 21160 550 21166 584
rect 21200 564 21206 584
rect 21790 578 21798 612
rect 21832 578 21838 612
rect 22062 711 22074 745
rect 22062 677 22108 711
rect 22062 643 22074 677
rect 22062 597 22108 643
rect 22142 745 22208 757
rect 22142 694 22158 745
rect 22192 694 22208 745
rect 22478 739 22512 790
rect 22142 677 22208 694
rect 22142 643 22158 677
rect 22192 643 22208 677
rect 22142 631 22208 643
rect 22379 705 22512 739
rect 22567 730 22603 802
rect 22754 798 22768 832
rect 22802 821 22820 832
rect 22754 787 22770 798
rect 22804 787 22820 821
rect 22379 684 22413 705
rect 22551 701 22603 730
rect 22379 629 22413 650
rect 22449 637 22465 671
rect 22499 637 22515 671
rect 21200 550 21210 564
rect 17798 420 17832 454
rect 17798 368 17832 384
rect 19190 444 19322 480
rect 19494 490 19528 506
rect 19590 490 19624 506
rect 19528 454 19529 455
rect 19190 396 19226 444
rect 19494 420 19529 454
rect 19528 418 19529 420
rect 19590 420 19624 454
rect 19374 396 19494 418
rect 19190 384 19494 396
rect 19528 384 19530 418
rect 19190 382 19530 384
rect 19190 360 19410 382
rect 19494 368 19528 382
rect 19590 368 19624 384
rect 19686 490 19720 506
rect 21160 480 21210 550
rect 21510 540 21526 574
rect 21560 540 21576 574
rect 21790 566 21838 578
rect 21998 563 22027 597
rect 22061 563 22119 597
rect 22153 563 22211 597
rect 22245 563 22274 597
rect 22449 595 22515 637
rect 22585 667 22603 701
rect 22551 629 22603 667
rect 22754 737 22800 753
rect 22854 749 22900 869
rect 23038 1047 23072 1066
rect 23124 1057 23329 1066
rect 23363 1089 23572 1091
rect 23363 1057 23448 1089
rect 23124 1055 23448 1057
rect 23482 1066 23572 1089
rect 23812 1066 23846 1424
rect 24756 1398 24790 1609
rect 24987 1306 25021 1609
rect 25072 1390 25106 2004
rect 25272 2002 25338 2004
rect 25589 2009 25605 2043
rect 25639 2009 25655 2043
rect 25589 1975 25655 2009
rect 25144 1943 25178 1962
rect 25144 1875 25178 1877
rect 25144 1839 25178 1841
rect 25144 1754 25178 1773
rect 25240 1943 25274 1962
rect 25240 1875 25274 1877
rect 25240 1839 25274 1841
rect 25240 1754 25274 1773
rect 25336 1943 25370 1962
rect 25589 1941 25605 1975
rect 25639 1959 25655 1975
rect 25761 2111 25827 2153
rect 25795 2077 25827 2111
rect 25761 2043 25827 2077
rect 25795 2009 25827 2043
rect 25761 1975 25827 2009
rect 25639 1941 25725 1959
rect 25589 1925 25725 1941
rect 25795 1941 25827 1975
rect 25761 1925 25827 1941
rect 26663 2111 26729 2116
rect 26663 2077 26679 2111
rect 26713 2077 26729 2111
rect 26663 2043 26729 2077
rect 26663 2009 26679 2043
rect 26713 2009 26729 2043
rect 26663 1975 26729 2009
rect 26663 1941 26679 1975
rect 26713 1959 26729 1975
rect 26835 2111 26901 2153
rect 26869 2077 26901 2111
rect 27068 2147 27350 2153
rect 27068 2113 27107 2147
rect 27141 2145 27350 2147
rect 27141 2113 27226 2145
rect 27068 2111 27226 2113
rect 27260 2111 27350 2145
rect 27068 2078 27350 2111
rect 27477 2111 27543 2116
rect 26835 2043 26901 2077
rect 26869 2009 26901 2043
rect 27477 2077 27493 2111
rect 27527 2077 27543 2111
rect 27477 2043 27543 2077
rect 26835 1975 26901 2009
rect 26713 1941 26799 1959
rect 26663 1925 26799 1941
rect 26869 1941 26901 1975
rect 26835 1925 26901 1941
rect 26960 2039 27226 2040
rect 26960 2005 27176 2039
rect 27210 2005 27226 2039
rect 26960 2004 27226 2005
rect 25336 1875 25370 1877
rect 25587 1882 25657 1891
rect 25587 1848 25603 1882
rect 25637 1875 25657 1882
rect 25587 1841 25607 1848
rect 25641 1841 25657 1875
rect 25336 1839 25370 1841
rect 25691 1805 25725 1925
rect 25759 1882 25829 1891
rect 25759 1875 25777 1882
rect 25759 1841 25775 1875
rect 25811 1848 25829 1882
rect 25809 1841 25829 1848
rect 26661 1884 26731 1891
rect 26661 1850 26679 1884
rect 26713 1875 26731 1884
rect 26661 1841 26681 1850
rect 26715 1841 26731 1875
rect 26765 1805 26799 1925
rect 26833 1880 26903 1891
rect 26833 1875 26852 1880
rect 26833 1841 26849 1875
rect 26886 1846 26903 1880
rect 26883 1841 26903 1846
rect 25336 1754 25370 1773
rect 25591 1789 25639 1805
rect 25591 1755 25605 1789
rect 25591 1721 25639 1755
rect 25176 1677 25192 1711
rect 25226 1677 25242 1711
rect 25591 1687 25605 1721
rect 25591 1643 25639 1687
rect 25673 1789 25739 1805
rect 25673 1755 25689 1789
rect 25723 1759 25739 1789
rect 25673 1725 25691 1755
rect 25725 1725 25739 1759
rect 25673 1721 25739 1725
rect 25673 1687 25689 1721
rect 25723 1687 25739 1721
rect 25673 1677 25739 1687
rect 25773 1789 25827 1805
rect 25807 1755 25827 1789
rect 25773 1721 25827 1755
rect 25807 1687 25827 1721
rect 25773 1643 25827 1687
rect 26665 1789 26713 1805
rect 26665 1755 26679 1789
rect 26665 1721 26713 1755
rect 26665 1687 26679 1721
rect 26665 1643 26713 1687
rect 26747 1789 26813 1805
rect 26747 1764 26763 1789
rect 26747 1730 26761 1764
rect 26797 1755 26813 1789
rect 26795 1730 26813 1755
rect 26747 1721 26813 1730
rect 26747 1687 26763 1721
rect 26797 1687 26813 1721
rect 26747 1677 26813 1687
rect 26847 1789 26901 1805
rect 26881 1755 26901 1789
rect 26847 1721 26901 1755
rect 26881 1687 26901 1721
rect 26847 1643 26901 1687
rect 25288 1596 25304 1630
rect 25338 1596 25354 1630
rect 25570 1609 25599 1643
rect 25633 1609 25691 1643
rect 25725 1609 25783 1643
rect 25817 1609 25846 1643
rect 26644 1609 26673 1643
rect 26707 1609 26765 1643
rect 26799 1609 26857 1643
rect 26891 1609 26920 1643
rect 25160 1546 25194 1562
rect 25160 1476 25194 1510
rect 25160 1424 25194 1440
rect 25256 1546 25290 1562
rect 25256 1476 25290 1510
rect 25256 1424 25290 1440
rect 25352 1546 25386 1562
rect 25352 1476 25386 1510
rect 25386 1440 25734 1464
rect 25352 1424 25734 1440
rect 25072 1356 25208 1390
rect 25242 1356 25258 1390
rect 24987 1286 25382 1306
rect 24987 1281 25249 1286
rect 24987 1272 25128 1281
rect 25112 1247 25128 1272
rect 25162 1252 25249 1281
rect 25283 1262 25382 1286
rect 25554 1264 25600 1266
rect 25554 1262 25558 1264
rect 25283 1252 25558 1262
rect 25162 1247 25558 1252
rect 25112 1230 25558 1247
rect 25592 1230 25600 1264
rect 25112 1228 25600 1230
rect 25554 1222 25600 1228
rect 23886 1107 23915 1141
rect 23949 1107 24007 1141
rect 24041 1107 24099 1141
rect 24133 1107 24162 1141
rect 23482 1055 23718 1066
rect 23124 1047 23718 1055
rect 23124 1022 23126 1047
rect 23038 979 23072 981
rect 23038 943 23072 945
rect 23038 858 23072 877
rect 23160 1022 23684 1047
rect 23770 1047 23846 1066
rect 23770 1026 23772 1047
rect 23126 979 23160 981
rect 23382 949 23398 983
rect 23432 949 23448 983
rect 23684 979 23718 981
rect 23126 943 23160 945
rect 23684 943 23718 945
rect 23126 858 23160 877
rect 23254 887 23288 906
rect 23254 819 23288 821
rect 23066 781 23082 815
rect 23116 781 23132 815
rect 23254 783 23288 785
rect 22754 703 22766 737
rect 22754 669 22800 703
rect 22754 635 22766 669
rect 22344 561 22373 595
rect 22407 561 22465 595
rect 22499 561 22557 595
rect 22591 561 22620 595
rect 22754 589 22800 635
rect 22834 737 22900 749
rect 22834 703 22850 737
rect 22884 703 22900 737
rect 22834 690 22900 703
rect 23254 698 23288 717
rect 23350 887 23384 906
rect 23350 819 23384 821
rect 23350 783 23384 785
rect 23350 698 23384 717
rect 23446 887 23480 906
rect 23684 858 23718 877
rect 23806 1026 23846 1047
rect 23954 1065 23996 1107
rect 24232 1105 24261 1139
rect 24295 1105 24353 1139
rect 24387 1105 24445 1139
rect 24479 1105 24508 1139
rect 24653 1133 24687 1140
rect 23954 1031 23962 1065
rect 23772 979 23806 981
rect 23772 943 23806 945
rect 23954 997 23996 1031
rect 23954 963 23962 997
rect 23954 929 23996 963
rect 23954 895 23962 929
rect 23954 879 23996 895
rect 24030 1065 24096 1073
rect 24030 1031 24046 1065
rect 24080 1031 24096 1065
rect 24030 997 24096 1031
rect 24030 963 24046 997
rect 24080 963 24096 997
rect 24030 929 24096 963
rect 24030 895 24046 929
rect 24080 895 24096 929
rect 24030 877 24096 895
rect 24265 1055 24301 1071
rect 24265 1021 24267 1055
rect 24265 987 24301 1021
rect 24265 953 24267 987
rect 24337 1055 24403 1105
rect 24578 1099 24607 1133
rect 24641 1099 24699 1133
rect 24733 1099 24791 1133
rect 24825 1099 24854 1133
rect 24954 1109 24970 1143
rect 25004 1109 25020 1143
rect 25178 1130 25292 1132
rect 24337 1021 24353 1055
rect 24387 1021 24403 1055
rect 24337 987 24403 1021
rect 24337 953 24353 987
rect 24387 953 24403 987
rect 24437 1055 24491 1071
rect 24437 1021 24439 1055
rect 24473 1021 24491 1055
rect 24437 974 24491 1021
rect 24265 919 24301 953
rect 24437 940 24439 974
rect 24473 940 24491 974
rect 24265 885 24400 919
rect 24437 890 24491 940
rect 23772 858 23806 877
rect 23446 819 23480 821
rect 23858 843 24002 844
rect 23858 829 24016 843
rect 23446 783 23480 785
rect 23712 816 23778 818
rect 23858 816 23966 829
rect 23712 815 23966 816
rect 23712 781 23728 815
rect 23762 802 23966 815
rect 23762 782 23898 802
rect 23950 795 23966 802
rect 24000 795 24016 829
rect 23762 781 23778 782
rect 23950 745 23996 761
rect 24050 757 24096 877
rect 24366 856 24400 885
rect 24253 827 24321 849
rect 24253 826 24269 827
rect 24253 792 24267 826
rect 24303 793 24321 827
rect 24301 792 24321 793
rect 24253 775 24321 792
rect 24366 840 24421 856
rect 24366 806 24387 840
rect 24366 790 24421 806
rect 24455 840 24491 890
rect 24646 1057 24688 1099
rect 25178 1091 25460 1130
rect 25600 1109 25616 1143
rect 25650 1109 25666 1143
rect 25178 1066 25217 1091
rect 24646 1023 24654 1057
rect 24646 989 24688 1023
rect 24646 955 24654 989
rect 24646 921 24688 955
rect 24646 887 24654 921
rect 24646 871 24688 887
rect 24722 1057 24788 1065
rect 24722 1023 24738 1057
rect 24772 1023 24788 1057
rect 24722 989 24788 1023
rect 24722 955 24738 989
rect 24772 955 24788 989
rect 24722 921 24788 955
rect 24722 887 24738 921
rect 24772 887 24788 921
rect 24722 869 24788 887
rect 24455 838 24496 840
rect 24455 804 24460 838
rect 24494 804 24496 838
rect 24455 802 24496 804
rect 24642 832 24708 835
rect 23480 717 23726 734
rect 23446 700 23726 717
rect 23446 698 23480 700
rect 22834 669 23176 690
rect 22834 635 22850 669
rect 22884 658 23176 669
rect 22884 655 23352 658
rect 22884 654 23302 655
rect 22884 635 22906 654
rect 22834 630 22906 635
rect 22834 623 22900 630
rect 23140 622 23302 654
rect 23286 621 23302 622
rect 23336 621 23352 655
rect 23678 612 23726 700
rect 22690 555 22719 589
rect 22753 555 22811 589
rect 22845 555 22903 589
rect 22937 555 22966 589
rect 23048 584 23094 594
rect 23048 550 23054 584
rect 23088 564 23094 584
rect 23678 578 23686 612
rect 23720 578 23726 612
rect 23950 711 23962 745
rect 23950 677 23996 711
rect 23950 643 23962 677
rect 23950 597 23996 643
rect 24030 745 24096 757
rect 24030 694 24046 745
rect 24080 694 24096 745
rect 24366 739 24400 790
rect 24030 677 24096 694
rect 24030 643 24046 677
rect 24080 643 24096 677
rect 24030 631 24096 643
rect 24267 705 24400 739
rect 24455 730 24491 802
rect 24642 798 24656 832
rect 24690 821 24708 832
rect 24642 787 24658 798
rect 24692 787 24708 821
rect 24267 684 24301 705
rect 24439 701 24491 730
rect 24267 629 24301 650
rect 24337 637 24353 671
rect 24387 637 24403 671
rect 23088 550 23098 564
rect 19686 420 19720 454
rect 19686 368 19720 384
rect 21078 444 21210 480
rect 21382 490 21416 506
rect 21478 490 21512 506
rect 21416 454 21417 455
rect 21078 396 21114 444
rect 21382 420 21417 454
rect 21416 418 21417 420
rect 21478 420 21512 454
rect 21262 396 21382 418
rect 21078 384 21382 396
rect 21416 384 21418 418
rect 21078 382 21418 384
rect 21078 360 21298 382
rect 21382 368 21416 382
rect 21478 368 21512 384
rect 21574 490 21608 506
rect 23048 480 23098 550
rect 23398 540 23414 574
rect 23448 540 23464 574
rect 23678 566 23726 578
rect 23886 563 23915 597
rect 23949 563 24007 597
rect 24041 563 24099 597
rect 24133 563 24162 597
rect 24337 595 24403 637
rect 24473 667 24491 701
rect 24439 629 24491 667
rect 24642 737 24688 753
rect 24742 749 24788 869
rect 24926 1047 24960 1066
rect 25012 1057 25217 1066
rect 25251 1089 25460 1091
rect 25251 1057 25336 1089
rect 25012 1055 25336 1057
rect 25370 1066 25460 1089
rect 25700 1066 25734 1424
rect 26644 1398 26678 1609
rect 26875 1306 26909 1609
rect 26960 1390 26994 2004
rect 27160 2002 27226 2004
rect 27477 2009 27493 2043
rect 27527 2009 27543 2043
rect 27477 1975 27543 2009
rect 27032 1943 27066 1962
rect 27032 1875 27066 1877
rect 27032 1839 27066 1841
rect 27032 1754 27066 1773
rect 27128 1943 27162 1962
rect 27128 1875 27162 1877
rect 27128 1839 27162 1841
rect 27128 1754 27162 1773
rect 27224 1943 27258 1962
rect 27477 1941 27493 1975
rect 27527 1959 27543 1975
rect 27649 2111 27715 2153
rect 27683 2077 27715 2111
rect 27649 2043 27715 2077
rect 27683 2009 27715 2043
rect 27649 1975 27715 2009
rect 27527 1941 27613 1959
rect 27477 1925 27613 1941
rect 27683 1941 27715 1975
rect 27649 1925 27715 1941
rect 28551 2111 28617 2116
rect 28551 2077 28567 2111
rect 28601 2077 28617 2111
rect 28551 2043 28617 2077
rect 28551 2009 28567 2043
rect 28601 2009 28617 2043
rect 28551 1975 28617 2009
rect 28551 1941 28567 1975
rect 28601 1959 28617 1975
rect 28723 2111 28789 2153
rect 28757 2077 28789 2111
rect 28956 2147 29238 2153
rect 28956 2113 28995 2147
rect 29029 2145 29238 2147
rect 29029 2113 29114 2145
rect 28956 2111 29114 2113
rect 29148 2111 29238 2145
rect 28956 2078 29238 2111
rect 29365 2111 29431 2116
rect 28723 2043 28789 2077
rect 28757 2009 28789 2043
rect 29365 2077 29381 2111
rect 29415 2077 29431 2111
rect 29365 2043 29431 2077
rect 28723 1975 28789 2009
rect 28601 1941 28687 1959
rect 28551 1925 28687 1941
rect 28757 1941 28789 1975
rect 28723 1925 28789 1941
rect 28848 2039 29114 2040
rect 28848 2005 29064 2039
rect 29098 2005 29114 2039
rect 28848 2004 29114 2005
rect 27224 1875 27258 1877
rect 27475 1882 27545 1891
rect 27475 1848 27491 1882
rect 27525 1875 27545 1882
rect 27475 1841 27495 1848
rect 27529 1841 27545 1875
rect 27224 1839 27258 1841
rect 27579 1805 27613 1925
rect 27647 1882 27717 1891
rect 27647 1875 27665 1882
rect 27647 1841 27663 1875
rect 27699 1848 27717 1882
rect 27697 1841 27717 1848
rect 28549 1884 28619 1891
rect 28549 1850 28567 1884
rect 28601 1875 28619 1884
rect 28549 1841 28569 1850
rect 28603 1841 28619 1875
rect 28653 1805 28687 1925
rect 28721 1880 28791 1891
rect 28721 1875 28740 1880
rect 28721 1841 28737 1875
rect 28774 1846 28791 1880
rect 28771 1841 28791 1846
rect 27224 1754 27258 1773
rect 27479 1789 27527 1805
rect 27479 1755 27493 1789
rect 27479 1721 27527 1755
rect 27064 1677 27080 1711
rect 27114 1677 27130 1711
rect 27479 1687 27493 1721
rect 27479 1643 27527 1687
rect 27561 1789 27627 1805
rect 27561 1755 27577 1789
rect 27611 1759 27627 1789
rect 27561 1725 27579 1755
rect 27613 1725 27627 1759
rect 27561 1721 27627 1725
rect 27561 1687 27577 1721
rect 27611 1687 27627 1721
rect 27561 1677 27627 1687
rect 27661 1789 27715 1805
rect 27695 1755 27715 1789
rect 27661 1721 27715 1755
rect 27695 1687 27715 1721
rect 27661 1643 27715 1687
rect 28553 1789 28601 1805
rect 28553 1755 28567 1789
rect 28553 1721 28601 1755
rect 28553 1687 28567 1721
rect 28553 1643 28601 1687
rect 28635 1789 28701 1805
rect 28635 1764 28651 1789
rect 28635 1730 28649 1764
rect 28685 1755 28701 1789
rect 28683 1730 28701 1755
rect 28635 1721 28701 1730
rect 28635 1687 28651 1721
rect 28685 1687 28701 1721
rect 28635 1677 28701 1687
rect 28735 1789 28789 1805
rect 28769 1755 28789 1789
rect 28735 1721 28789 1755
rect 28769 1687 28789 1721
rect 28735 1643 28789 1687
rect 27176 1596 27192 1630
rect 27226 1596 27242 1630
rect 27458 1609 27487 1643
rect 27521 1609 27579 1643
rect 27613 1609 27671 1643
rect 27705 1609 27734 1643
rect 28532 1609 28561 1643
rect 28595 1609 28653 1643
rect 28687 1609 28745 1643
rect 28779 1609 28808 1643
rect 27048 1546 27082 1562
rect 27048 1476 27082 1510
rect 27048 1424 27082 1440
rect 27144 1546 27178 1562
rect 27144 1476 27178 1510
rect 27144 1424 27178 1440
rect 27240 1546 27274 1562
rect 27240 1476 27274 1510
rect 27274 1440 27622 1464
rect 27240 1424 27622 1440
rect 26960 1356 27096 1390
rect 27130 1356 27146 1390
rect 26875 1286 27270 1306
rect 26875 1281 27137 1286
rect 26875 1272 27016 1281
rect 27000 1247 27016 1272
rect 27050 1252 27137 1281
rect 27171 1262 27270 1286
rect 27442 1264 27488 1266
rect 27442 1262 27446 1264
rect 27171 1252 27446 1262
rect 27050 1247 27446 1252
rect 27000 1230 27446 1247
rect 27480 1230 27488 1264
rect 27000 1228 27488 1230
rect 27442 1222 27488 1228
rect 25774 1107 25803 1141
rect 25837 1107 25895 1141
rect 25929 1107 25987 1141
rect 26021 1107 26050 1141
rect 25370 1055 25606 1066
rect 25012 1047 25606 1055
rect 25012 1022 25014 1047
rect 24926 979 24960 981
rect 24926 943 24960 945
rect 24926 858 24960 877
rect 25048 1022 25572 1047
rect 25658 1047 25734 1066
rect 25658 1026 25660 1047
rect 25014 979 25048 981
rect 25270 949 25286 983
rect 25320 949 25336 983
rect 25572 979 25606 981
rect 25014 943 25048 945
rect 25572 943 25606 945
rect 25014 858 25048 877
rect 25142 887 25176 906
rect 25142 819 25176 821
rect 24954 781 24970 815
rect 25004 781 25020 815
rect 25142 783 25176 785
rect 24642 703 24654 737
rect 24642 669 24688 703
rect 24642 635 24654 669
rect 24232 561 24261 595
rect 24295 561 24353 595
rect 24387 561 24445 595
rect 24479 561 24508 595
rect 24642 589 24688 635
rect 24722 737 24788 749
rect 24722 703 24738 737
rect 24772 703 24788 737
rect 24722 690 24788 703
rect 25142 698 25176 717
rect 25238 887 25272 906
rect 25238 819 25272 821
rect 25238 783 25272 785
rect 25238 698 25272 717
rect 25334 887 25368 906
rect 25572 858 25606 877
rect 25694 1026 25734 1047
rect 25842 1065 25884 1107
rect 26120 1105 26149 1139
rect 26183 1105 26241 1139
rect 26275 1105 26333 1139
rect 26367 1105 26396 1139
rect 26541 1133 26575 1140
rect 25842 1031 25850 1065
rect 25660 979 25694 981
rect 25660 943 25694 945
rect 25842 997 25884 1031
rect 25842 963 25850 997
rect 25842 929 25884 963
rect 25842 895 25850 929
rect 25842 879 25884 895
rect 25918 1065 25984 1073
rect 25918 1031 25934 1065
rect 25968 1031 25984 1065
rect 25918 997 25984 1031
rect 25918 963 25934 997
rect 25968 963 25984 997
rect 25918 929 25984 963
rect 25918 895 25934 929
rect 25968 895 25984 929
rect 25918 877 25984 895
rect 26153 1055 26189 1071
rect 26153 1021 26155 1055
rect 26153 987 26189 1021
rect 26153 953 26155 987
rect 26225 1055 26291 1105
rect 26466 1099 26495 1133
rect 26529 1099 26587 1133
rect 26621 1099 26679 1133
rect 26713 1099 26742 1133
rect 26842 1109 26858 1143
rect 26892 1109 26908 1143
rect 27066 1130 27180 1132
rect 26225 1021 26241 1055
rect 26275 1021 26291 1055
rect 26225 987 26291 1021
rect 26225 953 26241 987
rect 26275 953 26291 987
rect 26325 1055 26379 1071
rect 26325 1021 26327 1055
rect 26361 1021 26379 1055
rect 26325 974 26379 1021
rect 26153 919 26189 953
rect 26325 940 26327 974
rect 26361 940 26379 974
rect 26153 885 26288 919
rect 26325 890 26379 940
rect 25660 858 25694 877
rect 25334 819 25368 821
rect 25746 843 25890 844
rect 25746 829 25904 843
rect 25334 783 25368 785
rect 25600 816 25666 818
rect 25746 816 25854 829
rect 25600 815 25854 816
rect 25600 781 25616 815
rect 25650 802 25854 815
rect 25650 782 25786 802
rect 25838 795 25854 802
rect 25888 795 25904 829
rect 25650 781 25666 782
rect 25838 745 25884 761
rect 25938 757 25984 877
rect 26254 856 26288 885
rect 26141 827 26209 849
rect 26141 826 26157 827
rect 26141 792 26155 826
rect 26191 793 26209 827
rect 26189 792 26209 793
rect 26141 775 26209 792
rect 26254 840 26309 856
rect 26254 806 26275 840
rect 26254 790 26309 806
rect 26343 840 26379 890
rect 26534 1057 26576 1099
rect 27066 1091 27348 1130
rect 27488 1109 27504 1143
rect 27538 1109 27554 1143
rect 27066 1066 27105 1091
rect 26534 1023 26542 1057
rect 26534 989 26576 1023
rect 26534 955 26542 989
rect 26534 921 26576 955
rect 26534 887 26542 921
rect 26534 871 26576 887
rect 26610 1057 26676 1065
rect 26610 1023 26626 1057
rect 26660 1023 26676 1057
rect 26610 989 26676 1023
rect 26610 955 26626 989
rect 26660 955 26676 989
rect 26610 921 26676 955
rect 26610 887 26626 921
rect 26660 887 26676 921
rect 26610 869 26676 887
rect 26343 838 26384 840
rect 26343 804 26348 838
rect 26382 804 26384 838
rect 26343 802 26384 804
rect 26530 832 26596 835
rect 25368 717 25614 734
rect 25334 700 25614 717
rect 25334 698 25368 700
rect 24722 669 25064 690
rect 24722 635 24738 669
rect 24772 658 25064 669
rect 24772 655 25240 658
rect 24772 654 25190 655
rect 24772 635 24794 654
rect 24722 630 24794 635
rect 24722 623 24788 630
rect 25028 622 25190 654
rect 25174 621 25190 622
rect 25224 621 25240 655
rect 25566 612 25614 700
rect 24578 555 24607 589
rect 24641 555 24699 589
rect 24733 555 24791 589
rect 24825 555 24854 589
rect 24936 584 24982 594
rect 24936 550 24942 584
rect 24976 564 24982 584
rect 25566 578 25574 612
rect 25608 578 25614 612
rect 25838 711 25850 745
rect 25838 677 25884 711
rect 25838 643 25850 677
rect 25838 597 25884 643
rect 25918 745 25984 757
rect 25918 694 25934 745
rect 25968 694 25984 745
rect 26254 739 26288 790
rect 25918 677 25984 694
rect 25918 643 25934 677
rect 25968 643 25984 677
rect 25918 631 25984 643
rect 26155 705 26288 739
rect 26343 730 26379 802
rect 26530 798 26544 832
rect 26578 821 26596 832
rect 26530 787 26546 798
rect 26580 787 26596 821
rect 26155 684 26189 705
rect 26327 701 26379 730
rect 26155 629 26189 650
rect 26225 637 26241 671
rect 26275 637 26291 671
rect 24976 550 24986 564
rect 21574 420 21608 454
rect 21574 368 21608 384
rect 22966 444 23098 480
rect 23270 490 23304 506
rect 23366 490 23400 506
rect 23304 454 23305 455
rect 22966 396 23002 444
rect 23270 420 23305 454
rect 23304 418 23305 420
rect 23366 420 23400 454
rect 23150 396 23270 418
rect 22966 384 23270 396
rect 23304 384 23306 418
rect 22966 382 23306 384
rect 22966 360 23186 382
rect 23270 368 23304 382
rect 23366 368 23400 384
rect 23462 490 23496 506
rect 24936 480 24986 550
rect 25286 540 25302 574
rect 25336 540 25352 574
rect 25566 566 25614 578
rect 25774 563 25803 597
rect 25837 563 25895 597
rect 25929 563 25987 597
rect 26021 563 26050 597
rect 26225 595 26291 637
rect 26361 667 26379 701
rect 26327 629 26379 667
rect 26530 737 26576 753
rect 26630 749 26676 869
rect 26814 1047 26848 1066
rect 26900 1057 27105 1066
rect 27139 1089 27348 1091
rect 27139 1057 27224 1089
rect 26900 1055 27224 1057
rect 27258 1066 27348 1089
rect 27588 1066 27622 1424
rect 28532 1398 28566 1609
rect 28763 1306 28797 1609
rect 28848 1390 28882 2004
rect 29048 2002 29114 2004
rect 29365 2009 29381 2043
rect 29415 2009 29431 2043
rect 29365 1975 29431 2009
rect 28920 1943 28954 1962
rect 28920 1875 28954 1877
rect 28920 1839 28954 1841
rect 28920 1754 28954 1773
rect 29016 1943 29050 1962
rect 29016 1875 29050 1877
rect 29016 1839 29050 1841
rect 29016 1754 29050 1773
rect 29112 1943 29146 1962
rect 29365 1941 29381 1975
rect 29415 1959 29431 1975
rect 29537 2111 29603 2153
rect 29571 2077 29603 2111
rect 29537 2043 29603 2077
rect 29571 2009 29603 2043
rect 29537 1975 29603 2009
rect 29415 1941 29501 1959
rect 29365 1925 29501 1941
rect 29571 1941 29603 1975
rect 29537 1925 29603 1941
rect 30439 2111 30505 2116
rect 30439 2077 30455 2111
rect 30489 2077 30505 2111
rect 30439 2043 30505 2077
rect 30439 2009 30455 2043
rect 30489 2009 30505 2043
rect 30439 1975 30505 2009
rect 30439 1941 30455 1975
rect 30489 1959 30505 1975
rect 30611 2111 30677 2153
rect 30645 2077 30677 2111
rect 30844 2147 31126 2153
rect 30844 2113 30883 2147
rect 30917 2145 31126 2147
rect 30917 2113 31002 2145
rect 30844 2111 31002 2113
rect 31036 2111 31126 2145
rect 30844 2078 31126 2111
rect 31253 2111 31319 2116
rect 30611 2043 30677 2077
rect 30645 2009 30677 2043
rect 31253 2077 31269 2111
rect 31303 2077 31319 2111
rect 31253 2043 31319 2077
rect 30611 1975 30677 2009
rect 30489 1941 30575 1959
rect 30439 1925 30575 1941
rect 30645 1941 30677 1975
rect 30611 1925 30677 1941
rect 30736 2039 31002 2040
rect 30736 2005 30952 2039
rect 30986 2005 31002 2039
rect 30736 2004 31002 2005
rect 29112 1875 29146 1877
rect 29363 1882 29433 1891
rect 29363 1848 29379 1882
rect 29413 1875 29433 1882
rect 29363 1841 29383 1848
rect 29417 1841 29433 1875
rect 29112 1839 29146 1841
rect 29467 1805 29501 1925
rect 29535 1882 29605 1891
rect 29535 1875 29553 1882
rect 29535 1841 29551 1875
rect 29587 1848 29605 1882
rect 29585 1841 29605 1848
rect 30437 1884 30507 1891
rect 30437 1850 30455 1884
rect 30489 1875 30507 1884
rect 30437 1841 30457 1850
rect 30491 1841 30507 1875
rect 30541 1805 30575 1925
rect 30609 1880 30679 1891
rect 30609 1875 30628 1880
rect 30609 1841 30625 1875
rect 30662 1846 30679 1880
rect 30659 1841 30679 1846
rect 29112 1754 29146 1773
rect 29367 1789 29415 1805
rect 29367 1755 29381 1789
rect 29367 1721 29415 1755
rect 28952 1677 28968 1711
rect 29002 1677 29018 1711
rect 29367 1687 29381 1721
rect 29367 1643 29415 1687
rect 29449 1789 29515 1805
rect 29449 1755 29465 1789
rect 29499 1759 29515 1789
rect 29449 1725 29467 1755
rect 29501 1725 29515 1759
rect 29449 1721 29515 1725
rect 29449 1687 29465 1721
rect 29499 1687 29515 1721
rect 29449 1677 29515 1687
rect 29549 1789 29603 1805
rect 29583 1755 29603 1789
rect 29549 1721 29603 1755
rect 29583 1687 29603 1721
rect 29549 1643 29603 1687
rect 30441 1789 30489 1805
rect 30441 1755 30455 1789
rect 30441 1721 30489 1755
rect 30441 1687 30455 1721
rect 30441 1643 30489 1687
rect 30523 1789 30589 1805
rect 30523 1764 30539 1789
rect 30523 1730 30537 1764
rect 30573 1755 30589 1789
rect 30571 1730 30589 1755
rect 30523 1721 30589 1730
rect 30523 1687 30539 1721
rect 30573 1687 30589 1721
rect 30523 1677 30589 1687
rect 30623 1789 30677 1805
rect 30657 1755 30677 1789
rect 30623 1721 30677 1755
rect 30657 1687 30677 1721
rect 30623 1643 30677 1687
rect 29064 1596 29080 1630
rect 29114 1596 29130 1630
rect 29346 1609 29375 1643
rect 29409 1609 29467 1643
rect 29501 1609 29559 1643
rect 29593 1609 29622 1643
rect 30420 1609 30449 1643
rect 30483 1609 30541 1643
rect 30575 1609 30633 1643
rect 30667 1609 30696 1643
rect 28936 1546 28970 1562
rect 28936 1476 28970 1510
rect 28936 1424 28970 1440
rect 29032 1546 29066 1562
rect 29032 1476 29066 1510
rect 29032 1424 29066 1440
rect 29128 1546 29162 1562
rect 29128 1476 29162 1510
rect 29162 1440 29510 1464
rect 29128 1424 29510 1440
rect 28848 1356 28984 1390
rect 29018 1356 29034 1390
rect 28763 1286 29158 1306
rect 28763 1281 29025 1286
rect 28763 1272 28904 1281
rect 28888 1247 28904 1272
rect 28938 1252 29025 1281
rect 29059 1262 29158 1286
rect 29330 1264 29376 1266
rect 29330 1262 29334 1264
rect 29059 1252 29334 1262
rect 28938 1247 29334 1252
rect 28888 1230 29334 1247
rect 29368 1230 29376 1264
rect 28888 1228 29376 1230
rect 29330 1222 29376 1228
rect 27662 1107 27691 1141
rect 27725 1107 27783 1141
rect 27817 1107 27875 1141
rect 27909 1107 27938 1141
rect 27258 1055 27494 1066
rect 26900 1047 27494 1055
rect 26900 1022 26902 1047
rect 26814 979 26848 981
rect 26814 943 26848 945
rect 26814 858 26848 877
rect 26936 1022 27460 1047
rect 27546 1047 27622 1066
rect 27546 1026 27548 1047
rect 26902 979 26936 981
rect 27158 949 27174 983
rect 27208 949 27224 983
rect 27460 979 27494 981
rect 26902 943 26936 945
rect 27460 943 27494 945
rect 26902 858 26936 877
rect 27030 887 27064 906
rect 27030 819 27064 821
rect 26842 781 26858 815
rect 26892 781 26908 815
rect 27030 783 27064 785
rect 26530 703 26542 737
rect 26530 669 26576 703
rect 26530 635 26542 669
rect 26120 561 26149 595
rect 26183 561 26241 595
rect 26275 561 26333 595
rect 26367 561 26396 595
rect 26530 589 26576 635
rect 26610 737 26676 749
rect 26610 703 26626 737
rect 26660 703 26676 737
rect 26610 690 26676 703
rect 27030 698 27064 717
rect 27126 887 27160 906
rect 27126 819 27160 821
rect 27126 783 27160 785
rect 27126 698 27160 717
rect 27222 887 27256 906
rect 27460 858 27494 877
rect 27582 1026 27622 1047
rect 27730 1065 27772 1107
rect 28008 1105 28037 1139
rect 28071 1105 28129 1139
rect 28163 1105 28221 1139
rect 28255 1105 28284 1139
rect 28429 1133 28463 1140
rect 27730 1031 27738 1065
rect 27548 979 27582 981
rect 27548 943 27582 945
rect 27730 997 27772 1031
rect 27730 963 27738 997
rect 27730 929 27772 963
rect 27730 895 27738 929
rect 27730 879 27772 895
rect 27806 1065 27872 1073
rect 27806 1031 27822 1065
rect 27856 1031 27872 1065
rect 27806 997 27872 1031
rect 27806 963 27822 997
rect 27856 963 27872 997
rect 27806 929 27872 963
rect 27806 895 27822 929
rect 27856 895 27872 929
rect 27806 877 27872 895
rect 28041 1055 28077 1071
rect 28041 1021 28043 1055
rect 28041 987 28077 1021
rect 28041 953 28043 987
rect 28113 1055 28179 1105
rect 28354 1099 28383 1133
rect 28417 1099 28475 1133
rect 28509 1099 28567 1133
rect 28601 1099 28630 1133
rect 28730 1109 28746 1143
rect 28780 1109 28796 1143
rect 28954 1130 29068 1132
rect 28113 1021 28129 1055
rect 28163 1021 28179 1055
rect 28113 987 28179 1021
rect 28113 953 28129 987
rect 28163 953 28179 987
rect 28213 1055 28267 1071
rect 28213 1021 28215 1055
rect 28249 1021 28267 1055
rect 28213 974 28267 1021
rect 28041 919 28077 953
rect 28213 940 28215 974
rect 28249 940 28267 974
rect 28041 885 28176 919
rect 28213 890 28267 940
rect 27548 858 27582 877
rect 27222 819 27256 821
rect 27634 843 27778 844
rect 27634 829 27792 843
rect 27222 783 27256 785
rect 27488 816 27554 818
rect 27634 816 27742 829
rect 27488 815 27742 816
rect 27488 781 27504 815
rect 27538 802 27742 815
rect 27538 782 27674 802
rect 27726 795 27742 802
rect 27776 795 27792 829
rect 27538 781 27554 782
rect 27726 745 27772 761
rect 27826 757 27872 877
rect 28142 856 28176 885
rect 28029 827 28097 849
rect 28029 826 28045 827
rect 28029 792 28043 826
rect 28079 793 28097 827
rect 28077 792 28097 793
rect 28029 775 28097 792
rect 28142 840 28197 856
rect 28142 806 28163 840
rect 28142 790 28197 806
rect 28231 840 28267 890
rect 28422 1057 28464 1099
rect 28954 1091 29236 1130
rect 29376 1109 29392 1143
rect 29426 1109 29442 1143
rect 28954 1066 28993 1091
rect 28422 1023 28430 1057
rect 28422 989 28464 1023
rect 28422 955 28430 989
rect 28422 921 28464 955
rect 28422 887 28430 921
rect 28422 871 28464 887
rect 28498 1057 28564 1065
rect 28498 1023 28514 1057
rect 28548 1023 28564 1057
rect 28498 989 28564 1023
rect 28498 955 28514 989
rect 28548 955 28564 989
rect 28498 921 28564 955
rect 28498 887 28514 921
rect 28548 887 28564 921
rect 28498 869 28564 887
rect 28231 838 28272 840
rect 28231 804 28236 838
rect 28270 804 28272 838
rect 28231 802 28272 804
rect 28418 832 28484 835
rect 27256 717 27502 734
rect 27222 700 27502 717
rect 27222 698 27256 700
rect 26610 669 26952 690
rect 26610 635 26626 669
rect 26660 658 26952 669
rect 26660 655 27128 658
rect 26660 654 27078 655
rect 26660 635 26682 654
rect 26610 630 26682 635
rect 26610 623 26676 630
rect 26916 622 27078 654
rect 27062 621 27078 622
rect 27112 621 27128 655
rect 27454 612 27502 700
rect 26466 555 26495 589
rect 26529 555 26587 589
rect 26621 555 26679 589
rect 26713 555 26742 589
rect 26824 584 26870 594
rect 26824 550 26830 584
rect 26864 564 26870 584
rect 27454 578 27462 612
rect 27496 578 27502 612
rect 27726 711 27738 745
rect 27726 677 27772 711
rect 27726 643 27738 677
rect 27726 597 27772 643
rect 27806 745 27872 757
rect 27806 694 27822 745
rect 27856 694 27872 745
rect 28142 739 28176 790
rect 27806 677 27872 694
rect 27806 643 27822 677
rect 27856 643 27872 677
rect 27806 631 27872 643
rect 28043 705 28176 739
rect 28231 730 28267 802
rect 28418 798 28432 832
rect 28466 821 28484 832
rect 28418 787 28434 798
rect 28468 787 28484 821
rect 28043 684 28077 705
rect 28215 701 28267 730
rect 28043 629 28077 650
rect 28113 637 28129 671
rect 28163 637 28179 671
rect 26864 550 26874 564
rect 23462 420 23496 454
rect 23462 368 23496 384
rect 24854 444 24986 480
rect 25158 490 25192 506
rect 25254 490 25288 506
rect 25192 454 25193 455
rect 24854 396 24890 444
rect 25158 420 25193 454
rect 25192 418 25193 420
rect 25254 420 25288 454
rect 25038 396 25158 418
rect 24854 384 25158 396
rect 25192 384 25194 418
rect 24854 382 25194 384
rect 24854 360 25074 382
rect 25158 368 25192 382
rect 25254 368 25288 384
rect 25350 490 25384 506
rect 26824 480 26874 550
rect 27174 540 27190 574
rect 27224 540 27240 574
rect 27454 566 27502 578
rect 27662 563 27691 597
rect 27725 563 27783 597
rect 27817 563 27875 597
rect 27909 563 27938 597
rect 28113 595 28179 637
rect 28249 667 28267 701
rect 28215 629 28267 667
rect 28418 737 28464 753
rect 28518 749 28564 869
rect 28702 1047 28736 1066
rect 28788 1057 28993 1066
rect 29027 1089 29236 1091
rect 29027 1057 29112 1089
rect 28788 1055 29112 1057
rect 29146 1066 29236 1089
rect 29476 1066 29510 1424
rect 30420 1398 30454 1609
rect 30651 1306 30685 1609
rect 30736 1390 30770 2004
rect 30936 2002 31002 2004
rect 31253 2009 31269 2043
rect 31303 2009 31319 2043
rect 31253 1975 31319 2009
rect 30808 1943 30842 1962
rect 30808 1875 30842 1877
rect 30808 1839 30842 1841
rect 30808 1754 30842 1773
rect 30904 1943 30938 1962
rect 30904 1875 30938 1877
rect 30904 1839 30938 1841
rect 30904 1754 30938 1773
rect 31000 1943 31034 1962
rect 31253 1941 31269 1975
rect 31303 1959 31319 1975
rect 31425 2111 31491 2153
rect 31459 2077 31491 2111
rect 31425 2043 31491 2077
rect 31459 2009 31491 2043
rect 31425 1975 31491 2009
rect 31303 1941 31389 1959
rect 31253 1925 31389 1941
rect 31459 1941 31491 1975
rect 31425 1925 31491 1941
rect 32327 2111 32393 2116
rect 32327 2077 32343 2111
rect 32377 2077 32393 2111
rect 32327 2043 32393 2077
rect 32327 2009 32343 2043
rect 32377 2009 32393 2043
rect 32327 1975 32393 2009
rect 32327 1941 32343 1975
rect 32377 1959 32393 1975
rect 32499 2111 32565 2153
rect 32533 2077 32565 2111
rect 32732 2147 33014 2153
rect 32732 2113 32771 2147
rect 32805 2145 33014 2147
rect 32805 2113 32890 2145
rect 32732 2111 32890 2113
rect 32924 2111 33014 2145
rect 32732 2078 33014 2111
rect 33141 2111 33207 2116
rect 32499 2043 32565 2077
rect 32533 2009 32565 2043
rect 33141 2077 33157 2111
rect 33191 2077 33207 2111
rect 33141 2043 33207 2077
rect 32499 1975 32565 2009
rect 32377 1941 32463 1959
rect 32327 1925 32463 1941
rect 32533 1941 32565 1975
rect 32499 1925 32565 1941
rect 32624 2039 32890 2040
rect 32624 2005 32840 2039
rect 32874 2005 32890 2039
rect 32624 2004 32890 2005
rect 31000 1875 31034 1877
rect 31251 1882 31321 1891
rect 31251 1848 31267 1882
rect 31301 1875 31321 1882
rect 31251 1841 31271 1848
rect 31305 1841 31321 1875
rect 31000 1839 31034 1841
rect 31355 1805 31389 1925
rect 31423 1882 31493 1891
rect 31423 1875 31441 1882
rect 31423 1841 31439 1875
rect 31475 1848 31493 1882
rect 31473 1841 31493 1848
rect 32325 1884 32395 1891
rect 32325 1850 32343 1884
rect 32377 1875 32395 1884
rect 32325 1841 32345 1850
rect 32379 1841 32395 1875
rect 32429 1805 32463 1925
rect 32497 1880 32567 1891
rect 32497 1875 32516 1880
rect 32497 1841 32513 1875
rect 32550 1846 32567 1880
rect 32547 1841 32567 1846
rect 31000 1754 31034 1773
rect 31255 1789 31303 1805
rect 31255 1755 31269 1789
rect 31255 1721 31303 1755
rect 30840 1677 30856 1711
rect 30890 1677 30906 1711
rect 31255 1687 31269 1721
rect 31255 1643 31303 1687
rect 31337 1789 31403 1805
rect 31337 1755 31353 1789
rect 31387 1759 31403 1789
rect 31337 1725 31355 1755
rect 31389 1725 31403 1759
rect 31337 1721 31403 1725
rect 31337 1687 31353 1721
rect 31387 1687 31403 1721
rect 31337 1677 31403 1687
rect 31437 1789 31491 1805
rect 31471 1755 31491 1789
rect 31437 1721 31491 1755
rect 31471 1687 31491 1721
rect 31437 1643 31491 1687
rect 32329 1789 32377 1805
rect 32329 1755 32343 1789
rect 32329 1721 32377 1755
rect 32329 1687 32343 1721
rect 32329 1643 32377 1687
rect 32411 1789 32477 1805
rect 32411 1764 32427 1789
rect 32411 1730 32425 1764
rect 32461 1755 32477 1789
rect 32459 1730 32477 1755
rect 32411 1721 32477 1730
rect 32411 1687 32427 1721
rect 32461 1687 32477 1721
rect 32411 1677 32477 1687
rect 32511 1789 32565 1805
rect 32545 1755 32565 1789
rect 32511 1721 32565 1755
rect 32545 1687 32565 1721
rect 32511 1643 32565 1687
rect 30952 1596 30968 1630
rect 31002 1596 31018 1630
rect 31234 1609 31263 1643
rect 31297 1609 31355 1643
rect 31389 1609 31447 1643
rect 31481 1609 31510 1643
rect 32308 1609 32337 1643
rect 32371 1609 32429 1643
rect 32463 1609 32521 1643
rect 32555 1609 32584 1643
rect 30824 1546 30858 1562
rect 30824 1476 30858 1510
rect 30824 1424 30858 1440
rect 30920 1546 30954 1562
rect 30920 1476 30954 1510
rect 30920 1424 30954 1440
rect 31016 1546 31050 1562
rect 31016 1476 31050 1510
rect 31050 1440 31398 1464
rect 31016 1424 31398 1440
rect 30736 1356 30872 1390
rect 30906 1356 30922 1390
rect 30651 1286 31046 1306
rect 30651 1281 30913 1286
rect 30651 1272 30792 1281
rect 30776 1247 30792 1272
rect 30826 1252 30913 1281
rect 30947 1262 31046 1286
rect 31218 1264 31264 1266
rect 31218 1262 31222 1264
rect 30947 1252 31222 1262
rect 30826 1247 31222 1252
rect 30776 1230 31222 1247
rect 31256 1230 31264 1264
rect 30776 1228 31264 1230
rect 31218 1222 31264 1228
rect 29550 1107 29579 1141
rect 29613 1107 29671 1141
rect 29705 1107 29763 1141
rect 29797 1107 29826 1141
rect 29146 1055 29382 1066
rect 28788 1047 29382 1055
rect 28788 1022 28790 1047
rect 28702 979 28736 981
rect 28702 943 28736 945
rect 28702 858 28736 877
rect 28824 1022 29348 1047
rect 29434 1047 29510 1066
rect 29434 1026 29436 1047
rect 28790 979 28824 981
rect 29046 949 29062 983
rect 29096 949 29112 983
rect 29348 979 29382 981
rect 28790 943 28824 945
rect 29348 943 29382 945
rect 28790 858 28824 877
rect 28918 887 28952 906
rect 28918 819 28952 821
rect 28730 781 28746 815
rect 28780 781 28796 815
rect 28918 783 28952 785
rect 28418 703 28430 737
rect 28418 669 28464 703
rect 28418 635 28430 669
rect 28008 561 28037 595
rect 28071 561 28129 595
rect 28163 561 28221 595
rect 28255 561 28284 595
rect 28418 589 28464 635
rect 28498 737 28564 749
rect 28498 703 28514 737
rect 28548 703 28564 737
rect 28498 690 28564 703
rect 28918 698 28952 717
rect 29014 887 29048 906
rect 29014 819 29048 821
rect 29014 783 29048 785
rect 29014 698 29048 717
rect 29110 887 29144 906
rect 29348 858 29382 877
rect 29470 1026 29510 1047
rect 29618 1065 29660 1107
rect 29896 1105 29925 1139
rect 29959 1105 30017 1139
rect 30051 1105 30109 1139
rect 30143 1105 30172 1139
rect 30317 1133 30351 1140
rect 29618 1031 29626 1065
rect 29436 979 29470 981
rect 29436 943 29470 945
rect 29618 997 29660 1031
rect 29618 963 29626 997
rect 29618 929 29660 963
rect 29618 895 29626 929
rect 29618 879 29660 895
rect 29694 1065 29760 1073
rect 29694 1031 29710 1065
rect 29744 1031 29760 1065
rect 29694 997 29760 1031
rect 29694 963 29710 997
rect 29744 963 29760 997
rect 29694 929 29760 963
rect 29694 895 29710 929
rect 29744 895 29760 929
rect 29694 877 29760 895
rect 29929 1055 29965 1071
rect 29929 1021 29931 1055
rect 29929 987 29965 1021
rect 29929 953 29931 987
rect 30001 1055 30067 1105
rect 30242 1099 30271 1133
rect 30305 1099 30363 1133
rect 30397 1099 30455 1133
rect 30489 1099 30518 1133
rect 30618 1109 30634 1143
rect 30668 1109 30684 1143
rect 30842 1130 30956 1132
rect 30001 1021 30017 1055
rect 30051 1021 30067 1055
rect 30001 987 30067 1021
rect 30001 953 30017 987
rect 30051 953 30067 987
rect 30101 1055 30155 1071
rect 30101 1021 30103 1055
rect 30137 1021 30155 1055
rect 30101 974 30155 1021
rect 29929 919 29965 953
rect 30101 940 30103 974
rect 30137 940 30155 974
rect 29929 885 30064 919
rect 30101 890 30155 940
rect 29436 858 29470 877
rect 29110 819 29144 821
rect 29522 843 29666 844
rect 29522 829 29680 843
rect 29110 783 29144 785
rect 29376 816 29442 818
rect 29522 816 29630 829
rect 29376 815 29630 816
rect 29376 781 29392 815
rect 29426 802 29630 815
rect 29426 782 29562 802
rect 29614 795 29630 802
rect 29664 795 29680 829
rect 29426 781 29442 782
rect 29614 745 29660 761
rect 29714 757 29760 877
rect 30030 856 30064 885
rect 29917 827 29985 849
rect 29917 826 29933 827
rect 29917 792 29931 826
rect 29967 793 29985 827
rect 29965 792 29985 793
rect 29917 775 29985 792
rect 30030 840 30085 856
rect 30030 806 30051 840
rect 30030 790 30085 806
rect 30119 840 30155 890
rect 30310 1057 30352 1099
rect 30842 1091 31124 1130
rect 31264 1109 31280 1143
rect 31314 1109 31330 1143
rect 30842 1066 30881 1091
rect 30310 1023 30318 1057
rect 30310 989 30352 1023
rect 30310 955 30318 989
rect 30310 921 30352 955
rect 30310 887 30318 921
rect 30310 871 30352 887
rect 30386 1057 30452 1065
rect 30386 1023 30402 1057
rect 30436 1023 30452 1057
rect 30386 989 30452 1023
rect 30386 955 30402 989
rect 30436 955 30452 989
rect 30386 921 30452 955
rect 30386 887 30402 921
rect 30436 887 30452 921
rect 30386 869 30452 887
rect 30119 838 30160 840
rect 30119 804 30124 838
rect 30158 804 30160 838
rect 30119 802 30160 804
rect 30306 832 30372 835
rect 29144 717 29390 734
rect 29110 700 29390 717
rect 29110 698 29144 700
rect 28498 669 28840 690
rect 28498 635 28514 669
rect 28548 658 28840 669
rect 28548 655 29016 658
rect 28548 654 28966 655
rect 28548 635 28570 654
rect 28498 630 28570 635
rect 28498 623 28564 630
rect 28804 622 28966 654
rect 28950 621 28966 622
rect 29000 621 29016 655
rect 29342 612 29390 700
rect 28354 555 28383 589
rect 28417 555 28475 589
rect 28509 555 28567 589
rect 28601 555 28630 589
rect 28712 584 28758 594
rect 28712 550 28718 584
rect 28752 564 28758 584
rect 29342 578 29350 612
rect 29384 578 29390 612
rect 29614 711 29626 745
rect 29614 677 29660 711
rect 29614 643 29626 677
rect 29614 597 29660 643
rect 29694 745 29760 757
rect 29694 694 29710 745
rect 29744 694 29760 745
rect 30030 739 30064 790
rect 29694 677 29760 694
rect 29694 643 29710 677
rect 29744 643 29760 677
rect 29694 631 29760 643
rect 29931 705 30064 739
rect 30119 730 30155 802
rect 30306 798 30320 832
rect 30354 821 30372 832
rect 30306 787 30322 798
rect 30356 787 30372 821
rect 29931 684 29965 705
rect 30103 701 30155 730
rect 29931 629 29965 650
rect 30001 637 30017 671
rect 30051 637 30067 671
rect 28752 550 28762 564
rect 25350 420 25384 454
rect 25350 368 25384 384
rect 26742 444 26874 480
rect 27046 490 27080 506
rect 27142 490 27176 506
rect 27080 454 27081 455
rect 26742 396 26778 444
rect 27046 420 27081 454
rect 27080 418 27081 420
rect 27142 420 27176 454
rect 26926 396 27046 418
rect 26742 384 27046 396
rect 27080 384 27082 418
rect 26742 382 27082 384
rect 26742 360 26962 382
rect 27046 368 27080 382
rect 27142 368 27176 384
rect 27238 490 27272 506
rect 28712 480 28762 550
rect 29062 540 29078 574
rect 29112 540 29128 574
rect 29342 566 29390 578
rect 29550 563 29579 597
rect 29613 563 29671 597
rect 29705 563 29763 597
rect 29797 563 29826 597
rect 30001 595 30067 637
rect 30137 667 30155 701
rect 30103 629 30155 667
rect 30306 737 30352 753
rect 30406 749 30452 869
rect 30590 1047 30624 1066
rect 30676 1057 30881 1066
rect 30915 1089 31124 1091
rect 30915 1057 31000 1089
rect 30676 1055 31000 1057
rect 31034 1066 31124 1089
rect 31364 1066 31398 1424
rect 32308 1398 32342 1609
rect 32539 1306 32573 1609
rect 32624 1390 32658 2004
rect 32824 2002 32890 2004
rect 33141 2009 33157 2043
rect 33191 2009 33207 2043
rect 33141 1975 33207 2009
rect 32696 1943 32730 1962
rect 32696 1875 32730 1877
rect 32696 1839 32730 1841
rect 32696 1754 32730 1773
rect 32792 1943 32826 1962
rect 32792 1875 32826 1877
rect 32792 1839 32826 1841
rect 32792 1754 32826 1773
rect 32888 1943 32922 1962
rect 33141 1941 33157 1975
rect 33191 1959 33207 1975
rect 33313 2111 33379 2153
rect 33347 2077 33379 2111
rect 33313 2043 33379 2077
rect 33347 2009 33379 2043
rect 33313 1975 33379 2009
rect 33191 1941 33277 1959
rect 33141 1925 33277 1941
rect 33347 1941 33379 1975
rect 33313 1925 33379 1941
rect 34215 2111 34281 2116
rect 34215 2077 34231 2111
rect 34265 2077 34281 2111
rect 34215 2043 34281 2077
rect 34215 2009 34231 2043
rect 34265 2009 34281 2043
rect 34215 1975 34281 2009
rect 34215 1941 34231 1975
rect 34265 1959 34281 1975
rect 34387 2111 34453 2153
rect 34421 2077 34453 2111
rect 34620 2147 34902 2153
rect 34620 2113 34659 2147
rect 34693 2145 34902 2147
rect 34693 2113 34778 2145
rect 34620 2111 34778 2113
rect 34812 2111 34902 2145
rect 34620 2078 34902 2111
rect 35029 2111 35095 2116
rect 34387 2043 34453 2077
rect 34421 2009 34453 2043
rect 35029 2077 35045 2111
rect 35079 2077 35095 2111
rect 35029 2043 35095 2077
rect 34387 1975 34453 2009
rect 34265 1941 34351 1959
rect 34215 1925 34351 1941
rect 34421 1941 34453 1975
rect 34387 1925 34453 1941
rect 34512 2039 34778 2040
rect 34512 2005 34728 2039
rect 34762 2005 34778 2039
rect 34512 2004 34778 2005
rect 32888 1875 32922 1877
rect 33139 1882 33209 1891
rect 33139 1848 33155 1882
rect 33189 1875 33209 1882
rect 33139 1841 33159 1848
rect 33193 1841 33209 1875
rect 32888 1839 32922 1841
rect 33243 1805 33277 1925
rect 33311 1882 33381 1891
rect 33311 1875 33329 1882
rect 33311 1841 33327 1875
rect 33363 1848 33381 1882
rect 33361 1841 33381 1848
rect 34213 1884 34283 1891
rect 34213 1850 34231 1884
rect 34265 1875 34283 1884
rect 34213 1841 34233 1850
rect 34267 1841 34283 1875
rect 34317 1805 34351 1925
rect 34385 1880 34455 1891
rect 34385 1875 34404 1880
rect 34385 1841 34401 1875
rect 34438 1846 34455 1880
rect 34435 1841 34455 1846
rect 32888 1754 32922 1773
rect 33143 1789 33191 1805
rect 33143 1755 33157 1789
rect 33143 1721 33191 1755
rect 32728 1677 32744 1711
rect 32778 1677 32794 1711
rect 33143 1687 33157 1721
rect 33143 1643 33191 1687
rect 33225 1789 33291 1805
rect 33225 1755 33241 1789
rect 33275 1759 33291 1789
rect 33225 1725 33243 1755
rect 33277 1725 33291 1759
rect 33225 1721 33291 1725
rect 33225 1687 33241 1721
rect 33275 1687 33291 1721
rect 33225 1677 33291 1687
rect 33325 1789 33379 1805
rect 33359 1755 33379 1789
rect 33325 1721 33379 1755
rect 33359 1687 33379 1721
rect 33325 1643 33379 1687
rect 34217 1789 34265 1805
rect 34217 1755 34231 1789
rect 34217 1721 34265 1755
rect 34217 1687 34231 1721
rect 34217 1643 34265 1687
rect 34299 1789 34365 1805
rect 34299 1764 34315 1789
rect 34299 1730 34313 1764
rect 34349 1755 34365 1789
rect 34347 1730 34365 1755
rect 34299 1721 34365 1730
rect 34299 1687 34315 1721
rect 34349 1687 34365 1721
rect 34299 1677 34365 1687
rect 34399 1789 34453 1805
rect 34433 1755 34453 1789
rect 34399 1721 34453 1755
rect 34433 1687 34453 1721
rect 34399 1643 34453 1687
rect 32840 1596 32856 1630
rect 32890 1596 32906 1630
rect 33122 1609 33151 1643
rect 33185 1609 33243 1643
rect 33277 1609 33335 1643
rect 33369 1609 33398 1643
rect 34196 1609 34225 1643
rect 34259 1609 34317 1643
rect 34351 1609 34409 1643
rect 34443 1609 34472 1643
rect 32712 1546 32746 1562
rect 32712 1476 32746 1510
rect 32712 1424 32746 1440
rect 32808 1546 32842 1562
rect 32808 1476 32842 1510
rect 32808 1424 32842 1440
rect 32904 1546 32938 1562
rect 32904 1476 32938 1510
rect 32938 1440 33286 1464
rect 32904 1424 33286 1440
rect 32624 1356 32760 1390
rect 32794 1356 32810 1390
rect 32539 1286 32934 1306
rect 32539 1281 32801 1286
rect 32539 1272 32680 1281
rect 32664 1247 32680 1272
rect 32714 1252 32801 1281
rect 32835 1262 32934 1286
rect 33106 1264 33152 1266
rect 33106 1262 33110 1264
rect 32835 1252 33110 1262
rect 32714 1247 33110 1252
rect 32664 1230 33110 1247
rect 33144 1230 33152 1264
rect 32664 1228 33152 1230
rect 33106 1222 33152 1228
rect 31438 1107 31467 1141
rect 31501 1107 31559 1141
rect 31593 1107 31651 1141
rect 31685 1107 31714 1141
rect 31034 1055 31270 1066
rect 30676 1047 31270 1055
rect 30676 1022 30678 1047
rect 30590 979 30624 981
rect 30590 943 30624 945
rect 30590 858 30624 877
rect 30712 1022 31236 1047
rect 31322 1047 31398 1066
rect 31322 1026 31324 1047
rect 30678 979 30712 981
rect 30934 949 30950 983
rect 30984 949 31000 983
rect 31236 979 31270 981
rect 30678 943 30712 945
rect 31236 943 31270 945
rect 30678 858 30712 877
rect 30806 887 30840 906
rect 30806 819 30840 821
rect 30618 781 30634 815
rect 30668 781 30684 815
rect 30806 783 30840 785
rect 30306 703 30318 737
rect 30306 669 30352 703
rect 30306 635 30318 669
rect 29896 561 29925 595
rect 29959 561 30017 595
rect 30051 561 30109 595
rect 30143 561 30172 595
rect 30306 589 30352 635
rect 30386 737 30452 749
rect 30386 703 30402 737
rect 30436 703 30452 737
rect 30386 690 30452 703
rect 30806 698 30840 717
rect 30902 887 30936 906
rect 30902 819 30936 821
rect 30902 783 30936 785
rect 30902 698 30936 717
rect 30998 887 31032 906
rect 31236 858 31270 877
rect 31358 1026 31398 1047
rect 31506 1065 31548 1107
rect 31784 1105 31813 1139
rect 31847 1105 31905 1139
rect 31939 1105 31997 1139
rect 32031 1105 32060 1139
rect 32205 1133 32239 1140
rect 31506 1031 31514 1065
rect 31324 979 31358 981
rect 31324 943 31358 945
rect 31506 997 31548 1031
rect 31506 963 31514 997
rect 31506 929 31548 963
rect 31506 895 31514 929
rect 31506 879 31548 895
rect 31582 1065 31648 1073
rect 31582 1031 31598 1065
rect 31632 1031 31648 1065
rect 31582 997 31648 1031
rect 31582 963 31598 997
rect 31632 963 31648 997
rect 31582 929 31648 963
rect 31582 895 31598 929
rect 31632 895 31648 929
rect 31582 877 31648 895
rect 31817 1055 31853 1071
rect 31817 1021 31819 1055
rect 31817 987 31853 1021
rect 31817 953 31819 987
rect 31889 1055 31955 1105
rect 32130 1099 32159 1133
rect 32193 1099 32251 1133
rect 32285 1099 32343 1133
rect 32377 1099 32406 1133
rect 32506 1109 32522 1143
rect 32556 1109 32572 1143
rect 32730 1130 32844 1132
rect 31889 1021 31905 1055
rect 31939 1021 31955 1055
rect 31889 987 31955 1021
rect 31889 953 31905 987
rect 31939 953 31955 987
rect 31989 1055 32043 1071
rect 31989 1021 31991 1055
rect 32025 1021 32043 1055
rect 31989 974 32043 1021
rect 31817 919 31853 953
rect 31989 940 31991 974
rect 32025 940 32043 974
rect 31817 885 31952 919
rect 31989 890 32043 940
rect 31324 858 31358 877
rect 30998 819 31032 821
rect 31410 843 31554 844
rect 31410 829 31568 843
rect 30998 783 31032 785
rect 31264 816 31330 818
rect 31410 816 31518 829
rect 31264 815 31518 816
rect 31264 781 31280 815
rect 31314 802 31518 815
rect 31314 782 31450 802
rect 31502 795 31518 802
rect 31552 795 31568 829
rect 31314 781 31330 782
rect 31502 745 31548 761
rect 31602 757 31648 877
rect 31918 856 31952 885
rect 31805 827 31873 849
rect 31805 826 31821 827
rect 31805 792 31819 826
rect 31855 793 31873 827
rect 31853 792 31873 793
rect 31805 775 31873 792
rect 31918 840 31973 856
rect 31918 806 31939 840
rect 31918 790 31973 806
rect 32007 840 32043 890
rect 32198 1057 32240 1099
rect 32730 1091 33012 1130
rect 33152 1109 33168 1143
rect 33202 1109 33218 1143
rect 32730 1066 32769 1091
rect 32198 1023 32206 1057
rect 32198 989 32240 1023
rect 32198 955 32206 989
rect 32198 921 32240 955
rect 32198 887 32206 921
rect 32198 871 32240 887
rect 32274 1057 32340 1065
rect 32274 1023 32290 1057
rect 32324 1023 32340 1057
rect 32274 989 32340 1023
rect 32274 955 32290 989
rect 32324 955 32340 989
rect 32274 921 32340 955
rect 32274 887 32290 921
rect 32324 887 32340 921
rect 32274 869 32340 887
rect 32007 838 32048 840
rect 32007 804 32012 838
rect 32046 804 32048 838
rect 32007 802 32048 804
rect 32194 832 32260 835
rect 31032 717 31278 734
rect 30998 700 31278 717
rect 30998 698 31032 700
rect 30386 669 30728 690
rect 30386 635 30402 669
rect 30436 658 30728 669
rect 30436 655 30904 658
rect 30436 654 30854 655
rect 30436 635 30458 654
rect 30386 630 30458 635
rect 30386 623 30452 630
rect 30692 622 30854 654
rect 30838 621 30854 622
rect 30888 621 30904 655
rect 31230 612 31278 700
rect 30242 555 30271 589
rect 30305 555 30363 589
rect 30397 555 30455 589
rect 30489 555 30518 589
rect 30600 584 30646 594
rect 30600 550 30606 584
rect 30640 564 30646 584
rect 31230 578 31238 612
rect 31272 578 31278 612
rect 31502 711 31514 745
rect 31502 677 31548 711
rect 31502 643 31514 677
rect 31502 597 31548 643
rect 31582 745 31648 757
rect 31582 694 31598 745
rect 31632 694 31648 745
rect 31918 739 31952 790
rect 31582 677 31648 694
rect 31582 643 31598 677
rect 31632 643 31648 677
rect 31582 631 31648 643
rect 31819 705 31952 739
rect 32007 730 32043 802
rect 32194 798 32208 832
rect 32242 821 32260 832
rect 32194 787 32210 798
rect 32244 787 32260 821
rect 31819 684 31853 705
rect 31991 701 32043 730
rect 31819 629 31853 650
rect 31889 637 31905 671
rect 31939 637 31955 671
rect 30640 550 30650 564
rect 27238 420 27272 454
rect 27238 368 27272 384
rect 28630 444 28762 480
rect 28934 490 28968 506
rect 29030 490 29064 506
rect 28968 454 28969 455
rect 28630 396 28666 444
rect 28934 420 28969 454
rect 28968 418 28969 420
rect 29030 420 29064 454
rect 28814 396 28934 418
rect 28630 384 28934 396
rect 28968 384 28970 418
rect 28630 382 28970 384
rect 28630 360 28850 382
rect 28934 368 28968 382
rect 29030 368 29064 384
rect 29126 490 29160 506
rect 30600 480 30650 550
rect 30950 540 30966 574
rect 31000 540 31016 574
rect 31230 566 31278 578
rect 31438 563 31467 597
rect 31501 563 31559 597
rect 31593 563 31651 597
rect 31685 563 31714 597
rect 31889 595 31955 637
rect 32025 667 32043 701
rect 31991 629 32043 667
rect 32194 737 32240 753
rect 32294 749 32340 869
rect 32478 1047 32512 1066
rect 32564 1057 32769 1066
rect 32803 1089 33012 1091
rect 32803 1057 32888 1089
rect 32564 1055 32888 1057
rect 32922 1066 33012 1089
rect 33252 1066 33286 1424
rect 34196 1398 34230 1609
rect 34427 1306 34461 1609
rect 34512 1390 34546 2004
rect 34712 2002 34778 2004
rect 35029 2009 35045 2043
rect 35079 2009 35095 2043
rect 35029 1975 35095 2009
rect 34584 1943 34618 1962
rect 34584 1875 34618 1877
rect 34584 1839 34618 1841
rect 34584 1754 34618 1773
rect 34680 1943 34714 1962
rect 34680 1875 34714 1877
rect 34680 1839 34714 1841
rect 34680 1754 34714 1773
rect 34776 1943 34810 1962
rect 35029 1941 35045 1975
rect 35079 1959 35095 1975
rect 35201 2111 35267 2153
rect 35235 2077 35267 2111
rect 35201 2043 35267 2077
rect 35235 2009 35267 2043
rect 35201 1975 35267 2009
rect 35079 1941 35165 1959
rect 35029 1925 35165 1941
rect 35235 1941 35267 1975
rect 35201 1925 35267 1941
rect 36103 2111 36169 2116
rect 36103 2077 36119 2111
rect 36153 2077 36169 2111
rect 36103 2043 36169 2077
rect 36103 2009 36119 2043
rect 36153 2009 36169 2043
rect 36103 1975 36169 2009
rect 36103 1941 36119 1975
rect 36153 1959 36169 1975
rect 36275 2111 36341 2153
rect 36309 2077 36341 2111
rect 36508 2147 36790 2153
rect 36508 2113 36547 2147
rect 36581 2145 36790 2147
rect 36581 2113 36666 2145
rect 36508 2111 36666 2113
rect 36700 2111 36790 2145
rect 36508 2078 36790 2111
rect 36917 2111 36983 2116
rect 36275 2043 36341 2077
rect 36309 2009 36341 2043
rect 36917 2077 36933 2111
rect 36967 2077 36983 2111
rect 36917 2043 36983 2077
rect 36275 1975 36341 2009
rect 36153 1941 36239 1959
rect 36103 1925 36239 1941
rect 36309 1941 36341 1975
rect 36275 1925 36341 1941
rect 36400 2039 36666 2040
rect 36400 2005 36616 2039
rect 36650 2005 36666 2039
rect 36400 2004 36666 2005
rect 34776 1875 34810 1877
rect 35027 1882 35097 1891
rect 35027 1848 35043 1882
rect 35077 1875 35097 1882
rect 35027 1841 35047 1848
rect 35081 1841 35097 1875
rect 34776 1839 34810 1841
rect 35131 1805 35165 1925
rect 35199 1882 35269 1891
rect 35199 1875 35217 1882
rect 35199 1841 35215 1875
rect 35251 1848 35269 1882
rect 35249 1841 35269 1848
rect 36101 1884 36171 1891
rect 36101 1850 36119 1884
rect 36153 1875 36171 1884
rect 36101 1841 36121 1850
rect 36155 1841 36171 1875
rect 36205 1805 36239 1925
rect 36273 1880 36343 1891
rect 36273 1875 36292 1880
rect 36273 1841 36289 1875
rect 36326 1846 36343 1880
rect 36323 1841 36343 1846
rect 34776 1754 34810 1773
rect 35031 1789 35079 1805
rect 35031 1755 35045 1789
rect 35031 1721 35079 1755
rect 34616 1677 34632 1711
rect 34666 1677 34682 1711
rect 35031 1687 35045 1721
rect 35031 1643 35079 1687
rect 35113 1789 35179 1805
rect 35113 1755 35129 1789
rect 35163 1759 35179 1789
rect 35113 1725 35131 1755
rect 35165 1725 35179 1759
rect 35113 1721 35179 1725
rect 35113 1687 35129 1721
rect 35163 1687 35179 1721
rect 35113 1677 35179 1687
rect 35213 1789 35267 1805
rect 35247 1755 35267 1789
rect 35213 1721 35267 1755
rect 35247 1687 35267 1721
rect 35213 1643 35267 1687
rect 36105 1789 36153 1805
rect 36105 1755 36119 1789
rect 36105 1721 36153 1755
rect 36105 1687 36119 1721
rect 36105 1643 36153 1687
rect 36187 1789 36253 1805
rect 36187 1764 36203 1789
rect 36187 1730 36201 1764
rect 36237 1755 36253 1789
rect 36235 1730 36253 1755
rect 36187 1721 36253 1730
rect 36187 1687 36203 1721
rect 36237 1687 36253 1721
rect 36187 1677 36253 1687
rect 36287 1789 36341 1805
rect 36321 1755 36341 1789
rect 36287 1721 36341 1755
rect 36321 1687 36341 1721
rect 36287 1643 36341 1687
rect 34728 1596 34744 1630
rect 34778 1596 34794 1630
rect 35010 1609 35039 1643
rect 35073 1609 35131 1643
rect 35165 1609 35223 1643
rect 35257 1609 35286 1643
rect 36084 1609 36113 1643
rect 36147 1609 36205 1643
rect 36239 1609 36297 1643
rect 36331 1609 36360 1643
rect 34600 1546 34634 1562
rect 34600 1476 34634 1510
rect 34600 1424 34634 1440
rect 34696 1546 34730 1562
rect 34696 1476 34730 1510
rect 34696 1424 34730 1440
rect 34792 1546 34826 1562
rect 34792 1476 34826 1510
rect 34826 1440 35174 1464
rect 34792 1424 35174 1440
rect 34512 1356 34648 1390
rect 34682 1356 34698 1390
rect 34427 1286 34822 1306
rect 34427 1281 34689 1286
rect 34427 1272 34568 1281
rect 34552 1247 34568 1272
rect 34602 1252 34689 1281
rect 34723 1262 34822 1286
rect 34994 1264 35040 1266
rect 34994 1262 34998 1264
rect 34723 1252 34998 1262
rect 34602 1247 34998 1252
rect 34552 1230 34998 1247
rect 35032 1230 35040 1264
rect 34552 1228 35040 1230
rect 34994 1222 35040 1228
rect 33326 1107 33355 1141
rect 33389 1107 33447 1141
rect 33481 1107 33539 1141
rect 33573 1107 33602 1141
rect 32922 1055 33158 1066
rect 32564 1047 33158 1055
rect 32564 1022 32566 1047
rect 32478 979 32512 981
rect 32478 943 32512 945
rect 32478 858 32512 877
rect 32600 1022 33124 1047
rect 33210 1047 33286 1066
rect 33210 1026 33212 1047
rect 32566 979 32600 981
rect 32822 949 32838 983
rect 32872 949 32888 983
rect 33124 979 33158 981
rect 32566 943 32600 945
rect 33124 943 33158 945
rect 32566 858 32600 877
rect 32694 887 32728 906
rect 32694 819 32728 821
rect 32506 781 32522 815
rect 32556 781 32572 815
rect 32694 783 32728 785
rect 32194 703 32206 737
rect 32194 669 32240 703
rect 32194 635 32206 669
rect 31784 561 31813 595
rect 31847 561 31905 595
rect 31939 561 31997 595
rect 32031 561 32060 595
rect 32194 589 32240 635
rect 32274 737 32340 749
rect 32274 703 32290 737
rect 32324 703 32340 737
rect 32274 690 32340 703
rect 32694 698 32728 717
rect 32790 887 32824 906
rect 32790 819 32824 821
rect 32790 783 32824 785
rect 32790 698 32824 717
rect 32886 887 32920 906
rect 33124 858 33158 877
rect 33246 1026 33286 1047
rect 33394 1065 33436 1107
rect 33672 1105 33701 1139
rect 33735 1105 33793 1139
rect 33827 1105 33885 1139
rect 33919 1105 33948 1139
rect 34093 1133 34127 1140
rect 33394 1031 33402 1065
rect 33212 979 33246 981
rect 33212 943 33246 945
rect 33394 997 33436 1031
rect 33394 963 33402 997
rect 33394 929 33436 963
rect 33394 895 33402 929
rect 33394 879 33436 895
rect 33470 1065 33536 1073
rect 33470 1031 33486 1065
rect 33520 1031 33536 1065
rect 33470 997 33536 1031
rect 33470 963 33486 997
rect 33520 963 33536 997
rect 33470 929 33536 963
rect 33470 895 33486 929
rect 33520 895 33536 929
rect 33470 877 33536 895
rect 33705 1055 33741 1071
rect 33705 1021 33707 1055
rect 33705 987 33741 1021
rect 33705 953 33707 987
rect 33777 1055 33843 1105
rect 34018 1099 34047 1133
rect 34081 1099 34139 1133
rect 34173 1099 34231 1133
rect 34265 1099 34294 1133
rect 34394 1109 34410 1143
rect 34444 1109 34460 1143
rect 34618 1130 34732 1132
rect 33777 1021 33793 1055
rect 33827 1021 33843 1055
rect 33777 987 33843 1021
rect 33777 953 33793 987
rect 33827 953 33843 987
rect 33877 1055 33931 1071
rect 33877 1021 33879 1055
rect 33913 1021 33931 1055
rect 33877 974 33931 1021
rect 33705 919 33741 953
rect 33877 940 33879 974
rect 33913 940 33931 974
rect 33705 885 33840 919
rect 33877 890 33931 940
rect 33212 858 33246 877
rect 32886 819 32920 821
rect 33298 843 33442 844
rect 33298 829 33456 843
rect 32886 783 32920 785
rect 33152 816 33218 818
rect 33298 816 33406 829
rect 33152 815 33406 816
rect 33152 781 33168 815
rect 33202 802 33406 815
rect 33202 782 33338 802
rect 33390 795 33406 802
rect 33440 795 33456 829
rect 33202 781 33218 782
rect 33390 745 33436 761
rect 33490 757 33536 877
rect 33806 856 33840 885
rect 33693 827 33761 849
rect 33693 826 33709 827
rect 33693 792 33707 826
rect 33743 793 33761 827
rect 33741 792 33761 793
rect 33693 775 33761 792
rect 33806 840 33861 856
rect 33806 806 33827 840
rect 33806 790 33861 806
rect 33895 840 33931 890
rect 34086 1057 34128 1099
rect 34618 1091 34900 1130
rect 35040 1109 35056 1143
rect 35090 1109 35106 1143
rect 34618 1066 34657 1091
rect 34086 1023 34094 1057
rect 34086 989 34128 1023
rect 34086 955 34094 989
rect 34086 921 34128 955
rect 34086 887 34094 921
rect 34086 871 34128 887
rect 34162 1057 34228 1065
rect 34162 1023 34178 1057
rect 34212 1023 34228 1057
rect 34162 989 34228 1023
rect 34162 955 34178 989
rect 34212 955 34228 989
rect 34162 921 34228 955
rect 34162 887 34178 921
rect 34212 887 34228 921
rect 34162 869 34228 887
rect 33895 838 33936 840
rect 33895 804 33900 838
rect 33934 804 33936 838
rect 33895 802 33936 804
rect 34082 832 34148 835
rect 32920 717 33166 734
rect 32886 700 33166 717
rect 32886 698 32920 700
rect 32274 669 32616 690
rect 32274 635 32290 669
rect 32324 658 32616 669
rect 32324 655 32792 658
rect 32324 654 32742 655
rect 32324 635 32346 654
rect 32274 630 32346 635
rect 32274 623 32340 630
rect 32580 622 32742 654
rect 32726 621 32742 622
rect 32776 621 32792 655
rect 33118 612 33166 700
rect 32130 555 32159 589
rect 32193 555 32251 589
rect 32285 555 32343 589
rect 32377 555 32406 589
rect 32488 584 32534 594
rect 32488 550 32494 584
rect 32528 564 32534 584
rect 33118 578 33126 612
rect 33160 578 33166 612
rect 33390 711 33402 745
rect 33390 677 33436 711
rect 33390 643 33402 677
rect 33390 597 33436 643
rect 33470 745 33536 757
rect 33470 694 33486 745
rect 33520 694 33536 745
rect 33806 739 33840 790
rect 33470 677 33536 694
rect 33470 643 33486 677
rect 33520 643 33536 677
rect 33470 631 33536 643
rect 33707 705 33840 739
rect 33895 730 33931 802
rect 34082 798 34096 832
rect 34130 821 34148 832
rect 34082 787 34098 798
rect 34132 787 34148 821
rect 33707 684 33741 705
rect 33879 701 33931 730
rect 33707 629 33741 650
rect 33777 637 33793 671
rect 33827 637 33843 671
rect 32528 550 32538 564
rect 29126 420 29160 454
rect 29126 368 29160 384
rect 30518 444 30650 480
rect 30822 490 30856 506
rect 30918 490 30952 506
rect 30856 454 30857 455
rect 30518 396 30554 444
rect 30822 420 30857 454
rect 30856 418 30857 420
rect 30918 420 30952 454
rect 30702 396 30822 418
rect 30518 384 30822 396
rect 30856 384 30858 418
rect 30518 382 30858 384
rect 30518 360 30738 382
rect 30822 368 30856 382
rect 30918 368 30952 384
rect 31014 490 31048 506
rect 32488 480 32538 550
rect 32838 540 32854 574
rect 32888 540 32904 574
rect 33118 566 33166 578
rect 33326 563 33355 597
rect 33389 563 33447 597
rect 33481 563 33539 597
rect 33573 563 33602 597
rect 33777 595 33843 637
rect 33913 667 33931 701
rect 33879 629 33931 667
rect 34082 737 34128 753
rect 34182 749 34228 869
rect 34366 1047 34400 1066
rect 34452 1057 34657 1066
rect 34691 1089 34900 1091
rect 34691 1057 34776 1089
rect 34452 1055 34776 1057
rect 34810 1066 34900 1089
rect 35140 1066 35174 1424
rect 36084 1398 36118 1609
rect 36315 1306 36349 1609
rect 36400 1390 36434 2004
rect 36600 2002 36666 2004
rect 36917 2009 36933 2043
rect 36967 2009 36983 2043
rect 36917 1975 36983 2009
rect 36472 1943 36506 1962
rect 36472 1875 36506 1877
rect 36472 1839 36506 1841
rect 36472 1754 36506 1773
rect 36568 1943 36602 1962
rect 36568 1875 36602 1877
rect 36568 1839 36602 1841
rect 36568 1754 36602 1773
rect 36664 1943 36698 1962
rect 36917 1941 36933 1975
rect 36967 1959 36983 1975
rect 37089 2111 37155 2153
rect 37123 2077 37155 2111
rect 37089 2043 37155 2077
rect 37123 2009 37155 2043
rect 37089 1975 37155 2009
rect 36967 1941 37053 1959
rect 36917 1925 37053 1941
rect 37123 1941 37155 1975
rect 37089 1925 37155 1941
rect 37991 2111 38057 2116
rect 37991 2077 38007 2111
rect 38041 2077 38057 2111
rect 37991 2043 38057 2077
rect 37991 2009 38007 2043
rect 38041 2009 38057 2043
rect 37991 1975 38057 2009
rect 37991 1941 38007 1975
rect 38041 1959 38057 1975
rect 38163 2111 38229 2153
rect 38197 2077 38229 2111
rect 38396 2147 38678 2153
rect 38396 2113 38435 2147
rect 38469 2145 38678 2147
rect 38469 2113 38554 2145
rect 38396 2111 38554 2113
rect 38588 2111 38678 2145
rect 38396 2078 38678 2111
rect 38805 2111 38871 2116
rect 38163 2043 38229 2077
rect 38197 2009 38229 2043
rect 38805 2077 38821 2111
rect 38855 2077 38871 2111
rect 38805 2043 38871 2077
rect 38163 1975 38229 2009
rect 38041 1941 38127 1959
rect 37991 1925 38127 1941
rect 38197 1941 38229 1975
rect 38163 1925 38229 1941
rect 38288 2039 38554 2040
rect 38288 2005 38504 2039
rect 38538 2005 38554 2039
rect 38288 2004 38554 2005
rect 36664 1875 36698 1877
rect 36915 1882 36985 1891
rect 36915 1848 36931 1882
rect 36965 1875 36985 1882
rect 36915 1841 36935 1848
rect 36969 1841 36985 1875
rect 36664 1839 36698 1841
rect 37019 1805 37053 1925
rect 37087 1882 37157 1891
rect 37087 1875 37105 1882
rect 37087 1841 37103 1875
rect 37139 1848 37157 1882
rect 37137 1841 37157 1848
rect 37989 1884 38059 1891
rect 37989 1850 38007 1884
rect 38041 1875 38059 1884
rect 37989 1841 38009 1850
rect 38043 1841 38059 1875
rect 38093 1805 38127 1925
rect 38161 1880 38231 1891
rect 38161 1875 38180 1880
rect 38161 1841 38177 1875
rect 38214 1846 38231 1880
rect 38211 1841 38231 1846
rect 36664 1754 36698 1773
rect 36919 1789 36967 1805
rect 36919 1755 36933 1789
rect 36919 1721 36967 1755
rect 36504 1677 36520 1711
rect 36554 1677 36570 1711
rect 36919 1687 36933 1721
rect 36919 1643 36967 1687
rect 37001 1789 37067 1805
rect 37001 1755 37017 1789
rect 37051 1759 37067 1789
rect 37001 1725 37019 1755
rect 37053 1725 37067 1759
rect 37001 1721 37067 1725
rect 37001 1687 37017 1721
rect 37051 1687 37067 1721
rect 37001 1677 37067 1687
rect 37101 1789 37155 1805
rect 37135 1755 37155 1789
rect 37101 1721 37155 1755
rect 37135 1687 37155 1721
rect 37101 1643 37155 1687
rect 37993 1789 38041 1805
rect 37993 1755 38007 1789
rect 37993 1721 38041 1755
rect 37993 1687 38007 1721
rect 37993 1643 38041 1687
rect 38075 1789 38141 1805
rect 38075 1764 38091 1789
rect 38075 1730 38089 1764
rect 38125 1755 38141 1789
rect 38123 1730 38141 1755
rect 38075 1721 38141 1730
rect 38075 1687 38091 1721
rect 38125 1687 38141 1721
rect 38075 1677 38141 1687
rect 38175 1789 38229 1805
rect 38209 1755 38229 1789
rect 38175 1721 38229 1755
rect 38209 1687 38229 1721
rect 38175 1643 38229 1687
rect 36616 1596 36632 1630
rect 36666 1596 36682 1630
rect 36898 1609 36927 1643
rect 36961 1609 37019 1643
rect 37053 1609 37111 1643
rect 37145 1609 37174 1643
rect 37972 1609 38001 1643
rect 38035 1609 38093 1643
rect 38127 1609 38185 1643
rect 38219 1609 38248 1643
rect 36488 1546 36522 1562
rect 36488 1476 36522 1510
rect 36488 1424 36522 1440
rect 36584 1546 36618 1562
rect 36584 1476 36618 1510
rect 36584 1424 36618 1440
rect 36680 1546 36714 1562
rect 36680 1476 36714 1510
rect 36714 1440 37062 1464
rect 36680 1424 37062 1440
rect 36400 1356 36536 1390
rect 36570 1356 36586 1390
rect 36315 1286 36710 1306
rect 36315 1281 36577 1286
rect 36315 1272 36456 1281
rect 36440 1247 36456 1272
rect 36490 1252 36577 1281
rect 36611 1262 36710 1286
rect 36882 1264 36928 1266
rect 36882 1262 36886 1264
rect 36611 1252 36886 1262
rect 36490 1247 36886 1252
rect 36440 1230 36886 1247
rect 36920 1230 36928 1264
rect 36440 1228 36928 1230
rect 36882 1222 36928 1228
rect 35214 1107 35243 1141
rect 35277 1107 35335 1141
rect 35369 1107 35427 1141
rect 35461 1107 35490 1141
rect 34810 1055 35046 1066
rect 34452 1047 35046 1055
rect 34452 1022 34454 1047
rect 34366 979 34400 981
rect 34366 943 34400 945
rect 34366 858 34400 877
rect 34488 1022 35012 1047
rect 35098 1047 35174 1066
rect 35098 1026 35100 1047
rect 34454 979 34488 981
rect 34710 949 34726 983
rect 34760 949 34776 983
rect 35012 979 35046 981
rect 34454 943 34488 945
rect 35012 943 35046 945
rect 34454 858 34488 877
rect 34582 887 34616 906
rect 34582 819 34616 821
rect 34394 781 34410 815
rect 34444 781 34460 815
rect 34582 783 34616 785
rect 34082 703 34094 737
rect 34082 669 34128 703
rect 34082 635 34094 669
rect 33672 561 33701 595
rect 33735 561 33793 595
rect 33827 561 33885 595
rect 33919 561 33948 595
rect 34082 589 34128 635
rect 34162 737 34228 749
rect 34162 703 34178 737
rect 34212 703 34228 737
rect 34162 690 34228 703
rect 34582 698 34616 717
rect 34678 887 34712 906
rect 34678 819 34712 821
rect 34678 783 34712 785
rect 34678 698 34712 717
rect 34774 887 34808 906
rect 35012 858 35046 877
rect 35134 1026 35174 1047
rect 35282 1065 35324 1107
rect 35560 1105 35589 1139
rect 35623 1105 35681 1139
rect 35715 1105 35773 1139
rect 35807 1105 35836 1139
rect 35981 1133 36015 1140
rect 35282 1031 35290 1065
rect 35100 979 35134 981
rect 35100 943 35134 945
rect 35282 997 35324 1031
rect 35282 963 35290 997
rect 35282 929 35324 963
rect 35282 895 35290 929
rect 35282 879 35324 895
rect 35358 1065 35424 1073
rect 35358 1031 35374 1065
rect 35408 1031 35424 1065
rect 35358 997 35424 1031
rect 35358 963 35374 997
rect 35408 963 35424 997
rect 35358 929 35424 963
rect 35358 895 35374 929
rect 35408 895 35424 929
rect 35358 877 35424 895
rect 35593 1055 35629 1071
rect 35593 1021 35595 1055
rect 35593 987 35629 1021
rect 35593 953 35595 987
rect 35665 1055 35731 1105
rect 35906 1099 35935 1133
rect 35969 1099 36027 1133
rect 36061 1099 36119 1133
rect 36153 1099 36182 1133
rect 36282 1109 36298 1143
rect 36332 1109 36348 1143
rect 36506 1130 36620 1132
rect 35665 1021 35681 1055
rect 35715 1021 35731 1055
rect 35665 987 35731 1021
rect 35665 953 35681 987
rect 35715 953 35731 987
rect 35765 1055 35819 1071
rect 35765 1021 35767 1055
rect 35801 1021 35819 1055
rect 35765 974 35819 1021
rect 35593 919 35629 953
rect 35765 940 35767 974
rect 35801 940 35819 974
rect 35593 885 35728 919
rect 35765 890 35819 940
rect 35100 858 35134 877
rect 34774 819 34808 821
rect 35186 843 35330 844
rect 35186 829 35344 843
rect 34774 783 34808 785
rect 35040 816 35106 818
rect 35186 816 35294 829
rect 35040 815 35294 816
rect 35040 781 35056 815
rect 35090 802 35294 815
rect 35090 782 35226 802
rect 35278 795 35294 802
rect 35328 795 35344 829
rect 35090 781 35106 782
rect 35278 745 35324 761
rect 35378 757 35424 877
rect 35694 856 35728 885
rect 35581 827 35649 849
rect 35581 826 35597 827
rect 35581 792 35595 826
rect 35631 793 35649 827
rect 35629 792 35649 793
rect 35581 775 35649 792
rect 35694 840 35749 856
rect 35694 806 35715 840
rect 35694 790 35749 806
rect 35783 840 35819 890
rect 35974 1057 36016 1099
rect 36506 1091 36788 1130
rect 36928 1109 36944 1143
rect 36978 1109 36994 1143
rect 36506 1066 36545 1091
rect 35974 1023 35982 1057
rect 35974 989 36016 1023
rect 35974 955 35982 989
rect 35974 921 36016 955
rect 35974 887 35982 921
rect 35974 871 36016 887
rect 36050 1057 36116 1065
rect 36050 1023 36066 1057
rect 36100 1023 36116 1057
rect 36050 989 36116 1023
rect 36050 955 36066 989
rect 36100 955 36116 989
rect 36050 921 36116 955
rect 36050 887 36066 921
rect 36100 887 36116 921
rect 36050 869 36116 887
rect 35783 838 35824 840
rect 35783 804 35788 838
rect 35822 804 35824 838
rect 35783 802 35824 804
rect 35970 832 36036 835
rect 34808 717 35054 734
rect 34774 700 35054 717
rect 34774 698 34808 700
rect 34162 669 34504 690
rect 34162 635 34178 669
rect 34212 658 34504 669
rect 34212 655 34680 658
rect 34212 654 34630 655
rect 34212 635 34234 654
rect 34162 630 34234 635
rect 34162 623 34228 630
rect 34468 622 34630 654
rect 34614 621 34630 622
rect 34664 621 34680 655
rect 35006 612 35054 700
rect 34018 555 34047 589
rect 34081 555 34139 589
rect 34173 555 34231 589
rect 34265 555 34294 589
rect 34376 584 34422 594
rect 34376 550 34382 584
rect 34416 564 34422 584
rect 35006 578 35014 612
rect 35048 578 35054 612
rect 35278 711 35290 745
rect 35278 677 35324 711
rect 35278 643 35290 677
rect 35278 597 35324 643
rect 35358 745 35424 757
rect 35358 694 35374 745
rect 35408 694 35424 745
rect 35694 739 35728 790
rect 35358 677 35424 694
rect 35358 643 35374 677
rect 35408 643 35424 677
rect 35358 631 35424 643
rect 35595 705 35728 739
rect 35783 730 35819 802
rect 35970 798 35984 832
rect 36018 821 36036 832
rect 35970 787 35986 798
rect 36020 787 36036 821
rect 35595 684 35629 705
rect 35767 701 35819 730
rect 35595 629 35629 650
rect 35665 637 35681 671
rect 35715 637 35731 671
rect 34416 550 34426 564
rect 31014 420 31048 454
rect 31014 368 31048 384
rect 32406 444 32538 480
rect 32710 490 32744 506
rect 32806 490 32840 506
rect 32744 454 32745 455
rect 32406 396 32442 444
rect 32710 420 32745 454
rect 32744 418 32745 420
rect 32806 420 32840 454
rect 32590 396 32710 418
rect 32406 384 32710 396
rect 32744 384 32746 418
rect 32406 382 32746 384
rect 32406 360 32626 382
rect 32710 368 32744 382
rect 32806 368 32840 384
rect 32902 490 32936 506
rect 34376 480 34426 550
rect 34726 540 34742 574
rect 34776 540 34792 574
rect 35006 566 35054 578
rect 35214 563 35243 597
rect 35277 563 35335 597
rect 35369 563 35427 597
rect 35461 563 35490 597
rect 35665 595 35731 637
rect 35801 667 35819 701
rect 35767 629 35819 667
rect 35970 737 36016 753
rect 36070 749 36116 869
rect 36254 1047 36288 1066
rect 36340 1057 36545 1066
rect 36579 1089 36788 1091
rect 36579 1057 36664 1089
rect 36340 1055 36664 1057
rect 36698 1066 36788 1089
rect 37028 1066 37062 1424
rect 37972 1398 38006 1609
rect 38203 1306 38237 1609
rect 38288 1390 38322 2004
rect 38488 2002 38554 2004
rect 38805 2009 38821 2043
rect 38855 2009 38871 2043
rect 38805 1975 38871 2009
rect 38360 1943 38394 1962
rect 38360 1875 38394 1877
rect 38360 1839 38394 1841
rect 38360 1754 38394 1773
rect 38456 1943 38490 1962
rect 38456 1875 38490 1877
rect 38456 1839 38490 1841
rect 38456 1754 38490 1773
rect 38552 1943 38586 1962
rect 38805 1941 38821 1975
rect 38855 1959 38871 1975
rect 38977 2111 39043 2153
rect 39011 2077 39043 2111
rect 38977 2043 39043 2077
rect 39011 2009 39043 2043
rect 38977 1975 39043 2009
rect 38855 1941 38941 1959
rect 38805 1925 38941 1941
rect 39011 1941 39043 1975
rect 38977 1925 39043 1941
rect 39879 2111 39945 2116
rect 39879 2077 39895 2111
rect 39929 2077 39945 2111
rect 39879 2043 39945 2077
rect 39879 2009 39895 2043
rect 39929 2009 39945 2043
rect 39879 1975 39945 2009
rect 39879 1941 39895 1975
rect 39929 1959 39945 1975
rect 40051 2111 40117 2153
rect 40085 2077 40117 2111
rect 40284 2147 40566 2153
rect 40284 2113 40323 2147
rect 40357 2145 40566 2147
rect 40357 2113 40442 2145
rect 40284 2111 40442 2113
rect 40476 2111 40566 2145
rect 40284 2078 40566 2111
rect 40693 2111 40759 2116
rect 40051 2043 40117 2077
rect 40085 2009 40117 2043
rect 40693 2077 40709 2111
rect 40743 2077 40759 2111
rect 40693 2043 40759 2077
rect 40051 1975 40117 2009
rect 39929 1941 40015 1959
rect 39879 1925 40015 1941
rect 40085 1941 40117 1975
rect 40051 1925 40117 1941
rect 40176 2039 40442 2040
rect 40176 2005 40392 2039
rect 40426 2005 40442 2039
rect 40176 2004 40442 2005
rect 38552 1875 38586 1877
rect 38803 1882 38873 1891
rect 38803 1848 38819 1882
rect 38853 1875 38873 1882
rect 38803 1841 38823 1848
rect 38857 1841 38873 1875
rect 38552 1839 38586 1841
rect 38907 1805 38941 1925
rect 38975 1882 39045 1891
rect 38975 1875 38993 1882
rect 38975 1841 38991 1875
rect 39027 1848 39045 1882
rect 39025 1841 39045 1848
rect 39877 1884 39947 1891
rect 39877 1850 39895 1884
rect 39929 1875 39947 1884
rect 39877 1841 39897 1850
rect 39931 1841 39947 1875
rect 39981 1805 40015 1925
rect 40049 1880 40119 1891
rect 40049 1875 40068 1880
rect 40049 1841 40065 1875
rect 40102 1846 40119 1880
rect 40099 1841 40119 1846
rect 38552 1754 38586 1773
rect 38807 1789 38855 1805
rect 38807 1755 38821 1789
rect 38807 1721 38855 1755
rect 38392 1677 38408 1711
rect 38442 1677 38458 1711
rect 38807 1687 38821 1721
rect 38807 1643 38855 1687
rect 38889 1789 38955 1805
rect 38889 1755 38905 1789
rect 38939 1759 38955 1789
rect 38889 1725 38907 1755
rect 38941 1725 38955 1759
rect 38889 1721 38955 1725
rect 38889 1687 38905 1721
rect 38939 1687 38955 1721
rect 38889 1677 38955 1687
rect 38989 1789 39043 1805
rect 39023 1755 39043 1789
rect 38989 1721 39043 1755
rect 39023 1687 39043 1721
rect 38989 1643 39043 1687
rect 39881 1789 39929 1805
rect 39881 1755 39895 1789
rect 39881 1721 39929 1755
rect 39881 1687 39895 1721
rect 39881 1643 39929 1687
rect 39963 1789 40029 1805
rect 39963 1764 39979 1789
rect 39963 1730 39977 1764
rect 40013 1755 40029 1789
rect 40011 1730 40029 1755
rect 39963 1721 40029 1730
rect 39963 1687 39979 1721
rect 40013 1687 40029 1721
rect 39963 1677 40029 1687
rect 40063 1789 40117 1805
rect 40097 1755 40117 1789
rect 40063 1721 40117 1755
rect 40097 1687 40117 1721
rect 40063 1643 40117 1687
rect 38504 1596 38520 1630
rect 38554 1596 38570 1630
rect 38786 1609 38815 1643
rect 38849 1609 38907 1643
rect 38941 1609 38999 1643
rect 39033 1609 39062 1643
rect 39860 1609 39889 1643
rect 39923 1609 39981 1643
rect 40015 1609 40073 1643
rect 40107 1609 40136 1643
rect 38376 1546 38410 1562
rect 38376 1476 38410 1510
rect 38376 1424 38410 1440
rect 38472 1546 38506 1562
rect 38472 1476 38506 1510
rect 38472 1424 38506 1440
rect 38568 1546 38602 1562
rect 38568 1476 38602 1510
rect 38602 1440 38950 1464
rect 38568 1424 38950 1440
rect 38288 1356 38424 1390
rect 38458 1356 38474 1390
rect 38203 1286 38598 1306
rect 38203 1281 38465 1286
rect 38203 1272 38344 1281
rect 38328 1247 38344 1272
rect 38378 1252 38465 1281
rect 38499 1262 38598 1286
rect 38770 1264 38816 1266
rect 38770 1262 38774 1264
rect 38499 1252 38774 1262
rect 38378 1247 38774 1252
rect 38328 1230 38774 1247
rect 38808 1230 38816 1264
rect 38328 1228 38816 1230
rect 38770 1222 38816 1228
rect 37102 1107 37131 1141
rect 37165 1107 37223 1141
rect 37257 1107 37315 1141
rect 37349 1107 37378 1141
rect 36698 1055 36934 1066
rect 36340 1047 36934 1055
rect 36340 1022 36342 1047
rect 36254 979 36288 981
rect 36254 943 36288 945
rect 36254 858 36288 877
rect 36376 1022 36900 1047
rect 36986 1047 37062 1066
rect 36986 1026 36988 1047
rect 36342 979 36376 981
rect 36598 949 36614 983
rect 36648 949 36664 983
rect 36900 979 36934 981
rect 36342 943 36376 945
rect 36900 943 36934 945
rect 36342 858 36376 877
rect 36470 887 36504 906
rect 36470 819 36504 821
rect 36282 781 36298 815
rect 36332 781 36348 815
rect 36470 783 36504 785
rect 35970 703 35982 737
rect 35970 669 36016 703
rect 35970 635 35982 669
rect 35560 561 35589 595
rect 35623 561 35681 595
rect 35715 561 35773 595
rect 35807 561 35836 595
rect 35970 589 36016 635
rect 36050 737 36116 749
rect 36050 703 36066 737
rect 36100 703 36116 737
rect 36050 690 36116 703
rect 36470 698 36504 717
rect 36566 887 36600 906
rect 36566 819 36600 821
rect 36566 783 36600 785
rect 36566 698 36600 717
rect 36662 887 36696 906
rect 36900 858 36934 877
rect 37022 1026 37062 1047
rect 37170 1065 37212 1107
rect 37448 1105 37477 1139
rect 37511 1105 37569 1139
rect 37603 1105 37661 1139
rect 37695 1105 37724 1139
rect 37869 1133 37903 1140
rect 37170 1031 37178 1065
rect 36988 979 37022 981
rect 36988 943 37022 945
rect 37170 997 37212 1031
rect 37170 963 37178 997
rect 37170 929 37212 963
rect 37170 895 37178 929
rect 37170 879 37212 895
rect 37246 1065 37312 1073
rect 37246 1031 37262 1065
rect 37296 1031 37312 1065
rect 37246 997 37312 1031
rect 37246 963 37262 997
rect 37296 963 37312 997
rect 37246 929 37312 963
rect 37246 895 37262 929
rect 37296 895 37312 929
rect 37246 877 37312 895
rect 37481 1055 37517 1071
rect 37481 1021 37483 1055
rect 37481 987 37517 1021
rect 37481 953 37483 987
rect 37553 1055 37619 1105
rect 37794 1099 37823 1133
rect 37857 1099 37915 1133
rect 37949 1099 38007 1133
rect 38041 1099 38070 1133
rect 38170 1109 38186 1143
rect 38220 1109 38236 1143
rect 38394 1130 38508 1132
rect 37553 1021 37569 1055
rect 37603 1021 37619 1055
rect 37553 987 37619 1021
rect 37553 953 37569 987
rect 37603 953 37619 987
rect 37653 1055 37707 1071
rect 37653 1021 37655 1055
rect 37689 1021 37707 1055
rect 37653 974 37707 1021
rect 37481 919 37517 953
rect 37653 940 37655 974
rect 37689 940 37707 974
rect 37481 885 37616 919
rect 37653 890 37707 940
rect 36988 858 37022 877
rect 36662 819 36696 821
rect 37074 843 37218 844
rect 37074 829 37232 843
rect 36662 783 36696 785
rect 36928 816 36994 818
rect 37074 816 37182 829
rect 36928 815 37182 816
rect 36928 781 36944 815
rect 36978 802 37182 815
rect 36978 782 37114 802
rect 37166 795 37182 802
rect 37216 795 37232 829
rect 36978 781 36994 782
rect 37166 745 37212 761
rect 37266 757 37312 877
rect 37582 856 37616 885
rect 37469 827 37537 849
rect 37469 826 37485 827
rect 37469 792 37483 826
rect 37519 793 37537 827
rect 37517 792 37537 793
rect 37469 775 37537 792
rect 37582 840 37637 856
rect 37582 806 37603 840
rect 37582 790 37637 806
rect 37671 840 37707 890
rect 37862 1057 37904 1099
rect 38394 1091 38676 1130
rect 38816 1109 38832 1143
rect 38866 1109 38882 1143
rect 38394 1066 38433 1091
rect 37862 1023 37870 1057
rect 37862 989 37904 1023
rect 37862 955 37870 989
rect 37862 921 37904 955
rect 37862 887 37870 921
rect 37862 871 37904 887
rect 37938 1057 38004 1065
rect 37938 1023 37954 1057
rect 37988 1023 38004 1057
rect 37938 989 38004 1023
rect 37938 955 37954 989
rect 37988 955 38004 989
rect 37938 921 38004 955
rect 37938 887 37954 921
rect 37988 887 38004 921
rect 37938 869 38004 887
rect 37671 838 37712 840
rect 37671 804 37676 838
rect 37710 804 37712 838
rect 37671 802 37712 804
rect 37858 832 37924 835
rect 36696 717 36942 734
rect 36662 700 36942 717
rect 36662 698 36696 700
rect 36050 669 36392 690
rect 36050 635 36066 669
rect 36100 658 36392 669
rect 36100 655 36568 658
rect 36100 654 36518 655
rect 36100 635 36122 654
rect 36050 630 36122 635
rect 36050 623 36116 630
rect 36356 622 36518 654
rect 36502 621 36518 622
rect 36552 621 36568 655
rect 36894 612 36942 700
rect 35906 555 35935 589
rect 35969 555 36027 589
rect 36061 555 36119 589
rect 36153 555 36182 589
rect 36264 584 36310 594
rect 36264 550 36270 584
rect 36304 564 36310 584
rect 36894 578 36902 612
rect 36936 578 36942 612
rect 37166 711 37178 745
rect 37166 677 37212 711
rect 37166 643 37178 677
rect 37166 597 37212 643
rect 37246 745 37312 757
rect 37246 694 37262 745
rect 37296 694 37312 745
rect 37582 739 37616 790
rect 37246 677 37312 694
rect 37246 643 37262 677
rect 37296 643 37312 677
rect 37246 631 37312 643
rect 37483 705 37616 739
rect 37671 730 37707 802
rect 37858 798 37872 832
rect 37906 821 37924 832
rect 37858 787 37874 798
rect 37908 787 37924 821
rect 37483 684 37517 705
rect 37655 701 37707 730
rect 37483 629 37517 650
rect 37553 637 37569 671
rect 37603 637 37619 671
rect 36304 550 36314 564
rect 32902 420 32936 454
rect 32902 368 32936 384
rect 34294 444 34426 480
rect 34598 490 34632 506
rect 34694 490 34728 506
rect 34632 454 34633 455
rect 34294 396 34330 444
rect 34598 420 34633 454
rect 34632 418 34633 420
rect 34694 420 34728 454
rect 34478 396 34598 418
rect 34294 384 34598 396
rect 34632 384 34634 418
rect 34294 382 34634 384
rect 34294 360 34514 382
rect 34598 368 34632 382
rect 34694 368 34728 384
rect 34790 490 34824 506
rect 36264 480 36314 550
rect 36614 540 36630 574
rect 36664 540 36680 574
rect 36894 566 36942 578
rect 37102 563 37131 597
rect 37165 563 37223 597
rect 37257 563 37315 597
rect 37349 563 37378 597
rect 37553 595 37619 637
rect 37689 667 37707 701
rect 37655 629 37707 667
rect 37858 737 37904 753
rect 37958 749 38004 869
rect 38142 1047 38176 1066
rect 38228 1057 38433 1066
rect 38467 1089 38676 1091
rect 38467 1057 38552 1089
rect 38228 1055 38552 1057
rect 38586 1066 38676 1089
rect 38916 1066 38950 1424
rect 39860 1398 39894 1609
rect 40091 1306 40125 1609
rect 40176 1390 40210 2004
rect 40376 2002 40442 2004
rect 40693 2009 40709 2043
rect 40743 2009 40759 2043
rect 40693 1975 40759 2009
rect 40248 1943 40282 1962
rect 40248 1875 40282 1877
rect 40248 1839 40282 1841
rect 40248 1754 40282 1773
rect 40344 1943 40378 1962
rect 40344 1875 40378 1877
rect 40344 1839 40378 1841
rect 40344 1754 40378 1773
rect 40440 1943 40474 1962
rect 40693 1941 40709 1975
rect 40743 1959 40759 1975
rect 40865 2111 40931 2153
rect 40899 2077 40931 2111
rect 40865 2043 40931 2077
rect 40899 2009 40931 2043
rect 40865 1975 40931 2009
rect 40743 1941 40829 1959
rect 40693 1925 40829 1941
rect 40899 1941 40931 1975
rect 40865 1925 40931 1941
rect 41767 2111 41833 2116
rect 41767 2077 41783 2111
rect 41817 2077 41833 2111
rect 41767 2043 41833 2077
rect 41767 2009 41783 2043
rect 41817 2009 41833 2043
rect 41767 1975 41833 2009
rect 41767 1941 41783 1975
rect 41817 1959 41833 1975
rect 41939 2111 42005 2153
rect 41973 2077 42005 2111
rect 42172 2147 42454 2153
rect 42172 2113 42211 2147
rect 42245 2145 42454 2147
rect 42245 2113 42330 2145
rect 42172 2111 42330 2113
rect 42364 2111 42454 2145
rect 42172 2078 42454 2111
rect 42581 2111 42647 2116
rect 41939 2043 42005 2077
rect 41973 2009 42005 2043
rect 42581 2077 42597 2111
rect 42631 2077 42647 2111
rect 42581 2043 42647 2077
rect 41939 1975 42005 2009
rect 41817 1941 41903 1959
rect 41767 1925 41903 1941
rect 41973 1941 42005 1975
rect 41939 1925 42005 1941
rect 42064 2039 42330 2040
rect 42064 2005 42280 2039
rect 42314 2005 42330 2039
rect 42064 2004 42330 2005
rect 40440 1875 40474 1877
rect 40691 1882 40761 1891
rect 40691 1848 40707 1882
rect 40741 1875 40761 1882
rect 40691 1841 40711 1848
rect 40745 1841 40761 1875
rect 40440 1839 40474 1841
rect 40795 1805 40829 1925
rect 40863 1882 40933 1891
rect 40863 1875 40881 1882
rect 40863 1841 40879 1875
rect 40915 1848 40933 1882
rect 40913 1841 40933 1848
rect 41765 1884 41835 1891
rect 41765 1850 41783 1884
rect 41817 1875 41835 1884
rect 41765 1841 41785 1850
rect 41819 1841 41835 1875
rect 41869 1805 41903 1925
rect 41937 1880 42007 1891
rect 41937 1875 41956 1880
rect 41937 1841 41953 1875
rect 41990 1846 42007 1880
rect 41987 1841 42007 1846
rect 40440 1754 40474 1773
rect 40695 1789 40743 1805
rect 40695 1755 40709 1789
rect 40695 1721 40743 1755
rect 40280 1677 40296 1711
rect 40330 1677 40346 1711
rect 40695 1687 40709 1721
rect 40695 1643 40743 1687
rect 40777 1789 40843 1805
rect 40777 1755 40793 1789
rect 40827 1759 40843 1789
rect 40777 1725 40795 1755
rect 40829 1725 40843 1759
rect 40777 1721 40843 1725
rect 40777 1687 40793 1721
rect 40827 1687 40843 1721
rect 40777 1677 40843 1687
rect 40877 1789 40931 1805
rect 40911 1755 40931 1789
rect 40877 1721 40931 1755
rect 40911 1687 40931 1721
rect 40877 1643 40931 1687
rect 41769 1789 41817 1805
rect 41769 1755 41783 1789
rect 41769 1721 41817 1755
rect 41769 1687 41783 1721
rect 41769 1643 41817 1687
rect 41851 1789 41917 1805
rect 41851 1764 41867 1789
rect 41851 1730 41865 1764
rect 41901 1755 41917 1789
rect 41899 1730 41917 1755
rect 41851 1721 41917 1730
rect 41851 1687 41867 1721
rect 41901 1687 41917 1721
rect 41851 1677 41917 1687
rect 41951 1789 42005 1805
rect 41985 1755 42005 1789
rect 41951 1721 42005 1755
rect 41985 1687 42005 1721
rect 41951 1643 42005 1687
rect 40392 1596 40408 1630
rect 40442 1596 40458 1630
rect 40674 1609 40703 1643
rect 40737 1609 40795 1643
rect 40829 1609 40887 1643
rect 40921 1609 40950 1643
rect 41748 1609 41777 1643
rect 41811 1609 41869 1643
rect 41903 1609 41961 1643
rect 41995 1609 42024 1643
rect 40264 1546 40298 1562
rect 40264 1476 40298 1510
rect 40264 1424 40298 1440
rect 40360 1546 40394 1562
rect 40360 1476 40394 1510
rect 40360 1424 40394 1440
rect 40456 1546 40490 1562
rect 40456 1476 40490 1510
rect 40490 1440 40838 1464
rect 40456 1424 40838 1440
rect 40176 1356 40312 1390
rect 40346 1356 40362 1390
rect 40091 1286 40486 1306
rect 40091 1281 40353 1286
rect 40091 1272 40232 1281
rect 40216 1247 40232 1272
rect 40266 1252 40353 1281
rect 40387 1262 40486 1286
rect 40658 1264 40704 1266
rect 40658 1262 40662 1264
rect 40387 1252 40662 1262
rect 40266 1247 40662 1252
rect 40216 1230 40662 1247
rect 40696 1230 40704 1264
rect 40216 1228 40704 1230
rect 40658 1222 40704 1228
rect 38990 1107 39019 1141
rect 39053 1107 39111 1141
rect 39145 1107 39203 1141
rect 39237 1107 39266 1141
rect 38586 1055 38822 1066
rect 38228 1047 38822 1055
rect 38228 1022 38230 1047
rect 38142 979 38176 981
rect 38142 943 38176 945
rect 38142 858 38176 877
rect 38264 1022 38788 1047
rect 38874 1047 38950 1066
rect 38874 1026 38876 1047
rect 38230 979 38264 981
rect 38486 949 38502 983
rect 38536 949 38552 983
rect 38788 979 38822 981
rect 38230 943 38264 945
rect 38788 943 38822 945
rect 38230 858 38264 877
rect 38358 887 38392 906
rect 38358 819 38392 821
rect 38170 781 38186 815
rect 38220 781 38236 815
rect 38358 783 38392 785
rect 37858 703 37870 737
rect 37858 669 37904 703
rect 37858 635 37870 669
rect 37448 561 37477 595
rect 37511 561 37569 595
rect 37603 561 37661 595
rect 37695 561 37724 595
rect 37858 589 37904 635
rect 37938 737 38004 749
rect 37938 703 37954 737
rect 37988 703 38004 737
rect 37938 690 38004 703
rect 38358 698 38392 717
rect 38454 887 38488 906
rect 38454 819 38488 821
rect 38454 783 38488 785
rect 38454 698 38488 717
rect 38550 887 38584 906
rect 38788 858 38822 877
rect 38910 1026 38950 1047
rect 39058 1065 39100 1107
rect 39336 1105 39365 1139
rect 39399 1105 39457 1139
rect 39491 1105 39549 1139
rect 39583 1105 39612 1139
rect 39757 1133 39791 1140
rect 39058 1031 39066 1065
rect 38876 979 38910 981
rect 38876 943 38910 945
rect 39058 997 39100 1031
rect 39058 963 39066 997
rect 39058 929 39100 963
rect 39058 895 39066 929
rect 39058 879 39100 895
rect 39134 1065 39200 1073
rect 39134 1031 39150 1065
rect 39184 1031 39200 1065
rect 39134 997 39200 1031
rect 39134 963 39150 997
rect 39184 963 39200 997
rect 39134 929 39200 963
rect 39134 895 39150 929
rect 39184 895 39200 929
rect 39134 877 39200 895
rect 39369 1055 39405 1071
rect 39369 1021 39371 1055
rect 39369 987 39405 1021
rect 39369 953 39371 987
rect 39441 1055 39507 1105
rect 39682 1099 39711 1133
rect 39745 1099 39803 1133
rect 39837 1099 39895 1133
rect 39929 1099 39958 1133
rect 40058 1109 40074 1143
rect 40108 1109 40124 1143
rect 40282 1130 40396 1132
rect 39441 1021 39457 1055
rect 39491 1021 39507 1055
rect 39441 987 39507 1021
rect 39441 953 39457 987
rect 39491 953 39507 987
rect 39541 1055 39595 1071
rect 39541 1021 39543 1055
rect 39577 1021 39595 1055
rect 39541 974 39595 1021
rect 39369 919 39405 953
rect 39541 940 39543 974
rect 39577 940 39595 974
rect 39369 885 39504 919
rect 39541 890 39595 940
rect 38876 858 38910 877
rect 38550 819 38584 821
rect 38962 843 39106 844
rect 38962 829 39120 843
rect 38550 783 38584 785
rect 38816 816 38882 818
rect 38962 816 39070 829
rect 38816 815 39070 816
rect 38816 781 38832 815
rect 38866 802 39070 815
rect 38866 782 39002 802
rect 39054 795 39070 802
rect 39104 795 39120 829
rect 38866 781 38882 782
rect 39054 745 39100 761
rect 39154 757 39200 877
rect 39470 856 39504 885
rect 39357 827 39425 849
rect 39357 826 39373 827
rect 39357 792 39371 826
rect 39407 793 39425 827
rect 39405 792 39425 793
rect 39357 775 39425 792
rect 39470 840 39525 856
rect 39470 806 39491 840
rect 39470 790 39525 806
rect 39559 840 39595 890
rect 39750 1057 39792 1099
rect 40282 1091 40564 1130
rect 40704 1109 40720 1143
rect 40754 1109 40770 1143
rect 40282 1066 40321 1091
rect 39750 1023 39758 1057
rect 39750 989 39792 1023
rect 39750 955 39758 989
rect 39750 921 39792 955
rect 39750 887 39758 921
rect 39750 871 39792 887
rect 39826 1057 39892 1065
rect 39826 1023 39842 1057
rect 39876 1023 39892 1057
rect 39826 989 39892 1023
rect 39826 955 39842 989
rect 39876 955 39892 989
rect 39826 921 39892 955
rect 39826 887 39842 921
rect 39876 887 39892 921
rect 39826 869 39892 887
rect 39559 838 39600 840
rect 39559 804 39564 838
rect 39598 804 39600 838
rect 39559 802 39600 804
rect 39746 832 39812 835
rect 38584 717 38830 734
rect 38550 700 38830 717
rect 38550 698 38584 700
rect 37938 669 38280 690
rect 37938 635 37954 669
rect 37988 658 38280 669
rect 37988 655 38456 658
rect 37988 654 38406 655
rect 37988 635 38010 654
rect 37938 630 38010 635
rect 37938 623 38004 630
rect 38244 622 38406 654
rect 38390 621 38406 622
rect 38440 621 38456 655
rect 38782 612 38830 700
rect 37794 555 37823 589
rect 37857 555 37915 589
rect 37949 555 38007 589
rect 38041 555 38070 589
rect 38152 584 38198 594
rect 38152 550 38158 584
rect 38192 564 38198 584
rect 38782 578 38790 612
rect 38824 578 38830 612
rect 39054 711 39066 745
rect 39054 677 39100 711
rect 39054 643 39066 677
rect 39054 597 39100 643
rect 39134 745 39200 757
rect 39134 694 39150 745
rect 39184 694 39200 745
rect 39470 739 39504 790
rect 39134 677 39200 694
rect 39134 643 39150 677
rect 39184 643 39200 677
rect 39134 631 39200 643
rect 39371 705 39504 739
rect 39559 730 39595 802
rect 39746 798 39760 832
rect 39794 821 39812 832
rect 39746 787 39762 798
rect 39796 787 39812 821
rect 39371 684 39405 705
rect 39543 701 39595 730
rect 39371 629 39405 650
rect 39441 637 39457 671
rect 39491 637 39507 671
rect 38192 550 38202 564
rect 34790 420 34824 454
rect 34790 368 34824 384
rect 36182 444 36314 480
rect 36486 490 36520 506
rect 36582 490 36616 506
rect 36520 454 36521 455
rect 36182 396 36218 444
rect 36486 420 36521 454
rect 36520 418 36521 420
rect 36582 420 36616 454
rect 36366 396 36486 418
rect 36182 384 36486 396
rect 36520 384 36522 418
rect 36182 382 36522 384
rect 36182 360 36402 382
rect 36486 368 36520 382
rect 36582 368 36616 384
rect 36678 490 36712 506
rect 38152 480 38202 550
rect 38502 540 38518 574
rect 38552 540 38568 574
rect 38782 566 38830 578
rect 38990 563 39019 597
rect 39053 563 39111 597
rect 39145 563 39203 597
rect 39237 563 39266 597
rect 39441 595 39507 637
rect 39577 667 39595 701
rect 39543 629 39595 667
rect 39746 737 39792 753
rect 39846 749 39892 869
rect 40030 1047 40064 1066
rect 40116 1057 40321 1066
rect 40355 1089 40564 1091
rect 40355 1057 40440 1089
rect 40116 1055 40440 1057
rect 40474 1066 40564 1089
rect 40804 1066 40838 1424
rect 41748 1398 41782 1609
rect 41979 1306 42013 1609
rect 42064 1390 42098 2004
rect 42264 2002 42330 2004
rect 42581 2009 42597 2043
rect 42631 2009 42647 2043
rect 42581 1975 42647 2009
rect 42136 1943 42170 1962
rect 42136 1875 42170 1877
rect 42136 1839 42170 1841
rect 42136 1754 42170 1773
rect 42232 1943 42266 1962
rect 42232 1875 42266 1877
rect 42232 1839 42266 1841
rect 42232 1754 42266 1773
rect 42328 1943 42362 1962
rect 42581 1941 42597 1975
rect 42631 1959 42647 1975
rect 42753 2111 42819 2153
rect 42787 2077 42819 2111
rect 42753 2043 42819 2077
rect 42787 2009 42819 2043
rect 42753 1975 42819 2009
rect 42631 1941 42717 1959
rect 42581 1925 42717 1941
rect 42787 1941 42819 1975
rect 42753 1925 42819 1941
rect 43655 2111 43721 2116
rect 43655 2077 43671 2111
rect 43705 2077 43721 2111
rect 43655 2043 43721 2077
rect 43655 2009 43671 2043
rect 43705 2009 43721 2043
rect 43655 1975 43721 2009
rect 43655 1941 43671 1975
rect 43705 1959 43721 1975
rect 43827 2111 43893 2153
rect 43861 2077 43893 2111
rect 44060 2147 44342 2153
rect 44060 2113 44099 2147
rect 44133 2145 44342 2147
rect 44133 2113 44218 2145
rect 44060 2111 44218 2113
rect 44252 2111 44342 2145
rect 44060 2078 44342 2111
rect 44469 2111 44535 2116
rect 43827 2043 43893 2077
rect 43861 2009 43893 2043
rect 44469 2077 44485 2111
rect 44519 2077 44535 2111
rect 44469 2043 44535 2077
rect 43827 1975 43893 2009
rect 43705 1941 43791 1959
rect 43655 1925 43791 1941
rect 43861 1941 43893 1975
rect 43827 1925 43893 1941
rect 43952 2039 44218 2040
rect 43952 2005 44168 2039
rect 44202 2005 44218 2039
rect 43952 2004 44218 2005
rect 42328 1875 42362 1877
rect 42579 1882 42649 1891
rect 42579 1848 42595 1882
rect 42629 1875 42649 1882
rect 42579 1841 42599 1848
rect 42633 1841 42649 1875
rect 42328 1839 42362 1841
rect 42683 1805 42717 1925
rect 42751 1882 42821 1891
rect 42751 1875 42769 1882
rect 42751 1841 42767 1875
rect 42803 1848 42821 1882
rect 42801 1841 42821 1848
rect 43653 1884 43723 1891
rect 43653 1850 43671 1884
rect 43705 1875 43723 1884
rect 43653 1841 43673 1850
rect 43707 1841 43723 1875
rect 43757 1805 43791 1925
rect 43825 1880 43895 1891
rect 43825 1875 43844 1880
rect 43825 1841 43841 1875
rect 43878 1846 43895 1880
rect 43875 1841 43895 1846
rect 42328 1754 42362 1773
rect 42583 1789 42631 1805
rect 42583 1755 42597 1789
rect 42583 1721 42631 1755
rect 42168 1677 42184 1711
rect 42218 1677 42234 1711
rect 42583 1687 42597 1721
rect 42583 1643 42631 1687
rect 42665 1789 42731 1805
rect 42665 1755 42681 1789
rect 42715 1759 42731 1789
rect 42665 1725 42683 1755
rect 42717 1725 42731 1759
rect 42665 1721 42731 1725
rect 42665 1687 42681 1721
rect 42715 1687 42731 1721
rect 42665 1677 42731 1687
rect 42765 1789 42819 1805
rect 42799 1755 42819 1789
rect 42765 1721 42819 1755
rect 42799 1687 42819 1721
rect 42765 1643 42819 1687
rect 43657 1789 43705 1805
rect 43657 1755 43671 1789
rect 43657 1721 43705 1755
rect 43657 1687 43671 1721
rect 43657 1643 43705 1687
rect 43739 1789 43805 1805
rect 43739 1764 43755 1789
rect 43739 1730 43753 1764
rect 43789 1755 43805 1789
rect 43787 1730 43805 1755
rect 43739 1721 43805 1730
rect 43739 1687 43755 1721
rect 43789 1687 43805 1721
rect 43739 1677 43805 1687
rect 43839 1789 43893 1805
rect 43873 1755 43893 1789
rect 43839 1721 43893 1755
rect 43873 1687 43893 1721
rect 43839 1643 43893 1687
rect 42280 1596 42296 1630
rect 42330 1596 42346 1630
rect 42562 1609 42591 1643
rect 42625 1609 42683 1643
rect 42717 1609 42775 1643
rect 42809 1609 42838 1643
rect 43636 1609 43665 1643
rect 43699 1609 43757 1643
rect 43791 1609 43849 1643
rect 43883 1609 43912 1643
rect 42152 1546 42186 1562
rect 42152 1476 42186 1510
rect 42152 1424 42186 1440
rect 42248 1546 42282 1562
rect 42248 1476 42282 1510
rect 42248 1424 42282 1440
rect 42344 1546 42378 1562
rect 42344 1476 42378 1510
rect 42378 1440 42726 1464
rect 42344 1424 42726 1440
rect 42064 1356 42200 1390
rect 42234 1356 42250 1390
rect 41979 1286 42374 1306
rect 41979 1281 42241 1286
rect 41979 1272 42120 1281
rect 42104 1247 42120 1272
rect 42154 1252 42241 1281
rect 42275 1262 42374 1286
rect 42546 1264 42592 1266
rect 42546 1262 42550 1264
rect 42275 1252 42550 1262
rect 42154 1247 42550 1252
rect 42104 1230 42550 1247
rect 42584 1230 42592 1264
rect 42104 1228 42592 1230
rect 42546 1222 42592 1228
rect 40878 1107 40907 1141
rect 40941 1107 40999 1141
rect 41033 1107 41091 1141
rect 41125 1107 41154 1141
rect 40474 1055 40710 1066
rect 40116 1047 40710 1055
rect 40116 1022 40118 1047
rect 40030 979 40064 981
rect 40030 943 40064 945
rect 40030 858 40064 877
rect 40152 1022 40676 1047
rect 40762 1047 40838 1066
rect 40762 1026 40764 1047
rect 40118 979 40152 981
rect 40374 949 40390 983
rect 40424 949 40440 983
rect 40676 979 40710 981
rect 40118 943 40152 945
rect 40676 943 40710 945
rect 40118 858 40152 877
rect 40246 887 40280 906
rect 40246 819 40280 821
rect 40058 781 40074 815
rect 40108 781 40124 815
rect 40246 783 40280 785
rect 39746 703 39758 737
rect 39746 669 39792 703
rect 39746 635 39758 669
rect 39336 561 39365 595
rect 39399 561 39457 595
rect 39491 561 39549 595
rect 39583 561 39612 595
rect 39746 589 39792 635
rect 39826 737 39892 749
rect 39826 703 39842 737
rect 39876 703 39892 737
rect 39826 690 39892 703
rect 40246 698 40280 717
rect 40342 887 40376 906
rect 40342 819 40376 821
rect 40342 783 40376 785
rect 40342 698 40376 717
rect 40438 887 40472 906
rect 40676 858 40710 877
rect 40798 1026 40838 1047
rect 40946 1065 40988 1107
rect 41224 1105 41253 1139
rect 41287 1105 41345 1139
rect 41379 1105 41437 1139
rect 41471 1105 41500 1139
rect 41645 1133 41679 1140
rect 40946 1031 40954 1065
rect 40764 979 40798 981
rect 40764 943 40798 945
rect 40946 997 40988 1031
rect 40946 963 40954 997
rect 40946 929 40988 963
rect 40946 895 40954 929
rect 40946 879 40988 895
rect 41022 1065 41088 1073
rect 41022 1031 41038 1065
rect 41072 1031 41088 1065
rect 41022 997 41088 1031
rect 41022 963 41038 997
rect 41072 963 41088 997
rect 41022 929 41088 963
rect 41022 895 41038 929
rect 41072 895 41088 929
rect 41022 877 41088 895
rect 41257 1055 41293 1071
rect 41257 1021 41259 1055
rect 41257 987 41293 1021
rect 41257 953 41259 987
rect 41329 1055 41395 1105
rect 41570 1099 41599 1133
rect 41633 1099 41691 1133
rect 41725 1099 41783 1133
rect 41817 1099 41846 1133
rect 41946 1109 41962 1143
rect 41996 1109 42012 1143
rect 42170 1130 42284 1132
rect 41329 1021 41345 1055
rect 41379 1021 41395 1055
rect 41329 987 41395 1021
rect 41329 953 41345 987
rect 41379 953 41395 987
rect 41429 1055 41483 1071
rect 41429 1021 41431 1055
rect 41465 1021 41483 1055
rect 41429 974 41483 1021
rect 41257 919 41293 953
rect 41429 940 41431 974
rect 41465 940 41483 974
rect 41257 885 41392 919
rect 41429 890 41483 940
rect 40764 858 40798 877
rect 40438 819 40472 821
rect 40850 843 40994 844
rect 40850 829 41008 843
rect 40438 783 40472 785
rect 40704 816 40770 818
rect 40850 816 40958 829
rect 40704 815 40958 816
rect 40704 781 40720 815
rect 40754 802 40958 815
rect 40754 782 40890 802
rect 40942 795 40958 802
rect 40992 795 41008 829
rect 40754 781 40770 782
rect 40942 745 40988 761
rect 41042 757 41088 877
rect 41358 856 41392 885
rect 41245 827 41313 849
rect 41245 826 41261 827
rect 41245 792 41259 826
rect 41295 793 41313 827
rect 41293 792 41313 793
rect 41245 775 41313 792
rect 41358 840 41413 856
rect 41358 806 41379 840
rect 41358 790 41413 806
rect 41447 840 41483 890
rect 41638 1057 41680 1099
rect 42170 1091 42452 1130
rect 42592 1109 42608 1143
rect 42642 1109 42658 1143
rect 42170 1066 42209 1091
rect 41638 1023 41646 1057
rect 41638 989 41680 1023
rect 41638 955 41646 989
rect 41638 921 41680 955
rect 41638 887 41646 921
rect 41638 871 41680 887
rect 41714 1057 41780 1065
rect 41714 1023 41730 1057
rect 41764 1023 41780 1057
rect 41714 989 41780 1023
rect 41714 955 41730 989
rect 41764 955 41780 989
rect 41714 921 41780 955
rect 41714 887 41730 921
rect 41764 887 41780 921
rect 41714 869 41780 887
rect 41447 838 41488 840
rect 41447 804 41452 838
rect 41486 804 41488 838
rect 41447 802 41488 804
rect 41634 832 41700 835
rect 40472 717 40718 734
rect 40438 700 40718 717
rect 40438 698 40472 700
rect 39826 669 40168 690
rect 39826 635 39842 669
rect 39876 658 40168 669
rect 39876 655 40344 658
rect 39876 654 40294 655
rect 39876 635 39898 654
rect 39826 630 39898 635
rect 39826 623 39892 630
rect 40132 622 40294 654
rect 40278 621 40294 622
rect 40328 621 40344 655
rect 40670 612 40718 700
rect 39682 555 39711 589
rect 39745 555 39803 589
rect 39837 555 39895 589
rect 39929 555 39958 589
rect 40040 584 40086 594
rect 40040 550 40046 584
rect 40080 564 40086 584
rect 40670 578 40678 612
rect 40712 578 40718 612
rect 40942 711 40954 745
rect 40942 677 40988 711
rect 40942 643 40954 677
rect 40942 597 40988 643
rect 41022 745 41088 757
rect 41022 694 41038 745
rect 41072 694 41088 745
rect 41358 739 41392 790
rect 41022 677 41088 694
rect 41022 643 41038 677
rect 41072 643 41088 677
rect 41022 631 41088 643
rect 41259 705 41392 739
rect 41447 730 41483 802
rect 41634 798 41648 832
rect 41682 821 41700 832
rect 41634 787 41650 798
rect 41684 787 41700 821
rect 41259 684 41293 705
rect 41431 701 41483 730
rect 41259 629 41293 650
rect 41329 637 41345 671
rect 41379 637 41395 671
rect 40080 550 40090 564
rect 36678 420 36712 454
rect 36678 368 36712 384
rect 38070 444 38202 480
rect 38374 490 38408 506
rect 38470 490 38504 506
rect 38408 454 38409 455
rect 38070 396 38106 444
rect 38374 420 38409 454
rect 38408 418 38409 420
rect 38470 420 38504 454
rect 38254 396 38374 418
rect 38070 384 38374 396
rect 38408 384 38410 418
rect 38070 382 38410 384
rect 38070 360 38290 382
rect 38374 368 38408 382
rect 38470 368 38504 384
rect 38566 490 38600 506
rect 40040 480 40090 550
rect 40390 540 40406 574
rect 40440 540 40456 574
rect 40670 566 40718 578
rect 40878 563 40907 597
rect 40941 563 40999 597
rect 41033 563 41091 597
rect 41125 563 41154 597
rect 41329 595 41395 637
rect 41465 667 41483 701
rect 41431 629 41483 667
rect 41634 737 41680 753
rect 41734 749 41780 869
rect 41918 1047 41952 1066
rect 42004 1057 42209 1066
rect 42243 1089 42452 1091
rect 42243 1057 42328 1089
rect 42004 1055 42328 1057
rect 42362 1066 42452 1089
rect 42692 1066 42726 1424
rect 43636 1398 43670 1609
rect 43867 1306 43901 1609
rect 43952 1390 43986 2004
rect 44152 2002 44218 2004
rect 44469 2009 44485 2043
rect 44519 2009 44535 2043
rect 44469 1975 44535 2009
rect 44024 1943 44058 1962
rect 44024 1875 44058 1877
rect 44024 1839 44058 1841
rect 44024 1754 44058 1773
rect 44120 1943 44154 1962
rect 44120 1875 44154 1877
rect 44120 1839 44154 1841
rect 44120 1754 44154 1773
rect 44216 1943 44250 1962
rect 44469 1941 44485 1975
rect 44519 1959 44535 1975
rect 44641 2111 44707 2153
rect 44675 2077 44707 2111
rect 44641 2043 44707 2077
rect 44675 2009 44707 2043
rect 44641 1975 44707 2009
rect 44519 1941 44605 1959
rect 44469 1925 44605 1941
rect 44675 1941 44707 1975
rect 44641 1925 44707 1941
rect 45537 2111 45603 2116
rect 45537 2077 45553 2111
rect 45587 2077 45603 2111
rect 45537 2043 45603 2077
rect 45537 2009 45553 2043
rect 45587 2009 45603 2043
rect 45537 1975 45603 2009
rect 45537 1941 45553 1975
rect 45587 1959 45603 1975
rect 45709 2111 45775 2153
rect 45743 2077 45775 2111
rect 45942 2147 46224 2153
rect 45942 2113 45981 2147
rect 46015 2145 46224 2147
rect 46015 2113 46100 2145
rect 45942 2111 46100 2113
rect 46134 2111 46224 2145
rect 45942 2078 46224 2111
rect 46351 2111 46417 2116
rect 45709 2043 45775 2077
rect 45743 2009 45775 2043
rect 46351 2077 46367 2111
rect 46401 2077 46417 2111
rect 46351 2043 46417 2077
rect 45709 1975 45775 2009
rect 45587 1941 45673 1959
rect 45537 1925 45673 1941
rect 45743 1941 45775 1975
rect 45709 1925 45775 1941
rect 45834 2039 46100 2040
rect 45834 2005 46050 2039
rect 46084 2005 46100 2039
rect 45834 2004 46100 2005
rect 44216 1875 44250 1877
rect 44467 1882 44537 1891
rect 44467 1848 44483 1882
rect 44517 1875 44537 1882
rect 44467 1841 44487 1848
rect 44521 1841 44537 1875
rect 44216 1839 44250 1841
rect 44571 1805 44605 1925
rect 44639 1882 44709 1891
rect 44639 1875 44657 1882
rect 44639 1841 44655 1875
rect 44691 1848 44709 1882
rect 44689 1841 44709 1848
rect 45535 1884 45605 1891
rect 45535 1850 45553 1884
rect 45587 1875 45605 1884
rect 45535 1841 45555 1850
rect 45589 1841 45605 1875
rect 45639 1805 45673 1925
rect 45707 1880 45777 1891
rect 45707 1875 45726 1880
rect 45707 1841 45723 1875
rect 45760 1846 45777 1880
rect 45757 1841 45777 1846
rect 44216 1754 44250 1773
rect 44471 1789 44519 1805
rect 44471 1755 44485 1789
rect 44471 1721 44519 1755
rect 44056 1677 44072 1711
rect 44106 1677 44122 1711
rect 44471 1687 44485 1721
rect 44471 1643 44519 1687
rect 44553 1789 44619 1805
rect 44553 1755 44569 1789
rect 44603 1759 44619 1789
rect 44553 1725 44571 1755
rect 44605 1725 44619 1759
rect 44553 1721 44619 1725
rect 44553 1687 44569 1721
rect 44603 1687 44619 1721
rect 44553 1677 44619 1687
rect 44653 1789 44707 1805
rect 44687 1755 44707 1789
rect 44653 1721 44707 1755
rect 44687 1687 44707 1721
rect 44653 1643 44707 1687
rect 45539 1789 45587 1805
rect 45539 1755 45553 1789
rect 45539 1721 45587 1755
rect 45539 1687 45553 1721
rect 45539 1643 45587 1687
rect 45621 1789 45687 1805
rect 45621 1764 45637 1789
rect 45621 1730 45635 1764
rect 45671 1755 45687 1789
rect 45669 1730 45687 1755
rect 45621 1721 45687 1730
rect 45621 1687 45637 1721
rect 45671 1687 45687 1721
rect 45621 1677 45687 1687
rect 45721 1789 45775 1805
rect 45755 1755 45775 1789
rect 45721 1721 45775 1755
rect 45755 1687 45775 1721
rect 45721 1643 45775 1687
rect 44168 1596 44184 1630
rect 44218 1596 44234 1630
rect 44450 1609 44479 1643
rect 44513 1609 44571 1643
rect 44605 1609 44663 1643
rect 44697 1609 44726 1643
rect 45518 1609 45547 1643
rect 45581 1609 45639 1643
rect 45673 1609 45731 1643
rect 45765 1609 45794 1643
rect 44040 1546 44074 1562
rect 44040 1476 44074 1510
rect 44040 1424 44074 1440
rect 44136 1546 44170 1562
rect 44136 1476 44170 1510
rect 44136 1424 44170 1440
rect 44232 1546 44266 1562
rect 44232 1476 44266 1510
rect 44266 1440 44614 1464
rect 44232 1424 44614 1440
rect 43952 1356 44088 1390
rect 44122 1356 44138 1390
rect 43867 1286 44262 1306
rect 43867 1281 44129 1286
rect 43867 1272 44008 1281
rect 43992 1247 44008 1272
rect 44042 1252 44129 1281
rect 44163 1262 44262 1286
rect 44434 1264 44480 1266
rect 44434 1262 44438 1264
rect 44163 1252 44438 1262
rect 44042 1247 44438 1252
rect 43992 1230 44438 1247
rect 44472 1230 44480 1264
rect 43992 1228 44480 1230
rect 44434 1222 44480 1228
rect 42766 1107 42795 1141
rect 42829 1107 42887 1141
rect 42921 1107 42979 1141
rect 43013 1107 43042 1141
rect 42362 1055 42598 1066
rect 42004 1047 42598 1055
rect 42004 1022 42006 1047
rect 41918 979 41952 981
rect 41918 943 41952 945
rect 41918 858 41952 877
rect 42040 1022 42564 1047
rect 42650 1047 42726 1066
rect 42650 1026 42652 1047
rect 42006 979 42040 981
rect 42262 949 42278 983
rect 42312 949 42328 983
rect 42564 979 42598 981
rect 42006 943 42040 945
rect 42564 943 42598 945
rect 42006 858 42040 877
rect 42134 887 42168 906
rect 42134 819 42168 821
rect 41946 781 41962 815
rect 41996 781 42012 815
rect 42134 783 42168 785
rect 41634 703 41646 737
rect 41634 669 41680 703
rect 41634 635 41646 669
rect 41224 561 41253 595
rect 41287 561 41345 595
rect 41379 561 41437 595
rect 41471 561 41500 595
rect 41634 589 41680 635
rect 41714 737 41780 749
rect 41714 703 41730 737
rect 41764 703 41780 737
rect 41714 690 41780 703
rect 42134 698 42168 717
rect 42230 887 42264 906
rect 42230 819 42264 821
rect 42230 783 42264 785
rect 42230 698 42264 717
rect 42326 887 42360 906
rect 42564 858 42598 877
rect 42686 1026 42726 1047
rect 42834 1065 42876 1107
rect 43112 1105 43141 1139
rect 43175 1105 43233 1139
rect 43267 1105 43325 1139
rect 43359 1105 43388 1139
rect 43533 1133 43567 1140
rect 42834 1031 42842 1065
rect 42652 979 42686 981
rect 42652 943 42686 945
rect 42834 997 42876 1031
rect 42834 963 42842 997
rect 42834 929 42876 963
rect 42834 895 42842 929
rect 42834 879 42876 895
rect 42910 1065 42976 1073
rect 42910 1031 42926 1065
rect 42960 1031 42976 1065
rect 42910 997 42976 1031
rect 42910 963 42926 997
rect 42960 963 42976 997
rect 42910 929 42976 963
rect 42910 895 42926 929
rect 42960 895 42976 929
rect 42910 877 42976 895
rect 43145 1055 43181 1071
rect 43145 1021 43147 1055
rect 43145 987 43181 1021
rect 43145 953 43147 987
rect 43217 1055 43283 1105
rect 43458 1099 43487 1133
rect 43521 1099 43579 1133
rect 43613 1099 43671 1133
rect 43705 1099 43734 1133
rect 43834 1109 43850 1143
rect 43884 1109 43900 1143
rect 44058 1130 44172 1132
rect 43217 1021 43233 1055
rect 43267 1021 43283 1055
rect 43217 987 43283 1021
rect 43217 953 43233 987
rect 43267 953 43283 987
rect 43317 1055 43371 1071
rect 43317 1021 43319 1055
rect 43353 1021 43371 1055
rect 43317 974 43371 1021
rect 43145 919 43181 953
rect 43317 940 43319 974
rect 43353 940 43371 974
rect 43145 885 43280 919
rect 43317 890 43371 940
rect 42652 858 42686 877
rect 42326 819 42360 821
rect 42738 843 42882 844
rect 42738 829 42896 843
rect 42326 783 42360 785
rect 42592 816 42658 818
rect 42738 816 42846 829
rect 42592 815 42846 816
rect 42592 781 42608 815
rect 42642 802 42846 815
rect 42642 782 42778 802
rect 42830 795 42846 802
rect 42880 795 42896 829
rect 42642 781 42658 782
rect 42830 745 42876 761
rect 42930 757 42976 877
rect 43246 856 43280 885
rect 43133 827 43201 849
rect 43133 826 43149 827
rect 43133 792 43147 826
rect 43183 793 43201 827
rect 43181 792 43201 793
rect 43133 775 43201 792
rect 43246 840 43301 856
rect 43246 806 43267 840
rect 43246 790 43301 806
rect 43335 840 43371 890
rect 43526 1057 43568 1099
rect 44058 1091 44340 1130
rect 44480 1109 44496 1143
rect 44530 1109 44546 1143
rect 44058 1066 44097 1091
rect 43526 1023 43534 1057
rect 43526 989 43568 1023
rect 43526 955 43534 989
rect 43526 921 43568 955
rect 43526 887 43534 921
rect 43526 871 43568 887
rect 43602 1057 43668 1065
rect 43602 1023 43618 1057
rect 43652 1023 43668 1057
rect 43602 989 43668 1023
rect 43602 955 43618 989
rect 43652 955 43668 989
rect 43602 921 43668 955
rect 43602 887 43618 921
rect 43652 887 43668 921
rect 43602 869 43668 887
rect 43335 838 43376 840
rect 43335 804 43340 838
rect 43374 804 43376 838
rect 43335 802 43376 804
rect 43522 832 43588 835
rect 42360 717 42606 734
rect 42326 700 42606 717
rect 42326 698 42360 700
rect 41714 669 42056 690
rect 41714 635 41730 669
rect 41764 658 42056 669
rect 41764 655 42232 658
rect 41764 654 42182 655
rect 41764 635 41786 654
rect 41714 630 41786 635
rect 41714 623 41780 630
rect 42020 622 42182 654
rect 42166 621 42182 622
rect 42216 621 42232 655
rect 42558 612 42606 700
rect 41570 555 41599 589
rect 41633 555 41691 589
rect 41725 555 41783 589
rect 41817 555 41846 589
rect 41928 584 41974 594
rect 41928 550 41934 584
rect 41968 564 41974 584
rect 42558 578 42566 612
rect 42600 578 42606 612
rect 42830 711 42842 745
rect 42830 677 42876 711
rect 42830 643 42842 677
rect 42830 597 42876 643
rect 42910 745 42976 757
rect 42910 694 42926 745
rect 42960 694 42976 745
rect 43246 739 43280 790
rect 42910 677 42976 694
rect 42910 643 42926 677
rect 42960 643 42976 677
rect 42910 631 42976 643
rect 43147 705 43280 739
rect 43335 730 43371 802
rect 43522 798 43536 832
rect 43570 821 43588 832
rect 43522 787 43538 798
rect 43572 787 43588 821
rect 43147 684 43181 705
rect 43319 701 43371 730
rect 43147 629 43181 650
rect 43217 637 43233 671
rect 43267 637 43283 671
rect 41968 550 41978 564
rect 38566 420 38600 454
rect 38566 368 38600 384
rect 39958 444 40090 480
rect 40262 490 40296 506
rect 40358 490 40392 506
rect 40296 454 40297 455
rect 39958 396 39994 444
rect 40262 420 40297 454
rect 40296 418 40297 420
rect 40358 420 40392 454
rect 40142 396 40262 418
rect 39958 384 40262 396
rect 40296 384 40298 418
rect 39958 382 40298 384
rect 39958 360 40178 382
rect 40262 368 40296 382
rect 40358 368 40392 384
rect 40454 490 40488 506
rect 41928 480 41978 550
rect 42278 540 42294 574
rect 42328 540 42344 574
rect 42558 566 42606 578
rect 42766 563 42795 597
rect 42829 563 42887 597
rect 42921 563 42979 597
rect 43013 563 43042 597
rect 43217 595 43283 637
rect 43353 667 43371 701
rect 43319 629 43371 667
rect 43522 737 43568 753
rect 43622 749 43668 869
rect 43806 1047 43840 1066
rect 43892 1057 44097 1066
rect 44131 1089 44340 1091
rect 44131 1057 44216 1089
rect 43892 1055 44216 1057
rect 44250 1066 44340 1089
rect 44580 1066 44614 1424
rect 45518 1398 45552 1609
rect 45749 1306 45783 1609
rect 45834 1390 45868 2004
rect 46034 2002 46100 2004
rect 46351 2009 46367 2043
rect 46401 2009 46417 2043
rect 46351 1975 46417 2009
rect 45906 1943 45940 1962
rect 45906 1875 45940 1877
rect 45906 1839 45940 1841
rect 45906 1754 45940 1773
rect 46002 1943 46036 1962
rect 46002 1875 46036 1877
rect 46002 1839 46036 1841
rect 46002 1754 46036 1773
rect 46098 1943 46132 1962
rect 46351 1941 46367 1975
rect 46401 1959 46417 1975
rect 46523 2111 46589 2153
rect 46557 2077 46589 2111
rect 46523 2043 46589 2077
rect 46557 2009 46589 2043
rect 46523 1975 46589 2009
rect 46401 1941 46487 1959
rect 46351 1925 46487 1941
rect 46557 1941 46589 1975
rect 46523 1925 46589 1941
rect 47425 2111 47491 2116
rect 47425 2077 47441 2111
rect 47475 2077 47491 2111
rect 47425 2043 47491 2077
rect 47425 2009 47441 2043
rect 47475 2009 47491 2043
rect 47425 1975 47491 2009
rect 47425 1941 47441 1975
rect 47475 1959 47491 1975
rect 47597 2111 47663 2153
rect 47631 2077 47663 2111
rect 47830 2147 48112 2153
rect 47830 2113 47869 2147
rect 47903 2145 48112 2147
rect 47903 2113 47988 2145
rect 47830 2111 47988 2113
rect 48022 2111 48112 2145
rect 47830 2078 48112 2111
rect 48239 2111 48305 2116
rect 47597 2043 47663 2077
rect 47631 2009 47663 2043
rect 48239 2077 48255 2111
rect 48289 2077 48305 2111
rect 48239 2043 48305 2077
rect 47597 1975 47663 2009
rect 47475 1941 47561 1959
rect 47425 1925 47561 1941
rect 47631 1941 47663 1975
rect 47597 1925 47663 1941
rect 47722 2039 47988 2040
rect 47722 2005 47938 2039
rect 47972 2005 47988 2039
rect 47722 2004 47988 2005
rect 46098 1875 46132 1877
rect 46349 1882 46419 1891
rect 46349 1848 46365 1882
rect 46399 1875 46419 1882
rect 46349 1841 46369 1848
rect 46403 1841 46419 1875
rect 46098 1839 46132 1841
rect 46453 1805 46487 1925
rect 46521 1882 46591 1891
rect 46521 1875 46539 1882
rect 46521 1841 46537 1875
rect 46573 1848 46591 1882
rect 46571 1841 46591 1848
rect 47423 1884 47493 1891
rect 47423 1850 47441 1884
rect 47475 1875 47493 1884
rect 47423 1841 47443 1850
rect 47477 1841 47493 1875
rect 47527 1805 47561 1925
rect 47595 1880 47665 1891
rect 47595 1875 47614 1880
rect 47595 1841 47611 1875
rect 47648 1846 47665 1880
rect 47645 1841 47665 1846
rect 46098 1754 46132 1773
rect 46353 1789 46401 1805
rect 46353 1755 46367 1789
rect 46353 1721 46401 1755
rect 45938 1677 45954 1711
rect 45988 1677 46004 1711
rect 46353 1687 46367 1721
rect 46353 1643 46401 1687
rect 46435 1789 46501 1805
rect 46435 1755 46451 1789
rect 46485 1759 46501 1789
rect 46435 1725 46453 1755
rect 46487 1725 46501 1759
rect 46435 1721 46501 1725
rect 46435 1687 46451 1721
rect 46485 1687 46501 1721
rect 46435 1677 46501 1687
rect 46535 1789 46589 1805
rect 46569 1755 46589 1789
rect 46535 1721 46589 1755
rect 46569 1687 46589 1721
rect 46535 1643 46589 1687
rect 47427 1789 47475 1805
rect 47427 1755 47441 1789
rect 47427 1721 47475 1755
rect 47427 1687 47441 1721
rect 47427 1643 47475 1687
rect 47509 1789 47575 1805
rect 47509 1764 47525 1789
rect 47509 1730 47523 1764
rect 47559 1755 47575 1789
rect 47557 1730 47575 1755
rect 47509 1721 47575 1730
rect 47509 1687 47525 1721
rect 47559 1687 47575 1721
rect 47509 1677 47575 1687
rect 47609 1789 47663 1805
rect 47643 1755 47663 1789
rect 47609 1721 47663 1755
rect 47643 1687 47663 1721
rect 47609 1643 47663 1687
rect 46050 1596 46066 1630
rect 46100 1596 46116 1630
rect 46332 1609 46361 1643
rect 46395 1609 46453 1643
rect 46487 1609 46545 1643
rect 46579 1609 46608 1643
rect 47406 1609 47435 1643
rect 47469 1609 47527 1643
rect 47561 1609 47619 1643
rect 47653 1609 47682 1643
rect 45922 1546 45956 1562
rect 45922 1476 45956 1510
rect 45922 1424 45956 1440
rect 46018 1546 46052 1562
rect 46018 1476 46052 1510
rect 46018 1424 46052 1440
rect 46114 1546 46148 1562
rect 46114 1476 46148 1510
rect 46148 1440 46496 1464
rect 46114 1424 46496 1440
rect 45834 1356 45970 1390
rect 46004 1356 46020 1390
rect 45749 1286 46144 1306
rect 45749 1281 46011 1286
rect 45749 1272 45890 1281
rect 45874 1247 45890 1272
rect 45924 1252 46011 1281
rect 46045 1262 46144 1286
rect 46316 1264 46362 1266
rect 46316 1262 46320 1264
rect 46045 1252 46320 1262
rect 45924 1247 46320 1252
rect 45874 1230 46320 1247
rect 46354 1230 46362 1264
rect 45874 1228 46362 1230
rect 46316 1222 46362 1228
rect 44654 1107 44683 1141
rect 44717 1107 44775 1141
rect 44809 1107 44867 1141
rect 44901 1107 44930 1141
rect 44250 1055 44486 1066
rect 43892 1047 44486 1055
rect 43892 1022 43894 1047
rect 43806 979 43840 981
rect 43806 943 43840 945
rect 43806 858 43840 877
rect 43928 1022 44452 1047
rect 44538 1047 44614 1066
rect 44538 1026 44540 1047
rect 43894 979 43928 981
rect 44150 949 44166 983
rect 44200 949 44216 983
rect 44452 979 44486 981
rect 43894 943 43928 945
rect 44452 943 44486 945
rect 43894 858 43928 877
rect 44022 887 44056 906
rect 44022 819 44056 821
rect 43834 781 43850 815
rect 43884 781 43900 815
rect 44022 783 44056 785
rect 43522 703 43534 737
rect 43522 669 43568 703
rect 43522 635 43534 669
rect 43112 561 43141 595
rect 43175 561 43233 595
rect 43267 561 43325 595
rect 43359 561 43388 595
rect 43522 589 43568 635
rect 43602 737 43668 749
rect 43602 703 43618 737
rect 43652 703 43668 737
rect 43602 690 43668 703
rect 44022 698 44056 717
rect 44118 887 44152 906
rect 44118 819 44152 821
rect 44118 783 44152 785
rect 44118 698 44152 717
rect 44214 887 44248 906
rect 44452 858 44486 877
rect 44574 1026 44614 1047
rect 44722 1065 44764 1107
rect 45000 1105 45029 1139
rect 45063 1105 45121 1139
rect 45155 1105 45213 1139
rect 45247 1105 45276 1139
rect 45415 1133 45449 1140
rect 44722 1031 44730 1065
rect 44540 979 44574 981
rect 44540 943 44574 945
rect 44722 997 44764 1031
rect 44722 963 44730 997
rect 44722 929 44764 963
rect 44722 895 44730 929
rect 44722 879 44764 895
rect 44798 1065 44864 1073
rect 44798 1031 44814 1065
rect 44848 1031 44864 1065
rect 44798 997 44864 1031
rect 44798 963 44814 997
rect 44848 963 44864 997
rect 44798 929 44864 963
rect 44798 895 44814 929
rect 44848 895 44864 929
rect 44798 877 44864 895
rect 45033 1055 45069 1071
rect 45033 1021 45035 1055
rect 45033 987 45069 1021
rect 45033 953 45035 987
rect 45105 1055 45171 1105
rect 45340 1099 45369 1133
rect 45403 1099 45461 1133
rect 45495 1099 45553 1133
rect 45587 1099 45616 1133
rect 45716 1109 45732 1143
rect 45766 1109 45782 1143
rect 45940 1130 46054 1132
rect 45105 1021 45121 1055
rect 45155 1021 45171 1055
rect 45105 987 45171 1021
rect 45105 953 45121 987
rect 45155 953 45171 987
rect 45205 1055 45259 1071
rect 45205 1021 45207 1055
rect 45241 1021 45259 1055
rect 45205 974 45259 1021
rect 45033 919 45069 953
rect 45205 940 45207 974
rect 45241 940 45259 974
rect 45033 885 45168 919
rect 45205 890 45259 940
rect 44540 858 44574 877
rect 44214 819 44248 821
rect 44626 843 44770 844
rect 44626 829 44784 843
rect 44214 783 44248 785
rect 44480 816 44546 818
rect 44626 816 44734 829
rect 44480 815 44734 816
rect 44480 781 44496 815
rect 44530 802 44734 815
rect 44530 782 44666 802
rect 44718 795 44734 802
rect 44768 795 44784 829
rect 44530 781 44546 782
rect 44718 745 44764 761
rect 44818 757 44864 877
rect 45134 856 45168 885
rect 45021 827 45089 849
rect 45021 826 45037 827
rect 45021 792 45035 826
rect 45071 793 45089 827
rect 45069 792 45089 793
rect 45021 775 45089 792
rect 45134 840 45189 856
rect 45134 806 45155 840
rect 45134 790 45189 806
rect 45223 840 45259 890
rect 45408 1057 45450 1099
rect 45940 1091 46222 1130
rect 46362 1109 46378 1143
rect 46412 1109 46428 1143
rect 45940 1066 45979 1091
rect 45408 1023 45416 1057
rect 45408 989 45450 1023
rect 45408 955 45416 989
rect 45408 921 45450 955
rect 45408 887 45416 921
rect 45408 871 45450 887
rect 45484 1057 45550 1065
rect 45484 1023 45500 1057
rect 45534 1023 45550 1057
rect 45484 989 45550 1023
rect 45484 955 45500 989
rect 45534 955 45550 989
rect 45484 921 45550 955
rect 45484 887 45500 921
rect 45534 887 45550 921
rect 45484 869 45550 887
rect 45223 838 45264 840
rect 45223 804 45228 838
rect 45262 804 45264 838
rect 45223 802 45264 804
rect 45404 832 45470 835
rect 44248 717 44494 734
rect 44214 700 44494 717
rect 44214 698 44248 700
rect 43602 669 43944 690
rect 43602 635 43618 669
rect 43652 658 43944 669
rect 43652 655 44120 658
rect 43652 654 44070 655
rect 43652 635 43674 654
rect 43602 630 43674 635
rect 43602 623 43668 630
rect 43908 622 44070 654
rect 44054 621 44070 622
rect 44104 621 44120 655
rect 44446 612 44494 700
rect 43458 555 43487 589
rect 43521 555 43579 589
rect 43613 555 43671 589
rect 43705 555 43734 589
rect 43816 584 43862 594
rect 43816 550 43822 584
rect 43856 564 43862 584
rect 44446 578 44454 612
rect 44488 578 44494 612
rect 44718 711 44730 745
rect 44718 677 44764 711
rect 44718 643 44730 677
rect 44718 597 44764 643
rect 44798 745 44864 757
rect 44798 694 44814 745
rect 44848 694 44864 745
rect 45134 739 45168 790
rect 44798 677 44864 694
rect 44798 643 44814 677
rect 44848 643 44864 677
rect 44798 631 44864 643
rect 45035 705 45168 739
rect 45223 730 45259 802
rect 45404 798 45418 832
rect 45452 821 45470 832
rect 45404 787 45420 798
rect 45454 787 45470 821
rect 45035 684 45069 705
rect 45207 701 45259 730
rect 45035 629 45069 650
rect 45105 637 45121 671
rect 45155 637 45171 671
rect 43856 550 43866 564
rect 40454 420 40488 454
rect 40454 368 40488 384
rect 41846 444 41978 480
rect 42150 490 42184 506
rect 42246 490 42280 506
rect 42184 454 42185 455
rect 41846 396 41882 444
rect 42150 420 42185 454
rect 42184 418 42185 420
rect 42246 420 42280 454
rect 42030 396 42150 418
rect 41846 384 42150 396
rect 42184 384 42186 418
rect 41846 382 42186 384
rect 41846 360 42066 382
rect 42150 368 42184 382
rect 42246 368 42280 384
rect 42342 490 42376 506
rect 43816 480 43866 550
rect 44166 540 44182 574
rect 44216 540 44232 574
rect 44446 566 44494 578
rect 44654 563 44683 597
rect 44717 563 44775 597
rect 44809 563 44867 597
rect 44901 563 44930 597
rect 45105 595 45171 637
rect 45241 667 45259 701
rect 45207 629 45259 667
rect 45404 737 45450 753
rect 45504 749 45550 869
rect 45688 1047 45722 1066
rect 45774 1057 45979 1066
rect 46013 1089 46222 1091
rect 46013 1057 46098 1089
rect 45774 1055 46098 1057
rect 46132 1066 46222 1089
rect 46462 1066 46496 1424
rect 47406 1398 47440 1609
rect 47637 1306 47671 1609
rect 47722 1390 47756 2004
rect 47922 2002 47988 2004
rect 48239 2009 48255 2043
rect 48289 2009 48305 2043
rect 48239 1975 48305 2009
rect 47794 1943 47828 1962
rect 47794 1875 47828 1877
rect 47794 1839 47828 1841
rect 47794 1754 47828 1773
rect 47890 1943 47924 1962
rect 47890 1875 47924 1877
rect 47890 1839 47924 1841
rect 47890 1754 47924 1773
rect 47986 1943 48020 1962
rect 48239 1941 48255 1975
rect 48289 1959 48305 1975
rect 48411 2111 48477 2153
rect 48445 2077 48477 2111
rect 48411 2043 48477 2077
rect 48445 2009 48477 2043
rect 48411 1975 48477 2009
rect 48289 1941 48375 1959
rect 48239 1925 48375 1941
rect 48445 1941 48477 1975
rect 48411 1925 48477 1941
rect 49313 2111 49379 2116
rect 49313 2077 49329 2111
rect 49363 2077 49379 2111
rect 49313 2043 49379 2077
rect 49313 2009 49329 2043
rect 49363 2009 49379 2043
rect 49313 1975 49379 2009
rect 49313 1941 49329 1975
rect 49363 1959 49379 1975
rect 49485 2111 49551 2153
rect 49519 2077 49551 2111
rect 49718 2147 50000 2153
rect 49718 2113 49757 2147
rect 49791 2145 50000 2147
rect 49791 2113 49876 2145
rect 49718 2111 49876 2113
rect 49910 2111 50000 2145
rect 49718 2078 50000 2111
rect 50127 2111 50193 2116
rect 49485 2043 49551 2077
rect 49519 2009 49551 2043
rect 50127 2077 50143 2111
rect 50177 2077 50193 2111
rect 50127 2043 50193 2077
rect 49485 1975 49551 2009
rect 49363 1941 49449 1959
rect 49313 1925 49449 1941
rect 49519 1941 49551 1975
rect 49485 1925 49551 1941
rect 49610 2039 49876 2040
rect 49610 2005 49826 2039
rect 49860 2005 49876 2039
rect 49610 2004 49876 2005
rect 47986 1875 48020 1877
rect 48237 1882 48307 1891
rect 48237 1848 48253 1882
rect 48287 1875 48307 1882
rect 48237 1841 48257 1848
rect 48291 1841 48307 1875
rect 47986 1839 48020 1841
rect 48341 1805 48375 1925
rect 48409 1882 48479 1891
rect 48409 1875 48427 1882
rect 48409 1841 48425 1875
rect 48461 1848 48479 1882
rect 48459 1841 48479 1848
rect 49311 1884 49381 1891
rect 49311 1850 49329 1884
rect 49363 1875 49381 1884
rect 49311 1841 49331 1850
rect 49365 1841 49381 1875
rect 49415 1805 49449 1925
rect 49483 1880 49553 1891
rect 49483 1875 49502 1880
rect 49483 1841 49499 1875
rect 49536 1846 49553 1880
rect 49533 1841 49553 1846
rect 47986 1754 48020 1773
rect 48241 1789 48289 1805
rect 48241 1755 48255 1789
rect 48241 1721 48289 1755
rect 47826 1677 47842 1711
rect 47876 1677 47892 1711
rect 48241 1687 48255 1721
rect 48241 1643 48289 1687
rect 48323 1789 48389 1805
rect 48323 1755 48339 1789
rect 48373 1759 48389 1789
rect 48323 1725 48341 1755
rect 48375 1725 48389 1759
rect 48323 1721 48389 1725
rect 48323 1687 48339 1721
rect 48373 1687 48389 1721
rect 48323 1677 48389 1687
rect 48423 1789 48477 1805
rect 48457 1755 48477 1789
rect 48423 1721 48477 1755
rect 48457 1687 48477 1721
rect 48423 1643 48477 1687
rect 49315 1789 49363 1805
rect 49315 1755 49329 1789
rect 49315 1721 49363 1755
rect 49315 1687 49329 1721
rect 49315 1643 49363 1687
rect 49397 1789 49463 1805
rect 49397 1764 49413 1789
rect 49397 1730 49411 1764
rect 49447 1755 49463 1789
rect 49445 1730 49463 1755
rect 49397 1721 49463 1730
rect 49397 1687 49413 1721
rect 49447 1687 49463 1721
rect 49397 1677 49463 1687
rect 49497 1789 49551 1805
rect 49531 1755 49551 1789
rect 49497 1721 49551 1755
rect 49531 1687 49551 1721
rect 49497 1643 49551 1687
rect 47938 1596 47954 1630
rect 47988 1596 48004 1630
rect 48220 1609 48249 1643
rect 48283 1609 48341 1643
rect 48375 1609 48433 1643
rect 48467 1609 48496 1643
rect 49294 1609 49323 1643
rect 49357 1609 49415 1643
rect 49449 1609 49507 1643
rect 49541 1609 49570 1643
rect 47810 1546 47844 1562
rect 47810 1476 47844 1510
rect 47810 1424 47844 1440
rect 47906 1546 47940 1562
rect 47906 1476 47940 1510
rect 47906 1424 47940 1440
rect 48002 1546 48036 1562
rect 48002 1476 48036 1510
rect 48036 1440 48384 1464
rect 48002 1424 48384 1440
rect 47722 1356 47858 1390
rect 47892 1356 47908 1390
rect 47637 1286 48032 1306
rect 47637 1281 47899 1286
rect 47637 1272 47778 1281
rect 47762 1247 47778 1272
rect 47812 1252 47899 1281
rect 47933 1262 48032 1286
rect 48204 1264 48250 1266
rect 48204 1262 48208 1264
rect 47933 1252 48208 1262
rect 47812 1247 48208 1252
rect 47762 1230 48208 1247
rect 48242 1230 48250 1264
rect 47762 1228 48250 1230
rect 48204 1222 48250 1228
rect 46536 1107 46565 1141
rect 46599 1107 46657 1141
rect 46691 1107 46749 1141
rect 46783 1107 46812 1141
rect 46132 1055 46368 1066
rect 45774 1047 46368 1055
rect 45774 1022 45776 1047
rect 45688 979 45722 981
rect 45688 943 45722 945
rect 45688 858 45722 877
rect 45810 1022 46334 1047
rect 46420 1047 46496 1066
rect 46420 1026 46422 1047
rect 45776 979 45810 981
rect 46032 949 46048 983
rect 46082 949 46098 983
rect 46334 979 46368 981
rect 45776 943 45810 945
rect 46334 943 46368 945
rect 45776 858 45810 877
rect 45904 887 45938 906
rect 45904 819 45938 821
rect 45716 781 45732 815
rect 45766 781 45782 815
rect 45904 783 45938 785
rect 45404 703 45416 737
rect 45404 669 45450 703
rect 45404 635 45416 669
rect 45000 561 45029 595
rect 45063 561 45121 595
rect 45155 561 45213 595
rect 45247 561 45276 595
rect 45404 589 45450 635
rect 45484 737 45550 749
rect 45484 703 45500 737
rect 45534 703 45550 737
rect 45484 690 45550 703
rect 45904 698 45938 717
rect 46000 887 46034 906
rect 46000 819 46034 821
rect 46000 783 46034 785
rect 46000 698 46034 717
rect 46096 887 46130 906
rect 46334 858 46368 877
rect 46456 1026 46496 1047
rect 46604 1065 46646 1107
rect 46882 1105 46911 1139
rect 46945 1105 47003 1139
rect 47037 1105 47095 1139
rect 47129 1105 47158 1139
rect 47303 1133 47337 1140
rect 46604 1031 46612 1065
rect 46422 979 46456 981
rect 46422 943 46456 945
rect 46604 997 46646 1031
rect 46604 963 46612 997
rect 46604 929 46646 963
rect 46604 895 46612 929
rect 46604 879 46646 895
rect 46680 1065 46746 1073
rect 46680 1031 46696 1065
rect 46730 1031 46746 1065
rect 46680 997 46746 1031
rect 46680 963 46696 997
rect 46730 963 46746 997
rect 46680 929 46746 963
rect 46680 895 46696 929
rect 46730 895 46746 929
rect 46680 877 46746 895
rect 46915 1055 46951 1071
rect 46915 1021 46917 1055
rect 46915 987 46951 1021
rect 46915 953 46917 987
rect 46987 1055 47053 1105
rect 47228 1099 47257 1133
rect 47291 1099 47349 1133
rect 47383 1099 47441 1133
rect 47475 1099 47504 1133
rect 47604 1109 47620 1143
rect 47654 1109 47670 1143
rect 47828 1130 47942 1132
rect 46987 1021 47003 1055
rect 47037 1021 47053 1055
rect 46987 987 47053 1021
rect 46987 953 47003 987
rect 47037 953 47053 987
rect 47087 1055 47141 1071
rect 47087 1021 47089 1055
rect 47123 1021 47141 1055
rect 47087 974 47141 1021
rect 46915 919 46951 953
rect 47087 940 47089 974
rect 47123 940 47141 974
rect 46915 885 47050 919
rect 47087 890 47141 940
rect 46422 858 46456 877
rect 46096 819 46130 821
rect 46508 843 46652 844
rect 46508 829 46666 843
rect 46096 783 46130 785
rect 46362 816 46428 818
rect 46508 816 46616 829
rect 46362 815 46616 816
rect 46362 781 46378 815
rect 46412 802 46616 815
rect 46412 782 46548 802
rect 46600 795 46616 802
rect 46650 795 46666 829
rect 46412 781 46428 782
rect 46600 745 46646 761
rect 46700 757 46746 877
rect 47016 856 47050 885
rect 46903 827 46971 849
rect 46903 826 46919 827
rect 46903 792 46917 826
rect 46953 793 46971 827
rect 46951 792 46971 793
rect 46903 775 46971 792
rect 47016 840 47071 856
rect 47016 806 47037 840
rect 47016 790 47071 806
rect 47105 840 47141 890
rect 47296 1057 47338 1099
rect 47828 1091 48110 1130
rect 48250 1109 48266 1143
rect 48300 1109 48316 1143
rect 47828 1066 47867 1091
rect 47296 1023 47304 1057
rect 47296 989 47338 1023
rect 47296 955 47304 989
rect 47296 921 47338 955
rect 47296 887 47304 921
rect 47296 871 47338 887
rect 47372 1057 47438 1065
rect 47372 1023 47388 1057
rect 47422 1023 47438 1057
rect 47372 989 47438 1023
rect 47372 955 47388 989
rect 47422 955 47438 989
rect 47372 921 47438 955
rect 47372 887 47388 921
rect 47422 887 47438 921
rect 47372 869 47438 887
rect 47105 838 47146 840
rect 47105 804 47110 838
rect 47144 804 47146 838
rect 47105 802 47146 804
rect 47292 832 47358 835
rect 46130 717 46376 734
rect 46096 700 46376 717
rect 46096 698 46130 700
rect 45484 669 45826 690
rect 45484 635 45500 669
rect 45534 658 45826 669
rect 45534 655 46002 658
rect 45534 654 45952 655
rect 45534 635 45556 654
rect 45484 630 45556 635
rect 45484 623 45550 630
rect 45790 622 45952 654
rect 45936 621 45952 622
rect 45986 621 46002 655
rect 46328 612 46376 700
rect 45340 555 45369 589
rect 45403 555 45461 589
rect 45495 555 45553 589
rect 45587 555 45616 589
rect 45698 584 45744 594
rect 45698 550 45704 584
rect 45738 564 45744 584
rect 46328 578 46336 612
rect 46370 578 46376 612
rect 46600 711 46612 745
rect 46600 677 46646 711
rect 46600 643 46612 677
rect 46600 597 46646 643
rect 46680 745 46746 757
rect 46680 694 46696 745
rect 46730 694 46746 745
rect 47016 739 47050 790
rect 46680 677 46746 694
rect 46680 643 46696 677
rect 46730 643 46746 677
rect 46680 631 46746 643
rect 46917 705 47050 739
rect 47105 730 47141 802
rect 47292 798 47306 832
rect 47340 821 47358 832
rect 47292 787 47308 798
rect 47342 787 47358 821
rect 46917 684 46951 705
rect 47089 701 47141 730
rect 46917 629 46951 650
rect 46987 637 47003 671
rect 47037 637 47053 671
rect 45738 550 45748 564
rect 42342 420 42376 454
rect 42342 368 42376 384
rect 43734 444 43866 480
rect 44038 490 44072 506
rect 44134 490 44168 506
rect 44072 454 44073 455
rect 43734 396 43770 444
rect 44038 420 44073 454
rect 44072 418 44073 420
rect 44134 420 44168 454
rect 43918 396 44038 418
rect 43734 384 44038 396
rect 44072 384 44074 418
rect 43734 382 44074 384
rect 43734 360 43954 382
rect 44038 368 44072 382
rect 44134 368 44168 384
rect 44230 490 44264 506
rect 45698 480 45748 550
rect 46048 540 46064 574
rect 46098 540 46114 574
rect 46328 566 46376 578
rect 46536 563 46565 597
rect 46599 563 46657 597
rect 46691 563 46749 597
rect 46783 563 46812 597
rect 46987 595 47053 637
rect 47123 667 47141 701
rect 47089 629 47141 667
rect 47292 737 47338 753
rect 47392 749 47438 869
rect 47576 1047 47610 1066
rect 47662 1057 47867 1066
rect 47901 1089 48110 1091
rect 47901 1057 47986 1089
rect 47662 1055 47986 1057
rect 48020 1066 48110 1089
rect 48350 1066 48384 1424
rect 49294 1398 49328 1609
rect 49525 1306 49559 1609
rect 49610 1390 49644 2004
rect 49810 2002 49876 2004
rect 50127 2009 50143 2043
rect 50177 2009 50193 2043
rect 50127 1975 50193 2009
rect 49682 1943 49716 1962
rect 49682 1875 49716 1877
rect 49682 1839 49716 1841
rect 49682 1754 49716 1773
rect 49778 1943 49812 1962
rect 49778 1875 49812 1877
rect 49778 1839 49812 1841
rect 49778 1754 49812 1773
rect 49874 1943 49908 1962
rect 50127 1941 50143 1975
rect 50177 1959 50193 1975
rect 50299 2111 50365 2153
rect 50333 2077 50365 2111
rect 50299 2043 50365 2077
rect 50333 2009 50365 2043
rect 50299 1975 50365 2009
rect 50177 1941 50263 1959
rect 50127 1925 50263 1941
rect 50333 1941 50365 1975
rect 50299 1925 50365 1941
rect 51201 2111 51267 2116
rect 51201 2077 51217 2111
rect 51251 2077 51267 2111
rect 51201 2043 51267 2077
rect 51201 2009 51217 2043
rect 51251 2009 51267 2043
rect 51201 1975 51267 2009
rect 51201 1941 51217 1975
rect 51251 1959 51267 1975
rect 51373 2111 51439 2153
rect 51407 2077 51439 2111
rect 51606 2147 51888 2153
rect 51606 2113 51645 2147
rect 51679 2145 51888 2147
rect 51679 2113 51764 2145
rect 51606 2111 51764 2113
rect 51798 2111 51888 2145
rect 51606 2078 51888 2111
rect 52015 2111 52081 2116
rect 51373 2043 51439 2077
rect 51407 2009 51439 2043
rect 52015 2077 52031 2111
rect 52065 2077 52081 2111
rect 52015 2043 52081 2077
rect 51373 1975 51439 2009
rect 51251 1941 51337 1959
rect 51201 1925 51337 1941
rect 51407 1941 51439 1975
rect 51373 1925 51439 1941
rect 51498 2039 51764 2040
rect 51498 2005 51714 2039
rect 51748 2005 51764 2039
rect 51498 2004 51764 2005
rect 49874 1875 49908 1877
rect 50125 1882 50195 1891
rect 50125 1848 50141 1882
rect 50175 1875 50195 1882
rect 50125 1841 50145 1848
rect 50179 1841 50195 1875
rect 49874 1839 49908 1841
rect 50229 1805 50263 1925
rect 50297 1882 50367 1891
rect 50297 1875 50315 1882
rect 50297 1841 50313 1875
rect 50349 1848 50367 1882
rect 50347 1841 50367 1848
rect 51199 1884 51269 1891
rect 51199 1850 51217 1884
rect 51251 1875 51269 1884
rect 51199 1841 51219 1850
rect 51253 1841 51269 1875
rect 51303 1805 51337 1925
rect 51371 1880 51441 1891
rect 51371 1875 51390 1880
rect 51371 1841 51387 1875
rect 51424 1846 51441 1880
rect 51421 1841 51441 1846
rect 49874 1754 49908 1773
rect 50129 1789 50177 1805
rect 50129 1755 50143 1789
rect 50129 1721 50177 1755
rect 49714 1677 49730 1711
rect 49764 1677 49780 1711
rect 50129 1687 50143 1721
rect 50129 1643 50177 1687
rect 50211 1789 50277 1805
rect 50211 1755 50227 1789
rect 50261 1759 50277 1789
rect 50211 1725 50229 1755
rect 50263 1725 50277 1759
rect 50211 1721 50277 1725
rect 50211 1687 50227 1721
rect 50261 1687 50277 1721
rect 50211 1677 50277 1687
rect 50311 1789 50365 1805
rect 50345 1755 50365 1789
rect 50311 1721 50365 1755
rect 50345 1687 50365 1721
rect 50311 1643 50365 1687
rect 51203 1789 51251 1805
rect 51203 1755 51217 1789
rect 51203 1721 51251 1755
rect 51203 1687 51217 1721
rect 51203 1643 51251 1687
rect 51285 1789 51351 1805
rect 51285 1764 51301 1789
rect 51285 1730 51299 1764
rect 51335 1755 51351 1789
rect 51333 1730 51351 1755
rect 51285 1721 51351 1730
rect 51285 1687 51301 1721
rect 51335 1687 51351 1721
rect 51285 1677 51351 1687
rect 51385 1789 51439 1805
rect 51419 1755 51439 1789
rect 51385 1721 51439 1755
rect 51419 1687 51439 1721
rect 51385 1643 51439 1687
rect 49826 1596 49842 1630
rect 49876 1596 49892 1630
rect 50108 1609 50137 1643
rect 50171 1609 50229 1643
rect 50263 1609 50321 1643
rect 50355 1609 50384 1643
rect 51182 1609 51211 1643
rect 51245 1609 51303 1643
rect 51337 1609 51395 1643
rect 51429 1609 51458 1643
rect 49698 1546 49732 1562
rect 49698 1476 49732 1510
rect 49698 1424 49732 1440
rect 49794 1546 49828 1562
rect 49794 1476 49828 1510
rect 49794 1424 49828 1440
rect 49890 1546 49924 1562
rect 49890 1476 49924 1510
rect 49924 1440 50272 1464
rect 49890 1424 50272 1440
rect 49610 1356 49746 1390
rect 49780 1356 49796 1390
rect 49525 1286 49920 1306
rect 49525 1281 49787 1286
rect 49525 1272 49666 1281
rect 49650 1247 49666 1272
rect 49700 1252 49787 1281
rect 49821 1262 49920 1286
rect 50092 1264 50138 1266
rect 50092 1262 50096 1264
rect 49821 1252 50096 1262
rect 49700 1247 50096 1252
rect 49650 1230 50096 1247
rect 50130 1230 50138 1264
rect 49650 1228 50138 1230
rect 50092 1222 50138 1228
rect 48424 1107 48453 1141
rect 48487 1107 48545 1141
rect 48579 1107 48637 1141
rect 48671 1107 48700 1141
rect 48020 1055 48256 1066
rect 47662 1047 48256 1055
rect 47662 1022 47664 1047
rect 47576 979 47610 981
rect 47576 943 47610 945
rect 47576 858 47610 877
rect 47698 1022 48222 1047
rect 48308 1047 48384 1066
rect 48308 1026 48310 1047
rect 47664 979 47698 981
rect 47920 949 47936 983
rect 47970 949 47986 983
rect 48222 979 48256 981
rect 47664 943 47698 945
rect 48222 943 48256 945
rect 47664 858 47698 877
rect 47792 887 47826 906
rect 47792 819 47826 821
rect 47604 781 47620 815
rect 47654 781 47670 815
rect 47792 783 47826 785
rect 47292 703 47304 737
rect 47292 669 47338 703
rect 47292 635 47304 669
rect 46882 561 46911 595
rect 46945 561 47003 595
rect 47037 561 47095 595
rect 47129 561 47158 595
rect 47292 589 47338 635
rect 47372 737 47438 749
rect 47372 703 47388 737
rect 47422 703 47438 737
rect 47372 690 47438 703
rect 47792 698 47826 717
rect 47888 887 47922 906
rect 47888 819 47922 821
rect 47888 783 47922 785
rect 47888 698 47922 717
rect 47984 887 48018 906
rect 48222 858 48256 877
rect 48344 1026 48384 1047
rect 48492 1065 48534 1107
rect 48770 1105 48799 1139
rect 48833 1105 48891 1139
rect 48925 1105 48983 1139
rect 49017 1105 49046 1139
rect 49191 1133 49225 1140
rect 48492 1031 48500 1065
rect 48310 979 48344 981
rect 48310 943 48344 945
rect 48492 997 48534 1031
rect 48492 963 48500 997
rect 48492 929 48534 963
rect 48492 895 48500 929
rect 48492 879 48534 895
rect 48568 1065 48634 1073
rect 48568 1031 48584 1065
rect 48618 1031 48634 1065
rect 48568 997 48634 1031
rect 48568 963 48584 997
rect 48618 963 48634 997
rect 48568 929 48634 963
rect 48568 895 48584 929
rect 48618 895 48634 929
rect 48568 877 48634 895
rect 48803 1055 48839 1071
rect 48803 1021 48805 1055
rect 48803 987 48839 1021
rect 48803 953 48805 987
rect 48875 1055 48941 1105
rect 49116 1099 49145 1133
rect 49179 1099 49237 1133
rect 49271 1099 49329 1133
rect 49363 1099 49392 1133
rect 49492 1109 49508 1143
rect 49542 1109 49558 1143
rect 49716 1130 49830 1132
rect 48875 1021 48891 1055
rect 48925 1021 48941 1055
rect 48875 987 48941 1021
rect 48875 953 48891 987
rect 48925 953 48941 987
rect 48975 1055 49029 1071
rect 48975 1021 48977 1055
rect 49011 1021 49029 1055
rect 48975 974 49029 1021
rect 48803 919 48839 953
rect 48975 940 48977 974
rect 49011 940 49029 974
rect 48803 885 48938 919
rect 48975 890 49029 940
rect 48310 858 48344 877
rect 47984 819 48018 821
rect 48396 843 48540 844
rect 48396 829 48554 843
rect 47984 783 48018 785
rect 48250 816 48316 818
rect 48396 816 48504 829
rect 48250 815 48504 816
rect 48250 781 48266 815
rect 48300 802 48504 815
rect 48300 782 48436 802
rect 48488 795 48504 802
rect 48538 795 48554 829
rect 48300 781 48316 782
rect 48488 745 48534 761
rect 48588 757 48634 877
rect 48904 856 48938 885
rect 48791 827 48859 849
rect 48791 826 48807 827
rect 48791 792 48805 826
rect 48841 793 48859 827
rect 48839 792 48859 793
rect 48791 775 48859 792
rect 48904 840 48959 856
rect 48904 806 48925 840
rect 48904 790 48959 806
rect 48993 840 49029 890
rect 49184 1057 49226 1099
rect 49716 1091 49998 1130
rect 50138 1109 50154 1143
rect 50188 1109 50204 1143
rect 49716 1066 49755 1091
rect 49184 1023 49192 1057
rect 49184 989 49226 1023
rect 49184 955 49192 989
rect 49184 921 49226 955
rect 49184 887 49192 921
rect 49184 871 49226 887
rect 49260 1057 49326 1065
rect 49260 1023 49276 1057
rect 49310 1023 49326 1057
rect 49260 989 49326 1023
rect 49260 955 49276 989
rect 49310 955 49326 989
rect 49260 921 49326 955
rect 49260 887 49276 921
rect 49310 887 49326 921
rect 49260 869 49326 887
rect 48993 838 49034 840
rect 48993 804 48998 838
rect 49032 804 49034 838
rect 48993 802 49034 804
rect 49180 832 49246 835
rect 48018 717 48264 734
rect 47984 700 48264 717
rect 47984 698 48018 700
rect 47372 669 47714 690
rect 47372 635 47388 669
rect 47422 658 47714 669
rect 47422 655 47890 658
rect 47422 654 47840 655
rect 47422 635 47444 654
rect 47372 630 47444 635
rect 47372 623 47438 630
rect 47678 622 47840 654
rect 47824 621 47840 622
rect 47874 621 47890 655
rect 48216 612 48264 700
rect 47228 555 47257 589
rect 47291 555 47349 589
rect 47383 555 47441 589
rect 47475 555 47504 589
rect 47586 584 47632 594
rect 47586 550 47592 584
rect 47626 564 47632 584
rect 48216 578 48224 612
rect 48258 578 48264 612
rect 48488 711 48500 745
rect 48488 677 48534 711
rect 48488 643 48500 677
rect 48488 597 48534 643
rect 48568 745 48634 757
rect 48568 694 48584 745
rect 48618 694 48634 745
rect 48904 739 48938 790
rect 48568 677 48634 694
rect 48568 643 48584 677
rect 48618 643 48634 677
rect 48568 631 48634 643
rect 48805 705 48938 739
rect 48993 730 49029 802
rect 49180 798 49194 832
rect 49228 821 49246 832
rect 49180 787 49196 798
rect 49230 787 49246 821
rect 48805 684 48839 705
rect 48977 701 49029 730
rect 48805 629 48839 650
rect 48875 637 48891 671
rect 48925 637 48941 671
rect 47626 550 47636 564
rect 44230 420 44264 454
rect 44230 368 44264 384
rect 45616 444 45748 480
rect 45920 490 45954 506
rect 46016 490 46050 506
rect 45954 454 45955 455
rect 45616 396 45652 444
rect 45920 420 45955 454
rect 45954 418 45955 420
rect 46016 420 46050 454
rect 45800 396 45920 418
rect 45616 384 45920 396
rect 45954 384 45956 418
rect 45616 382 45956 384
rect 45616 360 45836 382
rect 45920 368 45954 382
rect 46016 368 46050 384
rect 46112 490 46146 506
rect 47586 480 47636 550
rect 47936 540 47952 574
rect 47986 540 48002 574
rect 48216 566 48264 578
rect 48424 563 48453 597
rect 48487 563 48545 597
rect 48579 563 48637 597
rect 48671 563 48700 597
rect 48875 595 48941 637
rect 49011 667 49029 701
rect 48977 629 49029 667
rect 49180 737 49226 753
rect 49280 749 49326 869
rect 49464 1047 49498 1066
rect 49550 1057 49755 1066
rect 49789 1089 49998 1091
rect 49789 1057 49874 1089
rect 49550 1055 49874 1057
rect 49908 1066 49998 1089
rect 50238 1066 50272 1424
rect 51182 1398 51216 1609
rect 51413 1306 51447 1609
rect 51498 1390 51532 2004
rect 51698 2002 51764 2004
rect 52015 2009 52031 2043
rect 52065 2009 52081 2043
rect 52015 1975 52081 2009
rect 51570 1943 51604 1962
rect 51570 1875 51604 1877
rect 51570 1839 51604 1841
rect 51570 1754 51604 1773
rect 51666 1943 51700 1962
rect 51666 1875 51700 1877
rect 51666 1839 51700 1841
rect 51666 1754 51700 1773
rect 51762 1943 51796 1962
rect 52015 1941 52031 1975
rect 52065 1959 52081 1975
rect 52187 2111 52253 2153
rect 52221 2077 52253 2111
rect 52187 2043 52253 2077
rect 52221 2009 52253 2043
rect 52187 1975 52253 2009
rect 52065 1941 52151 1959
rect 52015 1925 52151 1941
rect 52221 1941 52253 1975
rect 52187 1925 52253 1941
rect 53089 2111 53155 2116
rect 53089 2077 53105 2111
rect 53139 2077 53155 2111
rect 53089 2043 53155 2077
rect 53089 2009 53105 2043
rect 53139 2009 53155 2043
rect 53089 1975 53155 2009
rect 53089 1941 53105 1975
rect 53139 1959 53155 1975
rect 53261 2111 53327 2153
rect 53295 2077 53327 2111
rect 53494 2147 53776 2153
rect 53494 2113 53533 2147
rect 53567 2145 53776 2147
rect 53567 2113 53652 2145
rect 53494 2111 53652 2113
rect 53686 2111 53776 2145
rect 53494 2078 53776 2111
rect 53903 2111 53969 2116
rect 53261 2043 53327 2077
rect 53295 2009 53327 2043
rect 53903 2077 53919 2111
rect 53953 2077 53969 2111
rect 53903 2043 53969 2077
rect 53261 1975 53327 2009
rect 53139 1941 53225 1959
rect 53089 1925 53225 1941
rect 53295 1941 53327 1975
rect 53261 1925 53327 1941
rect 53386 2039 53652 2040
rect 53386 2005 53602 2039
rect 53636 2005 53652 2039
rect 53386 2004 53652 2005
rect 51762 1875 51796 1877
rect 52013 1882 52083 1891
rect 52013 1848 52029 1882
rect 52063 1875 52083 1882
rect 52013 1841 52033 1848
rect 52067 1841 52083 1875
rect 51762 1839 51796 1841
rect 52117 1805 52151 1925
rect 52185 1882 52255 1891
rect 52185 1875 52203 1882
rect 52185 1841 52201 1875
rect 52237 1848 52255 1882
rect 52235 1841 52255 1848
rect 53087 1884 53157 1891
rect 53087 1850 53105 1884
rect 53139 1875 53157 1884
rect 53087 1841 53107 1850
rect 53141 1841 53157 1875
rect 53191 1805 53225 1925
rect 53259 1880 53329 1891
rect 53259 1875 53278 1880
rect 53259 1841 53275 1875
rect 53312 1846 53329 1880
rect 53309 1841 53329 1846
rect 51762 1754 51796 1773
rect 52017 1789 52065 1805
rect 52017 1755 52031 1789
rect 52017 1721 52065 1755
rect 51602 1677 51618 1711
rect 51652 1677 51668 1711
rect 52017 1687 52031 1721
rect 52017 1643 52065 1687
rect 52099 1789 52165 1805
rect 52099 1755 52115 1789
rect 52149 1759 52165 1789
rect 52099 1725 52117 1755
rect 52151 1725 52165 1759
rect 52099 1721 52165 1725
rect 52099 1687 52115 1721
rect 52149 1687 52165 1721
rect 52099 1677 52165 1687
rect 52199 1789 52253 1805
rect 52233 1755 52253 1789
rect 52199 1721 52253 1755
rect 52233 1687 52253 1721
rect 52199 1643 52253 1687
rect 53091 1789 53139 1805
rect 53091 1755 53105 1789
rect 53091 1721 53139 1755
rect 53091 1687 53105 1721
rect 53091 1643 53139 1687
rect 53173 1789 53239 1805
rect 53173 1764 53189 1789
rect 53173 1730 53187 1764
rect 53223 1755 53239 1789
rect 53221 1730 53239 1755
rect 53173 1721 53239 1730
rect 53173 1687 53189 1721
rect 53223 1687 53239 1721
rect 53173 1677 53239 1687
rect 53273 1789 53327 1805
rect 53307 1755 53327 1789
rect 53273 1721 53327 1755
rect 53307 1687 53327 1721
rect 53273 1643 53327 1687
rect 51714 1596 51730 1630
rect 51764 1596 51780 1630
rect 51996 1609 52025 1643
rect 52059 1609 52117 1643
rect 52151 1609 52209 1643
rect 52243 1609 52272 1643
rect 53070 1609 53099 1643
rect 53133 1609 53191 1643
rect 53225 1609 53283 1643
rect 53317 1609 53346 1643
rect 51586 1546 51620 1562
rect 51586 1476 51620 1510
rect 51586 1424 51620 1440
rect 51682 1546 51716 1562
rect 51682 1476 51716 1510
rect 51682 1424 51716 1440
rect 51778 1546 51812 1562
rect 51778 1476 51812 1510
rect 51812 1440 52160 1464
rect 51778 1424 52160 1440
rect 51498 1356 51634 1390
rect 51668 1356 51684 1390
rect 51413 1286 51808 1306
rect 51413 1281 51675 1286
rect 51413 1272 51554 1281
rect 51538 1247 51554 1272
rect 51588 1252 51675 1281
rect 51709 1262 51808 1286
rect 51980 1264 52026 1266
rect 51980 1262 51984 1264
rect 51709 1252 51984 1262
rect 51588 1247 51984 1252
rect 51538 1230 51984 1247
rect 52018 1230 52026 1264
rect 51538 1228 52026 1230
rect 51980 1222 52026 1228
rect 50312 1107 50341 1141
rect 50375 1107 50433 1141
rect 50467 1107 50525 1141
rect 50559 1107 50588 1141
rect 49908 1055 50144 1066
rect 49550 1047 50144 1055
rect 49550 1022 49552 1047
rect 49464 979 49498 981
rect 49464 943 49498 945
rect 49464 858 49498 877
rect 49586 1022 50110 1047
rect 50196 1047 50272 1066
rect 50196 1026 50198 1047
rect 49552 979 49586 981
rect 49808 949 49824 983
rect 49858 949 49874 983
rect 50110 979 50144 981
rect 49552 943 49586 945
rect 50110 943 50144 945
rect 49552 858 49586 877
rect 49680 887 49714 906
rect 49680 819 49714 821
rect 49492 781 49508 815
rect 49542 781 49558 815
rect 49680 783 49714 785
rect 49180 703 49192 737
rect 49180 669 49226 703
rect 49180 635 49192 669
rect 48770 561 48799 595
rect 48833 561 48891 595
rect 48925 561 48983 595
rect 49017 561 49046 595
rect 49180 589 49226 635
rect 49260 737 49326 749
rect 49260 703 49276 737
rect 49310 703 49326 737
rect 49260 690 49326 703
rect 49680 698 49714 717
rect 49776 887 49810 906
rect 49776 819 49810 821
rect 49776 783 49810 785
rect 49776 698 49810 717
rect 49872 887 49906 906
rect 50110 858 50144 877
rect 50232 1026 50272 1047
rect 50380 1065 50422 1107
rect 50658 1105 50687 1139
rect 50721 1105 50779 1139
rect 50813 1105 50871 1139
rect 50905 1105 50934 1139
rect 51079 1133 51113 1140
rect 50380 1031 50388 1065
rect 50198 979 50232 981
rect 50198 943 50232 945
rect 50380 997 50422 1031
rect 50380 963 50388 997
rect 50380 929 50422 963
rect 50380 895 50388 929
rect 50380 879 50422 895
rect 50456 1065 50522 1073
rect 50456 1031 50472 1065
rect 50506 1031 50522 1065
rect 50456 997 50522 1031
rect 50456 963 50472 997
rect 50506 963 50522 997
rect 50456 929 50522 963
rect 50456 895 50472 929
rect 50506 895 50522 929
rect 50456 877 50522 895
rect 50691 1055 50727 1071
rect 50691 1021 50693 1055
rect 50691 987 50727 1021
rect 50691 953 50693 987
rect 50763 1055 50829 1105
rect 51004 1099 51033 1133
rect 51067 1099 51125 1133
rect 51159 1099 51217 1133
rect 51251 1099 51280 1133
rect 51380 1109 51396 1143
rect 51430 1109 51446 1143
rect 51604 1130 51718 1132
rect 50763 1021 50779 1055
rect 50813 1021 50829 1055
rect 50763 987 50829 1021
rect 50763 953 50779 987
rect 50813 953 50829 987
rect 50863 1055 50917 1071
rect 50863 1021 50865 1055
rect 50899 1021 50917 1055
rect 50863 974 50917 1021
rect 50691 919 50727 953
rect 50863 940 50865 974
rect 50899 940 50917 974
rect 50691 885 50826 919
rect 50863 890 50917 940
rect 50198 858 50232 877
rect 49872 819 49906 821
rect 50284 843 50428 844
rect 50284 829 50442 843
rect 49872 783 49906 785
rect 50138 816 50204 818
rect 50284 816 50392 829
rect 50138 815 50392 816
rect 50138 781 50154 815
rect 50188 802 50392 815
rect 50188 782 50324 802
rect 50376 795 50392 802
rect 50426 795 50442 829
rect 50188 781 50204 782
rect 50376 745 50422 761
rect 50476 757 50522 877
rect 50792 856 50826 885
rect 50679 827 50747 849
rect 50679 826 50695 827
rect 50679 792 50693 826
rect 50729 793 50747 827
rect 50727 792 50747 793
rect 50679 775 50747 792
rect 50792 840 50847 856
rect 50792 806 50813 840
rect 50792 790 50847 806
rect 50881 840 50917 890
rect 51072 1057 51114 1099
rect 51604 1091 51886 1130
rect 52026 1109 52042 1143
rect 52076 1109 52092 1143
rect 51604 1066 51643 1091
rect 51072 1023 51080 1057
rect 51072 989 51114 1023
rect 51072 955 51080 989
rect 51072 921 51114 955
rect 51072 887 51080 921
rect 51072 871 51114 887
rect 51148 1057 51214 1065
rect 51148 1023 51164 1057
rect 51198 1023 51214 1057
rect 51148 989 51214 1023
rect 51148 955 51164 989
rect 51198 955 51214 989
rect 51148 921 51214 955
rect 51148 887 51164 921
rect 51198 887 51214 921
rect 51148 869 51214 887
rect 50881 838 50922 840
rect 50881 804 50886 838
rect 50920 804 50922 838
rect 50881 802 50922 804
rect 51068 832 51134 835
rect 49906 717 50152 734
rect 49872 700 50152 717
rect 49872 698 49906 700
rect 49260 669 49602 690
rect 49260 635 49276 669
rect 49310 658 49602 669
rect 49310 655 49778 658
rect 49310 654 49728 655
rect 49310 635 49332 654
rect 49260 630 49332 635
rect 49260 623 49326 630
rect 49566 622 49728 654
rect 49712 621 49728 622
rect 49762 621 49778 655
rect 50104 612 50152 700
rect 49116 555 49145 589
rect 49179 555 49237 589
rect 49271 555 49329 589
rect 49363 555 49392 589
rect 49474 584 49520 594
rect 49474 550 49480 584
rect 49514 564 49520 584
rect 50104 578 50112 612
rect 50146 578 50152 612
rect 50376 711 50388 745
rect 50376 677 50422 711
rect 50376 643 50388 677
rect 50376 597 50422 643
rect 50456 745 50522 757
rect 50456 694 50472 745
rect 50506 694 50522 745
rect 50792 739 50826 790
rect 50456 677 50522 694
rect 50456 643 50472 677
rect 50506 643 50522 677
rect 50456 631 50522 643
rect 50693 705 50826 739
rect 50881 730 50917 802
rect 51068 798 51082 832
rect 51116 821 51134 832
rect 51068 787 51084 798
rect 51118 787 51134 821
rect 50693 684 50727 705
rect 50865 701 50917 730
rect 50693 629 50727 650
rect 50763 637 50779 671
rect 50813 637 50829 671
rect 49514 550 49524 564
rect 46112 420 46146 454
rect 46112 368 46146 384
rect 47504 444 47636 480
rect 47808 490 47842 506
rect 47904 490 47938 506
rect 47842 454 47843 455
rect 47504 396 47540 444
rect 47808 420 47843 454
rect 47842 418 47843 420
rect 47904 420 47938 454
rect 47688 396 47808 418
rect 47504 384 47808 396
rect 47842 384 47844 418
rect 47504 382 47844 384
rect 47504 360 47724 382
rect 47808 368 47842 382
rect 47904 368 47938 384
rect 48000 490 48034 506
rect 49474 480 49524 550
rect 49824 540 49840 574
rect 49874 540 49890 574
rect 50104 566 50152 578
rect 50312 563 50341 597
rect 50375 563 50433 597
rect 50467 563 50525 597
rect 50559 563 50588 597
rect 50763 595 50829 637
rect 50899 667 50917 701
rect 50865 629 50917 667
rect 51068 737 51114 753
rect 51168 749 51214 869
rect 51352 1047 51386 1066
rect 51438 1057 51643 1066
rect 51677 1089 51886 1091
rect 51677 1057 51762 1089
rect 51438 1055 51762 1057
rect 51796 1066 51886 1089
rect 52126 1066 52160 1424
rect 53070 1398 53104 1609
rect 53301 1306 53335 1609
rect 53386 1390 53420 2004
rect 53586 2002 53652 2004
rect 53903 2009 53919 2043
rect 53953 2009 53969 2043
rect 53903 1975 53969 2009
rect 53458 1943 53492 1962
rect 53458 1875 53492 1877
rect 53458 1839 53492 1841
rect 53458 1754 53492 1773
rect 53554 1943 53588 1962
rect 53554 1875 53588 1877
rect 53554 1839 53588 1841
rect 53554 1754 53588 1773
rect 53650 1943 53684 1962
rect 53903 1941 53919 1975
rect 53953 1959 53969 1975
rect 54075 2111 54141 2153
rect 54109 2077 54141 2111
rect 54075 2043 54141 2077
rect 54109 2009 54141 2043
rect 54075 1975 54141 2009
rect 53953 1941 54039 1959
rect 53903 1925 54039 1941
rect 54109 1941 54141 1975
rect 54075 1925 54141 1941
rect 54977 2111 55043 2116
rect 54977 2077 54993 2111
rect 55027 2077 55043 2111
rect 54977 2043 55043 2077
rect 54977 2009 54993 2043
rect 55027 2009 55043 2043
rect 54977 1975 55043 2009
rect 54977 1941 54993 1975
rect 55027 1959 55043 1975
rect 55149 2111 55215 2153
rect 55183 2077 55215 2111
rect 55382 2147 55664 2153
rect 55382 2113 55421 2147
rect 55455 2145 55664 2147
rect 55455 2113 55540 2145
rect 55382 2111 55540 2113
rect 55574 2111 55664 2145
rect 55382 2078 55664 2111
rect 55791 2111 55857 2116
rect 55149 2043 55215 2077
rect 55183 2009 55215 2043
rect 55791 2077 55807 2111
rect 55841 2077 55857 2111
rect 55791 2043 55857 2077
rect 55149 1975 55215 2009
rect 55027 1941 55113 1959
rect 54977 1925 55113 1941
rect 55183 1941 55215 1975
rect 55149 1925 55215 1941
rect 55274 2039 55540 2040
rect 55274 2005 55490 2039
rect 55524 2005 55540 2039
rect 55274 2004 55540 2005
rect 53650 1875 53684 1877
rect 53901 1882 53971 1891
rect 53901 1848 53917 1882
rect 53951 1875 53971 1882
rect 53901 1841 53921 1848
rect 53955 1841 53971 1875
rect 53650 1839 53684 1841
rect 54005 1805 54039 1925
rect 54073 1882 54143 1891
rect 54073 1875 54091 1882
rect 54073 1841 54089 1875
rect 54125 1848 54143 1882
rect 54123 1841 54143 1848
rect 54975 1884 55045 1891
rect 54975 1850 54993 1884
rect 55027 1875 55045 1884
rect 54975 1841 54995 1850
rect 55029 1841 55045 1875
rect 55079 1805 55113 1925
rect 55147 1880 55217 1891
rect 55147 1875 55166 1880
rect 55147 1841 55163 1875
rect 55200 1846 55217 1880
rect 55197 1841 55217 1846
rect 53650 1754 53684 1773
rect 53905 1789 53953 1805
rect 53905 1755 53919 1789
rect 53905 1721 53953 1755
rect 53490 1677 53506 1711
rect 53540 1677 53556 1711
rect 53905 1687 53919 1721
rect 53905 1643 53953 1687
rect 53987 1789 54053 1805
rect 53987 1755 54003 1789
rect 54037 1759 54053 1789
rect 53987 1725 54005 1755
rect 54039 1725 54053 1759
rect 53987 1721 54053 1725
rect 53987 1687 54003 1721
rect 54037 1687 54053 1721
rect 53987 1677 54053 1687
rect 54087 1789 54141 1805
rect 54121 1755 54141 1789
rect 54087 1721 54141 1755
rect 54121 1687 54141 1721
rect 54087 1643 54141 1687
rect 54979 1789 55027 1805
rect 54979 1755 54993 1789
rect 54979 1721 55027 1755
rect 54979 1687 54993 1721
rect 54979 1643 55027 1687
rect 55061 1789 55127 1805
rect 55061 1764 55077 1789
rect 55061 1730 55075 1764
rect 55111 1755 55127 1789
rect 55109 1730 55127 1755
rect 55061 1721 55127 1730
rect 55061 1687 55077 1721
rect 55111 1687 55127 1721
rect 55061 1677 55127 1687
rect 55161 1789 55215 1805
rect 55195 1755 55215 1789
rect 55161 1721 55215 1755
rect 55195 1687 55215 1721
rect 55161 1643 55215 1687
rect 53602 1596 53618 1630
rect 53652 1596 53668 1630
rect 53884 1609 53913 1643
rect 53947 1609 54005 1643
rect 54039 1609 54097 1643
rect 54131 1609 54160 1643
rect 54958 1609 54987 1643
rect 55021 1609 55079 1643
rect 55113 1609 55171 1643
rect 55205 1609 55234 1643
rect 53474 1546 53508 1562
rect 53474 1476 53508 1510
rect 53474 1424 53508 1440
rect 53570 1546 53604 1562
rect 53570 1476 53604 1510
rect 53570 1424 53604 1440
rect 53666 1546 53700 1562
rect 53666 1476 53700 1510
rect 53700 1440 54048 1464
rect 53666 1424 54048 1440
rect 53386 1356 53522 1390
rect 53556 1356 53572 1390
rect 53301 1286 53696 1306
rect 53301 1281 53563 1286
rect 53301 1272 53442 1281
rect 53426 1247 53442 1272
rect 53476 1252 53563 1281
rect 53597 1262 53696 1286
rect 53868 1264 53914 1266
rect 53868 1262 53872 1264
rect 53597 1252 53872 1262
rect 53476 1247 53872 1252
rect 53426 1230 53872 1247
rect 53906 1230 53914 1264
rect 53426 1228 53914 1230
rect 53868 1222 53914 1228
rect 52200 1107 52229 1141
rect 52263 1107 52321 1141
rect 52355 1107 52413 1141
rect 52447 1107 52476 1141
rect 51796 1055 52032 1066
rect 51438 1047 52032 1055
rect 51438 1022 51440 1047
rect 51352 979 51386 981
rect 51352 943 51386 945
rect 51352 858 51386 877
rect 51474 1022 51998 1047
rect 52084 1047 52160 1066
rect 52084 1026 52086 1047
rect 51440 979 51474 981
rect 51696 949 51712 983
rect 51746 949 51762 983
rect 51998 979 52032 981
rect 51440 943 51474 945
rect 51998 943 52032 945
rect 51440 858 51474 877
rect 51568 887 51602 906
rect 51568 819 51602 821
rect 51380 781 51396 815
rect 51430 781 51446 815
rect 51568 783 51602 785
rect 51068 703 51080 737
rect 51068 669 51114 703
rect 51068 635 51080 669
rect 50658 561 50687 595
rect 50721 561 50779 595
rect 50813 561 50871 595
rect 50905 561 50934 595
rect 51068 589 51114 635
rect 51148 737 51214 749
rect 51148 703 51164 737
rect 51198 703 51214 737
rect 51148 690 51214 703
rect 51568 698 51602 717
rect 51664 887 51698 906
rect 51664 819 51698 821
rect 51664 783 51698 785
rect 51664 698 51698 717
rect 51760 887 51794 906
rect 51998 858 52032 877
rect 52120 1026 52160 1047
rect 52268 1065 52310 1107
rect 52546 1105 52575 1139
rect 52609 1105 52667 1139
rect 52701 1105 52759 1139
rect 52793 1105 52822 1139
rect 52967 1133 53001 1140
rect 52268 1031 52276 1065
rect 52086 979 52120 981
rect 52086 943 52120 945
rect 52268 997 52310 1031
rect 52268 963 52276 997
rect 52268 929 52310 963
rect 52268 895 52276 929
rect 52268 879 52310 895
rect 52344 1065 52410 1073
rect 52344 1031 52360 1065
rect 52394 1031 52410 1065
rect 52344 997 52410 1031
rect 52344 963 52360 997
rect 52394 963 52410 997
rect 52344 929 52410 963
rect 52344 895 52360 929
rect 52394 895 52410 929
rect 52344 877 52410 895
rect 52579 1055 52615 1071
rect 52579 1021 52581 1055
rect 52579 987 52615 1021
rect 52579 953 52581 987
rect 52651 1055 52717 1105
rect 52892 1099 52921 1133
rect 52955 1099 53013 1133
rect 53047 1099 53105 1133
rect 53139 1099 53168 1133
rect 53268 1109 53284 1143
rect 53318 1109 53334 1143
rect 53492 1130 53606 1132
rect 52651 1021 52667 1055
rect 52701 1021 52717 1055
rect 52651 987 52717 1021
rect 52651 953 52667 987
rect 52701 953 52717 987
rect 52751 1055 52805 1071
rect 52751 1021 52753 1055
rect 52787 1021 52805 1055
rect 52751 974 52805 1021
rect 52579 919 52615 953
rect 52751 940 52753 974
rect 52787 940 52805 974
rect 52579 885 52714 919
rect 52751 890 52805 940
rect 52086 858 52120 877
rect 51760 819 51794 821
rect 52172 843 52316 844
rect 52172 829 52330 843
rect 51760 783 51794 785
rect 52026 816 52092 818
rect 52172 816 52280 829
rect 52026 815 52280 816
rect 52026 781 52042 815
rect 52076 802 52280 815
rect 52076 782 52212 802
rect 52264 795 52280 802
rect 52314 795 52330 829
rect 52076 781 52092 782
rect 52264 745 52310 761
rect 52364 757 52410 877
rect 52680 856 52714 885
rect 52567 827 52635 849
rect 52567 826 52583 827
rect 52567 792 52581 826
rect 52617 793 52635 827
rect 52615 792 52635 793
rect 52567 775 52635 792
rect 52680 840 52735 856
rect 52680 806 52701 840
rect 52680 790 52735 806
rect 52769 840 52805 890
rect 52960 1057 53002 1099
rect 53492 1091 53774 1130
rect 53914 1109 53930 1143
rect 53964 1109 53980 1143
rect 53492 1066 53531 1091
rect 52960 1023 52968 1057
rect 52960 989 53002 1023
rect 52960 955 52968 989
rect 52960 921 53002 955
rect 52960 887 52968 921
rect 52960 871 53002 887
rect 53036 1057 53102 1065
rect 53036 1023 53052 1057
rect 53086 1023 53102 1057
rect 53036 989 53102 1023
rect 53036 955 53052 989
rect 53086 955 53102 989
rect 53036 921 53102 955
rect 53036 887 53052 921
rect 53086 887 53102 921
rect 53036 869 53102 887
rect 52769 838 52810 840
rect 52769 804 52774 838
rect 52808 804 52810 838
rect 52769 802 52810 804
rect 52956 832 53022 835
rect 51794 717 52040 734
rect 51760 700 52040 717
rect 51760 698 51794 700
rect 51148 669 51490 690
rect 51148 635 51164 669
rect 51198 658 51490 669
rect 51198 655 51666 658
rect 51198 654 51616 655
rect 51198 635 51220 654
rect 51148 630 51220 635
rect 51148 623 51214 630
rect 51454 622 51616 654
rect 51600 621 51616 622
rect 51650 621 51666 655
rect 51992 612 52040 700
rect 51004 555 51033 589
rect 51067 555 51125 589
rect 51159 555 51217 589
rect 51251 555 51280 589
rect 51362 584 51408 594
rect 51362 550 51368 584
rect 51402 564 51408 584
rect 51992 578 52000 612
rect 52034 578 52040 612
rect 52264 711 52276 745
rect 52264 677 52310 711
rect 52264 643 52276 677
rect 52264 597 52310 643
rect 52344 745 52410 757
rect 52344 694 52360 745
rect 52394 694 52410 745
rect 52680 739 52714 790
rect 52344 677 52410 694
rect 52344 643 52360 677
rect 52394 643 52410 677
rect 52344 631 52410 643
rect 52581 705 52714 739
rect 52769 730 52805 802
rect 52956 798 52970 832
rect 53004 821 53022 832
rect 52956 787 52972 798
rect 53006 787 53022 821
rect 52581 684 52615 705
rect 52753 701 52805 730
rect 52581 629 52615 650
rect 52651 637 52667 671
rect 52701 637 52717 671
rect 51402 550 51412 564
rect 48000 420 48034 454
rect 48000 368 48034 384
rect 49392 444 49524 480
rect 49696 490 49730 506
rect 49792 490 49826 506
rect 49730 454 49731 455
rect 49392 396 49428 444
rect 49696 420 49731 454
rect 49730 418 49731 420
rect 49792 420 49826 454
rect 49576 396 49696 418
rect 49392 384 49696 396
rect 49730 384 49732 418
rect 49392 382 49732 384
rect 49392 360 49612 382
rect 49696 368 49730 382
rect 49792 368 49826 384
rect 49888 490 49922 506
rect 51362 480 51412 550
rect 51712 540 51728 574
rect 51762 540 51778 574
rect 51992 566 52040 578
rect 52200 563 52229 597
rect 52263 563 52321 597
rect 52355 563 52413 597
rect 52447 563 52476 597
rect 52651 595 52717 637
rect 52787 667 52805 701
rect 52753 629 52805 667
rect 52956 737 53002 753
rect 53056 749 53102 869
rect 53240 1047 53274 1066
rect 53326 1057 53531 1066
rect 53565 1089 53774 1091
rect 53565 1057 53650 1089
rect 53326 1055 53650 1057
rect 53684 1066 53774 1089
rect 54014 1066 54048 1424
rect 54958 1398 54992 1609
rect 55189 1306 55223 1609
rect 55274 1390 55308 2004
rect 55474 2002 55540 2004
rect 55791 2009 55807 2043
rect 55841 2009 55857 2043
rect 55791 1975 55857 2009
rect 55346 1943 55380 1962
rect 55346 1875 55380 1877
rect 55346 1839 55380 1841
rect 55346 1754 55380 1773
rect 55442 1943 55476 1962
rect 55442 1875 55476 1877
rect 55442 1839 55476 1841
rect 55442 1754 55476 1773
rect 55538 1943 55572 1962
rect 55791 1941 55807 1975
rect 55841 1959 55857 1975
rect 55963 2111 56029 2153
rect 55997 2077 56029 2111
rect 55963 2043 56029 2077
rect 55997 2009 56029 2043
rect 55963 1975 56029 2009
rect 55841 1941 55927 1959
rect 55791 1925 55927 1941
rect 55997 1941 56029 1975
rect 55963 1925 56029 1941
rect 56865 2111 56931 2116
rect 56865 2077 56881 2111
rect 56915 2077 56931 2111
rect 56865 2043 56931 2077
rect 56865 2009 56881 2043
rect 56915 2009 56931 2043
rect 56865 1975 56931 2009
rect 56865 1941 56881 1975
rect 56915 1959 56931 1975
rect 57037 2111 57103 2153
rect 57071 2077 57103 2111
rect 57270 2147 57552 2153
rect 57270 2113 57309 2147
rect 57343 2145 57552 2147
rect 57343 2113 57428 2145
rect 57270 2111 57428 2113
rect 57462 2111 57552 2145
rect 57270 2078 57552 2111
rect 57679 2111 57745 2116
rect 57037 2043 57103 2077
rect 57071 2009 57103 2043
rect 57679 2077 57695 2111
rect 57729 2077 57745 2111
rect 57679 2043 57745 2077
rect 57037 1975 57103 2009
rect 56915 1941 57001 1959
rect 56865 1925 57001 1941
rect 57071 1941 57103 1975
rect 57037 1925 57103 1941
rect 57162 2039 57428 2040
rect 57162 2005 57378 2039
rect 57412 2005 57428 2039
rect 57162 2004 57428 2005
rect 55538 1875 55572 1877
rect 55789 1882 55859 1891
rect 55789 1848 55805 1882
rect 55839 1875 55859 1882
rect 55789 1841 55809 1848
rect 55843 1841 55859 1875
rect 55538 1839 55572 1841
rect 55893 1805 55927 1925
rect 55961 1882 56031 1891
rect 55961 1875 55979 1882
rect 55961 1841 55977 1875
rect 56013 1848 56031 1882
rect 56011 1841 56031 1848
rect 56863 1884 56933 1891
rect 56863 1850 56881 1884
rect 56915 1875 56933 1884
rect 56863 1841 56883 1850
rect 56917 1841 56933 1875
rect 56967 1805 57001 1925
rect 57035 1880 57105 1891
rect 57035 1875 57054 1880
rect 57035 1841 57051 1875
rect 57088 1846 57105 1880
rect 57085 1841 57105 1846
rect 55538 1754 55572 1773
rect 55793 1789 55841 1805
rect 55793 1755 55807 1789
rect 55793 1721 55841 1755
rect 55378 1677 55394 1711
rect 55428 1677 55444 1711
rect 55793 1687 55807 1721
rect 55793 1643 55841 1687
rect 55875 1789 55941 1805
rect 55875 1755 55891 1789
rect 55925 1759 55941 1789
rect 55875 1725 55893 1755
rect 55927 1725 55941 1759
rect 55875 1721 55941 1725
rect 55875 1687 55891 1721
rect 55925 1687 55941 1721
rect 55875 1677 55941 1687
rect 55975 1789 56029 1805
rect 56009 1755 56029 1789
rect 55975 1721 56029 1755
rect 56009 1687 56029 1721
rect 55975 1643 56029 1687
rect 56867 1789 56915 1805
rect 56867 1755 56881 1789
rect 56867 1721 56915 1755
rect 56867 1687 56881 1721
rect 56867 1643 56915 1687
rect 56949 1789 57015 1805
rect 56949 1764 56965 1789
rect 56949 1730 56963 1764
rect 56999 1755 57015 1789
rect 56997 1730 57015 1755
rect 56949 1721 57015 1730
rect 56949 1687 56965 1721
rect 56999 1687 57015 1721
rect 56949 1677 57015 1687
rect 57049 1789 57103 1805
rect 57083 1755 57103 1789
rect 57049 1721 57103 1755
rect 57083 1687 57103 1721
rect 57049 1643 57103 1687
rect 55490 1596 55506 1630
rect 55540 1596 55556 1630
rect 55772 1609 55801 1643
rect 55835 1609 55893 1643
rect 55927 1609 55985 1643
rect 56019 1609 56048 1643
rect 56846 1609 56875 1643
rect 56909 1609 56967 1643
rect 57001 1609 57059 1643
rect 57093 1609 57122 1643
rect 55362 1546 55396 1562
rect 55362 1476 55396 1510
rect 55362 1424 55396 1440
rect 55458 1546 55492 1562
rect 55458 1476 55492 1510
rect 55458 1424 55492 1440
rect 55554 1546 55588 1562
rect 55554 1476 55588 1510
rect 55588 1440 55936 1464
rect 55554 1424 55936 1440
rect 55274 1356 55410 1390
rect 55444 1356 55460 1390
rect 55189 1286 55584 1306
rect 55189 1281 55451 1286
rect 55189 1272 55330 1281
rect 55314 1247 55330 1272
rect 55364 1252 55451 1281
rect 55485 1262 55584 1286
rect 55756 1264 55802 1266
rect 55756 1262 55760 1264
rect 55485 1252 55760 1262
rect 55364 1247 55760 1252
rect 55314 1230 55760 1247
rect 55794 1230 55802 1264
rect 55314 1228 55802 1230
rect 55756 1222 55802 1228
rect 54088 1107 54117 1141
rect 54151 1107 54209 1141
rect 54243 1107 54301 1141
rect 54335 1107 54364 1141
rect 53684 1055 53920 1066
rect 53326 1047 53920 1055
rect 53326 1022 53328 1047
rect 53240 979 53274 981
rect 53240 943 53274 945
rect 53240 858 53274 877
rect 53362 1022 53886 1047
rect 53972 1047 54048 1066
rect 53972 1026 53974 1047
rect 53328 979 53362 981
rect 53584 949 53600 983
rect 53634 949 53650 983
rect 53886 979 53920 981
rect 53328 943 53362 945
rect 53886 943 53920 945
rect 53328 858 53362 877
rect 53456 887 53490 906
rect 53456 819 53490 821
rect 53268 781 53284 815
rect 53318 781 53334 815
rect 53456 783 53490 785
rect 52956 703 52968 737
rect 52956 669 53002 703
rect 52956 635 52968 669
rect 52546 561 52575 595
rect 52609 561 52667 595
rect 52701 561 52759 595
rect 52793 561 52822 595
rect 52956 589 53002 635
rect 53036 737 53102 749
rect 53036 703 53052 737
rect 53086 703 53102 737
rect 53036 690 53102 703
rect 53456 698 53490 717
rect 53552 887 53586 906
rect 53552 819 53586 821
rect 53552 783 53586 785
rect 53552 698 53586 717
rect 53648 887 53682 906
rect 53886 858 53920 877
rect 54008 1026 54048 1047
rect 54156 1065 54198 1107
rect 54434 1105 54463 1139
rect 54497 1105 54555 1139
rect 54589 1105 54647 1139
rect 54681 1105 54710 1139
rect 54855 1133 54889 1140
rect 54156 1031 54164 1065
rect 53974 979 54008 981
rect 53974 943 54008 945
rect 54156 997 54198 1031
rect 54156 963 54164 997
rect 54156 929 54198 963
rect 54156 895 54164 929
rect 54156 879 54198 895
rect 54232 1065 54298 1073
rect 54232 1031 54248 1065
rect 54282 1031 54298 1065
rect 54232 997 54298 1031
rect 54232 963 54248 997
rect 54282 963 54298 997
rect 54232 929 54298 963
rect 54232 895 54248 929
rect 54282 895 54298 929
rect 54232 877 54298 895
rect 54467 1055 54503 1071
rect 54467 1021 54469 1055
rect 54467 987 54503 1021
rect 54467 953 54469 987
rect 54539 1055 54605 1105
rect 54780 1099 54809 1133
rect 54843 1099 54901 1133
rect 54935 1099 54993 1133
rect 55027 1099 55056 1133
rect 55156 1109 55172 1143
rect 55206 1109 55222 1143
rect 55380 1130 55494 1132
rect 54539 1021 54555 1055
rect 54589 1021 54605 1055
rect 54539 987 54605 1021
rect 54539 953 54555 987
rect 54589 953 54605 987
rect 54639 1055 54693 1071
rect 54639 1021 54641 1055
rect 54675 1021 54693 1055
rect 54639 974 54693 1021
rect 54467 919 54503 953
rect 54639 940 54641 974
rect 54675 940 54693 974
rect 54467 885 54602 919
rect 54639 890 54693 940
rect 53974 858 54008 877
rect 53648 819 53682 821
rect 54060 843 54204 844
rect 54060 829 54218 843
rect 53648 783 53682 785
rect 53914 816 53980 818
rect 54060 816 54168 829
rect 53914 815 54168 816
rect 53914 781 53930 815
rect 53964 802 54168 815
rect 53964 782 54100 802
rect 54152 795 54168 802
rect 54202 795 54218 829
rect 53964 781 53980 782
rect 54152 745 54198 761
rect 54252 757 54298 877
rect 54568 856 54602 885
rect 54455 827 54523 849
rect 54455 826 54471 827
rect 54455 792 54469 826
rect 54505 793 54523 827
rect 54503 792 54523 793
rect 54455 775 54523 792
rect 54568 840 54623 856
rect 54568 806 54589 840
rect 54568 790 54623 806
rect 54657 840 54693 890
rect 54848 1057 54890 1099
rect 55380 1091 55662 1130
rect 55802 1109 55818 1143
rect 55852 1109 55868 1143
rect 55380 1066 55419 1091
rect 54848 1023 54856 1057
rect 54848 989 54890 1023
rect 54848 955 54856 989
rect 54848 921 54890 955
rect 54848 887 54856 921
rect 54848 871 54890 887
rect 54924 1057 54990 1065
rect 54924 1023 54940 1057
rect 54974 1023 54990 1057
rect 54924 989 54990 1023
rect 54924 955 54940 989
rect 54974 955 54990 989
rect 54924 921 54990 955
rect 54924 887 54940 921
rect 54974 887 54990 921
rect 54924 869 54990 887
rect 54657 838 54698 840
rect 54657 804 54662 838
rect 54696 804 54698 838
rect 54657 802 54698 804
rect 54844 832 54910 835
rect 53682 717 53928 734
rect 53648 700 53928 717
rect 53648 698 53682 700
rect 53036 669 53378 690
rect 53036 635 53052 669
rect 53086 658 53378 669
rect 53086 655 53554 658
rect 53086 654 53504 655
rect 53086 635 53108 654
rect 53036 630 53108 635
rect 53036 623 53102 630
rect 53342 622 53504 654
rect 53488 621 53504 622
rect 53538 621 53554 655
rect 53880 612 53928 700
rect 52892 555 52921 589
rect 52955 555 53013 589
rect 53047 555 53105 589
rect 53139 555 53168 589
rect 53250 584 53296 594
rect 53250 550 53256 584
rect 53290 564 53296 584
rect 53880 578 53888 612
rect 53922 578 53928 612
rect 54152 711 54164 745
rect 54152 677 54198 711
rect 54152 643 54164 677
rect 54152 597 54198 643
rect 54232 745 54298 757
rect 54232 694 54248 745
rect 54282 694 54298 745
rect 54568 739 54602 790
rect 54232 677 54298 694
rect 54232 643 54248 677
rect 54282 643 54298 677
rect 54232 631 54298 643
rect 54469 705 54602 739
rect 54657 730 54693 802
rect 54844 798 54858 832
rect 54892 821 54910 832
rect 54844 787 54860 798
rect 54894 787 54910 821
rect 54469 684 54503 705
rect 54641 701 54693 730
rect 54469 629 54503 650
rect 54539 637 54555 671
rect 54589 637 54605 671
rect 53290 550 53300 564
rect 49888 420 49922 454
rect 49888 368 49922 384
rect 51280 444 51412 480
rect 51584 490 51618 506
rect 51680 490 51714 506
rect 51618 454 51619 455
rect 51280 396 51316 444
rect 51584 420 51619 454
rect 51618 418 51619 420
rect 51680 420 51714 454
rect 51464 396 51584 418
rect 51280 384 51584 396
rect 51618 384 51620 418
rect 51280 382 51620 384
rect 51280 360 51500 382
rect 51584 368 51618 382
rect 51680 368 51714 384
rect 51776 490 51810 506
rect 53250 480 53300 550
rect 53600 540 53616 574
rect 53650 540 53666 574
rect 53880 566 53928 578
rect 54088 563 54117 597
rect 54151 563 54209 597
rect 54243 563 54301 597
rect 54335 563 54364 597
rect 54539 595 54605 637
rect 54675 667 54693 701
rect 54641 629 54693 667
rect 54844 737 54890 753
rect 54944 749 54990 869
rect 55128 1047 55162 1066
rect 55214 1057 55419 1066
rect 55453 1089 55662 1091
rect 55453 1057 55538 1089
rect 55214 1055 55538 1057
rect 55572 1066 55662 1089
rect 55902 1066 55936 1424
rect 56846 1398 56880 1609
rect 57077 1306 57111 1609
rect 57162 1390 57196 2004
rect 57362 2002 57428 2004
rect 57679 2009 57695 2043
rect 57729 2009 57745 2043
rect 57679 1975 57745 2009
rect 57234 1943 57268 1962
rect 57234 1875 57268 1877
rect 57234 1839 57268 1841
rect 57234 1754 57268 1773
rect 57330 1943 57364 1962
rect 57330 1875 57364 1877
rect 57330 1839 57364 1841
rect 57330 1754 57364 1773
rect 57426 1943 57460 1962
rect 57679 1941 57695 1975
rect 57729 1959 57745 1975
rect 57851 2111 57917 2153
rect 57885 2077 57917 2111
rect 57851 2043 57917 2077
rect 57885 2009 57917 2043
rect 57851 1975 57917 2009
rect 57729 1941 57815 1959
rect 57679 1925 57815 1941
rect 57885 1941 57917 1975
rect 57851 1925 57917 1941
rect 58753 2111 58819 2116
rect 58753 2077 58769 2111
rect 58803 2077 58819 2111
rect 58753 2043 58819 2077
rect 58753 2009 58769 2043
rect 58803 2009 58819 2043
rect 58753 1975 58819 2009
rect 58753 1941 58769 1975
rect 58803 1959 58819 1975
rect 58925 2111 58991 2153
rect 58959 2077 58991 2111
rect 59158 2147 59440 2153
rect 59158 2113 59197 2147
rect 59231 2145 59440 2147
rect 59231 2113 59316 2145
rect 59158 2111 59316 2113
rect 59350 2111 59440 2145
rect 59158 2078 59440 2111
rect 59567 2111 59633 2116
rect 58925 2043 58991 2077
rect 58959 2009 58991 2043
rect 59567 2077 59583 2111
rect 59617 2077 59633 2111
rect 59567 2043 59633 2077
rect 58925 1975 58991 2009
rect 58803 1941 58889 1959
rect 58753 1925 58889 1941
rect 58959 1941 58991 1975
rect 58925 1925 58991 1941
rect 59050 2039 59316 2040
rect 59050 2005 59266 2039
rect 59300 2005 59316 2039
rect 59050 2004 59316 2005
rect 57426 1875 57460 1877
rect 57677 1882 57747 1891
rect 57677 1848 57693 1882
rect 57727 1875 57747 1882
rect 57677 1841 57697 1848
rect 57731 1841 57747 1875
rect 57426 1839 57460 1841
rect 57781 1805 57815 1925
rect 57849 1882 57919 1891
rect 57849 1875 57867 1882
rect 57849 1841 57865 1875
rect 57901 1848 57919 1882
rect 57899 1841 57919 1848
rect 58751 1884 58821 1891
rect 58751 1850 58769 1884
rect 58803 1875 58821 1884
rect 58751 1841 58771 1850
rect 58805 1841 58821 1875
rect 58855 1805 58889 1925
rect 58923 1880 58993 1891
rect 58923 1875 58942 1880
rect 58923 1841 58939 1875
rect 58976 1846 58993 1880
rect 58973 1841 58993 1846
rect 57426 1754 57460 1773
rect 57681 1789 57729 1805
rect 57681 1755 57695 1789
rect 57681 1721 57729 1755
rect 57266 1677 57282 1711
rect 57316 1677 57332 1711
rect 57681 1687 57695 1721
rect 57681 1643 57729 1687
rect 57763 1789 57829 1805
rect 57763 1755 57779 1789
rect 57813 1759 57829 1789
rect 57763 1725 57781 1755
rect 57815 1725 57829 1759
rect 57763 1721 57829 1725
rect 57763 1687 57779 1721
rect 57813 1687 57829 1721
rect 57763 1677 57829 1687
rect 57863 1789 57917 1805
rect 57897 1755 57917 1789
rect 57863 1721 57917 1755
rect 57897 1687 57917 1721
rect 57863 1643 57917 1687
rect 58755 1789 58803 1805
rect 58755 1755 58769 1789
rect 58755 1721 58803 1755
rect 58755 1687 58769 1721
rect 58755 1643 58803 1687
rect 58837 1789 58903 1805
rect 58837 1764 58853 1789
rect 58837 1730 58851 1764
rect 58887 1755 58903 1789
rect 58885 1730 58903 1755
rect 58837 1721 58903 1730
rect 58837 1687 58853 1721
rect 58887 1687 58903 1721
rect 58837 1677 58903 1687
rect 58937 1789 58991 1805
rect 58971 1755 58991 1789
rect 58937 1721 58991 1755
rect 58971 1687 58991 1721
rect 58937 1643 58991 1687
rect 57378 1596 57394 1630
rect 57428 1596 57444 1630
rect 57660 1609 57689 1643
rect 57723 1609 57781 1643
rect 57815 1609 57873 1643
rect 57907 1609 57936 1643
rect 58734 1609 58763 1643
rect 58797 1609 58855 1643
rect 58889 1609 58947 1643
rect 58981 1609 59010 1643
rect 57250 1546 57284 1562
rect 57250 1476 57284 1510
rect 57250 1424 57284 1440
rect 57346 1546 57380 1562
rect 57346 1476 57380 1510
rect 57346 1424 57380 1440
rect 57442 1546 57476 1562
rect 57442 1476 57476 1510
rect 57476 1440 57824 1464
rect 57442 1424 57824 1440
rect 57162 1356 57298 1390
rect 57332 1356 57348 1390
rect 57077 1286 57472 1306
rect 57077 1281 57339 1286
rect 57077 1272 57218 1281
rect 57202 1247 57218 1272
rect 57252 1252 57339 1281
rect 57373 1262 57472 1286
rect 57644 1264 57690 1266
rect 57644 1262 57648 1264
rect 57373 1252 57648 1262
rect 57252 1247 57648 1252
rect 57202 1230 57648 1247
rect 57682 1230 57690 1264
rect 57202 1228 57690 1230
rect 57644 1222 57690 1228
rect 55976 1107 56005 1141
rect 56039 1107 56097 1141
rect 56131 1107 56189 1141
rect 56223 1107 56252 1141
rect 55572 1055 55808 1066
rect 55214 1047 55808 1055
rect 55214 1022 55216 1047
rect 55128 979 55162 981
rect 55128 943 55162 945
rect 55128 858 55162 877
rect 55250 1022 55774 1047
rect 55860 1047 55936 1066
rect 55860 1026 55862 1047
rect 55216 979 55250 981
rect 55472 949 55488 983
rect 55522 949 55538 983
rect 55774 979 55808 981
rect 55216 943 55250 945
rect 55774 943 55808 945
rect 55216 858 55250 877
rect 55344 887 55378 906
rect 55344 819 55378 821
rect 55156 781 55172 815
rect 55206 781 55222 815
rect 55344 783 55378 785
rect 54844 703 54856 737
rect 54844 669 54890 703
rect 54844 635 54856 669
rect 54434 561 54463 595
rect 54497 561 54555 595
rect 54589 561 54647 595
rect 54681 561 54710 595
rect 54844 589 54890 635
rect 54924 737 54990 749
rect 54924 703 54940 737
rect 54974 703 54990 737
rect 54924 690 54990 703
rect 55344 698 55378 717
rect 55440 887 55474 906
rect 55440 819 55474 821
rect 55440 783 55474 785
rect 55440 698 55474 717
rect 55536 887 55570 906
rect 55774 858 55808 877
rect 55896 1026 55936 1047
rect 56044 1065 56086 1107
rect 56322 1105 56351 1139
rect 56385 1105 56443 1139
rect 56477 1105 56535 1139
rect 56569 1105 56598 1139
rect 56743 1133 56777 1140
rect 56044 1031 56052 1065
rect 55862 979 55896 981
rect 55862 943 55896 945
rect 56044 997 56086 1031
rect 56044 963 56052 997
rect 56044 929 56086 963
rect 56044 895 56052 929
rect 56044 879 56086 895
rect 56120 1065 56186 1073
rect 56120 1031 56136 1065
rect 56170 1031 56186 1065
rect 56120 997 56186 1031
rect 56120 963 56136 997
rect 56170 963 56186 997
rect 56120 929 56186 963
rect 56120 895 56136 929
rect 56170 895 56186 929
rect 56120 877 56186 895
rect 56355 1055 56391 1071
rect 56355 1021 56357 1055
rect 56355 987 56391 1021
rect 56355 953 56357 987
rect 56427 1055 56493 1105
rect 56668 1099 56697 1133
rect 56731 1099 56789 1133
rect 56823 1099 56881 1133
rect 56915 1099 56944 1133
rect 57044 1109 57060 1143
rect 57094 1109 57110 1143
rect 57268 1130 57382 1132
rect 56427 1021 56443 1055
rect 56477 1021 56493 1055
rect 56427 987 56493 1021
rect 56427 953 56443 987
rect 56477 953 56493 987
rect 56527 1055 56581 1071
rect 56527 1021 56529 1055
rect 56563 1021 56581 1055
rect 56527 974 56581 1021
rect 56355 919 56391 953
rect 56527 940 56529 974
rect 56563 940 56581 974
rect 56355 885 56490 919
rect 56527 890 56581 940
rect 55862 858 55896 877
rect 55536 819 55570 821
rect 55948 843 56092 844
rect 55948 829 56106 843
rect 55536 783 55570 785
rect 55802 816 55868 818
rect 55948 816 56056 829
rect 55802 815 56056 816
rect 55802 781 55818 815
rect 55852 802 56056 815
rect 55852 782 55988 802
rect 56040 795 56056 802
rect 56090 795 56106 829
rect 55852 781 55868 782
rect 56040 745 56086 761
rect 56140 757 56186 877
rect 56456 856 56490 885
rect 56343 827 56411 849
rect 56343 826 56359 827
rect 56343 792 56357 826
rect 56393 793 56411 827
rect 56391 792 56411 793
rect 56343 775 56411 792
rect 56456 840 56511 856
rect 56456 806 56477 840
rect 56456 790 56511 806
rect 56545 840 56581 890
rect 56736 1057 56778 1099
rect 57268 1091 57550 1130
rect 57690 1109 57706 1143
rect 57740 1109 57756 1143
rect 57268 1066 57307 1091
rect 56736 1023 56744 1057
rect 56736 989 56778 1023
rect 56736 955 56744 989
rect 56736 921 56778 955
rect 56736 887 56744 921
rect 56736 871 56778 887
rect 56812 1057 56878 1065
rect 56812 1023 56828 1057
rect 56862 1023 56878 1057
rect 56812 989 56878 1023
rect 56812 955 56828 989
rect 56862 955 56878 989
rect 56812 921 56878 955
rect 56812 887 56828 921
rect 56862 887 56878 921
rect 56812 869 56878 887
rect 56545 838 56586 840
rect 56545 804 56550 838
rect 56584 804 56586 838
rect 56545 802 56586 804
rect 56732 832 56798 835
rect 55570 717 55816 734
rect 55536 700 55816 717
rect 55536 698 55570 700
rect 54924 669 55266 690
rect 54924 635 54940 669
rect 54974 658 55266 669
rect 54974 655 55442 658
rect 54974 654 55392 655
rect 54974 635 54996 654
rect 54924 630 54996 635
rect 54924 623 54990 630
rect 55230 622 55392 654
rect 55376 621 55392 622
rect 55426 621 55442 655
rect 55768 612 55816 700
rect 54780 555 54809 589
rect 54843 555 54901 589
rect 54935 555 54993 589
rect 55027 555 55056 589
rect 55138 584 55184 594
rect 55138 550 55144 584
rect 55178 564 55184 584
rect 55768 578 55776 612
rect 55810 578 55816 612
rect 56040 711 56052 745
rect 56040 677 56086 711
rect 56040 643 56052 677
rect 56040 597 56086 643
rect 56120 745 56186 757
rect 56120 694 56136 745
rect 56170 694 56186 745
rect 56456 739 56490 790
rect 56120 677 56186 694
rect 56120 643 56136 677
rect 56170 643 56186 677
rect 56120 631 56186 643
rect 56357 705 56490 739
rect 56545 730 56581 802
rect 56732 798 56746 832
rect 56780 821 56798 832
rect 56732 787 56748 798
rect 56782 787 56798 821
rect 56357 684 56391 705
rect 56529 701 56581 730
rect 56357 629 56391 650
rect 56427 637 56443 671
rect 56477 637 56493 671
rect 55178 550 55188 564
rect 51776 420 51810 454
rect 51776 368 51810 384
rect 53168 444 53300 480
rect 53472 490 53506 506
rect 53568 490 53602 506
rect 53506 454 53507 455
rect 53168 396 53204 444
rect 53472 420 53507 454
rect 53506 418 53507 420
rect 53568 420 53602 454
rect 53352 396 53472 418
rect 53168 384 53472 396
rect 53506 384 53508 418
rect 53168 382 53508 384
rect 53168 360 53388 382
rect 53472 368 53506 382
rect 53568 368 53602 384
rect 53664 490 53698 506
rect 55138 480 55188 550
rect 55488 540 55504 574
rect 55538 540 55554 574
rect 55768 566 55816 578
rect 55976 563 56005 597
rect 56039 563 56097 597
rect 56131 563 56189 597
rect 56223 563 56252 597
rect 56427 595 56493 637
rect 56563 667 56581 701
rect 56529 629 56581 667
rect 56732 737 56778 753
rect 56832 749 56878 869
rect 57016 1047 57050 1066
rect 57102 1057 57307 1066
rect 57341 1089 57550 1091
rect 57341 1057 57426 1089
rect 57102 1055 57426 1057
rect 57460 1066 57550 1089
rect 57790 1066 57824 1424
rect 58734 1398 58768 1609
rect 58965 1306 58999 1609
rect 59050 1390 59084 2004
rect 59250 2002 59316 2004
rect 59567 2009 59583 2043
rect 59617 2009 59633 2043
rect 59567 1975 59633 2009
rect 59122 1943 59156 1962
rect 59122 1875 59156 1877
rect 59122 1839 59156 1841
rect 59122 1754 59156 1773
rect 59218 1943 59252 1962
rect 59218 1875 59252 1877
rect 59218 1839 59252 1841
rect 59218 1754 59252 1773
rect 59314 1943 59348 1962
rect 59567 1941 59583 1975
rect 59617 1959 59633 1975
rect 59739 2111 59805 2153
rect 59773 2077 59805 2111
rect 59739 2043 59805 2077
rect 59773 2009 59805 2043
rect 59739 1975 59805 2009
rect 59617 1941 59703 1959
rect 59567 1925 59703 1941
rect 59773 1941 59805 1975
rect 59739 1925 59805 1941
rect 59314 1875 59348 1877
rect 59565 1882 59635 1891
rect 59565 1848 59581 1882
rect 59615 1875 59635 1882
rect 59565 1841 59585 1848
rect 59619 1841 59635 1875
rect 59314 1839 59348 1841
rect 59669 1805 59703 1925
rect 59737 1882 59807 1891
rect 59737 1875 59755 1882
rect 59737 1841 59753 1875
rect 59789 1848 59807 1882
rect 59787 1841 59807 1848
rect 59314 1754 59348 1773
rect 59569 1789 59617 1805
rect 59569 1755 59583 1789
rect 59569 1721 59617 1755
rect 59154 1677 59170 1711
rect 59204 1677 59220 1711
rect 59569 1687 59583 1721
rect 59569 1643 59617 1687
rect 59651 1789 59717 1805
rect 59651 1755 59667 1789
rect 59701 1759 59717 1789
rect 59651 1725 59669 1755
rect 59703 1725 59717 1759
rect 59651 1721 59717 1725
rect 59651 1687 59667 1721
rect 59701 1687 59717 1721
rect 59651 1677 59717 1687
rect 59751 1789 59805 1805
rect 59785 1755 59805 1789
rect 59751 1721 59805 1755
rect 59785 1687 59805 1721
rect 59751 1643 59805 1687
rect 59266 1596 59282 1630
rect 59316 1596 59332 1630
rect 59548 1609 59577 1643
rect 59611 1609 59669 1643
rect 59703 1609 59761 1643
rect 59795 1609 59824 1643
rect 59138 1546 59172 1562
rect 59138 1476 59172 1510
rect 59138 1424 59172 1440
rect 59234 1546 59268 1562
rect 59234 1476 59268 1510
rect 59234 1424 59268 1440
rect 59330 1546 59364 1562
rect 59330 1476 59364 1510
rect 59364 1440 59712 1464
rect 59330 1424 59712 1440
rect 59050 1356 59186 1390
rect 59220 1356 59236 1390
rect 58965 1286 59360 1306
rect 58965 1281 59227 1286
rect 58965 1272 59106 1281
rect 59090 1247 59106 1272
rect 59140 1252 59227 1281
rect 59261 1262 59360 1286
rect 59532 1264 59578 1266
rect 59532 1262 59536 1264
rect 59261 1252 59536 1262
rect 59140 1247 59536 1252
rect 59090 1230 59536 1247
rect 59570 1230 59578 1264
rect 59090 1228 59578 1230
rect 59532 1222 59578 1228
rect 57864 1107 57893 1141
rect 57927 1107 57985 1141
rect 58019 1107 58077 1141
rect 58111 1107 58140 1141
rect 57460 1055 57696 1066
rect 57102 1047 57696 1055
rect 57102 1022 57104 1047
rect 57016 979 57050 981
rect 57016 943 57050 945
rect 57016 858 57050 877
rect 57138 1022 57662 1047
rect 57748 1047 57824 1066
rect 57748 1026 57750 1047
rect 57104 979 57138 981
rect 57360 949 57376 983
rect 57410 949 57426 983
rect 57662 979 57696 981
rect 57104 943 57138 945
rect 57662 943 57696 945
rect 57104 858 57138 877
rect 57232 887 57266 906
rect 57232 819 57266 821
rect 57044 781 57060 815
rect 57094 781 57110 815
rect 57232 783 57266 785
rect 56732 703 56744 737
rect 56732 669 56778 703
rect 56732 635 56744 669
rect 56322 561 56351 595
rect 56385 561 56443 595
rect 56477 561 56535 595
rect 56569 561 56598 595
rect 56732 589 56778 635
rect 56812 737 56878 749
rect 56812 703 56828 737
rect 56862 703 56878 737
rect 56812 690 56878 703
rect 57232 698 57266 717
rect 57328 887 57362 906
rect 57328 819 57362 821
rect 57328 783 57362 785
rect 57328 698 57362 717
rect 57424 887 57458 906
rect 57662 858 57696 877
rect 57784 1026 57824 1047
rect 57932 1065 57974 1107
rect 58210 1105 58239 1139
rect 58273 1105 58331 1139
rect 58365 1105 58423 1139
rect 58457 1105 58486 1139
rect 58631 1133 58665 1140
rect 57932 1031 57940 1065
rect 57750 979 57784 981
rect 57750 943 57784 945
rect 57932 997 57974 1031
rect 57932 963 57940 997
rect 57932 929 57974 963
rect 57932 895 57940 929
rect 57932 879 57974 895
rect 58008 1065 58074 1073
rect 58008 1031 58024 1065
rect 58058 1031 58074 1065
rect 58008 997 58074 1031
rect 58008 963 58024 997
rect 58058 963 58074 997
rect 58008 929 58074 963
rect 58008 895 58024 929
rect 58058 895 58074 929
rect 58008 877 58074 895
rect 58243 1055 58279 1071
rect 58243 1021 58245 1055
rect 58243 987 58279 1021
rect 58243 953 58245 987
rect 58315 1055 58381 1105
rect 58556 1099 58585 1133
rect 58619 1099 58677 1133
rect 58711 1099 58769 1133
rect 58803 1099 58832 1133
rect 58932 1109 58948 1143
rect 58982 1109 58998 1143
rect 59156 1130 59270 1132
rect 58315 1021 58331 1055
rect 58365 1021 58381 1055
rect 58315 987 58381 1021
rect 58315 953 58331 987
rect 58365 953 58381 987
rect 58415 1055 58469 1071
rect 58415 1021 58417 1055
rect 58451 1021 58469 1055
rect 58415 974 58469 1021
rect 58243 919 58279 953
rect 58415 940 58417 974
rect 58451 940 58469 974
rect 58243 885 58378 919
rect 58415 890 58469 940
rect 57750 858 57784 877
rect 57424 819 57458 821
rect 57836 843 57980 844
rect 57836 829 57994 843
rect 57424 783 57458 785
rect 57690 816 57756 818
rect 57836 816 57944 829
rect 57690 815 57944 816
rect 57690 781 57706 815
rect 57740 802 57944 815
rect 57740 782 57876 802
rect 57928 795 57944 802
rect 57978 795 57994 829
rect 57740 781 57756 782
rect 57928 745 57974 761
rect 58028 757 58074 877
rect 58344 856 58378 885
rect 58231 827 58299 849
rect 58231 826 58247 827
rect 58231 792 58245 826
rect 58281 793 58299 827
rect 58279 792 58299 793
rect 58231 775 58299 792
rect 58344 840 58399 856
rect 58344 806 58365 840
rect 58344 790 58399 806
rect 58433 840 58469 890
rect 58624 1057 58666 1099
rect 59156 1091 59438 1130
rect 59578 1109 59594 1143
rect 59628 1109 59644 1143
rect 59156 1066 59195 1091
rect 58624 1023 58632 1057
rect 58624 989 58666 1023
rect 58624 955 58632 989
rect 58624 921 58666 955
rect 58624 887 58632 921
rect 58624 871 58666 887
rect 58700 1057 58766 1065
rect 58700 1023 58716 1057
rect 58750 1023 58766 1057
rect 58700 989 58766 1023
rect 58700 955 58716 989
rect 58750 955 58766 989
rect 58700 921 58766 955
rect 58700 887 58716 921
rect 58750 887 58766 921
rect 58700 869 58766 887
rect 58433 838 58474 840
rect 58433 804 58438 838
rect 58472 804 58474 838
rect 58433 802 58474 804
rect 58620 832 58686 835
rect 57458 717 57704 734
rect 57424 700 57704 717
rect 57424 698 57458 700
rect 56812 669 57154 690
rect 56812 635 56828 669
rect 56862 658 57154 669
rect 56862 655 57330 658
rect 56862 654 57280 655
rect 56862 635 56884 654
rect 56812 630 56884 635
rect 56812 623 56878 630
rect 57118 622 57280 654
rect 57264 621 57280 622
rect 57314 621 57330 655
rect 57656 612 57704 700
rect 56668 555 56697 589
rect 56731 555 56789 589
rect 56823 555 56881 589
rect 56915 555 56944 589
rect 57026 584 57072 594
rect 57026 550 57032 584
rect 57066 564 57072 584
rect 57656 578 57664 612
rect 57698 578 57704 612
rect 57928 711 57940 745
rect 57928 677 57974 711
rect 57928 643 57940 677
rect 57928 597 57974 643
rect 58008 745 58074 757
rect 58008 694 58024 745
rect 58058 694 58074 745
rect 58344 739 58378 790
rect 58008 677 58074 694
rect 58008 643 58024 677
rect 58058 643 58074 677
rect 58008 631 58074 643
rect 58245 705 58378 739
rect 58433 730 58469 802
rect 58620 798 58634 832
rect 58668 821 58686 832
rect 58620 787 58636 798
rect 58670 787 58686 821
rect 58245 684 58279 705
rect 58417 701 58469 730
rect 58245 629 58279 650
rect 58315 637 58331 671
rect 58365 637 58381 671
rect 57066 550 57076 564
rect 53664 420 53698 454
rect 53664 368 53698 384
rect 55056 444 55188 480
rect 55360 490 55394 506
rect 55456 490 55490 506
rect 55394 454 55395 455
rect 55056 396 55092 444
rect 55360 420 55395 454
rect 55394 418 55395 420
rect 55456 420 55490 454
rect 55240 396 55360 418
rect 55056 384 55360 396
rect 55394 384 55396 418
rect 55056 382 55396 384
rect 55056 360 55276 382
rect 55360 368 55394 382
rect 55456 368 55490 384
rect 55552 490 55586 506
rect 57026 480 57076 550
rect 57376 540 57392 574
rect 57426 540 57442 574
rect 57656 566 57704 578
rect 57864 563 57893 597
rect 57927 563 57985 597
rect 58019 563 58077 597
rect 58111 563 58140 597
rect 58315 595 58381 637
rect 58451 667 58469 701
rect 58417 629 58469 667
rect 58620 737 58666 753
rect 58720 749 58766 869
rect 58904 1047 58938 1066
rect 58990 1057 59195 1066
rect 59229 1089 59438 1091
rect 59229 1057 59314 1089
rect 58990 1055 59314 1057
rect 59348 1066 59438 1089
rect 59678 1066 59712 1424
rect 59752 1107 59781 1141
rect 59815 1107 59873 1141
rect 59907 1107 59965 1141
rect 59999 1107 60028 1141
rect 59348 1055 59584 1066
rect 58990 1047 59584 1055
rect 58990 1022 58992 1047
rect 58904 979 58938 981
rect 58904 943 58938 945
rect 58904 858 58938 877
rect 59026 1022 59550 1047
rect 59636 1047 59712 1066
rect 59636 1026 59638 1047
rect 58992 979 59026 981
rect 59248 949 59264 983
rect 59298 949 59314 983
rect 59550 979 59584 981
rect 58992 943 59026 945
rect 59550 943 59584 945
rect 58992 858 59026 877
rect 59120 887 59154 906
rect 59120 819 59154 821
rect 58932 781 58948 815
rect 58982 781 58998 815
rect 59120 783 59154 785
rect 58620 703 58632 737
rect 58620 669 58666 703
rect 58620 635 58632 669
rect 58210 561 58239 595
rect 58273 561 58331 595
rect 58365 561 58423 595
rect 58457 561 58486 595
rect 58620 589 58666 635
rect 58700 737 58766 749
rect 58700 703 58716 737
rect 58750 703 58766 737
rect 58700 690 58766 703
rect 59120 698 59154 717
rect 59216 887 59250 906
rect 59216 819 59250 821
rect 59216 783 59250 785
rect 59216 698 59250 717
rect 59312 887 59346 906
rect 59550 858 59584 877
rect 59672 1026 59712 1047
rect 59820 1065 59862 1107
rect 60098 1105 60127 1139
rect 60161 1105 60219 1139
rect 60253 1105 60311 1139
rect 60345 1105 60374 1139
rect 59820 1031 59828 1065
rect 59638 979 59672 981
rect 59638 943 59672 945
rect 59820 997 59862 1031
rect 59820 963 59828 997
rect 59820 929 59862 963
rect 59820 895 59828 929
rect 59820 879 59862 895
rect 59896 1065 59962 1073
rect 59896 1031 59912 1065
rect 59946 1031 59962 1065
rect 59896 997 59962 1031
rect 59896 963 59912 997
rect 59946 963 59962 997
rect 59896 929 59962 963
rect 59896 895 59912 929
rect 59946 895 59962 929
rect 59896 877 59962 895
rect 60131 1055 60167 1071
rect 60131 1021 60133 1055
rect 60131 987 60167 1021
rect 60131 953 60133 987
rect 60203 1055 60269 1105
rect 60203 1021 60219 1055
rect 60253 1021 60269 1055
rect 60203 987 60269 1021
rect 60203 953 60219 987
rect 60253 953 60269 987
rect 60303 1055 60357 1071
rect 60303 1021 60305 1055
rect 60339 1021 60357 1055
rect 60303 974 60357 1021
rect 60131 919 60167 953
rect 60303 940 60305 974
rect 60339 940 60357 974
rect 60131 885 60266 919
rect 60303 890 60357 940
rect 59638 858 59672 877
rect 59312 819 59346 821
rect 59724 843 59868 844
rect 59724 829 59882 843
rect 59312 783 59346 785
rect 59578 816 59644 818
rect 59724 816 59832 829
rect 59578 815 59832 816
rect 59578 781 59594 815
rect 59628 802 59832 815
rect 59628 782 59764 802
rect 59816 795 59832 802
rect 59866 795 59882 829
rect 59628 781 59644 782
rect 59816 745 59862 761
rect 59916 757 59962 877
rect 60232 856 60266 885
rect 60119 827 60187 849
rect 60119 826 60135 827
rect 60119 792 60133 826
rect 60169 793 60187 827
rect 60167 792 60187 793
rect 60119 775 60187 792
rect 60232 840 60287 856
rect 60232 806 60253 840
rect 60232 790 60287 806
rect 60321 840 60357 890
rect 60321 838 60362 840
rect 60321 804 60326 838
rect 60360 804 60362 838
rect 60321 802 60362 804
rect 59346 717 59592 734
rect 59312 700 59592 717
rect 59312 698 59346 700
rect 58700 669 59042 690
rect 58700 635 58716 669
rect 58750 658 59042 669
rect 58750 655 59218 658
rect 58750 654 59168 655
rect 58750 635 58772 654
rect 58700 630 58772 635
rect 58700 623 58766 630
rect 59006 622 59168 654
rect 59152 621 59168 622
rect 59202 621 59218 655
rect 59544 612 59592 700
rect 58556 555 58585 589
rect 58619 555 58677 589
rect 58711 555 58769 589
rect 58803 555 58832 589
rect 58914 584 58960 594
rect 58914 550 58920 584
rect 58954 564 58960 584
rect 59544 578 59552 612
rect 59586 578 59592 612
rect 59816 711 59828 745
rect 59816 677 59862 711
rect 59816 643 59828 677
rect 59816 597 59862 643
rect 59896 745 59962 757
rect 59896 694 59912 745
rect 59946 694 59962 745
rect 60232 739 60266 790
rect 59896 677 59962 694
rect 59896 643 59912 677
rect 59946 643 59962 677
rect 59896 631 59962 643
rect 60133 705 60266 739
rect 60321 730 60357 802
rect 60133 684 60167 705
rect 60305 701 60357 730
rect 60133 629 60167 650
rect 60203 637 60219 671
rect 60253 637 60269 671
rect 58954 550 58964 564
rect 55552 420 55586 454
rect 55552 368 55586 384
rect 56944 444 57076 480
rect 57248 490 57282 506
rect 57344 490 57378 506
rect 57282 454 57283 455
rect 56944 396 56980 444
rect 57248 420 57283 454
rect 57282 418 57283 420
rect 57344 420 57378 454
rect 57128 396 57248 418
rect 56944 384 57248 396
rect 57282 384 57284 418
rect 56944 382 57284 384
rect 56944 360 57164 382
rect 57248 368 57282 382
rect 57344 368 57378 384
rect 57440 490 57474 506
rect 58914 480 58964 550
rect 59264 540 59280 574
rect 59314 540 59330 574
rect 59544 566 59592 578
rect 59752 563 59781 597
rect 59815 563 59873 597
rect 59907 563 59965 597
rect 59999 563 60028 597
rect 60203 595 60269 637
rect 60339 667 60357 701
rect 60305 629 60357 667
rect 60098 561 60127 595
rect 60161 561 60219 595
rect 60253 561 60311 595
rect 60345 561 60374 595
rect 57440 420 57474 454
rect 57440 368 57474 384
rect 58832 444 58964 480
rect 59136 490 59170 506
rect 59232 490 59266 506
rect 59170 454 59171 455
rect 58832 396 58868 444
rect 59136 420 59171 454
rect 59170 418 59171 420
rect 59232 420 59266 454
rect 59016 396 59136 418
rect 58832 384 59136 396
rect 59170 384 59172 418
rect 58832 382 59172 384
rect 58832 360 59052 382
rect 59136 368 59170 382
rect 59232 368 59266 384
rect 59328 490 59362 506
rect 59328 420 59362 454
rect 59328 368 59362 384
rect 652 300 668 334
rect 702 300 718 334
rect 2540 300 2556 334
rect 2590 300 2606 334
rect 4428 300 4444 334
rect 4478 300 4494 334
rect 6316 300 6332 334
rect 6366 300 6382 334
rect 8204 300 8220 334
rect 8254 300 8270 334
rect 10092 300 10108 334
rect 10142 300 10158 334
rect 11980 300 11996 334
rect 12030 300 12046 334
rect 13868 300 13884 334
rect 13918 300 13934 334
rect 15750 300 15766 334
rect 15800 300 15816 334
rect 17638 300 17654 334
rect 17688 300 17704 334
rect 19526 300 19542 334
rect 19576 300 19592 334
rect 21414 300 21430 334
rect 21464 300 21480 334
rect 23302 300 23318 334
rect 23352 300 23368 334
rect 25190 300 25206 334
rect 25240 300 25256 334
rect 27078 300 27094 334
rect 27128 300 27144 334
rect 28966 300 28982 334
rect 29016 300 29032 334
rect 30854 300 30870 334
rect 30904 300 30920 334
rect 32742 300 32758 334
rect 32792 300 32808 334
rect 34630 300 34646 334
rect 34680 300 34696 334
rect 36518 300 36534 334
rect 36568 300 36584 334
rect 38406 300 38422 334
rect 38456 300 38472 334
rect 40294 300 40310 334
rect 40344 300 40360 334
rect 42182 300 42198 334
rect 42232 300 42248 334
rect 44070 300 44086 334
rect 44120 300 44136 334
rect 45952 300 45968 334
rect 46002 300 46018 334
rect 47840 300 47856 334
rect 47890 300 47906 334
rect 49728 300 49744 334
rect 49778 300 49794 334
rect 51616 300 51632 334
rect 51666 300 51682 334
rect 53504 300 53520 334
rect 53554 300 53570 334
rect 55392 300 55408 334
rect 55442 300 55458 334
rect 57280 300 57296 334
rect 57330 300 57346 334
rect 59168 300 59184 334
rect 59218 300 59234 334
rect 572 230 842 250
rect 572 225 709 230
rect 572 191 588 225
rect 622 196 709 225
rect 743 196 842 230
rect 622 191 842 196
rect 572 172 842 191
rect 2460 230 2730 250
rect 2460 225 2597 230
rect 2460 191 2476 225
rect 2510 196 2597 225
rect 2631 196 2730 230
rect 2510 191 2730 196
rect 2460 172 2730 191
rect 4348 230 4618 250
rect 4348 225 4485 230
rect 4348 191 4364 225
rect 4398 196 4485 225
rect 4519 196 4618 230
rect 4398 191 4618 196
rect 4348 172 4618 191
rect 6236 230 6506 250
rect 6236 225 6373 230
rect 6236 191 6252 225
rect 6286 196 6373 225
rect 6407 196 6506 230
rect 6286 191 6506 196
rect 6236 172 6506 191
rect 8124 230 8394 250
rect 8124 225 8261 230
rect 8124 191 8140 225
rect 8174 196 8261 225
rect 8295 196 8394 230
rect 8174 191 8394 196
rect 8124 172 8394 191
rect 10012 230 10282 250
rect 10012 225 10149 230
rect 10012 191 10028 225
rect 10062 196 10149 225
rect 10183 196 10282 230
rect 10062 191 10282 196
rect 10012 172 10282 191
rect 11900 230 12170 250
rect 11900 225 12037 230
rect 11900 191 11916 225
rect 11950 196 12037 225
rect 12071 196 12170 230
rect 11950 191 12170 196
rect 11900 172 12170 191
rect 13788 230 14058 250
rect 13788 225 13925 230
rect 13788 191 13804 225
rect 13838 196 13925 225
rect 13959 196 14058 230
rect 13838 191 14058 196
rect 13788 172 14058 191
rect 15670 230 15940 250
rect 15670 225 15807 230
rect 15670 191 15686 225
rect 15720 196 15807 225
rect 15841 196 15940 230
rect 15720 191 15940 196
rect 15670 172 15940 191
rect 17558 230 17828 250
rect 17558 225 17695 230
rect 17558 191 17574 225
rect 17608 196 17695 225
rect 17729 196 17828 230
rect 17608 191 17828 196
rect 17558 172 17828 191
rect 19446 230 19716 250
rect 19446 225 19583 230
rect 19446 191 19462 225
rect 19496 196 19583 225
rect 19617 196 19716 230
rect 19496 191 19716 196
rect 19446 172 19716 191
rect 21334 230 21604 250
rect 21334 225 21471 230
rect 21334 191 21350 225
rect 21384 196 21471 225
rect 21505 196 21604 230
rect 21384 191 21604 196
rect 21334 172 21604 191
rect 23222 230 23492 250
rect 23222 225 23359 230
rect 23222 191 23238 225
rect 23272 196 23359 225
rect 23393 196 23492 230
rect 23272 191 23492 196
rect 23222 172 23492 191
rect 25110 230 25380 250
rect 25110 225 25247 230
rect 25110 191 25126 225
rect 25160 196 25247 225
rect 25281 196 25380 230
rect 25160 191 25380 196
rect 25110 172 25380 191
rect 26998 230 27268 250
rect 26998 225 27135 230
rect 26998 191 27014 225
rect 27048 196 27135 225
rect 27169 196 27268 230
rect 27048 191 27268 196
rect 26998 172 27268 191
rect 28886 230 29156 250
rect 28886 225 29023 230
rect 28886 191 28902 225
rect 28936 196 29023 225
rect 29057 196 29156 230
rect 28936 191 29156 196
rect 28886 172 29156 191
rect 30774 230 31044 250
rect 30774 225 30911 230
rect 30774 191 30790 225
rect 30824 196 30911 225
rect 30945 196 31044 230
rect 30824 191 31044 196
rect 30774 172 31044 191
rect 32662 230 32932 250
rect 32662 225 32799 230
rect 32662 191 32678 225
rect 32712 196 32799 225
rect 32833 196 32932 230
rect 32712 191 32932 196
rect 32662 172 32932 191
rect 34550 230 34820 250
rect 34550 225 34687 230
rect 34550 191 34566 225
rect 34600 196 34687 225
rect 34721 196 34820 230
rect 34600 191 34820 196
rect 34550 172 34820 191
rect 36438 230 36708 250
rect 36438 225 36575 230
rect 36438 191 36454 225
rect 36488 196 36575 225
rect 36609 196 36708 230
rect 36488 191 36708 196
rect 36438 172 36708 191
rect 38326 230 38596 250
rect 38326 225 38463 230
rect 38326 191 38342 225
rect 38376 196 38463 225
rect 38497 196 38596 230
rect 38376 191 38596 196
rect 38326 172 38596 191
rect 40214 230 40484 250
rect 40214 225 40351 230
rect 40214 191 40230 225
rect 40264 196 40351 225
rect 40385 196 40484 230
rect 40264 191 40484 196
rect 40214 172 40484 191
rect 42102 230 42372 250
rect 42102 225 42239 230
rect 42102 191 42118 225
rect 42152 196 42239 225
rect 42273 196 42372 230
rect 42152 191 42372 196
rect 42102 172 42372 191
rect 43990 230 44260 250
rect 43990 225 44127 230
rect 43990 191 44006 225
rect 44040 196 44127 225
rect 44161 196 44260 230
rect 44040 191 44260 196
rect 43990 172 44260 191
rect 45872 230 46142 250
rect 45872 225 46009 230
rect 45872 191 45888 225
rect 45922 196 46009 225
rect 46043 196 46142 230
rect 45922 191 46142 196
rect 45872 172 46142 191
rect 47760 230 48030 250
rect 47760 225 47897 230
rect 47760 191 47776 225
rect 47810 196 47897 225
rect 47931 196 48030 230
rect 47810 191 48030 196
rect 47760 172 48030 191
rect 49648 230 49918 250
rect 49648 225 49785 230
rect 49648 191 49664 225
rect 49698 196 49785 225
rect 49819 196 49918 230
rect 49698 191 49918 196
rect 49648 172 49918 191
rect 51536 230 51806 250
rect 51536 225 51673 230
rect 51536 191 51552 225
rect 51586 196 51673 225
rect 51707 196 51806 230
rect 51586 191 51806 196
rect 51536 172 51806 191
rect 53424 230 53694 250
rect 53424 225 53561 230
rect 53424 191 53440 225
rect 53474 196 53561 225
rect 53595 196 53694 230
rect 53474 191 53694 196
rect 53424 172 53694 191
rect 55312 230 55582 250
rect 55312 225 55449 230
rect 55312 191 55328 225
rect 55362 196 55449 225
rect 55483 196 55582 230
rect 55362 191 55582 196
rect 55312 172 55582 191
rect 57200 230 57470 250
rect 57200 225 57337 230
rect 57200 191 57216 225
rect 57250 196 57337 225
rect 57371 196 57470 230
rect 57250 191 57470 196
rect 57200 172 57470 191
rect 59088 230 59358 250
rect 59088 225 59225 230
rect 59088 191 59104 225
rect 59138 196 59225 225
rect 59259 196 59358 230
rect 59138 191 59358 196
rect 59088 172 59358 191
<< viali >>
rect 844 7215 878 7249
rect 2732 7215 2766 7249
rect 4620 7215 4654 7249
rect 6508 7215 6542 7249
rect 8396 7215 8430 7249
rect 10284 7215 10318 7249
rect 12172 7215 12206 7249
rect 14060 7215 14094 7249
rect 15942 7215 15976 7249
rect 17830 7215 17864 7249
rect 19718 7215 19752 7249
rect 21606 7215 21640 7249
rect 23494 7215 23528 7249
rect 25382 7215 25416 7249
rect 27270 7215 27304 7249
rect 29158 7215 29192 7249
rect 31046 7215 31080 7249
rect 32934 7215 32968 7249
rect 34822 7215 34856 7249
rect 36710 7215 36744 7249
rect 38598 7215 38632 7249
rect 40486 7215 40520 7249
rect 42374 7215 42408 7249
rect 44262 7215 44296 7249
rect 46144 7215 46178 7249
rect 48032 7215 48066 7249
rect 49920 7215 49954 7249
rect 51808 7215 51842 7249
rect 53696 7215 53730 7249
rect 55584 7215 55618 7249
rect 57472 7215 57506 7249
rect 59360 7215 59394 7249
rect 764 7106 798 7140
rect 2652 7106 2686 7140
rect 4540 7106 4574 7140
rect 6428 7106 6462 7140
rect 8316 7106 8350 7140
rect 10204 7106 10238 7140
rect 12092 7106 12126 7140
rect 13980 7106 14014 7140
rect 15862 7106 15896 7140
rect 17750 7106 17784 7140
rect 19638 7106 19672 7140
rect 21526 7106 21560 7140
rect 23414 7106 23448 7140
rect 25302 7106 25336 7140
rect 27190 7106 27224 7140
rect 29078 7106 29112 7140
rect 30966 7106 31000 7140
rect 32854 7106 32888 7140
rect 34742 7106 34776 7140
rect 36630 7106 36664 7140
rect 38518 7106 38552 7140
rect 40406 7106 40440 7140
rect 42294 7106 42328 7140
rect 44182 7106 44216 7140
rect 46064 7106 46098 7140
rect 47952 7106 47986 7140
rect 49840 7106 49874 7140
rect 51728 7106 51762 7140
rect 53616 7106 53650 7140
rect 55504 7106 55538 7140
rect 57392 7106 57426 7140
rect 59280 7106 59314 7140
rect 620 7054 654 7056
rect 620 7022 654 7054
rect 620 6952 654 6984
rect 620 6950 654 6952
rect 716 7054 750 7056
rect 716 7022 750 7054
rect 812 7054 846 7056
rect 812 7022 846 7054
rect 716 6952 750 6984
rect 716 6950 750 6952
rect 812 6952 846 6984
rect 812 6950 846 6952
rect 2508 7054 2542 7056
rect 2508 7022 2542 7054
rect -363 6845 -329 6879
rect -271 6845 -237 6879
rect -179 6845 -145 6879
rect -17 6843 17 6877
rect 75 6843 109 6877
rect 167 6843 201 6877
rect 668 6866 702 6900
rect 2508 6952 2542 6984
rect 2508 6950 2542 6952
rect 2604 7054 2638 7056
rect 2604 7022 2638 7054
rect 2700 7054 2734 7056
rect 2700 7022 2734 7054
rect 2604 6952 2638 6984
rect 2604 6950 2638 6952
rect 2700 6952 2734 6984
rect 2700 6950 2734 6952
rect 4396 7054 4430 7056
rect 4396 7022 4430 7054
rect 36 6729 70 6746
rect 36 6712 70 6729
rect 396 6828 430 6862
rect 1028 6856 1062 6890
rect 1179 6851 1213 6885
rect 1271 6851 1305 6885
rect 1363 6851 1397 6885
rect 780 6785 814 6819
rect -378 6602 -344 6636
rect -185 6647 -151 6648
rect -185 6614 -153 6647
rect -153 6614 -151 6647
rect 636 6689 670 6691
rect 354 6625 388 6659
rect 636 6657 670 6689
rect 636 6587 670 6619
rect 636 6585 670 6587
rect 310 6529 344 6531
rect 310 6497 344 6529
rect 310 6427 344 6459
rect 310 6425 344 6427
rect -363 6301 -329 6335
rect -271 6301 -237 6335
rect -179 6301 -145 6335
rect 732 6689 766 6691
rect 732 6657 766 6689
rect 732 6587 766 6619
rect 732 6585 766 6587
rect 828 6689 862 6691
rect 828 6657 862 6689
rect 1525 6845 1559 6879
rect 1617 6845 1651 6879
rect 1709 6845 1743 6879
rect 1000 6625 1034 6659
rect 828 6587 862 6619
rect 828 6585 862 6587
rect 398 6529 432 6531
rect 398 6497 432 6529
rect 956 6529 990 6531
rect 956 6497 990 6529
rect 398 6427 432 6459
rect 684 6457 718 6491
rect 398 6425 432 6427
rect 956 6427 990 6459
rect 956 6425 990 6427
rect 1044 6529 1078 6531
rect 1044 6497 1078 6529
rect 1044 6427 1078 6459
rect 1044 6425 1078 6427
rect -17 6299 17 6333
rect 75 6299 109 6333
rect 167 6299 201 6333
rect 753 6349 787 6383
rect 1871 6843 1905 6877
rect 1963 6843 1997 6877
rect 2055 6843 2089 6877
rect 2556 6866 2590 6900
rect 4396 6952 4430 6984
rect 4396 6950 4430 6952
rect 4492 7054 4526 7056
rect 4492 7022 4526 7054
rect 4588 7054 4622 7056
rect 4588 7022 4622 7054
rect 4492 6952 4526 6984
rect 4492 6950 4526 6952
rect 4588 6952 4622 6984
rect 4588 6950 4622 6952
rect 6284 7054 6318 7056
rect 6284 7022 6318 7054
rect 1314 6619 1346 6642
rect 1346 6619 1348 6642
rect 1314 6608 1348 6619
rect 1924 6729 1958 6746
rect 1924 6712 1958 6729
rect 2284 6828 2318 6862
rect 2916 6856 2950 6890
rect 3067 6851 3101 6885
rect 3159 6851 3193 6885
rect 3251 6851 3285 6885
rect 2668 6785 2702 6819
rect 1510 6602 1544 6636
rect 354 6297 388 6331
rect 1703 6647 1737 6648
rect 1703 6614 1735 6647
rect 1735 6614 1737 6647
rect 2524 6689 2558 6691
rect 2242 6625 2276 6659
rect 2524 6657 2558 6689
rect 2524 6587 2558 6619
rect 2524 6585 2558 6587
rect 1000 6297 1034 6331
rect 1179 6307 1213 6341
rect 1271 6307 1305 6341
rect 1363 6307 1397 6341
rect 2198 6529 2232 6531
rect 2198 6497 2232 6529
rect 2198 6427 2232 6459
rect 2198 6425 2232 6427
rect 1525 6301 1559 6335
rect 1617 6301 1651 6335
rect 1709 6301 1743 6335
rect 2620 6689 2654 6691
rect 2620 6657 2654 6689
rect 2620 6587 2654 6619
rect 2620 6585 2654 6587
rect 2716 6689 2750 6691
rect 2716 6657 2750 6689
rect 3413 6845 3447 6879
rect 3505 6845 3539 6879
rect 3597 6845 3631 6879
rect 2888 6625 2922 6659
rect 2716 6587 2750 6619
rect 2716 6585 2750 6587
rect 2286 6529 2320 6531
rect 2286 6497 2320 6529
rect 2844 6529 2878 6531
rect 2844 6497 2878 6529
rect 2286 6427 2320 6459
rect 2572 6457 2606 6491
rect 2286 6425 2320 6427
rect 2844 6427 2878 6459
rect 2844 6425 2878 6427
rect 2932 6529 2966 6531
rect 2932 6497 2966 6529
rect 2932 6427 2966 6459
rect 2932 6425 2966 6427
rect 1871 6299 1905 6333
rect 1963 6299 1997 6333
rect 2055 6299 2089 6333
rect 412 6176 446 6210
rect 842 6159 876 6193
rect 762 6050 796 6084
rect 618 5998 652 6000
rect 618 5966 652 5998
rect 618 5896 652 5928
rect 618 5894 652 5896
rect 714 5998 748 6000
rect 714 5966 748 5998
rect 714 5896 748 5928
rect 714 5894 748 5896
rect 810 5998 844 6000
rect 810 5966 844 5998
rect 810 5896 844 5928
rect 810 5894 844 5896
rect 187 5797 221 5831
rect 279 5797 313 5831
rect 371 5797 405 5831
rect 666 5810 700 5844
rect 279 5685 313 5715
rect 279 5681 281 5685
rect 281 5681 313 5685
rect 778 5729 812 5763
rect 193 5565 195 5592
rect 195 5565 227 5592
rect 193 5558 227 5565
rect 634 5633 668 5635
rect 634 5601 668 5633
rect 367 5565 397 5592
rect 397 5565 401 5592
rect 367 5558 401 5565
rect 634 5531 668 5563
rect 634 5529 668 5531
rect 730 5633 764 5635
rect 730 5601 764 5633
rect 730 5531 764 5563
rect 730 5529 764 5531
rect 826 5633 860 5635
rect 826 5601 860 5633
rect 826 5531 860 5563
rect 826 5529 860 5531
rect 1214 6042 1248 6076
rect 2641 6349 2675 6383
rect 3759 6843 3793 6877
rect 3851 6843 3885 6877
rect 3943 6843 3977 6877
rect 4444 6866 4478 6900
rect 6284 6952 6318 6984
rect 6284 6950 6318 6952
rect 6380 7054 6414 7056
rect 6380 7022 6414 7054
rect 6476 7054 6510 7056
rect 6476 7022 6510 7054
rect 6380 6952 6414 6984
rect 6380 6950 6414 6952
rect 6476 6952 6510 6984
rect 6476 6950 6510 6952
rect 8172 7054 8206 7056
rect 8172 7022 8206 7054
rect 3202 6619 3234 6642
rect 3234 6619 3236 6642
rect 3202 6608 3236 6619
rect 3812 6729 3846 6746
rect 3812 6712 3846 6729
rect 4172 6828 4206 6862
rect 4804 6856 4838 6890
rect 4955 6851 4989 6885
rect 5047 6851 5081 6885
rect 5139 6851 5173 6885
rect 4556 6785 4590 6819
rect 3398 6602 3432 6636
rect 2242 6297 2276 6331
rect 3591 6647 3625 6648
rect 3591 6614 3623 6647
rect 3623 6614 3625 6647
rect 4412 6689 4446 6691
rect 4130 6625 4164 6659
rect 4412 6657 4446 6689
rect 4412 6587 4446 6619
rect 4412 6585 4446 6587
rect 2888 6297 2922 6331
rect 3067 6307 3101 6341
rect 3159 6307 3193 6341
rect 3251 6307 3285 6341
rect 4086 6529 4120 6531
rect 4086 6497 4120 6529
rect 4086 6427 4120 6459
rect 4086 6425 4120 6427
rect 3413 6301 3447 6335
rect 3505 6301 3539 6335
rect 3597 6301 3631 6335
rect 4508 6689 4542 6691
rect 4508 6657 4542 6689
rect 4508 6587 4542 6619
rect 4508 6585 4542 6587
rect 4604 6689 4638 6691
rect 4604 6657 4638 6689
rect 5301 6845 5335 6879
rect 5393 6845 5427 6879
rect 5485 6845 5519 6879
rect 4776 6625 4810 6659
rect 4604 6587 4638 6619
rect 4604 6585 4638 6587
rect 4174 6529 4208 6531
rect 4174 6497 4208 6529
rect 4732 6529 4766 6531
rect 4732 6497 4766 6529
rect 4174 6427 4208 6459
rect 4460 6457 4494 6491
rect 4174 6425 4208 6427
rect 4732 6427 4766 6459
rect 4732 6425 4766 6427
rect 4820 6529 4854 6531
rect 4820 6497 4854 6529
rect 4820 6427 4854 6459
rect 4820 6425 4854 6427
rect 3759 6299 3793 6333
rect 3851 6299 3885 6333
rect 3943 6299 3977 6333
rect 2300 6176 2334 6210
rect 2730 6159 2764 6193
rect 2650 6050 2684 6084
rect 2506 5998 2540 6000
rect 2506 5966 2540 5998
rect 2506 5896 2540 5928
rect 2506 5894 2540 5896
rect 2602 5998 2636 6000
rect 2602 5966 2636 5998
rect 2602 5896 2636 5928
rect 2602 5894 2636 5896
rect 2698 5998 2732 6000
rect 2698 5966 2732 5998
rect 2698 5896 2732 5928
rect 2698 5894 2732 5896
rect 1001 5797 1035 5831
rect 1093 5797 1127 5831
rect 1185 5797 1219 5831
rect 2075 5797 2109 5831
rect 2167 5797 2201 5831
rect 2259 5797 2293 5831
rect 2554 5810 2588 5844
rect 1097 5685 1131 5710
rect 1097 5676 1129 5685
rect 1129 5676 1131 5685
rect 2167 5685 2201 5715
rect 2167 5681 2169 5685
rect 2169 5681 2201 5685
rect 2666 5729 2700 5763
rect 1006 5565 1009 5594
rect 1009 5565 1040 5594
rect 1006 5560 1040 5565
rect 1179 5565 1211 5590
rect 1211 5565 1213 5590
rect 1179 5556 1213 5565
rect 2081 5565 2083 5592
rect 2083 5565 2115 5592
rect 2081 5558 2115 5565
rect 2522 5633 2556 5635
rect 2522 5601 2556 5633
rect 2255 5565 2285 5592
rect 2285 5565 2289 5592
rect 2255 5558 2289 5565
rect 2522 5531 2556 5563
rect 2522 5529 2556 5531
rect 682 5401 716 5435
rect 751 5293 785 5327
rect 2618 5633 2652 5635
rect 2618 5601 2652 5633
rect 2618 5531 2652 5563
rect 2618 5529 2652 5531
rect 2714 5633 2748 5635
rect 2714 5601 2748 5633
rect 2714 5531 2748 5563
rect 2714 5529 2748 5531
rect 3102 6042 3136 6076
rect 4529 6349 4563 6383
rect 5647 6843 5681 6877
rect 5739 6843 5773 6877
rect 5831 6843 5865 6877
rect 6332 6866 6366 6900
rect 8172 6952 8206 6984
rect 8172 6950 8206 6952
rect 8268 7054 8302 7056
rect 8268 7022 8302 7054
rect 8364 7054 8398 7056
rect 8364 7022 8398 7054
rect 8268 6952 8302 6984
rect 8268 6950 8302 6952
rect 8364 6952 8398 6984
rect 8364 6950 8398 6952
rect 10060 7054 10094 7056
rect 10060 7022 10094 7054
rect 5090 6619 5122 6642
rect 5122 6619 5124 6642
rect 5090 6608 5124 6619
rect 5700 6729 5734 6746
rect 5700 6712 5734 6729
rect 6060 6828 6094 6862
rect 6692 6856 6726 6890
rect 6843 6851 6877 6885
rect 6935 6851 6969 6885
rect 7027 6851 7061 6885
rect 6444 6785 6478 6819
rect 5286 6602 5320 6636
rect 4130 6297 4164 6331
rect 5479 6647 5513 6648
rect 5479 6614 5511 6647
rect 5511 6614 5513 6647
rect 6300 6689 6334 6691
rect 6018 6625 6052 6659
rect 6300 6657 6334 6689
rect 6300 6587 6334 6619
rect 6300 6585 6334 6587
rect 4776 6297 4810 6331
rect 4955 6307 4989 6341
rect 5047 6307 5081 6341
rect 5139 6307 5173 6341
rect 5974 6529 6008 6531
rect 5974 6497 6008 6529
rect 5974 6427 6008 6459
rect 5974 6425 6008 6427
rect 5301 6301 5335 6335
rect 5393 6301 5427 6335
rect 5485 6301 5519 6335
rect 6396 6689 6430 6691
rect 6396 6657 6430 6689
rect 6396 6587 6430 6619
rect 6396 6585 6430 6587
rect 6492 6689 6526 6691
rect 6492 6657 6526 6689
rect 7189 6845 7223 6879
rect 7281 6845 7315 6879
rect 7373 6845 7407 6879
rect 6664 6625 6698 6659
rect 6492 6587 6526 6619
rect 6492 6585 6526 6587
rect 6062 6529 6096 6531
rect 6062 6497 6096 6529
rect 6620 6529 6654 6531
rect 6620 6497 6654 6529
rect 6062 6427 6096 6459
rect 6348 6457 6382 6491
rect 6062 6425 6096 6427
rect 6620 6427 6654 6459
rect 6620 6425 6654 6427
rect 6708 6529 6742 6531
rect 6708 6497 6742 6529
rect 6708 6427 6742 6459
rect 6708 6425 6742 6427
rect 5647 6299 5681 6333
rect 5739 6299 5773 6333
rect 5831 6299 5865 6333
rect 4188 6176 4222 6210
rect 4618 6159 4652 6193
rect 4538 6050 4572 6084
rect 4394 5998 4428 6000
rect 4394 5966 4428 5998
rect 4394 5896 4428 5928
rect 4394 5894 4428 5896
rect 4490 5998 4524 6000
rect 4490 5966 4524 5998
rect 4490 5896 4524 5928
rect 4490 5894 4524 5896
rect 4586 5998 4620 6000
rect 4586 5966 4620 5998
rect 4586 5896 4620 5928
rect 4586 5894 4620 5896
rect 2889 5797 2923 5831
rect 2981 5797 3015 5831
rect 3073 5797 3107 5831
rect 3963 5797 3997 5831
rect 4055 5797 4089 5831
rect 4147 5797 4181 5831
rect 4442 5810 4476 5844
rect 2985 5685 3019 5710
rect 2985 5676 3017 5685
rect 3017 5676 3019 5685
rect 4055 5685 4089 5715
rect 4055 5681 4057 5685
rect 4057 5681 4089 5685
rect 4554 5729 4588 5763
rect 2894 5565 2897 5594
rect 2897 5565 2928 5594
rect 2894 5560 2928 5565
rect 3067 5565 3099 5590
rect 3099 5565 3101 5590
rect 3067 5556 3101 5565
rect 3969 5565 3971 5592
rect 3971 5565 4003 5592
rect 3969 5558 4003 5565
rect 4410 5633 4444 5635
rect 4410 5601 4444 5633
rect 4143 5565 4173 5592
rect 4173 5565 4177 5592
rect 4143 5558 4177 5565
rect 4410 5531 4444 5563
rect 4410 5529 4444 5531
rect 2570 5401 2604 5435
rect 2639 5293 2673 5327
rect 4506 5633 4540 5635
rect 4506 5601 4540 5633
rect 4506 5531 4540 5563
rect 4506 5529 4540 5531
rect 4602 5633 4636 5635
rect 4602 5601 4636 5633
rect 4602 5531 4636 5563
rect 4602 5529 4636 5531
rect 4990 6042 5024 6076
rect 6417 6349 6451 6383
rect 7535 6843 7569 6877
rect 7627 6843 7661 6877
rect 7719 6843 7753 6877
rect 8220 6866 8254 6900
rect 10060 6952 10094 6984
rect 10060 6950 10094 6952
rect 10156 7054 10190 7056
rect 10156 7022 10190 7054
rect 10252 7054 10286 7056
rect 10252 7022 10286 7054
rect 10156 6952 10190 6984
rect 10156 6950 10190 6952
rect 10252 6952 10286 6984
rect 10252 6950 10286 6952
rect 11948 7054 11982 7056
rect 11948 7022 11982 7054
rect 6978 6619 7010 6642
rect 7010 6619 7012 6642
rect 6978 6608 7012 6619
rect 7588 6729 7622 6746
rect 7588 6712 7622 6729
rect 7948 6828 7982 6862
rect 8580 6856 8614 6890
rect 8731 6851 8765 6885
rect 8823 6851 8857 6885
rect 8915 6851 8949 6885
rect 8332 6785 8366 6819
rect 7174 6602 7208 6636
rect 6018 6297 6052 6331
rect 7367 6647 7401 6648
rect 7367 6614 7399 6647
rect 7399 6614 7401 6647
rect 8188 6689 8222 6691
rect 7906 6625 7940 6659
rect 8188 6657 8222 6689
rect 8188 6587 8222 6619
rect 8188 6585 8222 6587
rect 6664 6297 6698 6331
rect 6843 6307 6877 6341
rect 6935 6307 6969 6341
rect 7027 6307 7061 6341
rect 7862 6529 7896 6531
rect 7862 6497 7896 6529
rect 7862 6427 7896 6459
rect 7862 6425 7896 6427
rect 7189 6301 7223 6335
rect 7281 6301 7315 6335
rect 7373 6301 7407 6335
rect 8284 6689 8318 6691
rect 8284 6657 8318 6689
rect 8284 6587 8318 6619
rect 8284 6585 8318 6587
rect 8380 6689 8414 6691
rect 8380 6657 8414 6689
rect 9077 6845 9111 6879
rect 9169 6845 9203 6879
rect 9261 6845 9295 6879
rect 8552 6625 8586 6659
rect 8380 6587 8414 6619
rect 8380 6585 8414 6587
rect 7950 6529 7984 6531
rect 7950 6497 7984 6529
rect 8508 6529 8542 6531
rect 8508 6497 8542 6529
rect 7950 6427 7984 6459
rect 8236 6457 8270 6491
rect 7950 6425 7984 6427
rect 8508 6427 8542 6459
rect 8508 6425 8542 6427
rect 8596 6529 8630 6531
rect 8596 6497 8630 6529
rect 8596 6427 8630 6459
rect 8596 6425 8630 6427
rect 7535 6299 7569 6333
rect 7627 6299 7661 6333
rect 7719 6299 7753 6333
rect 6076 6176 6110 6210
rect 6506 6159 6540 6193
rect 6426 6050 6460 6084
rect 6282 5998 6316 6000
rect 6282 5966 6316 5998
rect 6282 5896 6316 5928
rect 6282 5894 6316 5896
rect 6378 5998 6412 6000
rect 6378 5966 6412 5998
rect 6378 5896 6412 5928
rect 6378 5894 6412 5896
rect 6474 5998 6508 6000
rect 6474 5966 6508 5998
rect 6474 5896 6508 5928
rect 6474 5894 6508 5896
rect 4777 5797 4811 5831
rect 4869 5797 4903 5831
rect 4961 5797 4995 5831
rect 5851 5797 5885 5831
rect 5943 5797 5977 5831
rect 6035 5797 6069 5831
rect 6330 5810 6364 5844
rect 4873 5685 4907 5710
rect 4873 5676 4905 5685
rect 4905 5676 4907 5685
rect 5943 5685 5977 5715
rect 5943 5681 5945 5685
rect 5945 5681 5977 5685
rect 6442 5729 6476 5763
rect 4782 5565 4785 5594
rect 4785 5565 4816 5594
rect 4782 5560 4816 5565
rect 4955 5565 4987 5590
rect 4987 5565 4989 5590
rect 4955 5556 4989 5565
rect 5857 5565 5859 5592
rect 5859 5565 5891 5592
rect 5857 5558 5891 5565
rect 6298 5633 6332 5635
rect 6298 5601 6332 5633
rect 6031 5565 6061 5592
rect 6061 5565 6065 5592
rect 6031 5558 6065 5565
rect 6298 5531 6332 5563
rect 6298 5529 6332 5531
rect 4458 5401 4492 5435
rect 4527 5293 4561 5327
rect 6394 5633 6428 5635
rect 6394 5601 6428 5633
rect 6394 5531 6428 5563
rect 6394 5529 6428 5531
rect 6490 5633 6524 5635
rect 6490 5601 6524 5633
rect 6490 5531 6524 5563
rect 6490 5529 6524 5531
rect 6878 6042 6912 6076
rect 8305 6349 8339 6383
rect 9423 6843 9457 6877
rect 9515 6843 9549 6877
rect 9607 6843 9641 6877
rect 10108 6866 10142 6900
rect 11948 6952 11982 6984
rect 11948 6950 11982 6952
rect 12044 7054 12078 7056
rect 12044 7022 12078 7054
rect 12140 7054 12174 7056
rect 12140 7022 12174 7054
rect 12044 6952 12078 6984
rect 12044 6950 12078 6952
rect 12140 6952 12174 6984
rect 12140 6950 12174 6952
rect 13836 7054 13870 7056
rect 13836 7022 13870 7054
rect 8866 6619 8898 6642
rect 8898 6619 8900 6642
rect 8866 6608 8900 6619
rect 9476 6729 9510 6746
rect 9476 6712 9510 6729
rect 9836 6828 9870 6862
rect 10468 6856 10502 6890
rect 10619 6851 10653 6885
rect 10711 6851 10745 6885
rect 10803 6851 10837 6885
rect 10220 6785 10254 6819
rect 9062 6602 9096 6636
rect 7906 6297 7940 6331
rect 9255 6647 9289 6648
rect 9255 6614 9287 6647
rect 9287 6614 9289 6647
rect 10076 6689 10110 6691
rect 9794 6625 9828 6659
rect 10076 6657 10110 6689
rect 10076 6587 10110 6619
rect 10076 6585 10110 6587
rect 8552 6297 8586 6331
rect 8731 6307 8765 6341
rect 8823 6307 8857 6341
rect 8915 6307 8949 6341
rect 9750 6529 9784 6531
rect 9750 6497 9784 6529
rect 9750 6427 9784 6459
rect 9750 6425 9784 6427
rect 9077 6301 9111 6335
rect 9169 6301 9203 6335
rect 9261 6301 9295 6335
rect 10172 6689 10206 6691
rect 10172 6657 10206 6689
rect 10172 6587 10206 6619
rect 10172 6585 10206 6587
rect 10268 6689 10302 6691
rect 10268 6657 10302 6689
rect 10965 6845 10999 6879
rect 11057 6845 11091 6879
rect 11149 6845 11183 6879
rect 10440 6625 10474 6659
rect 10268 6587 10302 6619
rect 10268 6585 10302 6587
rect 9838 6529 9872 6531
rect 9838 6497 9872 6529
rect 10396 6529 10430 6531
rect 10396 6497 10430 6529
rect 9838 6427 9872 6459
rect 10124 6457 10158 6491
rect 9838 6425 9872 6427
rect 10396 6427 10430 6459
rect 10396 6425 10430 6427
rect 10484 6529 10518 6531
rect 10484 6497 10518 6529
rect 10484 6427 10518 6459
rect 10484 6425 10518 6427
rect 9423 6299 9457 6333
rect 9515 6299 9549 6333
rect 9607 6299 9641 6333
rect 7964 6176 7998 6210
rect 8394 6159 8428 6193
rect 8314 6050 8348 6084
rect 8170 5998 8204 6000
rect 8170 5966 8204 5998
rect 8170 5896 8204 5928
rect 8170 5894 8204 5896
rect 8266 5998 8300 6000
rect 8266 5966 8300 5998
rect 8266 5896 8300 5928
rect 8266 5894 8300 5896
rect 8362 5998 8396 6000
rect 8362 5966 8396 5998
rect 8362 5896 8396 5928
rect 8362 5894 8396 5896
rect 6665 5797 6699 5831
rect 6757 5797 6791 5831
rect 6849 5797 6883 5831
rect 7739 5797 7773 5831
rect 7831 5797 7865 5831
rect 7923 5797 7957 5831
rect 8218 5810 8252 5844
rect 6761 5685 6795 5710
rect 6761 5676 6793 5685
rect 6793 5676 6795 5685
rect 7831 5685 7865 5715
rect 7831 5681 7833 5685
rect 7833 5681 7865 5685
rect 8330 5729 8364 5763
rect 6670 5565 6673 5594
rect 6673 5565 6704 5594
rect 6670 5560 6704 5565
rect 6843 5565 6875 5590
rect 6875 5565 6877 5590
rect 6843 5556 6877 5565
rect 7745 5565 7747 5592
rect 7747 5565 7779 5592
rect 7745 5558 7779 5565
rect 8186 5633 8220 5635
rect 8186 5601 8220 5633
rect 7919 5565 7949 5592
rect 7949 5565 7953 5592
rect 7919 5558 7953 5565
rect 8186 5531 8220 5563
rect 8186 5529 8220 5531
rect 6346 5401 6380 5435
rect 6415 5293 6449 5327
rect 8282 5633 8316 5635
rect 8282 5601 8316 5633
rect 8282 5531 8316 5563
rect 8282 5529 8316 5531
rect 8378 5633 8412 5635
rect 8378 5601 8412 5633
rect 8378 5531 8412 5563
rect 8378 5529 8412 5531
rect 8766 6042 8800 6076
rect 10193 6349 10227 6383
rect 11311 6843 11345 6877
rect 11403 6843 11437 6877
rect 11495 6843 11529 6877
rect 11996 6866 12030 6900
rect 13836 6952 13870 6984
rect 13836 6950 13870 6952
rect 13932 7054 13966 7056
rect 13932 7022 13966 7054
rect 14028 7054 14062 7056
rect 14028 7022 14062 7054
rect 13932 6952 13966 6984
rect 13932 6950 13966 6952
rect 14028 6952 14062 6984
rect 14028 6950 14062 6952
rect 15718 7054 15752 7056
rect 15718 7022 15752 7054
rect 10754 6619 10786 6642
rect 10786 6619 10788 6642
rect 10754 6608 10788 6619
rect 11364 6729 11398 6746
rect 11364 6712 11398 6729
rect 11724 6828 11758 6862
rect 12356 6856 12390 6890
rect 12507 6851 12541 6885
rect 12599 6851 12633 6885
rect 12691 6851 12725 6885
rect 12108 6785 12142 6819
rect 10950 6602 10984 6636
rect 9794 6297 9828 6331
rect 11143 6647 11177 6648
rect 11143 6614 11175 6647
rect 11175 6614 11177 6647
rect 11964 6689 11998 6691
rect 11682 6625 11716 6659
rect 11964 6657 11998 6689
rect 11964 6587 11998 6619
rect 11964 6585 11998 6587
rect 10440 6297 10474 6331
rect 10619 6307 10653 6341
rect 10711 6307 10745 6341
rect 10803 6307 10837 6341
rect 11638 6529 11672 6531
rect 11638 6497 11672 6529
rect 11638 6427 11672 6459
rect 11638 6425 11672 6427
rect 10965 6301 10999 6335
rect 11057 6301 11091 6335
rect 11149 6301 11183 6335
rect 12060 6689 12094 6691
rect 12060 6657 12094 6689
rect 12060 6587 12094 6619
rect 12060 6585 12094 6587
rect 12156 6689 12190 6691
rect 12156 6657 12190 6689
rect 12853 6845 12887 6879
rect 12945 6845 12979 6879
rect 13037 6845 13071 6879
rect 12328 6625 12362 6659
rect 12156 6587 12190 6619
rect 12156 6585 12190 6587
rect 11726 6529 11760 6531
rect 11726 6497 11760 6529
rect 12284 6529 12318 6531
rect 12284 6497 12318 6529
rect 11726 6427 11760 6459
rect 12012 6457 12046 6491
rect 11726 6425 11760 6427
rect 12284 6427 12318 6459
rect 12284 6425 12318 6427
rect 12372 6529 12406 6531
rect 12372 6497 12406 6529
rect 12372 6427 12406 6459
rect 12372 6425 12406 6427
rect 11311 6299 11345 6333
rect 11403 6299 11437 6333
rect 11495 6299 11529 6333
rect 9852 6176 9886 6210
rect 10282 6159 10316 6193
rect 10202 6050 10236 6084
rect 10058 5998 10092 6000
rect 10058 5966 10092 5998
rect 10058 5896 10092 5928
rect 10058 5894 10092 5896
rect 10154 5998 10188 6000
rect 10154 5966 10188 5998
rect 10154 5896 10188 5928
rect 10154 5894 10188 5896
rect 10250 5998 10284 6000
rect 10250 5966 10284 5998
rect 10250 5896 10284 5928
rect 10250 5894 10284 5896
rect 8553 5797 8587 5831
rect 8645 5797 8679 5831
rect 8737 5797 8771 5831
rect 9627 5797 9661 5831
rect 9719 5797 9753 5831
rect 9811 5797 9845 5831
rect 10106 5810 10140 5844
rect 8649 5685 8683 5710
rect 8649 5676 8681 5685
rect 8681 5676 8683 5685
rect 9719 5685 9753 5715
rect 9719 5681 9721 5685
rect 9721 5681 9753 5685
rect 10218 5729 10252 5763
rect 8558 5565 8561 5594
rect 8561 5565 8592 5594
rect 8558 5560 8592 5565
rect 8731 5565 8763 5590
rect 8763 5565 8765 5590
rect 8731 5556 8765 5565
rect 9633 5565 9635 5592
rect 9635 5565 9667 5592
rect 9633 5558 9667 5565
rect 10074 5633 10108 5635
rect 10074 5601 10108 5633
rect 9807 5565 9837 5592
rect 9837 5565 9841 5592
rect 9807 5558 9841 5565
rect 10074 5531 10108 5563
rect 10074 5529 10108 5531
rect 8234 5401 8268 5435
rect 8303 5293 8337 5327
rect 10170 5633 10204 5635
rect 10170 5601 10204 5633
rect 10170 5531 10204 5563
rect 10170 5529 10204 5531
rect 10266 5633 10300 5635
rect 10266 5601 10300 5633
rect 10266 5531 10300 5563
rect 10266 5529 10300 5531
rect 10654 6042 10688 6076
rect 12081 6349 12115 6383
rect 13199 6843 13233 6877
rect 13291 6843 13325 6877
rect 13383 6843 13417 6877
rect 13884 6866 13918 6900
rect 15718 6952 15752 6984
rect 15718 6950 15752 6952
rect 15814 7054 15848 7056
rect 15814 7022 15848 7054
rect 15910 7054 15944 7056
rect 15910 7022 15944 7054
rect 15814 6952 15848 6984
rect 15814 6950 15848 6952
rect 15910 6952 15944 6984
rect 15910 6950 15944 6952
rect 17606 7054 17640 7056
rect 17606 7022 17640 7054
rect 12642 6619 12674 6642
rect 12674 6619 12676 6642
rect 12642 6608 12676 6619
rect 13252 6729 13286 6746
rect 13252 6712 13286 6729
rect 13612 6828 13646 6862
rect 14244 6856 14278 6890
rect 14395 6851 14429 6885
rect 14487 6851 14521 6885
rect 14579 6851 14613 6885
rect 13996 6785 14030 6819
rect 12838 6602 12872 6636
rect 11682 6297 11716 6331
rect 13031 6647 13065 6648
rect 13031 6614 13063 6647
rect 13063 6614 13065 6647
rect 13852 6689 13886 6691
rect 13570 6625 13604 6659
rect 13852 6657 13886 6689
rect 13852 6587 13886 6619
rect 13852 6585 13886 6587
rect 12328 6297 12362 6331
rect 12507 6307 12541 6341
rect 12599 6307 12633 6341
rect 12691 6307 12725 6341
rect 13526 6529 13560 6531
rect 13526 6497 13560 6529
rect 13526 6427 13560 6459
rect 13526 6425 13560 6427
rect 12853 6301 12887 6335
rect 12945 6301 12979 6335
rect 13037 6301 13071 6335
rect 13948 6689 13982 6691
rect 13948 6657 13982 6689
rect 13948 6587 13982 6619
rect 13948 6585 13982 6587
rect 14044 6689 14078 6691
rect 14044 6657 14078 6689
rect 14735 6845 14769 6879
rect 14827 6845 14861 6879
rect 14919 6845 14953 6879
rect 14216 6625 14250 6659
rect 14044 6587 14078 6619
rect 14044 6585 14078 6587
rect 13614 6529 13648 6531
rect 13614 6497 13648 6529
rect 14172 6529 14206 6531
rect 14172 6497 14206 6529
rect 13614 6427 13648 6459
rect 13900 6457 13934 6491
rect 13614 6425 13648 6427
rect 14172 6427 14206 6459
rect 14172 6425 14206 6427
rect 14260 6529 14294 6531
rect 14260 6497 14294 6529
rect 14260 6427 14294 6459
rect 14260 6425 14294 6427
rect 13199 6299 13233 6333
rect 13291 6299 13325 6333
rect 13383 6299 13417 6333
rect 11740 6176 11774 6210
rect 12170 6159 12204 6193
rect 12090 6050 12124 6084
rect 11946 5998 11980 6000
rect 11946 5966 11980 5998
rect 11946 5896 11980 5928
rect 11946 5894 11980 5896
rect 12042 5998 12076 6000
rect 12042 5966 12076 5998
rect 12042 5896 12076 5928
rect 12042 5894 12076 5896
rect 12138 5998 12172 6000
rect 12138 5966 12172 5998
rect 12138 5896 12172 5928
rect 12138 5894 12172 5896
rect 10441 5797 10475 5831
rect 10533 5797 10567 5831
rect 10625 5797 10659 5831
rect 11515 5797 11549 5831
rect 11607 5797 11641 5831
rect 11699 5797 11733 5831
rect 11994 5810 12028 5844
rect 10537 5685 10571 5710
rect 10537 5676 10569 5685
rect 10569 5676 10571 5685
rect 11607 5685 11641 5715
rect 11607 5681 11609 5685
rect 11609 5681 11641 5685
rect 12106 5729 12140 5763
rect 10446 5565 10449 5594
rect 10449 5565 10480 5594
rect 10446 5560 10480 5565
rect 10619 5565 10651 5590
rect 10651 5565 10653 5590
rect 10619 5556 10653 5565
rect 11521 5565 11523 5592
rect 11523 5565 11555 5592
rect 11521 5558 11555 5565
rect 11962 5633 11996 5635
rect 11962 5601 11996 5633
rect 11695 5565 11725 5592
rect 11725 5565 11729 5592
rect 11695 5558 11729 5565
rect 11962 5531 11996 5563
rect 11962 5529 11996 5531
rect 10122 5401 10156 5435
rect 10191 5293 10225 5327
rect 12058 5633 12092 5635
rect 12058 5601 12092 5633
rect 12058 5531 12092 5563
rect 12058 5529 12092 5531
rect 12154 5633 12188 5635
rect 12154 5601 12188 5633
rect 12154 5531 12188 5563
rect 12154 5529 12188 5531
rect 12542 6042 12576 6076
rect 13969 6349 14003 6383
rect 15081 6843 15115 6877
rect 15173 6843 15207 6877
rect 15265 6843 15299 6877
rect 15766 6866 15800 6900
rect 17606 6952 17640 6984
rect 17606 6950 17640 6952
rect 17702 7054 17736 7056
rect 17702 7022 17736 7054
rect 17798 7054 17832 7056
rect 17798 7022 17832 7054
rect 17702 6952 17736 6984
rect 17702 6950 17736 6952
rect 17798 6952 17832 6984
rect 17798 6950 17832 6952
rect 19494 7054 19528 7056
rect 19494 7022 19528 7054
rect 14530 6619 14562 6642
rect 14562 6619 14564 6642
rect 14530 6608 14564 6619
rect 15134 6729 15168 6746
rect 15134 6712 15168 6729
rect 15494 6828 15528 6862
rect 16126 6856 16160 6890
rect 16277 6851 16311 6885
rect 16369 6851 16403 6885
rect 16461 6851 16495 6885
rect 15878 6785 15912 6819
rect 14720 6602 14754 6636
rect 13570 6297 13604 6331
rect 14913 6647 14947 6648
rect 14913 6614 14945 6647
rect 14945 6614 14947 6647
rect 15734 6689 15768 6691
rect 15452 6625 15486 6659
rect 15734 6657 15768 6689
rect 15734 6587 15768 6619
rect 15734 6585 15768 6587
rect 14216 6297 14250 6331
rect 14395 6307 14429 6341
rect 14487 6307 14521 6341
rect 14579 6307 14613 6341
rect 15408 6529 15442 6531
rect 15408 6497 15442 6529
rect 15408 6427 15442 6459
rect 15408 6425 15442 6427
rect 14735 6301 14769 6335
rect 14827 6301 14861 6335
rect 14919 6301 14953 6335
rect 15830 6689 15864 6691
rect 15830 6657 15864 6689
rect 15830 6587 15864 6619
rect 15830 6585 15864 6587
rect 15926 6689 15960 6691
rect 15926 6657 15960 6689
rect 16623 6845 16657 6879
rect 16715 6845 16749 6879
rect 16807 6845 16841 6879
rect 16098 6625 16132 6659
rect 15926 6587 15960 6619
rect 15926 6585 15960 6587
rect 15496 6529 15530 6531
rect 15496 6497 15530 6529
rect 16054 6529 16088 6531
rect 16054 6497 16088 6529
rect 15496 6427 15530 6459
rect 15782 6457 15816 6491
rect 15496 6425 15530 6427
rect 16054 6427 16088 6459
rect 16054 6425 16088 6427
rect 16142 6529 16176 6531
rect 16142 6497 16176 6529
rect 16142 6427 16176 6459
rect 16142 6425 16176 6427
rect 15081 6299 15115 6333
rect 15173 6299 15207 6333
rect 15265 6299 15299 6333
rect 13628 6176 13662 6210
rect 14058 6159 14092 6193
rect 13978 6050 14012 6084
rect 13834 5998 13868 6000
rect 13834 5966 13868 5998
rect 13834 5896 13868 5928
rect 13834 5894 13868 5896
rect 13930 5998 13964 6000
rect 13930 5966 13964 5998
rect 13930 5896 13964 5928
rect 13930 5894 13964 5896
rect 14026 5998 14060 6000
rect 14026 5966 14060 5998
rect 14026 5896 14060 5928
rect 14026 5894 14060 5896
rect 12329 5797 12363 5831
rect 12421 5797 12455 5831
rect 12513 5797 12547 5831
rect 13403 5797 13437 5831
rect 13495 5797 13529 5831
rect 13587 5797 13621 5831
rect 13882 5810 13916 5844
rect 12425 5685 12459 5710
rect 12425 5676 12457 5685
rect 12457 5676 12459 5685
rect 13495 5685 13529 5715
rect 13495 5681 13497 5685
rect 13497 5681 13529 5685
rect 13994 5729 14028 5763
rect 12334 5565 12337 5594
rect 12337 5565 12368 5594
rect 12334 5560 12368 5565
rect 12507 5565 12539 5590
rect 12539 5565 12541 5590
rect 12507 5556 12541 5565
rect 13409 5565 13411 5592
rect 13411 5565 13443 5592
rect 13409 5558 13443 5565
rect 13850 5633 13884 5635
rect 13850 5601 13884 5633
rect 13583 5565 13613 5592
rect 13613 5565 13617 5592
rect 13583 5558 13617 5565
rect 13850 5531 13884 5563
rect 13850 5529 13884 5531
rect 12010 5401 12044 5435
rect 12079 5293 12113 5327
rect 13946 5633 13980 5635
rect 13946 5601 13980 5633
rect 13946 5531 13980 5563
rect 13946 5529 13980 5531
rect 14042 5633 14076 5635
rect 14042 5601 14076 5633
rect 14042 5531 14076 5563
rect 14042 5529 14076 5531
rect 14430 6042 14464 6076
rect 15851 6349 15885 6383
rect 16969 6843 17003 6877
rect 17061 6843 17095 6877
rect 17153 6843 17187 6877
rect 17654 6866 17688 6900
rect 19494 6952 19528 6984
rect 19494 6950 19528 6952
rect 19590 7054 19624 7056
rect 19590 7022 19624 7054
rect 19686 7054 19720 7056
rect 19686 7022 19720 7054
rect 19590 6952 19624 6984
rect 19590 6950 19624 6952
rect 19686 6952 19720 6984
rect 19686 6950 19720 6952
rect 21382 7054 21416 7056
rect 21382 7022 21416 7054
rect 16412 6619 16444 6642
rect 16444 6619 16446 6642
rect 16412 6608 16446 6619
rect 17022 6729 17056 6746
rect 17022 6712 17056 6729
rect 17382 6828 17416 6862
rect 18014 6856 18048 6890
rect 18165 6851 18199 6885
rect 18257 6851 18291 6885
rect 18349 6851 18383 6885
rect 17766 6785 17800 6819
rect 16608 6602 16642 6636
rect 15452 6297 15486 6331
rect 16801 6647 16835 6648
rect 16801 6614 16833 6647
rect 16833 6614 16835 6647
rect 17622 6689 17656 6691
rect 17340 6625 17374 6659
rect 17622 6657 17656 6689
rect 17622 6587 17656 6619
rect 17622 6585 17656 6587
rect 16098 6297 16132 6331
rect 16277 6307 16311 6341
rect 16369 6307 16403 6341
rect 16461 6307 16495 6341
rect 17296 6529 17330 6531
rect 17296 6497 17330 6529
rect 17296 6427 17330 6459
rect 17296 6425 17330 6427
rect 16623 6301 16657 6335
rect 16715 6301 16749 6335
rect 16807 6301 16841 6335
rect 17718 6689 17752 6691
rect 17718 6657 17752 6689
rect 17718 6587 17752 6619
rect 17718 6585 17752 6587
rect 17814 6689 17848 6691
rect 17814 6657 17848 6689
rect 18511 6845 18545 6879
rect 18603 6845 18637 6879
rect 18695 6845 18729 6879
rect 17986 6625 18020 6659
rect 17814 6587 17848 6619
rect 17814 6585 17848 6587
rect 17384 6529 17418 6531
rect 17384 6497 17418 6529
rect 17942 6529 17976 6531
rect 17942 6497 17976 6529
rect 17384 6427 17418 6459
rect 17670 6457 17704 6491
rect 17384 6425 17418 6427
rect 17942 6427 17976 6459
rect 17942 6425 17976 6427
rect 18030 6529 18064 6531
rect 18030 6497 18064 6529
rect 18030 6427 18064 6459
rect 18030 6425 18064 6427
rect 16969 6299 17003 6333
rect 17061 6299 17095 6333
rect 17153 6299 17187 6333
rect 15510 6176 15544 6210
rect 15940 6159 15974 6193
rect 15860 6050 15894 6084
rect 15716 5998 15750 6000
rect 15716 5966 15750 5998
rect 15716 5896 15750 5928
rect 15716 5894 15750 5896
rect 15812 5998 15846 6000
rect 15812 5966 15846 5998
rect 15812 5896 15846 5928
rect 15812 5894 15846 5896
rect 15908 5998 15942 6000
rect 15908 5966 15942 5998
rect 15908 5896 15942 5928
rect 15908 5894 15942 5896
rect 14217 5797 14251 5831
rect 14309 5797 14343 5831
rect 14401 5797 14435 5831
rect 15285 5797 15319 5831
rect 15377 5797 15411 5831
rect 15469 5797 15503 5831
rect 15764 5810 15798 5844
rect 14313 5685 14347 5710
rect 14313 5676 14345 5685
rect 14345 5676 14347 5685
rect 15377 5685 15411 5715
rect 15377 5681 15379 5685
rect 15379 5681 15411 5685
rect 15876 5729 15910 5763
rect 14222 5565 14225 5594
rect 14225 5565 14256 5594
rect 14222 5560 14256 5565
rect 14395 5565 14427 5590
rect 14427 5565 14429 5590
rect 14395 5556 14429 5565
rect 15291 5565 15293 5592
rect 15293 5565 15325 5592
rect 15291 5558 15325 5565
rect 15732 5633 15766 5635
rect 15732 5601 15766 5633
rect 15465 5565 15495 5592
rect 15495 5565 15499 5592
rect 15465 5558 15499 5565
rect 15732 5531 15766 5563
rect 15732 5529 15766 5531
rect 13898 5401 13932 5435
rect 13967 5293 14001 5327
rect 15828 5633 15862 5635
rect 15828 5601 15862 5633
rect 15828 5531 15862 5563
rect 15828 5529 15862 5531
rect 15924 5633 15958 5635
rect 15924 5601 15958 5633
rect 15924 5531 15958 5563
rect 15924 5529 15958 5531
rect 16312 6042 16346 6076
rect 17739 6349 17773 6383
rect 18857 6843 18891 6877
rect 18949 6843 18983 6877
rect 19041 6843 19075 6877
rect 19542 6866 19576 6900
rect 21382 6952 21416 6984
rect 21382 6950 21416 6952
rect 21478 7054 21512 7056
rect 21478 7022 21512 7054
rect 21574 7054 21608 7056
rect 21574 7022 21608 7054
rect 21478 6952 21512 6984
rect 21478 6950 21512 6952
rect 21574 6952 21608 6984
rect 21574 6950 21608 6952
rect 23270 7054 23304 7056
rect 23270 7022 23304 7054
rect 18300 6619 18332 6642
rect 18332 6619 18334 6642
rect 18300 6608 18334 6619
rect 18910 6729 18944 6746
rect 18910 6712 18944 6729
rect 19270 6828 19304 6862
rect 19902 6856 19936 6890
rect 20053 6851 20087 6885
rect 20145 6851 20179 6885
rect 20237 6851 20271 6885
rect 19654 6785 19688 6819
rect 18496 6602 18530 6636
rect 17340 6297 17374 6331
rect 18689 6647 18723 6648
rect 18689 6614 18721 6647
rect 18721 6614 18723 6647
rect 19510 6689 19544 6691
rect 19228 6625 19262 6659
rect 19510 6657 19544 6689
rect 19510 6587 19544 6619
rect 19510 6585 19544 6587
rect 17986 6297 18020 6331
rect 18165 6307 18199 6341
rect 18257 6307 18291 6341
rect 18349 6307 18383 6341
rect 19184 6529 19218 6531
rect 19184 6497 19218 6529
rect 19184 6427 19218 6459
rect 19184 6425 19218 6427
rect 18511 6301 18545 6335
rect 18603 6301 18637 6335
rect 18695 6301 18729 6335
rect 19606 6689 19640 6691
rect 19606 6657 19640 6689
rect 19606 6587 19640 6619
rect 19606 6585 19640 6587
rect 19702 6689 19736 6691
rect 19702 6657 19736 6689
rect 20399 6845 20433 6879
rect 20491 6845 20525 6879
rect 20583 6845 20617 6879
rect 19874 6625 19908 6659
rect 19702 6587 19736 6619
rect 19702 6585 19736 6587
rect 19272 6529 19306 6531
rect 19272 6497 19306 6529
rect 19830 6529 19864 6531
rect 19830 6497 19864 6529
rect 19272 6427 19306 6459
rect 19558 6457 19592 6491
rect 19272 6425 19306 6427
rect 19830 6427 19864 6459
rect 19830 6425 19864 6427
rect 19918 6529 19952 6531
rect 19918 6497 19952 6529
rect 19918 6427 19952 6459
rect 19918 6425 19952 6427
rect 18857 6299 18891 6333
rect 18949 6299 18983 6333
rect 19041 6299 19075 6333
rect 17398 6176 17432 6210
rect 17828 6159 17862 6193
rect 17748 6050 17782 6084
rect 17604 5998 17638 6000
rect 17604 5966 17638 5998
rect 17604 5896 17638 5928
rect 17604 5894 17638 5896
rect 17700 5998 17734 6000
rect 17700 5966 17734 5998
rect 17700 5896 17734 5928
rect 17700 5894 17734 5896
rect 17796 5998 17830 6000
rect 17796 5966 17830 5998
rect 17796 5896 17830 5928
rect 17796 5894 17830 5896
rect 16099 5797 16133 5831
rect 16191 5797 16225 5831
rect 16283 5797 16317 5831
rect 17173 5797 17207 5831
rect 17265 5797 17299 5831
rect 17357 5797 17391 5831
rect 17652 5810 17686 5844
rect 16195 5685 16229 5710
rect 16195 5676 16227 5685
rect 16227 5676 16229 5685
rect 17265 5685 17299 5715
rect 17265 5681 17267 5685
rect 17267 5681 17299 5685
rect 17764 5729 17798 5763
rect 16104 5565 16107 5594
rect 16107 5565 16138 5594
rect 16104 5560 16138 5565
rect 16277 5565 16309 5590
rect 16309 5565 16311 5590
rect 16277 5556 16311 5565
rect 17179 5565 17181 5592
rect 17181 5565 17213 5592
rect 17179 5558 17213 5565
rect 17620 5633 17654 5635
rect 17620 5601 17654 5633
rect 17353 5565 17383 5592
rect 17383 5565 17387 5592
rect 17353 5558 17387 5565
rect 17620 5531 17654 5563
rect 17620 5529 17654 5531
rect 15780 5401 15814 5435
rect 15849 5293 15883 5327
rect 17716 5633 17750 5635
rect 17716 5601 17750 5633
rect 17716 5531 17750 5563
rect 17716 5529 17750 5531
rect 17812 5633 17846 5635
rect 17812 5601 17846 5633
rect 17812 5531 17846 5563
rect 17812 5529 17846 5531
rect 18200 6042 18234 6076
rect 19627 6349 19661 6383
rect 20745 6843 20779 6877
rect 20837 6843 20871 6877
rect 20929 6843 20963 6877
rect 21430 6866 21464 6900
rect 23270 6952 23304 6984
rect 23270 6950 23304 6952
rect 23366 7054 23400 7056
rect 23366 7022 23400 7054
rect 23462 7054 23496 7056
rect 23462 7022 23496 7054
rect 23366 6952 23400 6984
rect 23366 6950 23400 6952
rect 23462 6952 23496 6984
rect 23462 6950 23496 6952
rect 25158 7054 25192 7056
rect 25158 7022 25192 7054
rect 20188 6619 20220 6642
rect 20220 6619 20222 6642
rect 20188 6608 20222 6619
rect 20798 6729 20832 6746
rect 20798 6712 20832 6729
rect 21158 6828 21192 6862
rect 21790 6856 21824 6890
rect 21941 6851 21975 6885
rect 22033 6851 22067 6885
rect 22125 6851 22159 6885
rect 21542 6785 21576 6819
rect 20384 6602 20418 6636
rect 19228 6297 19262 6331
rect 20577 6647 20611 6648
rect 20577 6614 20609 6647
rect 20609 6614 20611 6647
rect 21398 6689 21432 6691
rect 21116 6625 21150 6659
rect 21398 6657 21432 6689
rect 21398 6587 21432 6619
rect 21398 6585 21432 6587
rect 19874 6297 19908 6331
rect 20053 6307 20087 6341
rect 20145 6307 20179 6341
rect 20237 6307 20271 6341
rect 21072 6529 21106 6531
rect 21072 6497 21106 6529
rect 21072 6427 21106 6459
rect 21072 6425 21106 6427
rect 20399 6301 20433 6335
rect 20491 6301 20525 6335
rect 20583 6301 20617 6335
rect 21494 6689 21528 6691
rect 21494 6657 21528 6689
rect 21494 6587 21528 6619
rect 21494 6585 21528 6587
rect 21590 6689 21624 6691
rect 21590 6657 21624 6689
rect 22287 6845 22321 6879
rect 22379 6845 22413 6879
rect 22471 6845 22505 6879
rect 21762 6625 21796 6659
rect 21590 6587 21624 6619
rect 21590 6585 21624 6587
rect 21160 6529 21194 6531
rect 21160 6497 21194 6529
rect 21718 6529 21752 6531
rect 21718 6497 21752 6529
rect 21160 6427 21194 6459
rect 21446 6457 21480 6491
rect 21160 6425 21194 6427
rect 21718 6427 21752 6459
rect 21718 6425 21752 6427
rect 21806 6529 21840 6531
rect 21806 6497 21840 6529
rect 21806 6427 21840 6459
rect 21806 6425 21840 6427
rect 20745 6299 20779 6333
rect 20837 6299 20871 6333
rect 20929 6299 20963 6333
rect 19286 6176 19320 6210
rect 19716 6159 19750 6193
rect 19636 6050 19670 6084
rect 19492 5998 19526 6000
rect 19492 5966 19526 5998
rect 19492 5896 19526 5928
rect 19492 5894 19526 5896
rect 19588 5998 19622 6000
rect 19588 5966 19622 5998
rect 19588 5896 19622 5928
rect 19588 5894 19622 5896
rect 19684 5998 19718 6000
rect 19684 5966 19718 5998
rect 19684 5896 19718 5928
rect 19684 5894 19718 5896
rect 17987 5797 18021 5831
rect 18079 5797 18113 5831
rect 18171 5797 18205 5831
rect 19061 5797 19095 5831
rect 19153 5797 19187 5831
rect 19245 5797 19279 5831
rect 19540 5810 19574 5844
rect 18083 5685 18117 5710
rect 18083 5676 18115 5685
rect 18115 5676 18117 5685
rect 19153 5685 19187 5715
rect 19153 5681 19155 5685
rect 19155 5681 19187 5685
rect 19652 5729 19686 5763
rect 17992 5565 17995 5594
rect 17995 5565 18026 5594
rect 17992 5560 18026 5565
rect 18165 5565 18197 5590
rect 18197 5565 18199 5590
rect 18165 5556 18199 5565
rect 19067 5565 19069 5592
rect 19069 5565 19101 5592
rect 19067 5558 19101 5565
rect 19508 5633 19542 5635
rect 19508 5601 19542 5633
rect 19241 5565 19271 5592
rect 19271 5565 19275 5592
rect 19241 5558 19275 5565
rect 19508 5531 19542 5563
rect 19508 5529 19542 5531
rect 17668 5401 17702 5435
rect 17737 5293 17771 5327
rect 19604 5633 19638 5635
rect 19604 5601 19638 5633
rect 19604 5531 19638 5563
rect 19604 5529 19638 5531
rect 19700 5633 19734 5635
rect 19700 5601 19734 5633
rect 19700 5531 19734 5563
rect 19700 5529 19734 5531
rect 20088 6042 20122 6076
rect 21515 6349 21549 6383
rect 22633 6843 22667 6877
rect 22725 6843 22759 6877
rect 22817 6843 22851 6877
rect 23318 6866 23352 6900
rect 25158 6952 25192 6984
rect 25158 6950 25192 6952
rect 25254 7054 25288 7056
rect 25254 7022 25288 7054
rect 25350 7054 25384 7056
rect 25350 7022 25384 7054
rect 25254 6952 25288 6984
rect 25254 6950 25288 6952
rect 25350 6952 25384 6984
rect 25350 6950 25384 6952
rect 27046 7054 27080 7056
rect 27046 7022 27080 7054
rect 22076 6619 22108 6642
rect 22108 6619 22110 6642
rect 22076 6608 22110 6619
rect 22686 6729 22720 6746
rect 22686 6712 22720 6729
rect 23046 6828 23080 6862
rect 23678 6856 23712 6890
rect 23829 6851 23863 6885
rect 23921 6851 23955 6885
rect 24013 6851 24047 6885
rect 23430 6785 23464 6819
rect 22272 6602 22306 6636
rect 21116 6297 21150 6331
rect 22465 6647 22499 6648
rect 22465 6614 22497 6647
rect 22497 6614 22499 6647
rect 23286 6689 23320 6691
rect 23004 6625 23038 6659
rect 23286 6657 23320 6689
rect 23286 6587 23320 6619
rect 23286 6585 23320 6587
rect 21762 6297 21796 6331
rect 21941 6307 21975 6341
rect 22033 6307 22067 6341
rect 22125 6307 22159 6341
rect 22960 6529 22994 6531
rect 22960 6497 22994 6529
rect 22960 6427 22994 6459
rect 22960 6425 22994 6427
rect 22287 6301 22321 6335
rect 22379 6301 22413 6335
rect 22471 6301 22505 6335
rect 23382 6689 23416 6691
rect 23382 6657 23416 6689
rect 23382 6587 23416 6619
rect 23382 6585 23416 6587
rect 23478 6689 23512 6691
rect 23478 6657 23512 6689
rect 24175 6845 24209 6879
rect 24267 6845 24301 6879
rect 24359 6845 24393 6879
rect 23650 6625 23684 6659
rect 23478 6587 23512 6619
rect 23478 6585 23512 6587
rect 23048 6529 23082 6531
rect 23048 6497 23082 6529
rect 23606 6529 23640 6531
rect 23606 6497 23640 6529
rect 23048 6427 23082 6459
rect 23334 6457 23368 6491
rect 23048 6425 23082 6427
rect 23606 6427 23640 6459
rect 23606 6425 23640 6427
rect 23694 6529 23728 6531
rect 23694 6497 23728 6529
rect 23694 6427 23728 6459
rect 23694 6425 23728 6427
rect 22633 6299 22667 6333
rect 22725 6299 22759 6333
rect 22817 6299 22851 6333
rect 21174 6176 21208 6210
rect 21604 6159 21638 6193
rect 21524 6050 21558 6084
rect 21380 5998 21414 6000
rect 21380 5966 21414 5998
rect 21380 5896 21414 5928
rect 21380 5894 21414 5896
rect 21476 5998 21510 6000
rect 21476 5966 21510 5998
rect 21476 5896 21510 5928
rect 21476 5894 21510 5896
rect 21572 5998 21606 6000
rect 21572 5966 21606 5998
rect 21572 5896 21606 5928
rect 21572 5894 21606 5896
rect 19875 5797 19909 5831
rect 19967 5797 20001 5831
rect 20059 5797 20093 5831
rect 20949 5797 20983 5831
rect 21041 5797 21075 5831
rect 21133 5797 21167 5831
rect 21428 5810 21462 5844
rect 19971 5685 20005 5710
rect 19971 5676 20003 5685
rect 20003 5676 20005 5685
rect 21041 5685 21075 5715
rect 21041 5681 21043 5685
rect 21043 5681 21075 5685
rect 21540 5729 21574 5763
rect 19880 5565 19883 5594
rect 19883 5565 19914 5594
rect 19880 5560 19914 5565
rect 20053 5565 20085 5590
rect 20085 5565 20087 5590
rect 20053 5556 20087 5565
rect 20955 5565 20957 5592
rect 20957 5565 20989 5592
rect 20955 5558 20989 5565
rect 21396 5633 21430 5635
rect 21396 5601 21430 5633
rect 21129 5565 21159 5592
rect 21159 5565 21163 5592
rect 21129 5558 21163 5565
rect 21396 5531 21430 5563
rect 21396 5529 21430 5531
rect 19556 5401 19590 5435
rect 19625 5293 19659 5327
rect 21492 5633 21526 5635
rect 21492 5601 21526 5633
rect 21492 5531 21526 5563
rect 21492 5529 21526 5531
rect 21588 5633 21622 5635
rect 21588 5601 21622 5633
rect 21588 5531 21622 5563
rect 21588 5529 21622 5531
rect 21976 6042 22010 6076
rect 23403 6349 23437 6383
rect 24521 6843 24555 6877
rect 24613 6843 24647 6877
rect 24705 6843 24739 6877
rect 25206 6866 25240 6900
rect 27046 6952 27080 6984
rect 27046 6950 27080 6952
rect 27142 7054 27176 7056
rect 27142 7022 27176 7054
rect 27238 7054 27272 7056
rect 27238 7022 27272 7054
rect 27142 6952 27176 6984
rect 27142 6950 27176 6952
rect 27238 6952 27272 6984
rect 27238 6950 27272 6952
rect 28934 7054 28968 7056
rect 28934 7022 28968 7054
rect 23964 6619 23996 6642
rect 23996 6619 23998 6642
rect 23964 6608 23998 6619
rect 24574 6729 24608 6746
rect 24574 6712 24608 6729
rect 24934 6828 24968 6862
rect 25566 6856 25600 6890
rect 25717 6851 25751 6885
rect 25809 6851 25843 6885
rect 25901 6851 25935 6885
rect 25318 6785 25352 6819
rect 24160 6602 24194 6636
rect 23004 6297 23038 6331
rect 24353 6647 24387 6648
rect 24353 6614 24385 6647
rect 24385 6614 24387 6647
rect 25174 6689 25208 6691
rect 24892 6625 24926 6659
rect 25174 6657 25208 6689
rect 25174 6587 25208 6619
rect 25174 6585 25208 6587
rect 23650 6297 23684 6331
rect 23829 6307 23863 6341
rect 23921 6307 23955 6341
rect 24013 6307 24047 6341
rect 24848 6529 24882 6531
rect 24848 6497 24882 6529
rect 24848 6427 24882 6459
rect 24848 6425 24882 6427
rect 24175 6301 24209 6335
rect 24267 6301 24301 6335
rect 24359 6301 24393 6335
rect 25270 6689 25304 6691
rect 25270 6657 25304 6689
rect 25270 6587 25304 6619
rect 25270 6585 25304 6587
rect 25366 6689 25400 6691
rect 25366 6657 25400 6689
rect 26063 6845 26097 6879
rect 26155 6845 26189 6879
rect 26247 6845 26281 6879
rect 25538 6625 25572 6659
rect 25366 6587 25400 6619
rect 25366 6585 25400 6587
rect 24936 6529 24970 6531
rect 24936 6497 24970 6529
rect 25494 6529 25528 6531
rect 25494 6497 25528 6529
rect 24936 6427 24970 6459
rect 25222 6457 25256 6491
rect 24936 6425 24970 6427
rect 25494 6427 25528 6459
rect 25494 6425 25528 6427
rect 25582 6529 25616 6531
rect 25582 6497 25616 6529
rect 25582 6427 25616 6459
rect 25582 6425 25616 6427
rect 24521 6299 24555 6333
rect 24613 6299 24647 6333
rect 24705 6299 24739 6333
rect 23062 6176 23096 6210
rect 23492 6159 23526 6193
rect 23412 6050 23446 6084
rect 23268 5998 23302 6000
rect 23268 5966 23302 5998
rect 23268 5896 23302 5928
rect 23268 5894 23302 5896
rect 23364 5998 23398 6000
rect 23364 5966 23398 5998
rect 23364 5896 23398 5928
rect 23364 5894 23398 5896
rect 23460 5998 23494 6000
rect 23460 5966 23494 5998
rect 23460 5896 23494 5928
rect 23460 5894 23494 5896
rect 21763 5797 21797 5831
rect 21855 5797 21889 5831
rect 21947 5797 21981 5831
rect 22837 5797 22871 5831
rect 22929 5797 22963 5831
rect 23021 5797 23055 5831
rect 23316 5810 23350 5844
rect 21859 5685 21893 5710
rect 21859 5676 21891 5685
rect 21891 5676 21893 5685
rect 22929 5685 22963 5715
rect 22929 5681 22931 5685
rect 22931 5681 22963 5685
rect 23428 5729 23462 5763
rect 21768 5565 21771 5594
rect 21771 5565 21802 5594
rect 21768 5560 21802 5565
rect 21941 5565 21973 5590
rect 21973 5565 21975 5590
rect 21941 5556 21975 5565
rect 22843 5565 22845 5592
rect 22845 5565 22877 5592
rect 22843 5558 22877 5565
rect 23284 5633 23318 5635
rect 23284 5601 23318 5633
rect 23017 5565 23047 5592
rect 23047 5565 23051 5592
rect 23017 5558 23051 5565
rect 23284 5531 23318 5563
rect 23284 5529 23318 5531
rect 21444 5401 21478 5435
rect 21513 5293 21547 5327
rect 23380 5633 23414 5635
rect 23380 5601 23414 5633
rect 23380 5531 23414 5563
rect 23380 5529 23414 5531
rect 23476 5633 23510 5635
rect 23476 5601 23510 5633
rect 23476 5531 23510 5563
rect 23476 5529 23510 5531
rect 23864 6042 23898 6076
rect 25291 6349 25325 6383
rect 26409 6843 26443 6877
rect 26501 6843 26535 6877
rect 26593 6843 26627 6877
rect 27094 6866 27128 6900
rect 28934 6952 28968 6984
rect 28934 6950 28968 6952
rect 29030 7054 29064 7056
rect 29030 7022 29064 7054
rect 29126 7054 29160 7056
rect 29126 7022 29160 7054
rect 29030 6952 29064 6984
rect 29030 6950 29064 6952
rect 29126 6952 29160 6984
rect 29126 6950 29160 6952
rect 30822 7054 30856 7056
rect 30822 7022 30856 7054
rect 25852 6619 25884 6642
rect 25884 6619 25886 6642
rect 25852 6608 25886 6619
rect 26462 6729 26496 6746
rect 26462 6712 26496 6729
rect 26822 6828 26856 6862
rect 27454 6856 27488 6890
rect 27605 6851 27639 6885
rect 27697 6851 27731 6885
rect 27789 6851 27823 6885
rect 27206 6785 27240 6819
rect 26048 6602 26082 6636
rect 24892 6297 24926 6331
rect 26241 6647 26275 6648
rect 26241 6614 26273 6647
rect 26273 6614 26275 6647
rect 27062 6689 27096 6691
rect 26780 6625 26814 6659
rect 27062 6657 27096 6689
rect 27062 6587 27096 6619
rect 27062 6585 27096 6587
rect 25538 6297 25572 6331
rect 25717 6307 25751 6341
rect 25809 6307 25843 6341
rect 25901 6307 25935 6341
rect 26736 6529 26770 6531
rect 26736 6497 26770 6529
rect 26736 6427 26770 6459
rect 26736 6425 26770 6427
rect 26063 6301 26097 6335
rect 26155 6301 26189 6335
rect 26247 6301 26281 6335
rect 27158 6689 27192 6691
rect 27158 6657 27192 6689
rect 27158 6587 27192 6619
rect 27158 6585 27192 6587
rect 27254 6689 27288 6691
rect 27254 6657 27288 6689
rect 27951 6845 27985 6879
rect 28043 6845 28077 6879
rect 28135 6845 28169 6879
rect 27426 6625 27460 6659
rect 27254 6587 27288 6619
rect 27254 6585 27288 6587
rect 26824 6529 26858 6531
rect 26824 6497 26858 6529
rect 27382 6529 27416 6531
rect 27382 6497 27416 6529
rect 26824 6427 26858 6459
rect 27110 6457 27144 6491
rect 26824 6425 26858 6427
rect 27382 6427 27416 6459
rect 27382 6425 27416 6427
rect 27470 6529 27504 6531
rect 27470 6497 27504 6529
rect 27470 6427 27504 6459
rect 27470 6425 27504 6427
rect 26409 6299 26443 6333
rect 26501 6299 26535 6333
rect 26593 6299 26627 6333
rect 24950 6176 24984 6210
rect 25380 6159 25414 6193
rect 25300 6050 25334 6084
rect 25156 5998 25190 6000
rect 25156 5966 25190 5998
rect 25156 5896 25190 5928
rect 25156 5894 25190 5896
rect 25252 5998 25286 6000
rect 25252 5966 25286 5998
rect 25252 5896 25286 5928
rect 25252 5894 25286 5896
rect 25348 5998 25382 6000
rect 25348 5966 25382 5998
rect 25348 5896 25382 5928
rect 25348 5894 25382 5896
rect 23651 5797 23685 5831
rect 23743 5797 23777 5831
rect 23835 5797 23869 5831
rect 24725 5797 24759 5831
rect 24817 5797 24851 5831
rect 24909 5797 24943 5831
rect 25204 5810 25238 5844
rect 23747 5685 23781 5710
rect 23747 5676 23779 5685
rect 23779 5676 23781 5685
rect 24817 5685 24851 5715
rect 24817 5681 24819 5685
rect 24819 5681 24851 5685
rect 25316 5729 25350 5763
rect 23656 5565 23659 5594
rect 23659 5565 23690 5594
rect 23656 5560 23690 5565
rect 23829 5565 23861 5590
rect 23861 5565 23863 5590
rect 23829 5556 23863 5565
rect 24731 5565 24733 5592
rect 24733 5565 24765 5592
rect 24731 5558 24765 5565
rect 25172 5633 25206 5635
rect 25172 5601 25206 5633
rect 24905 5565 24935 5592
rect 24935 5565 24939 5592
rect 24905 5558 24939 5565
rect 25172 5531 25206 5563
rect 25172 5529 25206 5531
rect 23332 5401 23366 5435
rect 23401 5293 23435 5327
rect 25268 5633 25302 5635
rect 25268 5601 25302 5633
rect 25268 5531 25302 5563
rect 25268 5529 25302 5531
rect 25364 5633 25398 5635
rect 25364 5601 25398 5633
rect 25364 5531 25398 5563
rect 25364 5529 25398 5531
rect 25752 6042 25786 6076
rect 27179 6349 27213 6383
rect 28297 6843 28331 6877
rect 28389 6843 28423 6877
rect 28481 6843 28515 6877
rect 28982 6866 29016 6900
rect 30822 6952 30856 6984
rect 30822 6950 30856 6952
rect 30918 7054 30952 7056
rect 30918 7022 30952 7054
rect 31014 7054 31048 7056
rect 31014 7022 31048 7054
rect 30918 6952 30952 6984
rect 30918 6950 30952 6952
rect 31014 6952 31048 6984
rect 31014 6950 31048 6952
rect 32710 7054 32744 7056
rect 32710 7022 32744 7054
rect 27740 6619 27772 6642
rect 27772 6619 27774 6642
rect 27740 6608 27774 6619
rect 28350 6729 28384 6746
rect 28350 6712 28384 6729
rect 28710 6828 28744 6862
rect 29342 6856 29376 6890
rect 29493 6851 29527 6885
rect 29585 6851 29619 6885
rect 29677 6851 29711 6885
rect 29094 6785 29128 6819
rect 27936 6602 27970 6636
rect 26780 6297 26814 6331
rect 28129 6647 28163 6648
rect 28129 6614 28161 6647
rect 28161 6614 28163 6647
rect 28950 6689 28984 6691
rect 28668 6625 28702 6659
rect 28950 6657 28984 6689
rect 28950 6587 28984 6619
rect 28950 6585 28984 6587
rect 27426 6297 27460 6331
rect 27605 6307 27639 6341
rect 27697 6307 27731 6341
rect 27789 6307 27823 6341
rect 28624 6529 28658 6531
rect 28624 6497 28658 6529
rect 28624 6427 28658 6459
rect 28624 6425 28658 6427
rect 27951 6301 27985 6335
rect 28043 6301 28077 6335
rect 28135 6301 28169 6335
rect 29046 6689 29080 6691
rect 29046 6657 29080 6689
rect 29046 6587 29080 6619
rect 29046 6585 29080 6587
rect 29142 6689 29176 6691
rect 29142 6657 29176 6689
rect 29839 6845 29873 6879
rect 29931 6845 29965 6879
rect 30023 6845 30057 6879
rect 29314 6625 29348 6659
rect 29142 6587 29176 6619
rect 29142 6585 29176 6587
rect 28712 6529 28746 6531
rect 28712 6497 28746 6529
rect 29270 6529 29304 6531
rect 29270 6497 29304 6529
rect 28712 6427 28746 6459
rect 28998 6457 29032 6491
rect 28712 6425 28746 6427
rect 29270 6427 29304 6459
rect 29270 6425 29304 6427
rect 29358 6529 29392 6531
rect 29358 6497 29392 6529
rect 29358 6427 29392 6459
rect 29358 6425 29392 6427
rect 28297 6299 28331 6333
rect 28389 6299 28423 6333
rect 28481 6299 28515 6333
rect 26838 6176 26872 6210
rect 27268 6159 27302 6193
rect 27188 6050 27222 6084
rect 27044 5998 27078 6000
rect 27044 5966 27078 5998
rect 27044 5896 27078 5928
rect 27044 5894 27078 5896
rect 27140 5998 27174 6000
rect 27140 5966 27174 5998
rect 27140 5896 27174 5928
rect 27140 5894 27174 5896
rect 27236 5998 27270 6000
rect 27236 5966 27270 5998
rect 27236 5896 27270 5928
rect 27236 5894 27270 5896
rect 25539 5797 25573 5831
rect 25631 5797 25665 5831
rect 25723 5797 25757 5831
rect 26613 5797 26647 5831
rect 26705 5797 26739 5831
rect 26797 5797 26831 5831
rect 27092 5810 27126 5844
rect 25635 5685 25669 5710
rect 25635 5676 25667 5685
rect 25667 5676 25669 5685
rect 26705 5685 26739 5715
rect 26705 5681 26707 5685
rect 26707 5681 26739 5685
rect 27204 5729 27238 5763
rect 25544 5565 25547 5594
rect 25547 5565 25578 5594
rect 25544 5560 25578 5565
rect 25717 5565 25749 5590
rect 25749 5565 25751 5590
rect 25717 5556 25751 5565
rect 26619 5565 26621 5592
rect 26621 5565 26653 5592
rect 26619 5558 26653 5565
rect 27060 5633 27094 5635
rect 27060 5601 27094 5633
rect 26793 5565 26823 5592
rect 26823 5565 26827 5592
rect 26793 5558 26827 5565
rect 27060 5531 27094 5563
rect 27060 5529 27094 5531
rect 25220 5401 25254 5435
rect 25289 5293 25323 5327
rect 27156 5633 27190 5635
rect 27156 5601 27190 5633
rect 27156 5531 27190 5563
rect 27156 5529 27190 5531
rect 27252 5633 27286 5635
rect 27252 5601 27286 5633
rect 27252 5531 27286 5563
rect 27252 5529 27286 5531
rect 27640 6042 27674 6076
rect 29067 6349 29101 6383
rect 30185 6843 30219 6877
rect 30277 6843 30311 6877
rect 30369 6843 30403 6877
rect 30870 6866 30904 6900
rect 32710 6952 32744 6984
rect 32710 6950 32744 6952
rect 32806 7054 32840 7056
rect 32806 7022 32840 7054
rect 32902 7054 32936 7056
rect 32902 7022 32936 7054
rect 32806 6952 32840 6984
rect 32806 6950 32840 6952
rect 32902 6952 32936 6984
rect 32902 6950 32936 6952
rect 34598 7054 34632 7056
rect 34598 7022 34632 7054
rect 29628 6619 29660 6642
rect 29660 6619 29662 6642
rect 29628 6608 29662 6619
rect 30238 6729 30272 6746
rect 30238 6712 30272 6729
rect 30598 6828 30632 6862
rect 31230 6856 31264 6890
rect 31381 6851 31415 6885
rect 31473 6851 31507 6885
rect 31565 6851 31599 6885
rect 30982 6785 31016 6819
rect 29824 6602 29858 6636
rect 28668 6297 28702 6331
rect 30017 6647 30051 6648
rect 30017 6614 30049 6647
rect 30049 6614 30051 6647
rect 30838 6689 30872 6691
rect 30556 6625 30590 6659
rect 30838 6657 30872 6689
rect 30838 6587 30872 6619
rect 30838 6585 30872 6587
rect 29314 6297 29348 6331
rect 29493 6307 29527 6341
rect 29585 6307 29619 6341
rect 29677 6307 29711 6341
rect 30512 6529 30546 6531
rect 30512 6497 30546 6529
rect 30512 6427 30546 6459
rect 30512 6425 30546 6427
rect 29839 6301 29873 6335
rect 29931 6301 29965 6335
rect 30023 6301 30057 6335
rect 30934 6689 30968 6691
rect 30934 6657 30968 6689
rect 30934 6587 30968 6619
rect 30934 6585 30968 6587
rect 31030 6689 31064 6691
rect 31030 6657 31064 6689
rect 31727 6845 31761 6879
rect 31819 6845 31853 6879
rect 31911 6845 31945 6879
rect 31202 6625 31236 6659
rect 31030 6587 31064 6619
rect 31030 6585 31064 6587
rect 30600 6529 30634 6531
rect 30600 6497 30634 6529
rect 31158 6529 31192 6531
rect 31158 6497 31192 6529
rect 30600 6427 30634 6459
rect 30886 6457 30920 6491
rect 30600 6425 30634 6427
rect 31158 6427 31192 6459
rect 31158 6425 31192 6427
rect 31246 6529 31280 6531
rect 31246 6497 31280 6529
rect 31246 6427 31280 6459
rect 31246 6425 31280 6427
rect 30185 6299 30219 6333
rect 30277 6299 30311 6333
rect 30369 6299 30403 6333
rect 28726 6176 28760 6210
rect 29156 6159 29190 6193
rect 29076 6050 29110 6084
rect 28932 5998 28966 6000
rect 28932 5966 28966 5998
rect 28932 5896 28966 5928
rect 28932 5894 28966 5896
rect 29028 5998 29062 6000
rect 29028 5966 29062 5998
rect 29028 5896 29062 5928
rect 29028 5894 29062 5896
rect 29124 5998 29158 6000
rect 29124 5966 29158 5998
rect 29124 5896 29158 5928
rect 29124 5894 29158 5896
rect 27427 5797 27461 5831
rect 27519 5797 27553 5831
rect 27611 5797 27645 5831
rect 28501 5797 28535 5831
rect 28593 5797 28627 5831
rect 28685 5797 28719 5831
rect 28980 5810 29014 5844
rect 27523 5685 27557 5710
rect 27523 5676 27555 5685
rect 27555 5676 27557 5685
rect 28593 5685 28627 5715
rect 28593 5681 28595 5685
rect 28595 5681 28627 5685
rect 29092 5729 29126 5763
rect 27432 5565 27435 5594
rect 27435 5565 27466 5594
rect 27432 5560 27466 5565
rect 27605 5565 27637 5590
rect 27637 5565 27639 5590
rect 27605 5556 27639 5565
rect 28507 5565 28509 5592
rect 28509 5565 28541 5592
rect 28507 5558 28541 5565
rect 28948 5633 28982 5635
rect 28948 5601 28982 5633
rect 28681 5565 28711 5592
rect 28711 5565 28715 5592
rect 28681 5558 28715 5565
rect 28948 5531 28982 5563
rect 28948 5529 28982 5531
rect 27108 5401 27142 5435
rect 27177 5293 27211 5327
rect 29044 5633 29078 5635
rect 29044 5601 29078 5633
rect 29044 5531 29078 5563
rect 29044 5529 29078 5531
rect 29140 5633 29174 5635
rect 29140 5601 29174 5633
rect 29140 5531 29174 5563
rect 29140 5529 29174 5531
rect 29528 6042 29562 6076
rect 30955 6349 30989 6383
rect 32073 6843 32107 6877
rect 32165 6843 32199 6877
rect 32257 6843 32291 6877
rect 32758 6866 32792 6900
rect 34598 6952 34632 6984
rect 34598 6950 34632 6952
rect 34694 7054 34728 7056
rect 34694 7022 34728 7054
rect 34790 7054 34824 7056
rect 34790 7022 34824 7054
rect 34694 6952 34728 6984
rect 34694 6950 34728 6952
rect 34790 6952 34824 6984
rect 34790 6950 34824 6952
rect 36486 7054 36520 7056
rect 36486 7022 36520 7054
rect 31516 6619 31548 6642
rect 31548 6619 31550 6642
rect 31516 6608 31550 6619
rect 32126 6729 32160 6746
rect 32126 6712 32160 6729
rect 32486 6828 32520 6862
rect 33118 6856 33152 6890
rect 33269 6851 33303 6885
rect 33361 6851 33395 6885
rect 33453 6851 33487 6885
rect 32870 6785 32904 6819
rect 31712 6602 31746 6636
rect 30556 6297 30590 6331
rect 31905 6647 31939 6648
rect 31905 6614 31937 6647
rect 31937 6614 31939 6647
rect 32726 6689 32760 6691
rect 32444 6625 32478 6659
rect 32726 6657 32760 6689
rect 32726 6587 32760 6619
rect 32726 6585 32760 6587
rect 31202 6297 31236 6331
rect 31381 6307 31415 6341
rect 31473 6307 31507 6341
rect 31565 6307 31599 6341
rect 32400 6529 32434 6531
rect 32400 6497 32434 6529
rect 32400 6427 32434 6459
rect 32400 6425 32434 6427
rect 31727 6301 31761 6335
rect 31819 6301 31853 6335
rect 31911 6301 31945 6335
rect 32822 6689 32856 6691
rect 32822 6657 32856 6689
rect 32822 6587 32856 6619
rect 32822 6585 32856 6587
rect 32918 6689 32952 6691
rect 32918 6657 32952 6689
rect 33615 6845 33649 6879
rect 33707 6845 33741 6879
rect 33799 6845 33833 6879
rect 33090 6625 33124 6659
rect 32918 6587 32952 6619
rect 32918 6585 32952 6587
rect 32488 6529 32522 6531
rect 32488 6497 32522 6529
rect 33046 6529 33080 6531
rect 33046 6497 33080 6529
rect 32488 6427 32522 6459
rect 32774 6457 32808 6491
rect 32488 6425 32522 6427
rect 33046 6427 33080 6459
rect 33046 6425 33080 6427
rect 33134 6529 33168 6531
rect 33134 6497 33168 6529
rect 33134 6427 33168 6459
rect 33134 6425 33168 6427
rect 32073 6299 32107 6333
rect 32165 6299 32199 6333
rect 32257 6299 32291 6333
rect 30614 6176 30648 6210
rect 31044 6159 31078 6193
rect 30964 6050 30998 6084
rect 30820 5998 30854 6000
rect 30820 5966 30854 5998
rect 30820 5896 30854 5928
rect 30820 5894 30854 5896
rect 30916 5998 30950 6000
rect 30916 5966 30950 5998
rect 30916 5896 30950 5928
rect 30916 5894 30950 5896
rect 31012 5998 31046 6000
rect 31012 5966 31046 5998
rect 31012 5896 31046 5928
rect 31012 5894 31046 5896
rect 29315 5797 29349 5831
rect 29407 5797 29441 5831
rect 29499 5797 29533 5831
rect 30389 5797 30423 5831
rect 30481 5797 30515 5831
rect 30573 5797 30607 5831
rect 30868 5810 30902 5844
rect 29411 5685 29445 5710
rect 29411 5676 29443 5685
rect 29443 5676 29445 5685
rect 30481 5685 30515 5715
rect 30481 5681 30483 5685
rect 30483 5681 30515 5685
rect 30980 5729 31014 5763
rect 29320 5565 29323 5594
rect 29323 5565 29354 5594
rect 29320 5560 29354 5565
rect 29493 5565 29525 5590
rect 29525 5565 29527 5590
rect 29493 5556 29527 5565
rect 30395 5565 30397 5592
rect 30397 5565 30429 5592
rect 30395 5558 30429 5565
rect 30836 5633 30870 5635
rect 30836 5601 30870 5633
rect 30569 5565 30599 5592
rect 30599 5565 30603 5592
rect 30569 5558 30603 5565
rect 30836 5531 30870 5563
rect 30836 5529 30870 5531
rect 28996 5401 29030 5435
rect 29065 5293 29099 5327
rect 30932 5633 30966 5635
rect 30932 5601 30966 5633
rect 30932 5531 30966 5563
rect 30932 5529 30966 5531
rect 31028 5633 31062 5635
rect 31028 5601 31062 5633
rect 31028 5531 31062 5563
rect 31028 5529 31062 5531
rect 31416 6042 31450 6076
rect 32843 6349 32877 6383
rect 33961 6843 33995 6877
rect 34053 6843 34087 6877
rect 34145 6843 34179 6877
rect 34646 6866 34680 6900
rect 36486 6952 36520 6984
rect 36486 6950 36520 6952
rect 36582 7054 36616 7056
rect 36582 7022 36616 7054
rect 36678 7054 36712 7056
rect 36678 7022 36712 7054
rect 36582 6952 36616 6984
rect 36582 6950 36616 6952
rect 36678 6952 36712 6984
rect 36678 6950 36712 6952
rect 38374 7054 38408 7056
rect 38374 7022 38408 7054
rect 33404 6619 33436 6642
rect 33436 6619 33438 6642
rect 33404 6608 33438 6619
rect 34014 6729 34048 6746
rect 34014 6712 34048 6729
rect 34374 6828 34408 6862
rect 35006 6856 35040 6890
rect 35157 6851 35191 6885
rect 35249 6851 35283 6885
rect 35341 6851 35375 6885
rect 34758 6785 34792 6819
rect 33600 6602 33634 6636
rect 32444 6297 32478 6331
rect 33793 6647 33827 6648
rect 33793 6614 33825 6647
rect 33825 6614 33827 6647
rect 34614 6689 34648 6691
rect 34332 6625 34366 6659
rect 34614 6657 34648 6689
rect 34614 6587 34648 6619
rect 34614 6585 34648 6587
rect 33090 6297 33124 6331
rect 33269 6307 33303 6341
rect 33361 6307 33395 6341
rect 33453 6307 33487 6341
rect 34288 6529 34322 6531
rect 34288 6497 34322 6529
rect 34288 6427 34322 6459
rect 34288 6425 34322 6427
rect 33615 6301 33649 6335
rect 33707 6301 33741 6335
rect 33799 6301 33833 6335
rect 34710 6689 34744 6691
rect 34710 6657 34744 6689
rect 34710 6587 34744 6619
rect 34710 6585 34744 6587
rect 34806 6689 34840 6691
rect 34806 6657 34840 6689
rect 35503 6845 35537 6879
rect 35595 6845 35629 6879
rect 35687 6845 35721 6879
rect 34978 6625 35012 6659
rect 34806 6587 34840 6619
rect 34806 6585 34840 6587
rect 34376 6529 34410 6531
rect 34376 6497 34410 6529
rect 34934 6529 34968 6531
rect 34934 6497 34968 6529
rect 34376 6427 34410 6459
rect 34662 6457 34696 6491
rect 34376 6425 34410 6427
rect 34934 6427 34968 6459
rect 34934 6425 34968 6427
rect 35022 6529 35056 6531
rect 35022 6497 35056 6529
rect 35022 6427 35056 6459
rect 35022 6425 35056 6427
rect 33961 6299 33995 6333
rect 34053 6299 34087 6333
rect 34145 6299 34179 6333
rect 32502 6176 32536 6210
rect 32932 6159 32966 6193
rect 32852 6050 32886 6084
rect 32708 5998 32742 6000
rect 32708 5966 32742 5998
rect 32708 5896 32742 5928
rect 32708 5894 32742 5896
rect 32804 5998 32838 6000
rect 32804 5966 32838 5998
rect 32804 5896 32838 5928
rect 32804 5894 32838 5896
rect 32900 5998 32934 6000
rect 32900 5966 32934 5998
rect 32900 5896 32934 5928
rect 32900 5894 32934 5896
rect 31203 5797 31237 5831
rect 31295 5797 31329 5831
rect 31387 5797 31421 5831
rect 32277 5797 32311 5831
rect 32369 5797 32403 5831
rect 32461 5797 32495 5831
rect 32756 5810 32790 5844
rect 31299 5685 31333 5710
rect 31299 5676 31331 5685
rect 31331 5676 31333 5685
rect 32369 5685 32403 5715
rect 32369 5681 32371 5685
rect 32371 5681 32403 5685
rect 32868 5729 32902 5763
rect 31208 5565 31211 5594
rect 31211 5565 31242 5594
rect 31208 5560 31242 5565
rect 31381 5565 31413 5590
rect 31413 5565 31415 5590
rect 31381 5556 31415 5565
rect 32283 5565 32285 5592
rect 32285 5565 32317 5592
rect 32283 5558 32317 5565
rect 32724 5633 32758 5635
rect 32724 5601 32758 5633
rect 32457 5565 32487 5592
rect 32487 5565 32491 5592
rect 32457 5558 32491 5565
rect 32724 5531 32758 5563
rect 32724 5529 32758 5531
rect 30884 5401 30918 5435
rect 30953 5293 30987 5327
rect 32820 5633 32854 5635
rect 32820 5601 32854 5633
rect 32820 5531 32854 5563
rect 32820 5529 32854 5531
rect 32916 5633 32950 5635
rect 32916 5601 32950 5633
rect 32916 5531 32950 5563
rect 32916 5529 32950 5531
rect 33304 6042 33338 6076
rect 34731 6349 34765 6383
rect 35849 6843 35883 6877
rect 35941 6843 35975 6877
rect 36033 6843 36067 6877
rect 36534 6866 36568 6900
rect 38374 6952 38408 6984
rect 38374 6950 38408 6952
rect 38470 7054 38504 7056
rect 38470 7022 38504 7054
rect 38566 7054 38600 7056
rect 38566 7022 38600 7054
rect 38470 6952 38504 6984
rect 38470 6950 38504 6952
rect 38566 6952 38600 6984
rect 38566 6950 38600 6952
rect 40262 7054 40296 7056
rect 40262 7022 40296 7054
rect 35292 6619 35324 6642
rect 35324 6619 35326 6642
rect 35292 6608 35326 6619
rect 35902 6729 35936 6746
rect 35902 6712 35936 6729
rect 36262 6828 36296 6862
rect 36894 6856 36928 6890
rect 37045 6851 37079 6885
rect 37137 6851 37171 6885
rect 37229 6851 37263 6885
rect 36646 6785 36680 6819
rect 35488 6602 35522 6636
rect 34332 6297 34366 6331
rect 35681 6647 35715 6648
rect 35681 6614 35713 6647
rect 35713 6614 35715 6647
rect 36502 6689 36536 6691
rect 36220 6625 36254 6659
rect 36502 6657 36536 6689
rect 36502 6587 36536 6619
rect 36502 6585 36536 6587
rect 34978 6297 35012 6331
rect 35157 6307 35191 6341
rect 35249 6307 35283 6341
rect 35341 6307 35375 6341
rect 36176 6529 36210 6531
rect 36176 6497 36210 6529
rect 36176 6427 36210 6459
rect 36176 6425 36210 6427
rect 35503 6301 35537 6335
rect 35595 6301 35629 6335
rect 35687 6301 35721 6335
rect 36598 6689 36632 6691
rect 36598 6657 36632 6689
rect 36598 6587 36632 6619
rect 36598 6585 36632 6587
rect 36694 6689 36728 6691
rect 36694 6657 36728 6689
rect 37391 6845 37425 6879
rect 37483 6845 37517 6879
rect 37575 6845 37609 6879
rect 36866 6625 36900 6659
rect 36694 6587 36728 6619
rect 36694 6585 36728 6587
rect 36264 6529 36298 6531
rect 36264 6497 36298 6529
rect 36822 6529 36856 6531
rect 36822 6497 36856 6529
rect 36264 6427 36298 6459
rect 36550 6457 36584 6491
rect 36264 6425 36298 6427
rect 36822 6427 36856 6459
rect 36822 6425 36856 6427
rect 36910 6529 36944 6531
rect 36910 6497 36944 6529
rect 36910 6427 36944 6459
rect 36910 6425 36944 6427
rect 35849 6299 35883 6333
rect 35941 6299 35975 6333
rect 36033 6299 36067 6333
rect 34390 6176 34424 6210
rect 34820 6159 34854 6193
rect 34740 6050 34774 6084
rect 34596 5998 34630 6000
rect 34596 5966 34630 5998
rect 34596 5896 34630 5928
rect 34596 5894 34630 5896
rect 34692 5998 34726 6000
rect 34692 5966 34726 5998
rect 34692 5896 34726 5928
rect 34692 5894 34726 5896
rect 34788 5998 34822 6000
rect 34788 5966 34822 5998
rect 34788 5896 34822 5928
rect 34788 5894 34822 5896
rect 33091 5797 33125 5831
rect 33183 5797 33217 5831
rect 33275 5797 33309 5831
rect 34165 5797 34199 5831
rect 34257 5797 34291 5831
rect 34349 5797 34383 5831
rect 34644 5810 34678 5844
rect 33187 5685 33221 5710
rect 33187 5676 33219 5685
rect 33219 5676 33221 5685
rect 34257 5685 34291 5715
rect 34257 5681 34259 5685
rect 34259 5681 34291 5685
rect 34756 5729 34790 5763
rect 33096 5565 33099 5594
rect 33099 5565 33130 5594
rect 33096 5560 33130 5565
rect 33269 5565 33301 5590
rect 33301 5565 33303 5590
rect 33269 5556 33303 5565
rect 34171 5565 34173 5592
rect 34173 5565 34205 5592
rect 34171 5558 34205 5565
rect 34612 5633 34646 5635
rect 34612 5601 34646 5633
rect 34345 5565 34375 5592
rect 34375 5565 34379 5592
rect 34345 5558 34379 5565
rect 34612 5531 34646 5563
rect 34612 5529 34646 5531
rect 32772 5401 32806 5435
rect 32841 5293 32875 5327
rect 34708 5633 34742 5635
rect 34708 5601 34742 5633
rect 34708 5531 34742 5563
rect 34708 5529 34742 5531
rect 34804 5633 34838 5635
rect 34804 5601 34838 5633
rect 34804 5531 34838 5563
rect 34804 5529 34838 5531
rect 35192 6042 35226 6076
rect 36619 6349 36653 6383
rect 37737 6843 37771 6877
rect 37829 6843 37863 6877
rect 37921 6843 37955 6877
rect 38422 6866 38456 6900
rect 40262 6952 40296 6984
rect 40262 6950 40296 6952
rect 40358 7054 40392 7056
rect 40358 7022 40392 7054
rect 40454 7054 40488 7056
rect 40454 7022 40488 7054
rect 40358 6952 40392 6984
rect 40358 6950 40392 6952
rect 40454 6952 40488 6984
rect 40454 6950 40488 6952
rect 42150 7054 42184 7056
rect 42150 7022 42184 7054
rect 37180 6619 37212 6642
rect 37212 6619 37214 6642
rect 37180 6608 37214 6619
rect 37790 6729 37824 6746
rect 37790 6712 37824 6729
rect 38150 6828 38184 6862
rect 38782 6856 38816 6890
rect 38933 6851 38967 6885
rect 39025 6851 39059 6885
rect 39117 6851 39151 6885
rect 38534 6785 38568 6819
rect 37376 6602 37410 6636
rect 36220 6297 36254 6331
rect 37569 6647 37603 6648
rect 37569 6614 37601 6647
rect 37601 6614 37603 6647
rect 38390 6689 38424 6691
rect 38108 6625 38142 6659
rect 38390 6657 38424 6689
rect 38390 6587 38424 6619
rect 38390 6585 38424 6587
rect 36866 6297 36900 6331
rect 37045 6307 37079 6341
rect 37137 6307 37171 6341
rect 37229 6307 37263 6341
rect 38064 6529 38098 6531
rect 38064 6497 38098 6529
rect 38064 6427 38098 6459
rect 38064 6425 38098 6427
rect 37391 6301 37425 6335
rect 37483 6301 37517 6335
rect 37575 6301 37609 6335
rect 38486 6689 38520 6691
rect 38486 6657 38520 6689
rect 38486 6587 38520 6619
rect 38486 6585 38520 6587
rect 38582 6689 38616 6691
rect 38582 6657 38616 6689
rect 39279 6845 39313 6879
rect 39371 6845 39405 6879
rect 39463 6845 39497 6879
rect 38754 6625 38788 6659
rect 38582 6587 38616 6619
rect 38582 6585 38616 6587
rect 38152 6529 38186 6531
rect 38152 6497 38186 6529
rect 38710 6529 38744 6531
rect 38710 6497 38744 6529
rect 38152 6427 38186 6459
rect 38438 6457 38472 6491
rect 38152 6425 38186 6427
rect 38710 6427 38744 6459
rect 38710 6425 38744 6427
rect 38798 6529 38832 6531
rect 38798 6497 38832 6529
rect 38798 6427 38832 6459
rect 38798 6425 38832 6427
rect 37737 6299 37771 6333
rect 37829 6299 37863 6333
rect 37921 6299 37955 6333
rect 36278 6176 36312 6210
rect 36708 6159 36742 6193
rect 36628 6050 36662 6084
rect 36484 5998 36518 6000
rect 36484 5966 36518 5998
rect 36484 5896 36518 5928
rect 36484 5894 36518 5896
rect 36580 5998 36614 6000
rect 36580 5966 36614 5998
rect 36580 5896 36614 5928
rect 36580 5894 36614 5896
rect 36676 5998 36710 6000
rect 36676 5966 36710 5998
rect 36676 5896 36710 5928
rect 36676 5894 36710 5896
rect 34979 5797 35013 5831
rect 35071 5797 35105 5831
rect 35163 5797 35197 5831
rect 36053 5797 36087 5831
rect 36145 5797 36179 5831
rect 36237 5797 36271 5831
rect 36532 5810 36566 5844
rect 35075 5685 35109 5710
rect 35075 5676 35107 5685
rect 35107 5676 35109 5685
rect 36145 5685 36179 5715
rect 36145 5681 36147 5685
rect 36147 5681 36179 5685
rect 36644 5729 36678 5763
rect 34984 5565 34987 5594
rect 34987 5565 35018 5594
rect 34984 5560 35018 5565
rect 35157 5565 35189 5590
rect 35189 5565 35191 5590
rect 35157 5556 35191 5565
rect 36059 5565 36061 5592
rect 36061 5565 36093 5592
rect 36059 5558 36093 5565
rect 36500 5633 36534 5635
rect 36500 5601 36534 5633
rect 36233 5565 36263 5592
rect 36263 5565 36267 5592
rect 36233 5558 36267 5565
rect 36500 5531 36534 5563
rect 36500 5529 36534 5531
rect 34660 5401 34694 5435
rect 34729 5293 34763 5327
rect 36596 5633 36630 5635
rect 36596 5601 36630 5633
rect 36596 5531 36630 5563
rect 36596 5529 36630 5531
rect 36692 5633 36726 5635
rect 36692 5601 36726 5633
rect 36692 5531 36726 5563
rect 36692 5529 36726 5531
rect 37080 6042 37114 6076
rect 38507 6349 38541 6383
rect 39625 6843 39659 6877
rect 39717 6843 39751 6877
rect 39809 6843 39843 6877
rect 40310 6866 40344 6900
rect 42150 6952 42184 6984
rect 42150 6950 42184 6952
rect 42246 7054 42280 7056
rect 42246 7022 42280 7054
rect 42342 7054 42376 7056
rect 42342 7022 42376 7054
rect 42246 6952 42280 6984
rect 42246 6950 42280 6952
rect 42342 6952 42376 6984
rect 42342 6950 42376 6952
rect 44038 7054 44072 7056
rect 44038 7022 44072 7054
rect 39068 6619 39100 6642
rect 39100 6619 39102 6642
rect 39068 6608 39102 6619
rect 39678 6729 39712 6746
rect 39678 6712 39712 6729
rect 40038 6828 40072 6862
rect 40670 6856 40704 6890
rect 40821 6851 40855 6885
rect 40913 6851 40947 6885
rect 41005 6851 41039 6885
rect 40422 6785 40456 6819
rect 39264 6602 39298 6636
rect 38108 6297 38142 6331
rect 39457 6647 39491 6648
rect 39457 6614 39489 6647
rect 39489 6614 39491 6647
rect 40278 6689 40312 6691
rect 39996 6625 40030 6659
rect 40278 6657 40312 6689
rect 40278 6587 40312 6619
rect 40278 6585 40312 6587
rect 38754 6297 38788 6331
rect 38933 6307 38967 6341
rect 39025 6307 39059 6341
rect 39117 6307 39151 6341
rect 39952 6529 39986 6531
rect 39952 6497 39986 6529
rect 39952 6427 39986 6459
rect 39952 6425 39986 6427
rect 39279 6301 39313 6335
rect 39371 6301 39405 6335
rect 39463 6301 39497 6335
rect 40374 6689 40408 6691
rect 40374 6657 40408 6689
rect 40374 6587 40408 6619
rect 40374 6585 40408 6587
rect 40470 6689 40504 6691
rect 40470 6657 40504 6689
rect 41167 6845 41201 6879
rect 41259 6845 41293 6879
rect 41351 6845 41385 6879
rect 40642 6625 40676 6659
rect 40470 6587 40504 6619
rect 40470 6585 40504 6587
rect 40040 6529 40074 6531
rect 40040 6497 40074 6529
rect 40598 6529 40632 6531
rect 40598 6497 40632 6529
rect 40040 6427 40074 6459
rect 40326 6457 40360 6491
rect 40040 6425 40074 6427
rect 40598 6427 40632 6459
rect 40598 6425 40632 6427
rect 40686 6529 40720 6531
rect 40686 6497 40720 6529
rect 40686 6427 40720 6459
rect 40686 6425 40720 6427
rect 39625 6299 39659 6333
rect 39717 6299 39751 6333
rect 39809 6299 39843 6333
rect 38166 6176 38200 6210
rect 38596 6159 38630 6193
rect 38516 6050 38550 6084
rect 38372 5998 38406 6000
rect 38372 5966 38406 5998
rect 38372 5896 38406 5928
rect 38372 5894 38406 5896
rect 38468 5998 38502 6000
rect 38468 5966 38502 5998
rect 38468 5896 38502 5928
rect 38468 5894 38502 5896
rect 38564 5998 38598 6000
rect 38564 5966 38598 5998
rect 38564 5896 38598 5928
rect 38564 5894 38598 5896
rect 36867 5797 36901 5831
rect 36959 5797 36993 5831
rect 37051 5797 37085 5831
rect 37941 5797 37975 5831
rect 38033 5797 38067 5831
rect 38125 5797 38159 5831
rect 38420 5810 38454 5844
rect 36963 5685 36997 5710
rect 36963 5676 36995 5685
rect 36995 5676 36997 5685
rect 38033 5685 38067 5715
rect 38033 5681 38035 5685
rect 38035 5681 38067 5685
rect 38532 5729 38566 5763
rect 36872 5565 36875 5594
rect 36875 5565 36906 5594
rect 36872 5560 36906 5565
rect 37045 5565 37077 5590
rect 37077 5565 37079 5590
rect 37045 5556 37079 5565
rect 37947 5565 37949 5592
rect 37949 5565 37981 5592
rect 37947 5558 37981 5565
rect 38388 5633 38422 5635
rect 38388 5601 38422 5633
rect 38121 5565 38151 5592
rect 38151 5565 38155 5592
rect 38121 5558 38155 5565
rect 38388 5531 38422 5563
rect 38388 5529 38422 5531
rect 36548 5401 36582 5435
rect 36617 5293 36651 5327
rect 38484 5633 38518 5635
rect 38484 5601 38518 5633
rect 38484 5531 38518 5563
rect 38484 5529 38518 5531
rect 38580 5633 38614 5635
rect 38580 5601 38614 5633
rect 38580 5531 38614 5563
rect 38580 5529 38614 5531
rect 38968 6042 39002 6076
rect 40395 6349 40429 6383
rect 41513 6843 41547 6877
rect 41605 6843 41639 6877
rect 41697 6843 41731 6877
rect 42198 6866 42232 6900
rect 44038 6952 44072 6984
rect 44038 6950 44072 6952
rect 44134 7054 44168 7056
rect 44134 7022 44168 7054
rect 44230 7054 44264 7056
rect 44230 7022 44264 7054
rect 44134 6952 44168 6984
rect 44134 6950 44168 6952
rect 44230 6952 44264 6984
rect 44230 6950 44264 6952
rect 45920 7054 45954 7056
rect 45920 7022 45954 7054
rect 40956 6619 40988 6642
rect 40988 6619 40990 6642
rect 40956 6608 40990 6619
rect 41566 6729 41600 6746
rect 41566 6712 41600 6729
rect 41926 6828 41960 6862
rect 42558 6856 42592 6890
rect 42709 6851 42743 6885
rect 42801 6851 42835 6885
rect 42893 6851 42927 6885
rect 42310 6785 42344 6819
rect 41152 6602 41186 6636
rect 39996 6297 40030 6331
rect 41345 6647 41379 6648
rect 41345 6614 41377 6647
rect 41377 6614 41379 6647
rect 42166 6689 42200 6691
rect 41884 6625 41918 6659
rect 42166 6657 42200 6689
rect 42166 6587 42200 6619
rect 42166 6585 42200 6587
rect 40642 6297 40676 6331
rect 40821 6307 40855 6341
rect 40913 6307 40947 6341
rect 41005 6307 41039 6341
rect 41840 6529 41874 6531
rect 41840 6497 41874 6529
rect 41840 6427 41874 6459
rect 41840 6425 41874 6427
rect 41167 6301 41201 6335
rect 41259 6301 41293 6335
rect 41351 6301 41385 6335
rect 42262 6689 42296 6691
rect 42262 6657 42296 6689
rect 42262 6587 42296 6619
rect 42262 6585 42296 6587
rect 42358 6689 42392 6691
rect 42358 6657 42392 6689
rect 43055 6845 43089 6879
rect 43147 6845 43181 6879
rect 43239 6845 43273 6879
rect 42530 6625 42564 6659
rect 42358 6587 42392 6619
rect 42358 6585 42392 6587
rect 41928 6529 41962 6531
rect 41928 6497 41962 6529
rect 42486 6529 42520 6531
rect 42486 6497 42520 6529
rect 41928 6427 41962 6459
rect 42214 6457 42248 6491
rect 41928 6425 41962 6427
rect 42486 6427 42520 6459
rect 42486 6425 42520 6427
rect 42574 6529 42608 6531
rect 42574 6497 42608 6529
rect 42574 6427 42608 6459
rect 42574 6425 42608 6427
rect 41513 6299 41547 6333
rect 41605 6299 41639 6333
rect 41697 6299 41731 6333
rect 40054 6176 40088 6210
rect 40484 6159 40518 6193
rect 40404 6050 40438 6084
rect 40260 5998 40294 6000
rect 40260 5966 40294 5998
rect 40260 5896 40294 5928
rect 40260 5894 40294 5896
rect 40356 5998 40390 6000
rect 40356 5966 40390 5998
rect 40356 5896 40390 5928
rect 40356 5894 40390 5896
rect 40452 5998 40486 6000
rect 40452 5966 40486 5998
rect 40452 5896 40486 5928
rect 40452 5894 40486 5896
rect 38755 5797 38789 5831
rect 38847 5797 38881 5831
rect 38939 5797 38973 5831
rect 39829 5797 39863 5831
rect 39921 5797 39955 5831
rect 40013 5797 40047 5831
rect 40308 5810 40342 5844
rect 38851 5685 38885 5710
rect 38851 5676 38883 5685
rect 38883 5676 38885 5685
rect 39921 5685 39955 5715
rect 39921 5681 39923 5685
rect 39923 5681 39955 5685
rect 40420 5729 40454 5763
rect 38760 5565 38763 5594
rect 38763 5565 38794 5594
rect 38760 5560 38794 5565
rect 38933 5565 38965 5590
rect 38965 5565 38967 5590
rect 38933 5556 38967 5565
rect 39835 5565 39837 5592
rect 39837 5565 39869 5592
rect 39835 5558 39869 5565
rect 40276 5633 40310 5635
rect 40276 5601 40310 5633
rect 40009 5565 40039 5592
rect 40039 5565 40043 5592
rect 40009 5558 40043 5565
rect 40276 5531 40310 5563
rect 40276 5529 40310 5531
rect 38436 5401 38470 5435
rect 38505 5293 38539 5327
rect 40372 5633 40406 5635
rect 40372 5601 40406 5633
rect 40372 5531 40406 5563
rect 40372 5529 40406 5531
rect 40468 5633 40502 5635
rect 40468 5601 40502 5633
rect 40468 5531 40502 5563
rect 40468 5529 40502 5531
rect 40856 6042 40890 6076
rect 42283 6349 42317 6383
rect 43401 6843 43435 6877
rect 43493 6843 43527 6877
rect 43585 6843 43619 6877
rect 44086 6866 44120 6900
rect 45920 6952 45954 6984
rect 45920 6950 45954 6952
rect 46016 7054 46050 7056
rect 46016 7022 46050 7054
rect 46112 7054 46146 7056
rect 46112 7022 46146 7054
rect 46016 6952 46050 6984
rect 46016 6950 46050 6952
rect 46112 6952 46146 6984
rect 46112 6950 46146 6952
rect 47808 7054 47842 7056
rect 47808 7022 47842 7054
rect 42844 6619 42876 6642
rect 42876 6619 42878 6642
rect 42844 6608 42878 6619
rect 43454 6729 43488 6746
rect 43454 6712 43488 6729
rect 43814 6828 43848 6862
rect 44446 6856 44480 6890
rect 44597 6851 44631 6885
rect 44689 6851 44723 6885
rect 44781 6851 44815 6885
rect 44198 6785 44232 6819
rect 43040 6602 43074 6636
rect 41884 6297 41918 6331
rect 43233 6647 43267 6648
rect 43233 6614 43265 6647
rect 43265 6614 43267 6647
rect 44054 6689 44088 6691
rect 43772 6625 43806 6659
rect 44054 6657 44088 6689
rect 44054 6587 44088 6619
rect 44054 6585 44088 6587
rect 42530 6297 42564 6331
rect 42709 6307 42743 6341
rect 42801 6307 42835 6341
rect 42893 6307 42927 6341
rect 43728 6529 43762 6531
rect 43728 6497 43762 6529
rect 43728 6427 43762 6459
rect 43728 6425 43762 6427
rect 43055 6301 43089 6335
rect 43147 6301 43181 6335
rect 43239 6301 43273 6335
rect 44150 6689 44184 6691
rect 44150 6657 44184 6689
rect 44150 6587 44184 6619
rect 44150 6585 44184 6587
rect 44246 6689 44280 6691
rect 44246 6657 44280 6689
rect 44937 6845 44971 6879
rect 45029 6845 45063 6879
rect 45121 6845 45155 6879
rect 44418 6625 44452 6659
rect 44246 6587 44280 6619
rect 44246 6585 44280 6587
rect 43816 6529 43850 6531
rect 43816 6497 43850 6529
rect 44374 6529 44408 6531
rect 44374 6497 44408 6529
rect 43816 6427 43850 6459
rect 44102 6457 44136 6491
rect 43816 6425 43850 6427
rect 44374 6427 44408 6459
rect 44374 6425 44408 6427
rect 44462 6529 44496 6531
rect 44462 6497 44496 6529
rect 44462 6427 44496 6459
rect 44462 6425 44496 6427
rect 43401 6299 43435 6333
rect 43493 6299 43527 6333
rect 43585 6299 43619 6333
rect 41942 6176 41976 6210
rect 42372 6159 42406 6193
rect 42292 6050 42326 6084
rect 42148 5998 42182 6000
rect 42148 5966 42182 5998
rect 42148 5896 42182 5928
rect 42148 5894 42182 5896
rect 42244 5998 42278 6000
rect 42244 5966 42278 5998
rect 42244 5896 42278 5928
rect 42244 5894 42278 5896
rect 42340 5998 42374 6000
rect 42340 5966 42374 5998
rect 42340 5896 42374 5928
rect 42340 5894 42374 5896
rect 40643 5797 40677 5831
rect 40735 5797 40769 5831
rect 40827 5797 40861 5831
rect 41717 5797 41751 5831
rect 41809 5797 41843 5831
rect 41901 5797 41935 5831
rect 42196 5810 42230 5844
rect 40739 5685 40773 5710
rect 40739 5676 40771 5685
rect 40771 5676 40773 5685
rect 41809 5685 41843 5715
rect 41809 5681 41811 5685
rect 41811 5681 41843 5685
rect 42308 5729 42342 5763
rect 40648 5565 40651 5594
rect 40651 5565 40682 5594
rect 40648 5560 40682 5565
rect 40821 5565 40853 5590
rect 40853 5565 40855 5590
rect 40821 5556 40855 5565
rect 41723 5565 41725 5592
rect 41725 5565 41757 5592
rect 41723 5558 41757 5565
rect 42164 5633 42198 5635
rect 42164 5601 42198 5633
rect 41897 5565 41927 5592
rect 41927 5565 41931 5592
rect 41897 5558 41931 5565
rect 42164 5531 42198 5563
rect 42164 5529 42198 5531
rect 40324 5401 40358 5435
rect 40393 5293 40427 5327
rect 42260 5633 42294 5635
rect 42260 5601 42294 5633
rect 42260 5531 42294 5563
rect 42260 5529 42294 5531
rect 42356 5633 42390 5635
rect 42356 5601 42390 5633
rect 42356 5531 42390 5563
rect 42356 5529 42390 5531
rect 42744 6042 42778 6076
rect 44171 6349 44205 6383
rect 45283 6843 45317 6877
rect 45375 6843 45409 6877
rect 45467 6843 45501 6877
rect 45968 6866 46002 6900
rect 47808 6952 47842 6984
rect 47808 6950 47842 6952
rect 47904 7054 47938 7056
rect 47904 7022 47938 7054
rect 48000 7054 48034 7056
rect 48000 7022 48034 7054
rect 47904 6952 47938 6984
rect 47904 6950 47938 6952
rect 48000 6952 48034 6984
rect 48000 6950 48034 6952
rect 49696 7054 49730 7056
rect 49696 7022 49730 7054
rect 44732 6619 44764 6642
rect 44764 6619 44766 6642
rect 44732 6608 44766 6619
rect 45336 6729 45370 6746
rect 45336 6712 45370 6729
rect 45696 6828 45730 6862
rect 46328 6856 46362 6890
rect 46479 6851 46513 6885
rect 46571 6851 46605 6885
rect 46663 6851 46697 6885
rect 46080 6785 46114 6819
rect 44922 6602 44956 6636
rect 43772 6297 43806 6331
rect 45115 6647 45149 6648
rect 45115 6614 45147 6647
rect 45147 6614 45149 6647
rect 45936 6689 45970 6691
rect 45654 6625 45688 6659
rect 45936 6657 45970 6689
rect 45936 6587 45970 6619
rect 45936 6585 45970 6587
rect 44418 6297 44452 6331
rect 44597 6307 44631 6341
rect 44689 6307 44723 6341
rect 44781 6307 44815 6341
rect 45610 6529 45644 6531
rect 45610 6497 45644 6529
rect 45610 6427 45644 6459
rect 45610 6425 45644 6427
rect 44937 6301 44971 6335
rect 45029 6301 45063 6335
rect 45121 6301 45155 6335
rect 46032 6689 46066 6691
rect 46032 6657 46066 6689
rect 46032 6587 46066 6619
rect 46032 6585 46066 6587
rect 46128 6689 46162 6691
rect 46128 6657 46162 6689
rect 46825 6845 46859 6879
rect 46917 6845 46951 6879
rect 47009 6845 47043 6879
rect 46300 6625 46334 6659
rect 46128 6587 46162 6619
rect 46128 6585 46162 6587
rect 45698 6529 45732 6531
rect 45698 6497 45732 6529
rect 46256 6529 46290 6531
rect 46256 6497 46290 6529
rect 45698 6427 45732 6459
rect 45984 6457 46018 6491
rect 45698 6425 45732 6427
rect 46256 6427 46290 6459
rect 46256 6425 46290 6427
rect 46344 6529 46378 6531
rect 46344 6497 46378 6529
rect 46344 6427 46378 6459
rect 46344 6425 46378 6427
rect 45283 6299 45317 6333
rect 45375 6299 45409 6333
rect 45467 6299 45501 6333
rect 43830 6176 43864 6210
rect 44260 6159 44294 6193
rect 44180 6050 44214 6084
rect 44036 5998 44070 6000
rect 44036 5966 44070 5998
rect 44036 5896 44070 5928
rect 44036 5894 44070 5896
rect 44132 5998 44166 6000
rect 44132 5966 44166 5998
rect 44132 5896 44166 5928
rect 44132 5894 44166 5896
rect 44228 5998 44262 6000
rect 44228 5966 44262 5998
rect 44228 5896 44262 5928
rect 44228 5894 44262 5896
rect 42531 5797 42565 5831
rect 42623 5797 42657 5831
rect 42715 5797 42749 5831
rect 43605 5797 43639 5831
rect 43697 5797 43731 5831
rect 43789 5797 43823 5831
rect 44084 5810 44118 5844
rect 42627 5685 42661 5710
rect 42627 5676 42659 5685
rect 42659 5676 42661 5685
rect 43697 5685 43731 5715
rect 43697 5681 43699 5685
rect 43699 5681 43731 5685
rect 44196 5729 44230 5763
rect 42536 5565 42539 5594
rect 42539 5565 42570 5594
rect 42536 5560 42570 5565
rect 42709 5565 42741 5590
rect 42741 5565 42743 5590
rect 42709 5556 42743 5565
rect 43611 5565 43613 5592
rect 43613 5565 43645 5592
rect 43611 5558 43645 5565
rect 44052 5633 44086 5635
rect 44052 5601 44086 5633
rect 43785 5565 43815 5592
rect 43815 5565 43819 5592
rect 43785 5558 43819 5565
rect 44052 5531 44086 5563
rect 44052 5529 44086 5531
rect 42212 5401 42246 5435
rect 42281 5293 42315 5327
rect 44148 5633 44182 5635
rect 44148 5601 44182 5633
rect 44148 5531 44182 5563
rect 44148 5529 44182 5531
rect 44244 5633 44278 5635
rect 44244 5601 44278 5633
rect 44244 5531 44278 5563
rect 44244 5529 44278 5531
rect 44632 6042 44666 6076
rect 46053 6349 46087 6383
rect 47171 6843 47205 6877
rect 47263 6843 47297 6877
rect 47355 6843 47389 6877
rect 47856 6866 47890 6900
rect 49696 6952 49730 6984
rect 49696 6950 49730 6952
rect 49792 7054 49826 7056
rect 49792 7022 49826 7054
rect 49888 7054 49922 7056
rect 49888 7022 49922 7054
rect 49792 6952 49826 6984
rect 49792 6950 49826 6952
rect 49888 6952 49922 6984
rect 49888 6950 49922 6952
rect 51584 7054 51618 7056
rect 51584 7022 51618 7054
rect 46614 6619 46646 6642
rect 46646 6619 46648 6642
rect 46614 6608 46648 6619
rect 47224 6729 47258 6746
rect 47224 6712 47258 6729
rect 47584 6828 47618 6862
rect 48216 6856 48250 6890
rect 48367 6851 48401 6885
rect 48459 6851 48493 6885
rect 48551 6851 48585 6885
rect 47968 6785 48002 6819
rect 46810 6602 46844 6636
rect 45654 6297 45688 6331
rect 47003 6647 47037 6648
rect 47003 6614 47035 6647
rect 47035 6614 47037 6647
rect 47824 6689 47858 6691
rect 47542 6625 47576 6659
rect 47824 6657 47858 6689
rect 47824 6587 47858 6619
rect 47824 6585 47858 6587
rect 46300 6297 46334 6331
rect 46479 6307 46513 6341
rect 46571 6307 46605 6341
rect 46663 6307 46697 6341
rect 47498 6529 47532 6531
rect 47498 6497 47532 6529
rect 47498 6427 47532 6459
rect 47498 6425 47532 6427
rect 46825 6301 46859 6335
rect 46917 6301 46951 6335
rect 47009 6301 47043 6335
rect 47920 6689 47954 6691
rect 47920 6657 47954 6689
rect 47920 6587 47954 6619
rect 47920 6585 47954 6587
rect 48016 6689 48050 6691
rect 48016 6657 48050 6689
rect 48713 6845 48747 6879
rect 48805 6845 48839 6879
rect 48897 6845 48931 6879
rect 48188 6625 48222 6659
rect 48016 6587 48050 6619
rect 48016 6585 48050 6587
rect 47586 6529 47620 6531
rect 47586 6497 47620 6529
rect 48144 6529 48178 6531
rect 48144 6497 48178 6529
rect 47586 6427 47620 6459
rect 47872 6457 47906 6491
rect 47586 6425 47620 6427
rect 48144 6427 48178 6459
rect 48144 6425 48178 6427
rect 48232 6529 48266 6531
rect 48232 6497 48266 6529
rect 48232 6427 48266 6459
rect 48232 6425 48266 6427
rect 47171 6299 47205 6333
rect 47263 6299 47297 6333
rect 47355 6299 47389 6333
rect 45712 6176 45746 6210
rect 46142 6159 46176 6193
rect 46062 6050 46096 6084
rect 45918 5998 45952 6000
rect 45918 5966 45952 5998
rect 45918 5896 45952 5928
rect 45918 5894 45952 5896
rect 46014 5998 46048 6000
rect 46014 5966 46048 5998
rect 46014 5896 46048 5928
rect 46014 5894 46048 5896
rect 46110 5998 46144 6000
rect 46110 5966 46144 5998
rect 46110 5896 46144 5928
rect 46110 5894 46144 5896
rect 44419 5797 44453 5831
rect 44511 5797 44545 5831
rect 44603 5797 44637 5831
rect 45487 5797 45521 5831
rect 45579 5797 45613 5831
rect 45671 5797 45705 5831
rect 45966 5810 46000 5844
rect 44515 5685 44549 5710
rect 44515 5676 44547 5685
rect 44547 5676 44549 5685
rect 45579 5685 45613 5715
rect 45579 5681 45581 5685
rect 45581 5681 45613 5685
rect 46078 5729 46112 5763
rect 44424 5565 44427 5594
rect 44427 5565 44458 5594
rect 44424 5560 44458 5565
rect 44597 5565 44629 5590
rect 44629 5565 44631 5590
rect 44597 5556 44631 5565
rect 45493 5565 45495 5592
rect 45495 5565 45527 5592
rect 45493 5558 45527 5565
rect 45934 5633 45968 5635
rect 45934 5601 45968 5633
rect 45667 5565 45697 5592
rect 45697 5565 45701 5592
rect 45667 5558 45701 5565
rect 45934 5531 45968 5563
rect 45934 5529 45968 5531
rect 44100 5401 44134 5435
rect 44169 5293 44203 5327
rect 46030 5633 46064 5635
rect 46030 5601 46064 5633
rect 46030 5531 46064 5563
rect 46030 5529 46064 5531
rect 46126 5633 46160 5635
rect 46126 5601 46160 5633
rect 46126 5531 46160 5563
rect 46126 5529 46160 5531
rect 46514 6042 46548 6076
rect 47941 6349 47975 6383
rect 49059 6843 49093 6877
rect 49151 6843 49185 6877
rect 49243 6843 49277 6877
rect 49744 6866 49778 6900
rect 51584 6952 51618 6984
rect 51584 6950 51618 6952
rect 51680 7054 51714 7056
rect 51680 7022 51714 7054
rect 51776 7054 51810 7056
rect 51776 7022 51810 7054
rect 51680 6952 51714 6984
rect 51680 6950 51714 6952
rect 51776 6952 51810 6984
rect 51776 6950 51810 6952
rect 53472 7054 53506 7056
rect 53472 7022 53506 7054
rect 48502 6619 48534 6642
rect 48534 6619 48536 6642
rect 48502 6608 48536 6619
rect 49112 6729 49146 6746
rect 49112 6712 49146 6729
rect 49472 6828 49506 6862
rect 50104 6856 50138 6890
rect 50255 6851 50289 6885
rect 50347 6851 50381 6885
rect 50439 6851 50473 6885
rect 49856 6785 49890 6819
rect 48698 6602 48732 6636
rect 47542 6297 47576 6331
rect 48891 6647 48925 6648
rect 48891 6614 48923 6647
rect 48923 6614 48925 6647
rect 49712 6689 49746 6691
rect 49430 6625 49464 6659
rect 49712 6657 49746 6689
rect 49712 6587 49746 6619
rect 49712 6585 49746 6587
rect 48188 6297 48222 6331
rect 48367 6307 48401 6341
rect 48459 6307 48493 6341
rect 48551 6307 48585 6341
rect 49386 6529 49420 6531
rect 49386 6497 49420 6529
rect 49386 6427 49420 6459
rect 49386 6425 49420 6427
rect 48713 6301 48747 6335
rect 48805 6301 48839 6335
rect 48897 6301 48931 6335
rect 49808 6689 49842 6691
rect 49808 6657 49842 6689
rect 49808 6587 49842 6619
rect 49808 6585 49842 6587
rect 49904 6689 49938 6691
rect 49904 6657 49938 6689
rect 50601 6845 50635 6879
rect 50693 6845 50727 6879
rect 50785 6845 50819 6879
rect 50076 6625 50110 6659
rect 49904 6587 49938 6619
rect 49904 6585 49938 6587
rect 49474 6529 49508 6531
rect 49474 6497 49508 6529
rect 50032 6529 50066 6531
rect 50032 6497 50066 6529
rect 49474 6427 49508 6459
rect 49760 6457 49794 6491
rect 49474 6425 49508 6427
rect 50032 6427 50066 6459
rect 50032 6425 50066 6427
rect 50120 6529 50154 6531
rect 50120 6497 50154 6529
rect 50120 6427 50154 6459
rect 50120 6425 50154 6427
rect 49059 6299 49093 6333
rect 49151 6299 49185 6333
rect 49243 6299 49277 6333
rect 47600 6176 47634 6210
rect 48030 6159 48064 6193
rect 47950 6050 47984 6084
rect 47806 5998 47840 6000
rect 47806 5966 47840 5998
rect 47806 5896 47840 5928
rect 47806 5894 47840 5896
rect 47902 5998 47936 6000
rect 47902 5966 47936 5998
rect 47902 5896 47936 5928
rect 47902 5894 47936 5896
rect 47998 5998 48032 6000
rect 47998 5966 48032 5998
rect 47998 5896 48032 5928
rect 47998 5894 48032 5896
rect 46301 5797 46335 5831
rect 46393 5797 46427 5831
rect 46485 5797 46519 5831
rect 47375 5797 47409 5831
rect 47467 5797 47501 5831
rect 47559 5797 47593 5831
rect 47854 5810 47888 5844
rect 46397 5685 46431 5710
rect 46397 5676 46429 5685
rect 46429 5676 46431 5685
rect 47467 5685 47501 5715
rect 47467 5681 47469 5685
rect 47469 5681 47501 5685
rect 47966 5729 48000 5763
rect 46306 5565 46309 5594
rect 46309 5565 46340 5594
rect 46306 5560 46340 5565
rect 46479 5565 46511 5590
rect 46511 5565 46513 5590
rect 46479 5556 46513 5565
rect 47381 5565 47383 5592
rect 47383 5565 47415 5592
rect 47381 5558 47415 5565
rect 47822 5633 47856 5635
rect 47822 5601 47856 5633
rect 47555 5565 47585 5592
rect 47585 5565 47589 5592
rect 47555 5558 47589 5565
rect 47822 5531 47856 5563
rect 47822 5529 47856 5531
rect 45982 5401 46016 5435
rect 46051 5293 46085 5327
rect 47918 5633 47952 5635
rect 47918 5601 47952 5633
rect 47918 5531 47952 5563
rect 47918 5529 47952 5531
rect 48014 5633 48048 5635
rect 48014 5601 48048 5633
rect 48014 5531 48048 5563
rect 48014 5529 48048 5531
rect 48402 6042 48436 6076
rect 49829 6349 49863 6383
rect 50947 6843 50981 6877
rect 51039 6843 51073 6877
rect 51131 6843 51165 6877
rect 51632 6866 51666 6900
rect 53472 6952 53506 6984
rect 53472 6950 53506 6952
rect 53568 7054 53602 7056
rect 53568 7022 53602 7054
rect 53664 7054 53698 7056
rect 53664 7022 53698 7054
rect 53568 6952 53602 6984
rect 53568 6950 53602 6952
rect 53664 6952 53698 6984
rect 53664 6950 53698 6952
rect 55360 7054 55394 7056
rect 55360 7022 55394 7054
rect 50390 6619 50422 6642
rect 50422 6619 50424 6642
rect 50390 6608 50424 6619
rect 51000 6729 51034 6746
rect 51000 6712 51034 6729
rect 51360 6828 51394 6862
rect 51992 6856 52026 6890
rect 52143 6851 52177 6885
rect 52235 6851 52269 6885
rect 52327 6851 52361 6885
rect 51744 6785 51778 6819
rect 50586 6602 50620 6636
rect 49430 6297 49464 6331
rect 50779 6647 50813 6648
rect 50779 6614 50811 6647
rect 50811 6614 50813 6647
rect 51600 6689 51634 6691
rect 51318 6625 51352 6659
rect 51600 6657 51634 6689
rect 51600 6587 51634 6619
rect 51600 6585 51634 6587
rect 50076 6297 50110 6331
rect 50255 6307 50289 6341
rect 50347 6307 50381 6341
rect 50439 6307 50473 6341
rect 51274 6529 51308 6531
rect 51274 6497 51308 6529
rect 51274 6427 51308 6459
rect 51274 6425 51308 6427
rect 50601 6301 50635 6335
rect 50693 6301 50727 6335
rect 50785 6301 50819 6335
rect 51696 6689 51730 6691
rect 51696 6657 51730 6689
rect 51696 6587 51730 6619
rect 51696 6585 51730 6587
rect 51792 6689 51826 6691
rect 51792 6657 51826 6689
rect 52489 6845 52523 6879
rect 52581 6845 52615 6879
rect 52673 6845 52707 6879
rect 51964 6625 51998 6659
rect 51792 6587 51826 6619
rect 51792 6585 51826 6587
rect 51362 6529 51396 6531
rect 51362 6497 51396 6529
rect 51920 6529 51954 6531
rect 51920 6497 51954 6529
rect 51362 6427 51396 6459
rect 51648 6457 51682 6491
rect 51362 6425 51396 6427
rect 51920 6427 51954 6459
rect 51920 6425 51954 6427
rect 52008 6529 52042 6531
rect 52008 6497 52042 6529
rect 52008 6427 52042 6459
rect 52008 6425 52042 6427
rect 50947 6299 50981 6333
rect 51039 6299 51073 6333
rect 51131 6299 51165 6333
rect 49488 6176 49522 6210
rect 49918 6159 49952 6193
rect 49838 6050 49872 6084
rect 49694 5998 49728 6000
rect 49694 5966 49728 5998
rect 49694 5896 49728 5928
rect 49694 5894 49728 5896
rect 49790 5998 49824 6000
rect 49790 5966 49824 5998
rect 49790 5896 49824 5928
rect 49790 5894 49824 5896
rect 49886 5998 49920 6000
rect 49886 5966 49920 5998
rect 49886 5896 49920 5928
rect 49886 5894 49920 5896
rect 48189 5797 48223 5831
rect 48281 5797 48315 5831
rect 48373 5797 48407 5831
rect 49263 5797 49297 5831
rect 49355 5797 49389 5831
rect 49447 5797 49481 5831
rect 49742 5810 49776 5844
rect 48285 5685 48319 5710
rect 48285 5676 48317 5685
rect 48317 5676 48319 5685
rect 49355 5685 49389 5715
rect 49355 5681 49357 5685
rect 49357 5681 49389 5685
rect 49854 5729 49888 5763
rect 48194 5565 48197 5594
rect 48197 5565 48228 5594
rect 48194 5560 48228 5565
rect 48367 5565 48399 5590
rect 48399 5565 48401 5590
rect 48367 5556 48401 5565
rect 49269 5565 49271 5592
rect 49271 5565 49303 5592
rect 49269 5558 49303 5565
rect 49710 5633 49744 5635
rect 49710 5601 49744 5633
rect 49443 5565 49473 5592
rect 49473 5565 49477 5592
rect 49443 5558 49477 5565
rect 49710 5531 49744 5563
rect 49710 5529 49744 5531
rect 47870 5401 47904 5435
rect 47939 5293 47973 5327
rect 49806 5633 49840 5635
rect 49806 5601 49840 5633
rect 49806 5531 49840 5563
rect 49806 5529 49840 5531
rect 49902 5633 49936 5635
rect 49902 5601 49936 5633
rect 49902 5531 49936 5563
rect 49902 5529 49936 5531
rect 50290 6042 50324 6076
rect 51717 6349 51751 6383
rect 52835 6843 52869 6877
rect 52927 6843 52961 6877
rect 53019 6843 53053 6877
rect 53520 6866 53554 6900
rect 55360 6952 55394 6984
rect 55360 6950 55394 6952
rect 55456 7054 55490 7056
rect 55456 7022 55490 7054
rect 55552 7054 55586 7056
rect 55552 7022 55586 7054
rect 55456 6952 55490 6984
rect 55456 6950 55490 6952
rect 55552 6952 55586 6984
rect 55552 6950 55586 6952
rect 57248 7054 57282 7056
rect 57248 7022 57282 7054
rect 52278 6619 52310 6642
rect 52310 6619 52312 6642
rect 52278 6608 52312 6619
rect 52888 6729 52922 6746
rect 52888 6712 52922 6729
rect 53248 6828 53282 6862
rect 53880 6856 53914 6890
rect 54031 6851 54065 6885
rect 54123 6851 54157 6885
rect 54215 6851 54249 6885
rect 53632 6785 53666 6819
rect 52474 6602 52508 6636
rect 51318 6297 51352 6331
rect 52667 6647 52701 6648
rect 52667 6614 52699 6647
rect 52699 6614 52701 6647
rect 53488 6689 53522 6691
rect 53206 6625 53240 6659
rect 53488 6657 53522 6689
rect 53488 6587 53522 6619
rect 53488 6585 53522 6587
rect 51964 6297 51998 6331
rect 52143 6307 52177 6341
rect 52235 6307 52269 6341
rect 52327 6307 52361 6341
rect 53162 6529 53196 6531
rect 53162 6497 53196 6529
rect 53162 6427 53196 6459
rect 53162 6425 53196 6427
rect 52489 6301 52523 6335
rect 52581 6301 52615 6335
rect 52673 6301 52707 6335
rect 53584 6689 53618 6691
rect 53584 6657 53618 6689
rect 53584 6587 53618 6619
rect 53584 6585 53618 6587
rect 53680 6689 53714 6691
rect 53680 6657 53714 6689
rect 54377 6845 54411 6879
rect 54469 6845 54503 6879
rect 54561 6845 54595 6879
rect 53852 6625 53886 6659
rect 53680 6587 53714 6619
rect 53680 6585 53714 6587
rect 53250 6529 53284 6531
rect 53250 6497 53284 6529
rect 53808 6529 53842 6531
rect 53808 6497 53842 6529
rect 53250 6427 53284 6459
rect 53536 6457 53570 6491
rect 53250 6425 53284 6427
rect 53808 6427 53842 6459
rect 53808 6425 53842 6427
rect 53896 6529 53930 6531
rect 53896 6497 53930 6529
rect 53896 6427 53930 6459
rect 53896 6425 53930 6427
rect 52835 6299 52869 6333
rect 52927 6299 52961 6333
rect 53019 6299 53053 6333
rect 51376 6176 51410 6210
rect 51806 6159 51840 6193
rect 51726 6050 51760 6084
rect 51582 5998 51616 6000
rect 51582 5966 51616 5998
rect 51582 5896 51616 5928
rect 51582 5894 51616 5896
rect 51678 5998 51712 6000
rect 51678 5966 51712 5998
rect 51678 5896 51712 5928
rect 51678 5894 51712 5896
rect 51774 5998 51808 6000
rect 51774 5966 51808 5998
rect 51774 5896 51808 5928
rect 51774 5894 51808 5896
rect 50077 5797 50111 5831
rect 50169 5797 50203 5831
rect 50261 5797 50295 5831
rect 51151 5797 51185 5831
rect 51243 5797 51277 5831
rect 51335 5797 51369 5831
rect 51630 5810 51664 5844
rect 50173 5685 50207 5710
rect 50173 5676 50205 5685
rect 50205 5676 50207 5685
rect 51243 5685 51277 5715
rect 51243 5681 51245 5685
rect 51245 5681 51277 5685
rect 51742 5729 51776 5763
rect 50082 5565 50085 5594
rect 50085 5565 50116 5594
rect 50082 5560 50116 5565
rect 50255 5565 50287 5590
rect 50287 5565 50289 5590
rect 50255 5556 50289 5565
rect 51157 5565 51159 5592
rect 51159 5565 51191 5592
rect 51157 5558 51191 5565
rect 51598 5633 51632 5635
rect 51598 5601 51632 5633
rect 51331 5565 51361 5592
rect 51361 5565 51365 5592
rect 51331 5558 51365 5565
rect 51598 5531 51632 5563
rect 51598 5529 51632 5531
rect 49758 5401 49792 5435
rect 49827 5293 49861 5327
rect 51694 5633 51728 5635
rect 51694 5601 51728 5633
rect 51694 5531 51728 5563
rect 51694 5529 51728 5531
rect 51790 5633 51824 5635
rect 51790 5601 51824 5633
rect 51790 5531 51824 5563
rect 51790 5529 51824 5531
rect 52178 6042 52212 6076
rect 53605 6349 53639 6383
rect 54723 6843 54757 6877
rect 54815 6843 54849 6877
rect 54907 6843 54941 6877
rect 55408 6866 55442 6900
rect 57248 6952 57282 6984
rect 57248 6950 57282 6952
rect 57344 7054 57378 7056
rect 57344 7022 57378 7054
rect 57440 7054 57474 7056
rect 57440 7022 57474 7054
rect 57344 6952 57378 6984
rect 57344 6950 57378 6952
rect 57440 6952 57474 6984
rect 57440 6950 57474 6952
rect 59136 7054 59170 7056
rect 59136 7022 59170 7054
rect 54166 6619 54198 6642
rect 54198 6619 54200 6642
rect 54166 6608 54200 6619
rect 54776 6729 54810 6746
rect 54776 6712 54810 6729
rect 55136 6828 55170 6862
rect 55768 6856 55802 6890
rect 55919 6851 55953 6885
rect 56011 6851 56045 6885
rect 56103 6851 56137 6885
rect 55520 6785 55554 6819
rect 54362 6602 54396 6636
rect 53206 6297 53240 6331
rect 54555 6647 54589 6648
rect 54555 6614 54587 6647
rect 54587 6614 54589 6647
rect 55376 6689 55410 6691
rect 55094 6625 55128 6659
rect 55376 6657 55410 6689
rect 55376 6587 55410 6619
rect 55376 6585 55410 6587
rect 53852 6297 53886 6331
rect 54031 6307 54065 6341
rect 54123 6307 54157 6341
rect 54215 6307 54249 6341
rect 55050 6529 55084 6531
rect 55050 6497 55084 6529
rect 55050 6427 55084 6459
rect 55050 6425 55084 6427
rect 54377 6301 54411 6335
rect 54469 6301 54503 6335
rect 54561 6301 54595 6335
rect 55472 6689 55506 6691
rect 55472 6657 55506 6689
rect 55472 6587 55506 6619
rect 55472 6585 55506 6587
rect 55568 6689 55602 6691
rect 55568 6657 55602 6689
rect 56265 6845 56299 6879
rect 56357 6845 56391 6879
rect 56449 6845 56483 6879
rect 55740 6625 55774 6659
rect 55568 6587 55602 6619
rect 55568 6585 55602 6587
rect 55138 6529 55172 6531
rect 55138 6497 55172 6529
rect 55696 6529 55730 6531
rect 55696 6497 55730 6529
rect 55138 6427 55172 6459
rect 55424 6457 55458 6491
rect 55138 6425 55172 6427
rect 55696 6427 55730 6459
rect 55696 6425 55730 6427
rect 55784 6529 55818 6531
rect 55784 6497 55818 6529
rect 55784 6427 55818 6459
rect 55784 6425 55818 6427
rect 54723 6299 54757 6333
rect 54815 6299 54849 6333
rect 54907 6299 54941 6333
rect 53264 6176 53298 6210
rect 53694 6159 53728 6193
rect 53614 6050 53648 6084
rect 53470 5998 53504 6000
rect 53470 5966 53504 5998
rect 53470 5896 53504 5928
rect 53470 5894 53504 5896
rect 53566 5998 53600 6000
rect 53566 5966 53600 5998
rect 53566 5896 53600 5928
rect 53566 5894 53600 5896
rect 53662 5998 53696 6000
rect 53662 5966 53696 5998
rect 53662 5896 53696 5928
rect 53662 5894 53696 5896
rect 51965 5797 51999 5831
rect 52057 5797 52091 5831
rect 52149 5797 52183 5831
rect 53039 5797 53073 5831
rect 53131 5797 53165 5831
rect 53223 5797 53257 5831
rect 53518 5810 53552 5844
rect 52061 5685 52095 5710
rect 52061 5676 52093 5685
rect 52093 5676 52095 5685
rect 53131 5685 53165 5715
rect 53131 5681 53133 5685
rect 53133 5681 53165 5685
rect 53630 5729 53664 5763
rect 51970 5565 51973 5594
rect 51973 5565 52004 5594
rect 51970 5560 52004 5565
rect 52143 5565 52175 5590
rect 52175 5565 52177 5590
rect 52143 5556 52177 5565
rect 53045 5565 53047 5592
rect 53047 5565 53079 5592
rect 53045 5558 53079 5565
rect 53486 5633 53520 5635
rect 53486 5601 53520 5633
rect 53219 5565 53249 5592
rect 53249 5565 53253 5592
rect 53219 5558 53253 5565
rect 53486 5531 53520 5563
rect 53486 5529 53520 5531
rect 51646 5401 51680 5435
rect 51715 5293 51749 5327
rect 53582 5633 53616 5635
rect 53582 5601 53616 5633
rect 53582 5531 53616 5563
rect 53582 5529 53616 5531
rect 53678 5633 53712 5635
rect 53678 5601 53712 5633
rect 53678 5531 53712 5563
rect 53678 5529 53712 5531
rect 54066 6042 54100 6076
rect 55493 6349 55527 6383
rect 56611 6843 56645 6877
rect 56703 6843 56737 6877
rect 56795 6843 56829 6877
rect 57296 6866 57330 6900
rect 59136 6952 59170 6984
rect 59136 6950 59170 6952
rect 59232 7054 59266 7056
rect 59232 7022 59266 7054
rect 59328 7054 59362 7056
rect 59328 7022 59362 7054
rect 59232 6952 59266 6984
rect 59232 6950 59266 6952
rect 59328 6952 59362 6984
rect 59328 6950 59362 6952
rect 56054 6619 56086 6642
rect 56086 6619 56088 6642
rect 56054 6608 56088 6619
rect 56664 6729 56698 6746
rect 56664 6712 56698 6729
rect 57024 6828 57058 6862
rect 57656 6856 57690 6890
rect 57807 6851 57841 6885
rect 57899 6851 57933 6885
rect 57991 6851 58025 6885
rect 57408 6785 57442 6819
rect 56250 6602 56284 6636
rect 55094 6297 55128 6331
rect 56443 6647 56477 6648
rect 56443 6614 56475 6647
rect 56475 6614 56477 6647
rect 57264 6689 57298 6691
rect 56982 6625 57016 6659
rect 57264 6657 57298 6689
rect 57264 6587 57298 6619
rect 57264 6585 57298 6587
rect 55740 6297 55774 6331
rect 55919 6307 55953 6341
rect 56011 6307 56045 6341
rect 56103 6307 56137 6341
rect 56938 6529 56972 6531
rect 56938 6497 56972 6529
rect 56938 6427 56972 6459
rect 56938 6425 56972 6427
rect 56265 6301 56299 6335
rect 56357 6301 56391 6335
rect 56449 6301 56483 6335
rect 57360 6689 57394 6691
rect 57360 6657 57394 6689
rect 57360 6587 57394 6619
rect 57360 6585 57394 6587
rect 57456 6689 57490 6691
rect 57456 6657 57490 6689
rect 58153 6845 58187 6879
rect 58245 6845 58279 6879
rect 58337 6845 58371 6879
rect 57628 6625 57662 6659
rect 57456 6587 57490 6619
rect 57456 6585 57490 6587
rect 57026 6529 57060 6531
rect 57026 6497 57060 6529
rect 57584 6529 57618 6531
rect 57584 6497 57618 6529
rect 57026 6427 57060 6459
rect 57312 6457 57346 6491
rect 57026 6425 57060 6427
rect 57584 6427 57618 6459
rect 57584 6425 57618 6427
rect 57672 6529 57706 6531
rect 57672 6497 57706 6529
rect 57672 6427 57706 6459
rect 57672 6425 57706 6427
rect 56611 6299 56645 6333
rect 56703 6299 56737 6333
rect 56795 6299 56829 6333
rect 55152 6176 55186 6210
rect 55582 6159 55616 6193
rect 55502 6050 55536 6084
rect 55358 5998 55392 6000
rect 55358 5966 55392 5998
rect 55358 5896 55392 5928
rect 55358 5894 55392 5896
rect 55454 5998 55488 6000
rect 55454 5966 55488 5998
rect 55454 5896 55488 5928
rect 55454 5894 55488 5896
rect 55550 5998 55584 6000
rect 55550 5966 55584 5998
rect 55550 5896 55584 5928
rect 55550 5894 55584 5896
rect 53853 5797 53887 5831
rect 53945 5797 53979 5831
rect 54037 5797 54071 5831
rect 54927 5797 54961 5831
rect 55019 5797 55053 5831
rect 55111 5797 55145 5831
rect 55406 5810 55440 5844
rect 53949 5685 53983 5710
rect 53949 5676 53981 5685
rect 53981 5676 53983 5685
rect 55019 5685 55053 5715
rect 55019 5681 55021 5685
rect 55021 5681 55053 5685
rect 55518 5729 55552 5763
rect 53858 5565 53861 5594
rect 53861 5565 53892 5594
rect 53858 5560 53892 5565
rect 54031 5565 54063 5590
rect 54063 5565 54065 5590
rect 54031 5556 54065 5565
rect 54933 5565 54935 5592
rect 54935 5565 54967 5592
rect 54933 5558 54967 5565
rect 55374 5633 55408 5635
rect 55374 5601 55408 5633
rect 55107 5565 55137 5592
rect 55137 5565 55141 5592
rect 55107 5558 55141 5565
rect 55374 5531 55408 5563
rect 55374 5529 55408 5531
rect 53534 5401 53568 5435
rect 53603 5293 53637 5327
rect 55470 5633 55504 5635
rect 55470 5601 55504 5633
rect 55470 5531 55504 5563
rect 55470 5529 55504 5531
rect 55566 5633 55600 5635
rect 55566 5601 55600 5633
rect 55566 5531 55600 5563
rect 55566 5529 55600 5531
rect 55954 6042 55988 6076
rect 57381 6349 57415 6383
rect 58499 6843 58533 6877
rect 58591 6843 58625 6877
rect 58683 6843 58717 6877
rect 59184 6866 59218 6900
rect 57942 6619 57974 6642
rect 57974 6619 57976 6642
rect 57942 6608 57976 6619
rect 58552 6729 58586 6746
rect 58552 6712 58586 6729
rect 58912 6828 58946 6862
rect 59544 6856 59578 6890
rect 59695 6851 59729 6885
rect 59787 6851 59821 6885
rect 59879 6851 59913 6885
rect 59296 6785 59330 6819
rect 58138 6602 58172 6636
rect 56982 6297 57016 6331
rect 58331 6647 58365 6648
rect 58331 6614 58363 6647
rect 58363 6614 58365 6647
rect 59152 6689 59186 6691
rect 58870 6625 58904 6659
rect 59152 6657 59186 6689
rect 59152 6587 59186 6619
rect 59152 6585 59186 6587
rect 57628 6297 57662 6331
rect 57807 6307 57841 6341
rect 57899 6307 57933 6341
rect 57991 6307 58025 6341
rect 58826 6529 58860 6531
rect 58826 6497 58860 6529
rect 58826 6427 58860 6459
rect 58826 6425 58860 6427
rect 58153 6301 58187 6335
rect 58245 6301 58279 6335
rect 58337 6301 58371 6335
rect 59248 6689 59282 6691
rect 59248 6657 59282 6689
rect 59248 6587 59282 6619
rect 59248 6585 59282 6587
rect 59344 6689 59378 6691
rect 59344 6657 59378 6689
rect 59516 6625 59550 6659
rect 59344 6587 59378 6619
rect 59344 6585 59378 6587
rect 58914 6529 58948 6531
rect 58914 6497 58948 6529
rect 59472 6529 59506 6531
rect 59472 6497 59506 6529
rect 58914 6427 58948 6459
rect 59200 6457 59234 6491
rect 58914 6425 58948 6427
rect 59472 6427 59506 6459
rect 59472 6425 59506 6427
rect 59560 6529 59594 6531
rect 59560 6497 59594 6529
rect 59560 6427 59594 6459
rect 59560 6425 59594 6427
rect 58499 6299 58533 6333
rect 58591 6299 58625 6333
rect 58683 6299 58717 6333
rect 57040 6176 57074 6210
rect 57470 6159 57504 6193
rect 57390 6050 57424 6084
rect 57246 5998 57280 6000
rect 57246 5966 57280 5998
rect 57246 5896 57280 5928
rect 57246 5894 57280 5896
rect 57342 5998 57376 6000
rect 57342 5966 57376 5998
rect 57342 5896 57376 5928
rect 57342 5894 57376 5896
rect 57438 5998 57472 6000
rect 57438 5966 57472 5998
rect 57438 5896 57472 5928
rect 57438 5894 57472 5896
rect 55741 5797 55775 5831
rect 55833 5797 55867 5831
rect 55925 5797 55959 5831
rect 56815 5797 56849 5831
rect 56907 5797 56941 5831
rect 56999 5797 57033 5831
rect 57294 5810 57328 5844
rect 55837 5685 55871 5710
rect 55837 5676 55869 5685
rect 55869 5676 55871 5685
rect 56907 5685 56941 5715
rect 56907 5681 56909 5685
rect 56909 5681 56941 5685
rect 57406 5729 57440 5763
rect 55746 5565 55749 5594
rect 55749 5565 55780 5594
rect 55746 5560 55780 5565
rect 55919 5565 55951 5590
rect 55951 5565 55953 5590
rect 55919 5556 55953 5565
rect 56821 5565 56823 5592
rect 56823 5565 56855 5592
rect 56821 5558 56855 5565
rect 57262 5633 57296 5635
rect 57262 5601 57296 5633
rect 56995 5565 57025 5592
rect 57025 5565 57029 5592
rect 56995 5558 57029 5565
rect 57262 5531 57296 5563
rect 57262 5529 57296 5531
rect 55422 5401 55456 5435
rect 55491 5293 55525 5327
rect 57358 5633 57392 5635
rect 57358 5601 57392 5633
rect 57358 5531 57392 5563
rect 57358 5529 57392 5531
rect 57454 5633 57488 5635
rect 57454 5601 57488 5633
rect 57454 5531 57488 5563
rect 57454 5529 57488 5531
rect 57842 6042 57876 6076
rect 59269 6349 59303 6383
rect 59830 6619 59862 6642
rect 59862 6619 59864 6642
rect 59830 6608 59864 6619
rect 58870 6297 58904 6331
rect 59516 6297 59550 6331
rect 59695 6307 59729 6341
rect 59787 6307 59821 6341
rect 59879 6307 59913 6341
rect 58928 6176 58962 6210
rect 59358 6159 59392 6193
rect 59278 6050 59312 6084
rect 59134 5998 59168 6000
rect 59134 5966 59168 5998
rect 59134 5896 59168 5928
rect 59134 5894 59168 5896
rect 59230 5998 59264 6000
rect 59230 5966 59264 5998
rect 59230 5896 59264 5928
rect 59230 5894 59264 5896
rect 59326 5998 59360 6000
rect 59326 5966 59360 5998
rect 59326 5896 59360 5928
rect 59326 5894 59360 5896
rect 57629 5797 57663 5831
rect 57721 5797 57755 5831
rect 57813 5797 57847 5831
rect 58703 5797 58737 5831
rect 58795 5797 58829 5831
rect 58887 5797 58921 5831
rect 59182 5810 59216 5844
rect 57725 5685 57759 5710
rect 57725 5676 57757 5685
rect 57757 5676 57759 5685
rect 58795 5685 58829 5715
rect 58795 5681 58797 5685
rect 58797 5681 58829 5685
rect 59294 5729 59328 5763
rect 57634 5565 57637 5594
rect 57637 5565 57668 5594
rect 57634 5560 57668 5565
rect 57807 5565 57839 5590
rect 57839 5565 57841 5590
rect 57807 5556 57841 5565
rect 58709 5565 58711 5592
rect 58711 5565 58743 5592
rect 58709 5558 58743 5565
rect 59150 5633 59184 5635
rect 59150 5601 59184 5633
rect 58883 5565 58913 5592
rect 58913 5565 58917 5592
rect 58883 5558 58917 5565
rect 59150 5531 59184 5563
rect 59150 5529 59184 5531
rect 57310 5401 57344 5435
rect 57379 5293 57413 5327
rect 59246 5633 59280 5635
rect 59246 5601 59280 5633
rect 59246 5531 59280 5563
rect 59246 5529 59280 5531
rect 59342 5633 59376 5635
rect 59342 5601 59376 5633
rect 59342 5531 59376 5563
rect 59342 5529 59376 5531
rect 59730 6042 59764 6076
rect 59517 5797 59551 5831
rect 59609 5797 59643 5831
rect 59701 5797 59735 5831
rect 59613 5685 59647 5710
rect 59613 5676 59645 5685
rect 59645 5676 59647 5685
rect 59522 5565 59525 5594
rect 59525 5565 59556 5594
rect 59522 5560 59556 5565
rect 59695 5565 59727 5590
rect 59727 5565 59729 5590
rect 59695 5556 59729 5565
rect 59198 5401 59232 5435
rect 59267 5293 59301 5327
rect 187 5253 221 5287
rect 279 5253 313 5287
rect 371 5253 405 5287
rect 1001 5253 1035 5287
rect 1093 5253 1127 5287
rect 1185 5253 1219 5287
rect 2075 5253 2109 5287
rect 2167 5253 2201 5287
rect 2259 5253 2293 5287
rect 2889 5253 2923 5287
rect 2981 5253 3015 5287
rect 3073 5253 3107 5287
rect 3963 5253 3997 5287
rect 4055 5253 4089 5287
rect 4147 5253 4181 5287
rect 4777 5253 4811 5287
rect 4869 5253 4903 5287
rect 4961 5253 4995 5287
rect 5851 5253 5885 5287
rect 5943 5253 5977 5287
rect 6035 5253 6069 5287
rect 6665 5253 6699 5287
rect 6757 5253 6791 5287
rect 6849 5253 6883 5287
rect 7739 5253 7773 5287
rect 7831 5253 7865 5287
rect 7923 5253 7957 5287
rect 8553 5253 8587 5287
rect 8645 5253 8679 5287
rect 8737 5253 8771 5287
rect 9627 5253 9661 5287
rect 9719 5253 9753 5287
rect 9811 5253 9845 5287
rect 10441 5253 10475 5287
rect 10533 5253 10567 5287
rect 10625 5253 10659 5287
rect 11515 5253 11549 5287
rect 11607 5253 11641 5287
rect 11699 5253 11733 5287
rect 12329 5253 12363 5287
rect 12421 5253 12455 5287
rect 12513 5253 12547 5287
rect 13403 5253 13437 5287
rect 13495 5253 13529 5287
rect 13587 5253 13621 5287
rect 14217 5253 14251 5287
rect 14309 5253 14343 5287
rect 14401 5253 14435 5287
rect 15285 5253 15319 5287
rect 15377 5253 15411 5287
rect 15469 5253 15503 5287
rect 16099 5253 16133 5287
rect 16191 5253 16225 5287
rect 16283 5253 16317 5287
rect 17173 5253 17207 5287
rect 17265 5253 17299 5287
rect 17357 5253 17391 5287
rect 17987 5253 18021 5287
rect 18079 5253 18113 5287
rect 18171 5253 18205 5287
rect 19061 5253 19095 5287
rect 19153 5253 19187 5287
rect 19245 5253 19279 5287
rect 19875 5253 19909 5287
rect 19967 5253 20001 5287
rect 20059 5253 20093 5287
rect 20949 5253 20983 5287
rect 21041 5253 21075 5287
rect 21133 5253 21167 5287
rect 21763 5253 21797 5287
rect 21855 5253 21889 5287
rect 21947 5253 21981 5287
rect 22837 5253 22871 5287
rect 22929 5253 22963 5287
rect 23021 5253 23055 5287
rect 23651 5253 23685 5287
rect 23743 5253 23777 5287
rect 23835 5253 23869 5287
rect 24725 5253 24759 5287
rect 24817 5253 24851 5287
rect 24909 5253 24943 5287
rect 25539 5253 25573 5287
rect 25631 5253 25665 5287
rect 25723 5253 25757 5287
rect 26613 5253 26647 5287
rect 26705 5253 26739 5287
rect 26797 5253 26831 5287
rect 27427 5253 27461 5287
rect 27519 5253 27553 5287
rect 27611 5253 27645 5287
rect 28501 5253 28535 5287
rect 28593 5253 28627 5287
rect 28685 5253 28719 5287
rect 29315 5253 29349 5287
rect 29407 5253 29441 5287
rect 29499 5253 29533 5287
rect 30389 5253 30423 5287
rect 30481 5253 30515 5287
rect 30573 5253 30607 5287
rect 31203 5253 31237 5287
rect 31295 5253 31329 5287
rect 31387 5253 31421 5287
rect 32277 5253 32311 5287
rect 32369 5253 32403 5287
rect 32461 5253 32495 5287
rect 33091 5253 33125 5287
rect 33183 5253 33217 5287
rect 33275 5253 33309 5287
rect 34165 5253 34199 5287
rect 34257 5253 34291 5287
rect 34349 5253 34383 5287
rect 34979 5253 35013 5287
rect 35071 5253 35105 5287
rect 35163 5253 35197 5287
rect 36053 5253 36087 5287
rect 36145 5253 36179 5287
rect 36237 5253 36271 5287
rect 36867 5253 36901 5287
rect 36959 5253 36993 5287
rect 37051 5253 37085 5287
rect 37941 5253 37975 5287
rect 38033 5253 38067 5287
rect 38125 5253 38159 5287
rect 38755 5253 38789 5287
rect 38847 5253 38881 5287
rect 38939 5253 38973 5287
rect 39829 5253 39863 5287
rect 39921 5253 39955 5287
rect 40013 5253 40047 5287
rect 40643 5253 40677 5287
rect 40735 5253 40769 5287
rect 40827 5253 40861 5287
rect 41717 5253 41751 5287
rect 41809 5253 41843 5287
rect 41901 5253 41935 5287
rect 42531 5253 42565 5287
rect 42623 5253 42657 5287
rect 42715 5253 42749 5287
rect 43605 5253 43639 5287
rect 43697 5253 43731 5287
rect 43789 5253 43823 5287
rect 44419 5253 44453 5287
rect 44511 5253 44545 5287
rect 44603 5253 44637 5287
rect 45487 5253 45521 5287
rect 45579 5253 45613 5287
rect 45671 5253 45705 5287
rect 46301 5253 46335 5287
rect 46393 5253 46427 5287
rect 46485 5253 46519 5287
rect 47375 5253 47409 5287
rect 47467 5253 47501 5287
rect 47559 5253 47593 5287
rect 48189 5253 48223 5287
rect 48281 5253 48315 5287
rect 48373 5253 48407 5287
rect 49263 5253 49297 5287
rect 49355 5253 49389 5287
rect 49447 5253 49481 5287
rect 50077 5253 50111 5287
rect 50169 5253 50203 5287
rect 50261 5253 50295 5287
rect 51151 5253 51185 5287
rect 51243 5253 51277 5287
rect 51335 5253 51369 5287
rect 51965 5253 51999 5287
rect 52057 5253 52091 5287
rect 52149 5253 52183 5287
rect 53039 5253 53073 5287
rect 53131 5253 53165 5287
rect 53223 5253 53257 5287
rect 53853 5253 53887 5287
rect 53945 5253 53979 5287
rect 54037 5253 54071 5287
rect 54927 5253 54961 5287
rect 55019 5253 55053 5287
rect 55111 5253 55145 5287
rect 55741 5253 55775 5287
rect 55833 5253 55867 5287
rect 55925 5253 55959 5287
rect 56815 5253 56849 5287
rect 56907 5253 56941 5287
rect 56999 5253 57033 5287
rect 57629 5253 57663 5287
rect 57721 5253 57755 5287
rect 57813 5253 57847 5287
rect 58703 5253 58737 5287
rect 58795 5253 58829 5287
rect 58887 5253 58921 5287
rect 59517 5253 59551 5287
rect 59609 5253 59643 5287
rect 59701 5253 59735 5287
rect 5693 5175 5727 5209
rect 5785 5175 5819 5209
rect 5877 5175 5911 5209
rect 5969 5175 6003 5209
rect 6061 5175 6095 5209
rect 6153 5175 6187 5209
rect 6245 5175 6279 5209
rect 6337 5175 6371 5209
rect 6429 5175 6463 5209
rect 6521 5175 6555 5209
rect 6613 5175 6647 5209
rect 6705 5175 6739 5209
rect 6797 5175 6831 5209
rect 6889 5175 6923 5209
rect 6981 5175 7015 5209
rect 7073 5175 7107 5209
rect 5799 4995 5833 5005
rect 5799 4971 5828 4995
rect 5828 4971 5833 4995
rect 5962 4995 5996 5009
rect 5962 4975 5996 4995
rect 6132 4995 6166 5007
rect 6132 4973 6164 4995
rect 6164 4973 6166 4995
rect 6297 4995 6331 5007
rect 6297 4973 6298 4995
rect 6298 4973 6331 4995
rect 6466 4961 6500 4993
rect 6637 4995 6671 4996
rect 6637 4962 6668 4995
rect 6668 4962 6671 4995
rect 6799 4995 6833 5001
rect 6799 4967 6802 4995
rect 6802 4967 6833 4995
rect 6972 4995 7006 5002
rect 6972 4968 7004 4995
rect 7004 4968 7006 4995
rect 6466 4959 6500 4961
rect 7575 5173 7609 5207
rect 7667 5173 7701 5207
rect 7759 5173 7793 5207
rect 7851 5173 7885 5207
rect 7943 5173 7977 5207
rect 8035 5173 8069 5207
rect 8127 5173 8161 5207
rect 8219 5173 8253 5207
rect 8311 5173 8345 5207
rect 8403 5173 8437 5207
rect 8495 5173 8529 5207
rect 8587 5173 8621 5207
rect 8679 5173 8713 5207
rect 8771 5173 8805 5207
rect 8863 5173 8897 5207
rect 8955 5173 8989 5207
rect 20791 5175 20825 5209
rect 20883 5175 20917 5209
rect 20975 5175 21009 5209
rect 21067 5175 21101 5209
rect 21159 5175 21193 5209
rect 21251 5175 21285 5209
rect 21343 5175 21377 5209
rect 21435 5175 21469 5209
rect 21527 5175 21561 5209
rect 21619 5175 21653 5209
rect 21711 5175 21745 5209
rect 21803 5175 21837 5209
rect 21895 5175 21929 5209
rect 21987 5175 22021 5209
rect 22079 5175 22113 5209
rect 22171 5175 22205 5209
rect 7845 4993 7879 5003
rect 7845 4969 7878 4993
rect 7878 4969 7879 4993
rect 8015 4993 8049 5012
rect 8015 4978 8046 4993
rect 8046 4978 8049 4993
rect 8183 4993 8217 5010
rect 8183 4976 8214 4993
rect 8214 4976 8217 4993
rect 8350 4993 8384 4997
rect 8350 4963 8382 4993
rect 8382 4963 8384 4993
rect 8515 4993 8549 5002
rect 8515 4968 8516 4993
rect 8516 4968 8549 4993
rect 8688 4993 8722 5006
rect 8688 4972 8718 4993
rect 8718 4972 8722 4993
rect 8851 4993 8885 5001
rect 8851 4967 8852 4993
rect 8852 4967 8885 4993
rect 6318 4866 6352 4900
rect 6426 4866 6460 4900
rect 6534 4897 6568 4900
rect 6534 4866 6549 4897
rect 6549 4866 6568 4897
rect 6642 4866 6676 4900
rect 6750 4897 6784 4900
rect 6750 4866 6752 4897
rect 6752 4866 6784 4897
rect 6858 4897 6892 4900
rect 6858 4866 6886 4897
rect 6886 4866 6892 4897
rect 6966 4866 7000 4900
rect 7074 4897 7108 4900
rect 7074 4866 7094 4897
rect 7094 4866 7108 4897
rect 20901 4995 20935 4996
rect 20901 4962 20926 4995
rect 20926 4962 20935 4995
rect 21060 4995 21094 4998
rect 21060 4964 21094 4995
rect 21230 4995 21264 5000
rect 21230 4966 21262 4995
rect 21262 4966 21264 4995
rect 21400 4995 21434 5006
rect 21400 4972 21430 4995
rect 21430 4972 21434 4995
rect 21564 4961 21598 4993
rect 21733 4995 21767 5003
rect 21733 4969 21766 4995
rect 21766 4969 21767 4995
rect 21900 4995 21934 4997
rect 21900 4963 21934 4995
rect 22060 4995 22094 4997
rect 22060 4963 22068 4995
rect 22068 4963 22094 4995
rect 21564 4959 21598 4961
rect 22673 5173 22707 5207
rect 22765 5173 22799 5207
rect 22857 5173 22891 5207
rect 22949 5173 22983 5207
rect 23041 5173 23075 5207
rect 23133 5173 23167 5207
rect 23225 5173 23259 5207
rect 23317 5173 23351 5207
rect 23409 5173 23443 5207
rect 23501 5173 23535 5207
rect 23593 5173 23627 5207
rect 23685 5173 23719 5207
rect 23777 5173 23811 5207
rect 23869 5173 23903 5207
rect 23961 5173 23995 5207
rect 24053 5173 24087 5207
rect 35895 5175 35929 5209
rect 35987 5175 36021 5209
rect 36079 5175 36113 5209
rect 36171 5175 36205 5209
rect 36263 5175 36297 5209
rect 36355 5175 36389 5209
rect 36447 5175 36481 5209
rect 36539 5175 36573 5209
rect 36631 5175 36665 5209
rect 36723 5175 36757 5209
rect 36815 5175 36849 5209
rect 36907 5175 36941 5209
rect 36999 5175 37033 5209
rect 37091 5175 37125 5209
rect 37183 5175 37217 5209
rect 37275 5175 37309 5209
rect 7930 4895 7964 4900
rect 7930 4866 7963 4895
rect 7963 4866 7964 4895
rect 8081 4895 8115 4900
rect 8081 4866 8096 4895
rect 8096 4866 8115 4895
rect 8178 4866 8212 4900
rect 8275 4895 8309 4900
rect 8275 4866 8298 4895
rect 8298 4866 8309 4895
rect 8372 4866 8406 4900
rect 8469 4866 8503 4900
rect 8566 4866 8600 4900
rect 8663 4866 8697 4900
rect 8760 4895 8794 4900
rect 8760 4866 8768 4895
rect 8768 4866 8794 4895
rect 22774 4993 22808 4994
rect 22774 4960 22808 4993
rect 22944 4993 22978 4996
rect 22944 4962 22976 4993
rect 22976 4962 22978 4993
rect 23110 4993 23144 5002
rect 23110 4968 23144 4993
rect 23279 4993 23313 5001
rect 23279 4967 23312 4993
rect 23312 4967 23313 4993
rect 23448 4993 23482 4997
rect 23448 4963 23480 4993
rect 23480 4963 23482 4993
rect 23619 4993 23653 4999
rect 23619 4965 23648 4993
rect 23648 4965 23653 4993
rect 23783 4993 23817 4997
rect 23783 4963 23816 4993
rect 23816 4963 23817 4993
rect 23949 4993 23983 4995
rect 23949 4961 23950 4993
rect 23950 4961 23983 4993
rect 21458 4897 21492 4900
rect 21458 4866 21480 4897
rect 21480 4866 21492 4897
rect 21577 4866 21611 4900
rect 21696 4866 21730 4900
rect 21815 4897 21849 4900
rect 21815 4866 21816 4897
rect 21816 4866 21849 4897
rect 21934 4866 21968 4900
rect 22053 4866 22087 4900
rect 22172 4897 22206 4900
rect 22172 4866 22192 4897
rect 22192 4866 22206 4897
rect 5693 4631 5727 4665
rect 5785 4631 5819 4665
rect 5877 4631 5911 4665
rect 5969 4631 6003 4665
rect 6061 4631 6095 4665
rect 6153 4631 6187 4665
rect 6245 4631 6279 4665
rect 6337 4631 6371 4665
rect 6429 4631 6463 4665
rect 6521 4631 6555 4665
rect 6613 4631 6647 4665
rect 6705 4631 6739 4665
rect 6797 4631 6831 4665
rect 6889 4631 6923 4665
rect 6981 4631 7015 4665
rect 7073 4631 7107 4665
rect 36001 4995 36035 5005
rect 36001 4971 36030 4995
rect 36030 4971 36035 4995
rect 36164 4995 36198 5009
rect 36164 4975 36198 4995
rect 36334 4995 36368 5007
rect 36334 4973 36366 4995
rect 36366 4973 36368 4995
rect 36499 4995 36533 5007
rect 36499 4973 36500 4995
rect 36500 4973 36533 4995
rect 36668 4961 36702 4993
rect 36839 4995 36873 4996
rect 36839 4962 36870 4995
rect 36870 4962 36873 4995
rect 37001 4995 37035 5001
rect 37001 4967 37004 4995
rect 37004 4967 37035 4995
rect 37174 4995 37208 5002
rect 37174 4968 37206 4995
rect 37206 4968 37208 4995
rect 36668 4959 36702 4961
rect 37777 5173 37811 5207
rect 37869 5173 37903 5207
rect 37961 5173 37995 5207
rect 38053 5173 38087 5207
rect 38145 5173 38179 5207
rect 38237 5173 38271 5207
rect 38329 5173 38363 5207
rect 38421 5173 38455 5207
rect 38513 5173 38547 5207
rect 38605 5173 38639 5207
rect 38697 5173 38731 5207
rect 38789 5173 38823 5207
rect 38881 5173 38915 5207
rect 38973 5173 39007 5207
rect 39065 5173 39099 5207
rect 39157 5173 39191 5207
rect 50993 5175 51027 5209
rect 51085 5175 51119 5209
rect 51177 5175 51211 5209
rect 51269 5175 51303 5209
rect 51361 5175 51395 5209
rect 51453 5175 51487 5209
rect 51545 5175 51579 5209
rect 51637 5175 51671 5209
rect 51729 5175 51763 5209
rect 51821 5175 51855 5209
rect 51913 5175 51947 5209
rect 52005 5175 52039 5209
rect 52097 5175 52131 5209
rect 52189 5175 52223 5209
rect 52281 5175 52315 5209
rect 52373 5175 52407 5209
rect 23028 4895 23062 4900
rect 23028 4866 23061 4895
rect 23061 4866 23062 4895
rect 23132 4866 23166 4900
rect 23248 4866 23282 4900
rect 23361 4895 23395 4900
rect 23361 4866 23362 4895
rect 23362 4866 23395 4895
rect 23474 4866 23508 4900
rect 23587 4866 23621 4900
rect 23700 4895 23734 4900
rect 23700 4866 23732 4895
rect 23732 4866 23734 4895
rect 23813 4866 23847 4900
rect 23926 4866 23960 4900
rect 38047 4993 38081 5003
rect 38047 4969 38080 4993
rect 38080 4969 38081 4993
rect 38217 4993 38251 5012
rect 38217 4978 38248 4993
rect 38248 4978 38251 4993
rect 38385 4993 38419 5010
rect 38385 4976 38416 4993
rect 38416 4976 38419 4993
rect 38552 4993 38586 4997
rect 38552 4963 38584 4993
rect 38584 4963 38586 4993
rect 38717 4993 38751 5002
rect 38717 4968 38718 4993
rect 38718 4968 38751 4993
rect 38890 4993 38924 5006
rect 38890 4972 38920 4993
rect 38920 4972 38924 4993
rect 39053 4993 39087 5001
rect 39053 4967 39054 4993
rect 39054 4967 39087 4993
rect 36520 4866 36554 4900
rect 36628 4866 36662 4900
rect 36736 4897 36770 4900
rect 36736 4866 36751 4897
rect 36751 4866 36770 4897
rect 36844 4866 36878 4900
rect 36952 4897 36986 4900
rect 36952 4866 36954 4897
rect 36954 4866 36986 4897
rect 37060 4897 37094 4900
rect 37060 4866 37088 4897
rect 37088 4866 37094 4897
rect 37168 4866 37202 4900
rect 37276 4897 37310 4900
rect 37276 4866 37296 4897
rect 37296 4866 37310 4897
rect 7575 4629 7609 4663
rect 7667 4629 7701 4663
rect 7759 4629 7793 4663
rect 7851 4629 7885 4663
rect 7943 4629 7977 4663
rect 8035 4629 8069 4663
rect 8127 4629 8161 4663
rect 8219 4629 8253 4663
rect 8311 4629 8345 4663
rect 8403 4629 8437 4663
rect 8495 4629 8529 4663
rect 8587 4629 8621 4663
rect 8679 4629 8713 4663
rect 8771 4629 8805 4663
rect 8863 4629 8897 4663
rect 8955 4629 8989 4663
rect 20791 4631 20825 4665
rect 20883 4631 20917 4665
rect 20975 4631 21009 4665
rect 21067 4631 21101 4665
rect 21159 4631 21193 4665
rect 21251 4631 21285 4665
rect 21343 4631 21377 4665
rect 21435 4631 21469 4665
rect 21527 4631 21561 4665
rect 21619 4631 21653 4665
rect 21711 4631 21745 4665
rect 21803 4631 21837 4665
rect 21895 4631 21929 4665
rect 21987 4631 22021 4665
rect 22079 4631 22113 4665
rect 22171 4631 22205 4665
rect 51103 4995 51137 4996
rect 51103 4962 51128 4995
rect 51128 4962 51137 4995
rect 51262 4995 51296 4998
rect 51262 4964 51296 4995
rect 51432 4995 51466 5000
rect 51432 4966 51464 4995
rect 51464 4966 51466 4995
rect 51602 4995 51636 5006
rect 51602 4972 51632 4995
rect 51632 4972 51636 4995
rect 51766 4961 51800 4993
rect 51935 4995 51969 5003
rect 51935 4969 51968 4995
rect 51968 4969 51969 4995
rect 52102 4995 52136 4997
rect 52102 4963 52136 4995
rect 52262 4995 52296 4997
rect 52262 4963 52270 4995
rect 52270 4963 52296 4995
rect 51766 4959 51800 4961
rect 52875 5173 52909 5207
rect 52967 5173 53001 5207
rect 53059 5173 53093 5207
rect 53151 5173 53185 5207
rect 53243 5173 53277 5207
rect 53335 5173 53369 5207
rect 53427 5173 53461 5207
rect 53519 5173 53553 5207
rect 53611 5173 53645 5207
rect 53703 5173 53737 5207
rect 53795 5173 53829 5207
rect 53887 5173 53921 5207
rect 53979 5173 54013 5207
rect 54071 5173 54105 5207
rect 54163 5173 54197 5207
rect 54255 5173 54289 5207
rect 38132 4895 38166 4900
rect 38132 4866 38165 4895
rect 38165 4866 38166 4895
rect 38283 4895 38317 4900
rect 38283 4866 38298 4895
rect 38298 4866 38317 4895
rect 38380 4866 38414 4900
rect 38477 4895 38511 4900
rect 38477 4866 38500 4895
rect 38500 4866 38511 4895
rect 38574 4866 38608 4900
rect 38671 4866 38705 4900
rect 38768 4866 38802 4900
rect 38865 4866 38899 4900
rect 38962 4895 38996 4900
rect 38962 4866 38970 4895
rect 38970 4866 38996 4895
rect 52976 4993 53010 4994
rect 52976 4960 53010 4993
rect 53146 4993 53180 4996
rect 53146 4962 53178 4993
rect 53178 4962 53180 4993
rect 53312 4993 53346 5002
rect 53312 4968 53346 4993
rect 53481 4993 53515 5001
rect 53481 4967 53514 4993
rect 53514 4967 53515 4993
rect 53650 4993 53684 4997
rect 53650 4963 53682 4993
rect 53682 4963 53684 4993
rect 53821 4993 53855 4999
rect 53821 4965 53850 4993
rect 53850 4965 53855 4993
rect 53985 4993 54019 4997
rect 53985 4963 54018 4993
rect 54018 4963 54019 4993
rect 54151 4993 54185 4995
rect 54151 4961 54152 4993
rect 54152 4961 54185 4993
rect 51660 4897 51694 4900
rect 51660 4866 51682 4897
rect 51682 4866 51694 4897
rect 51779 4866 51813 4900
rect 51898 4866 51932 4900
rect 52017 4897 52051 4900
rect 52017 4866 52018 4897
rect 52018 4866 52051 4897
rect 52136 4866 52170 4900
rect 52255 4866 52289 4900
rect 52374 4897 52408 4900
rect 52374 4866 52394 4897
rect 52394 4866 52408 4897
rect 22673 4629 22707 4663
rect 22765 4629 22799 4663
rect 22857 4629 22891 4663
rect 22949 4629 22983 4663
rect 23041 4629 23075 4663
rect 23133 4629 23167 4663
rect 23225 4629 23259 4663
rect 23317 4629 23351 4663
rect 23409 4629 23443 4663
rect 23501 4629 23535 4663
rect 23593 4629 23627 4663
rect 23685 4629 23719 4663
rect 23777 4629 23811 4663
rect 23869 4629 23903 4663
rect 23961 4629 23995 4663
rect 24053 4629 24087 4663
rect 35895 4631 35929 4665
rect 35987 4631 36021 4665
rect 36079 4631 36113 4665
rect 36171 4631 36205 4665
rect 36263 4631 36297 4665
rect 36355 4631 36389 4665
rect 36447 4631 36481 4665
rect 36539 4631 36573 4665
rect 36631 4631 36665 4665
rect 36723 4631 36757 4665
rect 36815 4631 36849 4665
rect 36907 4631 36941 4665
rect 36999 4631 37033 4665
rect 37091 4631 37125 4665
rect 37183 4631 37217 4665
rect 37275 4631 37309 4665
rect 53230 4895 53264 4900
rect 53230 4866 53263 4895
rect 53263 4866 53264 4895
rect 53334 4866 53368 4900
rect 53450 4866 53484 4900
rect 53563 4895 53597 4900
rect 53563 4866 53564 4895
rect 53564 4866 53597 4895
rect 53676 4866 53710 4900
rect 53789 4866 53823 4900
rect 53902 4895 53936 4900
rect 53902 4866 53934 4895
rect 53934 4866 53936 4895
rect 54015 4866 54049 4900
rect 54128 4866 54162 4900
rect 37777 4629 37811 4663
rect 37869 4629 37903 4663
rect 37961 4629 37995 4663
rect 38053 4629 38087 4663
rect 38145 4629 38179 4663
rect 38237 4629 38271 4663
rect 38329 4629 38363 4663
rect 38421 4629 38455 4663
rect 38513 4629 38547 4663
rect 38605 4629 38639 4663
rect 38697 4629 38731 4663
rect 38789 4629 38823 4663
rect 38881 4629 38915 4663
rect 38973 4629 39007 4663
rect 39065 4629 39099 4663
rect 39157 4629 39191 4663
rect 50993 4631 51027 4665
rect 51085 4631 51119 4665
rect 51177 4631 51211 4665
rect 51269 4631 51303 4665
rect 51361 4631 51395 4665
rect 51453 4631 51487 4665
rect 51545 4631 51579 4665
rect 51637 4631 51671 4665
rect 51729 4631 51763 4665
rect 51821 4631 51855 4665
rect 51913 4631 51947 4665
rect 52005 4631 52039 4665
rect 52097 4631 52131 4665
rect 52189 4631 52223 4665
rect 52281 4631 52315 4665
rect 52373 4631 52407 4665
rect 52875 4629 52909 4663
rect 52967 4629 53001 4663
rect 53059 4629 53093 4663
rect 53151 4629 53185 4663
rect 53243 4629 53277 4663
rect 53335 4629 53369 4663
rect 53427 4629 53461 4663
rect 53519 4629 53553 4663
rect 53611 4629 53645 4663
rect 53703 4629 53737 4663
rect 53795 4629 53829 4663
rect 53887 4629 53921 4663
rect 53979 4629 54013 4663
rect 54071 4629 54105 4663
rect 54163 4629 54197 4663
rect 54255 4629 54289 4663
rect 30056 4098 30090 4132
rect 30148 4098 30182 4132
rect 30240 4098 30274 4132
rect 30332 4098 30366 4132
rect 30424 4098 30458 4132
rect 30584 4098 30618 4132
rect 30676 4098 30710 4132
rect 30768 4098 30802 4132
rect 30860 4098 30894 4132
rect 30952 4098 30986 4132
rect 31044 4098 31078 4132
rect 31136 4098 31170 4132
rect 31228 4098 31262 4132
rect 31320 4098 31354 4132
rect 31412 4098 31446 4132
rect 31504 4098 31538 4132
rect 31596 4098 31630 4132
rect 31688 4098 31722 4132
rect 31780 4098 31814 4132
rect 31872 4098 31906 4132
rect 31964 4098 31998 4132
rect 43410 3882 43444 3916
rect 43502 3882 43536 3916
rect 43594 3882 43628 3916
rect 43686 3882 43720 3916
rect 43778 3882 43812 3916
rect 43870 3882 43904 3916
rect 43962 3882 43996 3916
rect 44054 3882 44088 3916
rect 44146 3882 44180 3916
rect 44238 3882 44272 3916
rect 44330 3882 44364 3916
rect 44422 3882 44456 3916
rect 44514 3882 44548 3916
rect 44606 3882 44640 3916
rect 44698 3882 44732 3916
rect 44790 3882 44824 3916
rect 45340 3882 45374 3916
rect 45432 3882 45466 3916
rect 45524 3882 45558 3916
rect 45616 3882 45650 3916
rect 45708 3882 45742 3916
rect 45800 3882 45834 3916
rect 45892 3882 45926 3916
rect 45984 3882 46018 3916
rect 46076 3882 46110 3916
rect 46168 3882 46202 3916
rect 46260 3882 46294 3916
rect 46352 3882 46386 3916
rect 46444 3882 46478 3916
rect 46536 3882 46570 3916
rect 46628 3882 46662 3916
rect 46720 3882 46754 3916
rect 30423 3828 30457 3862
rect 30606 3820 30640 3826
rect 30606 3792 30631 3820
rect 30631 3792 30640 3820
rect 30694 3792 30728 3826
rect 30782 3820 30816 3826
rect 30782 3792 30805 3820
rect 30805 3792 30816 3820
rect 30870 3792 30904 3826
rect 30958 3820 30992 3826
rect 30958 3792 30973 3820
rect 30973 3792 30992 3820
rect 31046 3792 31080 3826
rect 31134 3820 31168 3826
rect 31134 3792 31142 3820
rect 31142 3792 31168 3820
rect 31222 3792 31256 3826
rect 31310 3792 31344 3826
rect 13268 3722 13302 3756
rect 13360 3722 13394 3756
rect 13452 3722 13486 3756
rect 13544 3722 13578 3756
rect 13636 3722 13670 3756
rect 13728 3722 13762 3756
rect 13820 3722 13854 3756
rect 13912 3722 13946 3756
rect 14004 3722 14038 3756
rect 14096 3722 14130 3756
rect 14188 3722 14222 3756
rect 14280 3722 14314 3756
rect 14372 3722 14406 3756
rect 14464 3722 14498 3756
rect 14556 3722 14590 3756
rect 14648 3722 14682 3756
rect 15198 3722 15232 3756
rect 15290 3722 15324 3756
rect 15382 3722 15416 3756
rect 15474 3722 15508 3756
rect 15566 3722 15600 3756
rect 15658 3722 15692 3756
rect 15750 3722 15784 3756
rect 15842 3722 15876 3756
rect 15934 3722 15968 3756
rect 16026 3722 16060 3756
rect 16118 3722 16152 3756
rect 16210 3722 16244 3756
rect 16302 3722 16336 3756
rect 16394 3722 16428 3756
rect 16486 3722 16520 3756
rect 16578 3722 16612 3756
rect 30423 3748 30457 3782
rect 13372 3542 13406 3554
rect 13372 3509 13405 3542
rect 13405 3509 13406 3542
rect 13540 3542 13574 3561
rect 13540 3516 13573 3542
rect 13573 3516 13574 3542
rect 13708 3542 13742 3551
rect 13708 3508 13741 3542
rect 13741 3508 13742 3542
rect 13876 3542 13910 3563
rect 13876 3518 13909 3542
rect 13909 3518 13910 3542
rect 14042 3542 14076 3561
rect 14042 3516 14043 3542
rect 14043 3516 14076 3542
rect 14208 3542 14242 3563
rect 14208 3518 14211 3542
rect 14211 3518 14242 3542
rect 14376 3542 14410 3563
rect 14376 3518 14379 3542
rect 14379 3518 14410 3542
rect 14550 3542 14584 3561
rect 14550 3516 14581 3542
rect 14581 3516 14584 3542
rect 13708 3506 13742 3508
rect 13572 3418 13606 3452
rect 13672 3418 13706 3452
rect 13772 3444 13806 3452
rect 13772 3418 13792 3444
rect 13792 3418 13806 3444
rect 13872 3418 13906 3452
rect 13972 3444 14006 3452
rect 13972 3418 13993 3444
rect 13993 3418 14006 3444
rect 14072 3418 14106 3452
rect 14172 3418 14206 3452
rect 14272 3444 14306 3452
rect 14272 3418 14294 3444
rect 14294 3418 14306 3444
rect 15306 3542 15340 3555
rect 15306 3510 15335 3542
rect 15335 3510 15340 3542
rect 15468 3542 15502 3559
rect 15468 3514 15469 3542
rect 15469 3514 15502 3542
rect 15638 3542 15672 3563
rect 15638 3518 15671 3542
rect 15671 3518 15672 3542
rect 15802 3542 15836 3559
rect 15802 3514 15805 3542
rect 15805 3514 15836 3542
rect 15972 3542 16006 3559
rect 15972 3514 15973 3542
rect 15973 3514 16006 3542
rect 16140 3542 16174 3555
rect 16140 3510 16141 3542
rect 16141 3510 16174 3542
rect 16308 3542 16342 3559
rect 16308 3514 16309 3542
rect 16309 3514 16342 3542
rect 31029 3698 31057 3724
rect 31057 3698 31063 3724
rect 31029 3690 31063 3698
rect 31195 3698 31225 3720
rect 31225 3698 31229 3720
rect 31195 3686 31229 3698
rect 31363 3698 31393 3726
rect 31393 3698 31397 3726
rect 31363 3692 31397 3698
rect 31530 3698 31561 3724
rect 31561 3698 31564 3724
rect 31530 3690 31564 3698
rect 31700 3698 31729 3725
rect 31729 3698 31734 3725
rect 31700 3691 31734 3698
rect 31864 3698 31897 3726
rect 31897 3698 31898 3726
rect 31864 3692 31898 3698
rect 43514 3702 43548 3714
rect 43514 3669 43547 3702
rect 43547 3669 43548 3702
rect 43682 3702 43716 3721
rect 43682 3676 43715 3702
rect 43715 3676 43716 3702
rect 43850 3702 43884 3711
rect 43850 3668 43883 3702
rect 43883 3668 43884 3702
rect 44018 3702 44052 3723
rect 44018 3678 44051 3702
rect 44051 3678 44052 3702
rect 44184 3702 44218 3721
rect 44184 3676 44185 3702
rect 44185 3676 44218 3702
rect 44350 3702 44384 3723
rect 44350 3678 44353 3702
rect 44353 3678 44384 3702
rect 44518 3702 44552 3723
rect 44518 3678 44521 3702
rect 44521 3678 44552 3702
rect 44692 3702 44726 3721
rect 44692 3676 44723 3702
rect 44723 3676 44726 3702
rect 43850 3666 43884 3668
rect 16482 3542 16516 3555
rect 16482 3510 16511 3542
rect 16511 3510 16516 3542
rect 30056 3554 30090 3588
rect 30148 3554 30182 3588
rect 30240 3554 30274 3588
rect 30332 3554 30366 3588
rect 30424 3554 30458 3588
rect 30584 3554 30618 3588
rect 30676 3554 30710 3588
rect 30768 3554 30802 3588
rect 30860 3554 30894 3588
rect 30952 3554 30986 3588
rect 31044 3554 31078 3588
rect 31136 3554 31170 3588
rect 31228 3554 31262 3588
rect 31320 3554 31354 3588
rect 31412 3554 31446 3588
rect 31504 3554 31538 3588
rect 31596 3554 31630 3588
rect 31688 3554 31722 3588
rect 31780 3554 31814 3588
rect 31872 3554 31906 3588
rect 31964 3554 31998 3588
rect 43714 3578 43748 3612
rect 43814 3578 43848 3612
rect 43914 3604 43948 3612
rect 43914 3578 43934 3604
rect 43934 3578 43948 3604
rect 44014 3578 44048 3612
rect 44114 3604 44148 3612
rect 44114 3578 44135 3604
rect 44135 3578 44148 3604
rect 44214 3578 44248 3612
rect 44314 3578 44348 3612
rect 44414 3604 44448 3612
rect 44414 3578 44436 3604
rect 44436 3578 44448 3604
rect 45448 3702 45482 3715
rect 45448 3670 45477 3702
rect 45477 3670 45482 3702
rect 45610 3702 45644 3719
rect 45610 3674 45611 3702
rect 45611 3674 45644 3702
rect 45780 3702 45814 3723
rect 45780 3678 45813 3702
rect 45813 3678 45814 3702
rect 45944 3702 45978 3719
rect 45944 3674 45947 3702
rect 45947 3674 45978 3702
rect 46114 3702 46148 3719
rect 46114 3674 46115 3702
rect 46115 3674 46148 3702
rect 46282 3702 46316 3715
rect 46282 3670 46283 3702
rect 46283 3670 46316 3702
rect 46450 3702 46484 3719
rect 46450 3674 46451 3702
rect 46451 3674 46484 3702
rect 46624 3702 46658 3715
rect 46624 3670 46653 3702
rect 46653 3670 46658 3702
rect 45374 3604 45408 3612
rect 45374 3578 45387 3604
rect 45387 3578 45408 3604
rect 45474 3578 45508 3612
rect 45574 3578 45608 3612
rect 45674 3604 45708 3612
rect 45674 3578 45695 3604
rect 45695 3578 45708 3604
rect 45774 3578 45808 3612
rect 45874 3604 45908 3612
rect 45874 3578 45898 3604
rect 45898 3578 45908 3604
rect 45974 3578 46008 3612
rect 46074 3578 46108 3612
rect 15232 3444 15266 3452
rect 15232 3418 15245 3444
rect 15245 3418 15266 3444
rect 15332 3418 15366 3452
rect 15432 3418 15466 3452
rect 15532 3444 15566 3452
rect 15532 3418 15553 3444
rect 15553 3418 15566 3444
rect 15632 3418 15666 3452
rect 15732 3444 15766 3452
rect 15732 3418 15756 3444
rect 15756 3418 15766 3444
rect 15832 3418 15866 3452
rect 15932 3418 15966 3452
rect 43410 3338 43444 3372
rect 43502 3338 43536 3372
rect 43594 3338 43628 3372
rect 43686 3338 43720 3372
rect 43778 3338 43812 3372
rect 43870 3338 43904 3372
rect 43962 3338 43996 3372
rect 44054 3338 44088 3372
rect 44146 3338 44180 3372
rect 44238 3338 44272 3372
rect 44330 3338 44364 3372
rect 44422 3338 44456 3372
rect 44514 3338 44548 3372
rect 44606 3338 44640 3372
rect 44698 3338 44732 3372
rect 44790 3338 44824 3372
rect 45340 3338 45374 3372
rect 45432 3338 45466 3372
rect 45524 3338 45558 3372
rect 45616 3338 45650 3372
rect 45708 3338 45742 3372
rect 45800 3338 45834 3372
rect 45892 3338 45926 3372
rect 45984 3338 46018 3372
rect 46076 3338 46110 3372
rect 46168 3338 46202 3372
rect 46260 3338 46294 3372
rect 46352 3338 46386 3372
rect 46444 3338 46478 3372
rect 46536 3338 46570 3372
rect 46628 3338 46662 3372
rect 46720 3338 46754 3372
rect 13268 3178 13302 3212
rect 13360 3178 13394 3212
rect 13452 3178 13486 3212
rect 13544 3178 13578 3212
rect 13636 3178 13670 3212
rect 13728 3178 13762 3212
rect 13820 3178 13854 3212
rect 13912 3178 13946 3212
rect 14004 3178 14038 3212
rect 14096 3178 14130 3212
rect 14188 3178 14222 3212
rect 14280 3178 14314 3212
rect 14372 3178 14406 3212
rect 14464 3178 14498 3212
rect 14556 3178 14590 3212
rect 14648 3178 14682 3212
rect 15198 3178 15232 3212
rect 15290 3178 15324 3212
rect 15382 3178 15416 3212
rect 15474 3178 15508 3212
rect 15566 3178 15600 3212
rect 15658 3178 15692 3212
rect 15750 3178 15784 3212
rect 15842 3178 15876 3212
rect 15934 3178 15968 3212
rect 16026 3178 16060 3212
rect 16118 3178 16152 3212
rect 16210 3178 16244 3212
rect 16302 3178 16336 3212
rect 16394 3178 16428 3212
rect 16486 3178 16520 3212
rect 16578 3178 16612 3212
rect 5693 2777 5727 2811
rect 5785 2777 5819 2811
rect 5877 2777 5911 2811
rect 5969 2777 6003 2811
rect 6061 2777 6095 2811
rect 6153 2777 6187 2811
rect 6245 2777 6279 2811
rect 6337 2777 6371 2811
rect 6429 2777 6463 2811
rect 6521 2777 6555 2811
rect 6613 2777 6647 2811
rect 6705 2777 6739 2811
rect 6797 2777 6831 2811
rect 6889 2777 6923 2811
rect 6981 2777 7015 2811
rect 7073 2777 7107 2811
rect 7575 2775 7609 2809
rect 7667 2775 7701 2809
rect 7759 2775 7793 2809
rect 7851 2775 7885 2809
rect 7943 2775 7977 2809
rect 8035 2775 8069 2809
rect 8127 2775 8161 2809
rect 8219 2775 8253 2809
rect 8311 2775 8345 2809
rect 8403 2775 8437 2809
rect 8495 2775 8529 2809
rect 8587 2775 8621 2809
rect 8679 2775 8713 2809
rect 8771 2775 8805 2809
rect 8863 2775 8897 2809
rect 8955 2775 8989 2809
rect 20791 2777 20825 2811
rect 20883 2777 20917 2811
rect 20975 2777 21009 2811
rect 21067 2777 21101 2811
rect 21159 2777 21193 2811
rect 21251 2777 21285 2811
rect 21343 2777 21377 2811
rect 21435 2777 21469 2811
rect 21527 2777 21561 2811
rect 21619 2777 21653 2811
rect 21711 2777 21745 2811
rect 21803 2777 21837 2811
rect 21895 2777 21929 2811
rect 21987 2777 22021 2811
rect 22079 2777 22113 2811
rect 22171 2777 22205 2811
rect 5820 2540 5854 2574
rect 5933 2540 5967 2574
rect 6046 2545 6048 2574
rect 6048 2545 6080 2574
rect 6046 2540 6080 2545
rect 6159 2540 6193 2574
rect 6272 2540 6306 2574
rect 6385 2545 6418 2574
rect 6418 2545 6419 2574
rect 6385 2540 6419 2545
rect 6498 2540 6532 2574
rect 6614 2540 6648 2574
rect 6718 2545 6719 2574
rect 6719 2545 6752 2574
rect 6718 2540 6752 2545
rect 22673 2775 22707 2809
rect 22765 2775 22799 2809
rect 22857 2775 22891 2809
rect 22949 2775 22983 2809
rect 23041 2775 23075 2809
rect 23133 2775 23167 2809
rect 23225 2775 23259 2809
rect 23317 2775 23351 2809
rect 23409 2775 23443 2809
rect 23501 2775 23535 2809
rect 23593 2775 23627 2809
rect 23685 2775 23719 2809
rect 23777 2775 23811 2809
rect 23869 2775 23903 2809
rect 23961 2775 23995 2809
rect 24053 2775 24087 2809
rect 35895 2777 35929 2811
rect 35987 2777 36021 2811
rect 36079 2777 36113 2811
rect 36171 2777 36205 2811
rect 36263 2777 36297 2811
rect 36355 2777 36389 2811
rect 36447 2777 36481 2811
rect 36539 2777 36573 2811
rect 36631 2777 36665 2811
rect 36723 2777 36757 2811
rect 36815 2777 36849 2811
rect 36907 2777 36941 2811
rect 36999 2777 37033 2811
rect 37091 2777 37125 2811
rect 37183 2777 37217 2811
rect 37275 2777 37309 2811
rect 7574 2543 7588 2574
rect 7588 2543 7608 2574
rect 7574 2540 7608 2543
rect 7693 2540 7727 2574
rect 7812 2540 7846 2574
rect 7931 2543 7964 2574
rect 7964 2543 7965 2574
rect 7931 2540 7965 2543
rect 8050 2540 8084 2574
rect 8169 2540 8203 2574
rect 8288 2543 8300 2574
rect 8300 2543 8322 2574
rect 8288 2540 8322 2543
rect 5797 2447 5830 2479
rect 5830 2447 5831 2479
rect 5797 2445 5831 2447
rect 5963 2447 5964 2477
rect 5964 2447 5997 2477
rect 5963 2443 5997 2447
rect 6127 2447 6132 2475
rect 6132 2447 6161 2475
rect 6127 2441 6161 2447
rect 6298 2447 6300 2477
rect 6300 2447 6332 2477
rect 6298 2443 6332 2447
rect 6467 2447 6468 2473
rect 6468 2447 6501 2473
rect 6467 2439 6501 2447
rect 6636 2447 6670 2472
rect 6636 2438 6670 2447
rect 6802 2447 6804 2478
rect 6804 2447 6836 2478
rect 6802 2444 6836 2447
rect 6972 2447 7006 2480
rect 6972 2446 7006 2447
rect 20986 2545 21012 2574
rect 21012 2545 21020 2574
rect 20986 2540 21020 2545
rect 21083 2540 21117 2574
rect 21180 2540 21214 2574
rect 21277 2540 21311 2574
rect 21374 2540 21408 2574
rect 21471 2545 21482 2574
rect 21482 2545 21505 2574
rect 21471 2540 21505 2545
rect 21568 2540 21602 2574
rect 21665 2545 21684 2574
rect 21684 2545 21699 2574
rect 21665 2540 21699 2545
rect 21816 2545 21817 2574
rect 21817 2545 21850 2574
rect 21816 2540 21850 2545
rect 5693 2233 5727 2267
rect 5785 2233 5819 2267
rect 5877 2233 5911 2267
rect 5969 2233 6003 2267
rect 6061 2233 6095 2267
rect 6153 2233 6187 2267
rect 6245 2233 6279 2267
rect 6337 2233 6371 2267
rect 6429 2233 6463 2267
rect 6521 2233 6555 2267
rect 6613 2233 6647 2267
rect 6705 2233 6739 2267
rect 6797 2233 6831 2267
rect 6889 2233 6923 2267
rect 6981 2233 7015 2267
rect 7073 2233 7107 2267
rect 8182 2479 8216 2481
rect 7686 2445 7712 2477
rect 7712 2445 7720 2477
rect 7686 2443 7720 2445
rect 7846 2445 7880 2477
rect 7846 2443 7880 2445
rect 8013 2445 8014 2471
rect 8014 2445 8047 2471
rect 8013 2437 8047 2445
rect 8182 2447 8216 2479
rect 8346 2445 8350 2468
rect 8350 2445 8380 2468
rect 8346 2434 8380 2445
rect 8516 2445 8518 2474
rect 8518 2445 8550 2474
rect 8516 2440 8550 2445
rect 8686 2445 8720 2476
rect 8686 2442 8720 2445
rect 8845 2445 8854 2478
rect 8854 2445 8879 2478
rect 8845 2444 8879 2445
rect 37777 2775 37811 2809
rect 37869 2775 37903 2809
rect 37961 2775 37995 2809
rect 38053 2775 38087 2809
rect 38145 2775 38179 2809
rect 38237 2775 38271 2809
rect 38329 2775 38363 2809
rect 38421 2775 38455 2809
rect 38513 2775 38547 2809
rect 38605 2775 38639 2809
rect 38697 2775 38731 2809
rect 38789 2775 38823 2809
rect 38881 2775 38915 2809
rect 38973 2775 39007 2809
rect 39065 2775 39099 2809
rect 39157 2775 39191 2809
rect 50993 2777 51027 2811
rect 51085 2777 51119 2811
rect 51177 2777 51211 2811
rect 51269 2777 51303 2811
rect 51361 2777 51395 2811
rect 51453 2777 51487 2811
rect 51545 2777 51579 2811
rect 51637 2777 51671 2811
rect 51729 2777 51763 2811
rect 51821 2777 51855 2811
rect 51913 2777 51947 2811
rect 52005 2777 52039 2811
rect 52097 2777 52131 2811
rect 52189 2777 52223 2811
rect 52281 2777 52315 2811
rect 52373 2777 52407 2811
rect 22672 2543 22686 2574
rect 22686 2543 22706 2574
rect 22672 2540 22706 2543
rect 22780 2540 22814 2574
rect 22888 2543 22894 2574
rect 22894 2543 22922 2574
rect 22888 2540 22922 2543
rect 22996 2543 23028 2574
rect 23028 2543 23030 2574
rect 22996 2540 23030 2543
rect 23104 2540 23138 2574
rect 23212 2543 23231 2574
rect 23231 2543 23246 2574
rect 23212 2540 23246 2543
rect 23320 2540 23354 2574
rect 23428 2540 23462 2574
rect 20895 2447 20928 2473
rect 20928 2447 20929 2473
rect 20895 2439 20929 2447
rect 21058 2447 21062 2468
rect 21062 2447 21092 2468
rect 21058 2434 21092 2447
rect 21231 2447 21264 2472
rect 21264 2447 21265 2472
rect 21231 2438 21265 2447
rect 21396 2447 21398 2477
rect 21398 2447 21430 2477
rect 21396 2443 21430 2447
rect 21563 2447 21566 2464
rect 21566 2447 21597 2464
rect 21563 2430 21597 2447
rect 21731 2447 21734 2462
rect 21734 2447 21765 2462
rect 21731 2428 21765 2447
rect 21901 2447 21902 2471
rect 21902 2447 21935 2471
rect 21901 2437 21935 2447
rect 36022 2540 36056 2574
rect 36135 2540 36169 2574
rect 36248 2545 36250 2574
rect 36250 2545 36282 2574
rect 36248 2540 36282 2545
rect 36361 2540 36395 2574
rect 36474 2540 36508 2574
rect 36587 2545 36620 2574
rect 36620 2545 36621 2574
rect 36587 2540 36621 2545
rect 36700 2540 36734 2574
rect 36816 2540 36850 2574
rect 36920 2545 36921 2574
rect 36921 2545 36954 2574
rect 36920 2540 36954 2545
rect 7575 2231 7609 2265
rect 7667 2231 7701 2265
rect 7759 2231 7793 2265
rect 7851 2231 7885 2265
rect 7943 2231 7977 2265
rect 8035 2231 8069 2265
rect 8127 2231 8161 2265
rect 8219 2231 8253 2265
rect 8311 2231 8345 2265
rect 8403 2231 8437 2265
rect 8495 2231 8529 2265
rect 8587 2231 8621 2265
rect 8679 2231 8713 2265
rect 8771 2231 8805 2265
rect 8863 2231 8897 2265
rect 8955 2231 8989 2265
rect 20791 2233 20825 2267
rect 20883 2233 20917 2267
rect 20975 2233 21009 2267
rect 21067 2233 21101 2267
rect 21159 2233 21193 2267
rect 21251 2233 21285 2267
rect 21343 2233 21377 2267
rect 21435 2233 21469 2267
rect 21527 2233 21561 2267
rect 21619 2233 21653 2267
rect 21711 2233 21745 2267
rect 21803 2233 21837 2267
rect 21895 2233 21929 2267
rect 21987 2233 22021 2267
rect 22079 2233 22113 2267
rect 22171 2233 22205 2267
rect 23280 2479 23314 2481
rect 22774 2445 22776 2472
rect 22776 2445 22808 2472
rect 22774 2438 22808 2445
rect 22947 2445 22978 2473
rect 22978 2445 22981 2473
rect 22947 2439 22981 2445
rect 23109 2445 23112 2478
rect 23112 2445 23143 2478
rect 23109 2444 23143 2445
rect 23280 2447 23314 2479
rect 23449 2445 23482 2467
rect 23482 2445 23483 2467
rect 23449 2433 23483 2445
rect 23614 2445 23616 2467
rect 23616 2445 23648 2467
rect 23614 2433 23648 2445
rect 23784 2445 23818 2465
rect 23784 2431 23818 2445
rect 23947 2445 23952 2469
rect 23952 2445 23981 2469
rect 23947 2435 23981 2445
rect 52875 2775 52909 2809
rect 52967 2775 53001 2809
rect 53059 2775 53093 2809
rect 53151 2775 53185 2809
rect 53243 2775 53277 2809
rect 53335 2775 53369 2809
rect 53427 2775 53461 2809
rect 53519 2775 53553 2809
rect 53611 2775 53645 2809
rect 53703 2775 53737 2809
rect 53795 2775 53829 2809
rect 53887 2775 53921 2809
rect 53979 2775 54013 2809
rect 54071 2775 54105 2809
rect 54163 2775 54197 2809
rect 54255 2775 54289 2809
rect 37776 2543 37790 2574
rect 37790 2543 37810 2574
rect 37776 2540 37810 2543
rect 37895 2540 37929 2574
rect 38014 2540 38048 2574
rect 38133 2543 38166 2574
rect 38166 2543 38167 2574
rect 38133 2540 38167 2543
rect 38252 2540 38286 2574
rect 38371 2540 38405 2574
rect 38490 2543 38502 2574
rect 38502 2543 38524 2574
rect 38490 2540 38524 2543
rect 35999 2447 36032 2479
rect 36032 2447 36033 2479
rect 35999 2445 36033 2447
rect 36165 2447 36166 2477
rect 36166 2447 36199 2477
rect 36165 2443 36199 2447
rect 36329 2447 36334 2475
rect 36334 2447 36363 2475
rect 36329 2441 36363 2447
rect 36500 2447 36502 2477
rect 36502 2447 36534 2477
rect 36500 2443 36534 2447
rect 36669 2447 36670 2473
rect 36670 2447 36703 2473
rect 36669 2439 36703 2447
rect 36838 2447 36872 2472
rect 36838 2438 36872 2447
rect 37004 2447 37006 2478
rect 37006 2447 37038 2478
rect 37004 2444 37038 2447
rect 37174 2447 37208 2480
rect 37174 2446 37208 2447
rect 51188 2545 51214 2574
rect 51214 2545 51222 2574
rect 51188 2540 51222 2545
rect 51285 2540 51319 2574
rect 51382 2540 51416 2574
rect 51479 2540 51513 2574
rect 51576 2540 51610 2574
rect 51673 2545 51684 2574
rect 51684 2545 51707 2574
rect 51673 2540 51707 2545
rect 51770 2540 51804 2574
rect 51867 2545 51886 2574
rect 51886 2545 51901 2574
rect 51867 2540 51901 2545
rect 52018 2545 52019 2574
rect 52019 2545 52052 2574
rect 52018 2540 52052 2545
rect 22673 2231 22707 2265
rect 22765 2231 22799 2265
rect 22857 2231 22891 2265
rect 22949 2231 22983 2265
rect 23041 2231 23075 2265
rect 23133 2231 23167 2265
rect 23225 2231 23259 2265
rect 23317 2231 23351 2265
rect 23409 2231 23443 2265
rect 23501 2231 23535 2265
rect 23593 2231 23627 2265
rect 23685 2231 23719 2265
rect 23777 2231 23811 2265
rect 23869 2231 23903 2265
rect 23961 2231 23995 2265
rect 24053 2231 24087 2265
rect 35895 2233 35929 2267
rect 35987 2233 36021 2267
rect 36079 2233 36113 2267
rect 36171 2233 36205 2267
rect 36263 2233 36297 2267
rect 36355 2233 36389 2267
rect 36447 2233 36481 2267
rect 36539 2233 36573 2267
rect 36631 2233 36665 2267
rect 36723 2233 36757 2267
rect 36815 2233 36849 2267
rect 36907 2233 36941 2267
rect 36999 2233 37033 2267
rect 37091 2233 37125 2267
rect 37183 2233 37217 2267
rect 37275 2233 37309 2267
rect 38384 2479 38418 2481
rect 37888 2445 37914 2477
rect 37914 2445 37922 2477
rect 37888 2443 37922 2445
rect 38048 2445 38082 2477
rect 38048 2443 38082 2445
rect 38215 2445 38216 2471
rect 38216 2445 38249 2471
rect 38215 2437 38249 2445
rect 38384 2447 38418 2479
rect 38548 2445 38552 2468
rect 38552 2445 38582 2468
rect 38548 2434 38582 2445
rect 38718 2445 38720 2474
rect 38720 2445 38752 2474
rect 38718 2440 38752 2445
rect 38888 2445 38922 2476
rect 38888 2442 38922 2445
rect 39047 2445 39056 2478
rect 39056 2445 39081 2478
rect 39047 2444 39081 2445
rect 52874 2543 52888 2574
rect 52888 2543 52908 2574
rect 52874 2540 52908 2543
rect 52982 2540 53016 2574
rect 53090 2543 53096 2574
rect 53096 2543 53124 2574
rect 53090 2540 53124 2543
rect 53198 2543 53230 2574
rect 53230 2543 53232 2574
rect 53198 2540 53232 2543
rect 53306 2540 53340 2574
rect 53414 2543 53433 2574
rect 53433 2543 53448 2574
rect 53414 2540 53448 2543
rect 53522 2540 53556 2574
rect 53630 2540 53664 2574
rect 51097 2447 51130 2473
rect 51130 2447 51131 2473
rect 51097 2439 51131 2447
rect 51260 2447 51264 2468
rect 51264 2447 51294 2468
rect 51260 2434 51294 2447
rect 51433 2447 51466 2472
rect 51466 2447 51467 2472
rect 51433 2438 51467 2447
rect 51598 2447 51600 2477
rect 51600 2447 51632 2477
rect 51598 2443 51632 2447
rect 51765 2447 51768 2464
rect 51768 2447 51799 2464
rect 51765 2430 51799 2447
rect 51933 2447 51936 2462
rect 51936 2447 51967 2462
rect 51933 2428 51967 2447
rect 52103 2447 52104 2471
rect 52104 2447 52137 2471
rect 52103 2437 52137 2447
rect 37777 2231 37811 2265
rect 37869 2231 37903 2265
rect 37961 2231 37995 2265
rect 38053 2231 38087 2265
rect 38145 2231 38179 2265
rect 38237 2231 38271 2265
rect 38329 2231 38363 2265
rect 38421 2231 38455 2265
rect 38513 2231 38547 2265
rect 38605 2231 38639 2265
rect 38697 2231 38731 2265
rect 38789 2231 38823 2265
rect 38881 2231 38915 2265
rect 38973 2231 39007 2265
rect 39065 2231 39099 2265
rect 39157 2231 39191 2265
rect 50993 2233 51027 2267
rect 51085 2233 51119 2267
rect 51177 2233 51211 2267
rect 51269 2233 51303 2267
rect 51361 2233 51395 2267
rect 51453 2233 51487 2267
rect 51545 2233 51579 2267
rect 51637 2233 51671 2267
rect 51729 2233 51763 2267
rect 51821 2233 51855 2267
rect 51913 2233 51947 2267
rect 52005 2233 52039 2267
rect 52097 2233 52131 2267
rect 52189 2233 52223 2267
rect 52281 2233 52315 2267
rect 52373 2233 52407 2267
rect 53482 2479 53516 2481
rect 52976 2445 52978 2472
rect 52978 2445 53010 2472
rect 52976 2438 53010 2445
rect 53149 2445 53180 2473
rect 53180 2445 53183 2473
rect 53149 2439 53183 2445
rect 53311 2445 53314 2478
rect 53314 2445 53345 2478
rect 53311 2444 53345 2445
rect 53482 2447 53516 2479
rect 53651 2445 53684 2467
rect 53684 2445 53685 2467
rect 53651 2433 53685 2445
rect 53816 2445 53818 2467
rect 53818 2445 53850 2467
rect 53816 2433 53850 2445
rect 53986 2445 54020 2465
rect 53986 2431 54020 2445
rect 54149 2445 54154 2469
rect 54154 2445 54183 2469
rect 54149 2435 54183 2445
rect 52875 2231 52909 2265
rect 52967 2231 53001 2265
rect 53059 2231 53093 2265
rect 53151 2231 53185 2265
rect 53243 2231 53277 2265
rect 53335 2231 53369 2265
rect 53427 2231 53461 2265
rect 53519 2231 53553 2265
rect 53611 2231 53645 2265
rect 53703 2231 53737 2265
rect 53795 2231 53829 2265
rect 53887 2231 53921 2265
rect 53979 2231 54013 2265
rect 54071 2231 54105 2265
rect 54163 2231 54197 2265
rect 54255 2231 54289 2265
rect 247 2153 281 2187
rect 339 2153 373 2187
rect 431 2153 465 2187
rect 1061 2153 1095 2187
rect 1153 2153 1187 2187
rect 1245 2153 1279 2187
rect 2135 2153 2169 2187
rect 2227 2153 2261 2187
rect 2319 2153 2353 2187
rect 2949 2153 2983 2187
rect 3041 2153 3075 2187
rect 3133 2153 3167 2187
rect 4023 2153 4057 2187
rect 4115 2153 4149 2187
rect 4207 2153 4241 2187
rect 4837 2153 4871 2187
rect 4929 2153 4963 2187
rect 5021 2153 5055 2187
rect 5911 2153 5945 2187
rect 6003 2153 6037 2187
rect 6095 2153 6129 2187
rect 6725 2153 6759 2187
rect 6817 2153 6851 2187
rect 6909 2153 6943 2187
rect 7799 2153 7833 2187
rect 7891 2153 7925 2187
rect 7983 2153 8017 2187
rect 8613 2153 8647 2187
rect 8705 2153 8739 2187
rect 8797 2153 8831 2187
rect 9687 2153 9721 2187
rect 9779 2153 9813 2187
rect 9871 2153 9905 2187
rect 10501 2153 10535 2187
rect 10593 2153 10627 2187
rect 10685 2153 10719 2187
rect 11575 2153 11609 2187
rect 11667 2153 11701 2187
rect 11759 2153 11793 2187
rect 12389 2153 12423 2187
rect 12481 2153 12515 2187
rect 12573 2153 12607 2187
rect 13463 2153 13497 2187
rect 13555 2153 13589 2187
rect 13647 2153 13681 2187
rect 14277 2153 14311 2187
rect 14369 2153 14403 2187
rect 14461 2153 14495 2187
rect 15345 2153 15379 2187
rect 15437 2153 15471 2187
rect 15529 2153 15563 2187
rect 16159 2153 16193 2187
rect 16251 2153 16285 2187
rect 16343 2153 16377 2187
rect 17233 2153 17267 2187
rect 17325 2153 17359 2187
rect 17417 2153 17451 2187
rect 18047 2153 18081 2187
rect 18139 2153 18173 2187
rect 18231 2153 18265 2187
rect 19121 2153 19155 2187
rect 19213 2153 19247 2187
rect 19305 2153 19339 2187
rect 19935 2153 19969 2187
rect 20027 2153 20061 2187
rect 20119 2153 20153 2187
rect 21009 2153 21043 2187
rect 21101 2153 21135 2187
rect 21193 2153 21227 2187
rect 21823 2153 21857 2187
rect 21915 2153 21949 2187
rect 22007 2153 22041 2187
rect 22897 2153 22931 2187
rect 22989 2153 23023 2187
rect 23081 2153 23115 2187
rect 23711 2153 23745 2187
rect 23803 2153 23837 2187
rect 23895 2153 23929 2187
rect 24785 2153 24819 2187
rect 24877 2153 24911 2187
rect 24969 2153 25003 2187
rect 25599 2153 25633 2187
rect 25691 2153 25725 2187
rect 25783 2153 25817 2187
rect 26673 2153 26707 2187
rect 26765 2153 26799 2187
rect 26857 2153 26891 2187
rect 27487 2153 27521 2187
rect 27579 2153 27613 2187
rect 27671 2153 27705 2187
rect 28561 2153 28595 2187
rect 28653 2153 28687 2187
rect 28745 2153 28779 2187
rect 29375 2153 29409 2187
rect 29467 2153 29501 2187
rect 29559 2153 29593 2187
rect 30449 2153 30483 2187
rect 30541 2153 30575 2187
rect 30633 2153 30667 2187
rect 31263 2153 31297 2187
rect 31355 2153 31389 2187
rect 31447 2153 31481 2187
rect 32337 2153 32371 2187
rect 32429 2153 32463 2187
rect 32521 2153 32555 2187
rect 33151 2153 33185 2187
rect 33243 2153 33277 2187
rect 33335 2153 33369 2187
rect 34225 2153 34259 2187
rect 34317 2153 34351 2187
rect 34409 2153 34443 2187
rect 35039 2153 35073 2187
rect 35131 2153 35165 2187
rect 35223 2153 35257 2187
rect 36113 2153 36147 2187
rect 36205 2153 36239 2187
rect 36297 2153 36331 2187
rect 36927 2153 36961 2187
rect 37019 2153 37053 2187
rect 37111 2153 37145 2187
rect 38001 2153 38035 2187
rect 38093 2153 38127 2187
rect 38185 2153 38219 2187
rect 38815 2153 38849 2187
rect 38907 2153 38941 2187
rect 38999 2153 39033 2187
rect 39889 2153 39923 2187
rect 39981 2153 40015 2187
rect 40073 2153 40107 2187
rect 40703 2153 40737 2187
rect 40795 2153 40829 2187
rect 40887 2153 40921 2187
rect 41777 2153 41811 2187
rect 41869 2153 41903 2187
rect 41961 2153 41995 2187
rect 42591 2153 42625 2187
rect 42683 2153 42717 2187
rect 42775 2153 42809 2187
rect 43665 2153 43699 2187
rect 43757 2153 43791 2187
rect 43849 2153 43883 2187
rect 44479 2153 44513 2187
rect 44571 2153 44605 2187
rect 44663 2153 44697 2187
rect 45547 2153 45581 2187
rect 45639 2153 45673 2187
rect 45731 2153 45765 2187
rect 46361 2153 46395 2187
rect 46453 2153 46487 2187
rect 46545 2153 46579 2187
rect 47435 2153 47469 2187
rect 47527 2153 47561 2187
rect 47619 2153 47653 2187
rect 48249 2153 48283 2187
rect 48341 2153 48375 2187
rect 48433 2153 48467 2187
rect 49323 2153 49357 2187
rect 49415 2153 49449 2187
rect 49507 2153 49541 2187
rect 50137 2153 50171 2187
rect 50229 2153 50263 2187
rect 50321 2153 50355 2187
rect 51211 2153 51245 2187
rect 51303 2153 51337 2187
rect 51395 2153 51429 2187
rect 52025 2153 52059 2187
rect 52117 2153 52151 2187
rect 52209 2153 52243 2187
rect 53099 2153 53133 2187
rect 53191 2153 53225 2187
rect 53283 2153 53317 2187
rect 53913 2153 53947 2187
rect 54005 2153 54039 2187
rect 54097 2153 54131 2187
rect 54987 2153 55021 2187
rect 55079 2153 55113 2187
rect 55171 2153 55205 2187
rect 55801 2153 55835 2187
rect 55893 2153 55927 2187
rect 55985 2153 56019 2187
rect 56875 2153 56909 2187
rect 56967 2153 57001 2187
rect 57059 2153 57093 2187
rect 57689 2153 57723 2187
rect 57781 2153 57815 2187
rect 57873 2153 57907 2187
rect 58763 2153 58797 2187
rect 58855 2153 58889 2187
rect 58947 2153 58981 2187
rect 59577 2153 59611 2187
rect 59669 2153 59703 2187
rect 59761 2153 59795 2187
rect 681 2113 715 2147
rect 750 2005 784 2039
rect 253 1875 287 1884
rect 253 1850 255 1875
rect 255 1850 287 1875
rect 426 1875 460 1880
rect 426 1846 457 1875
rect 457 1846 460 1875
rect 335 1755 337 1764
rect 337 1755 369 1764
rect 335 1730 369 1755
rect 247 1609 281 1643
rect 339 1609 373 1643
rect 431 1609 465 1643
rect 218 1364 252 1398
rect 606 1909 640 1911
rect 606 1877 640 1909
rect 606 1807 640 1839
rect 606 1805 640 1807
rect 702 1909 736 1911
rect 702 1877 736 1909
rect 702 1807 736 1839
rect 702 1805 736 1807
rect 2569 2113 2603 2147
rect 2638 2005 2672 2039
rect 798 1909 832 1911
rect 798 1877 832 1909
rect 1065 1875 1099 1882
rect 1065 1848 1069 1875
rect 1069 1848 1099 1875
rect 798 1807 832 1839
rect 798 1805 832 1807
rect 1239 1875 1273 1882
rect 1239 1848 1271 1875
rect 1271 1848 1273 1875
rect 2141 1875 2175 1884
rect 2141 1850 2143 1875
rect 2143 1850 2175 1875
rect 2314 1875 2348 1880
rect 2314 1846 2345 1875
rect 2345 1846 2348 1875
rect 654 1677 688 1711
rect 1153 1755 1185 1759
rect 1185 1755 1187 1759
rect 1153 1725 1187 1755
rect 2223 1755 2225 1764
rect 2225 1755 2257 1764
rect 2223 1730 2257 1755
rect 766 1596 800 1630
rect 1061 1609 1095 1643
rect 1153 1609 1187 1643
rect 1245 1609 1279 1643
rect 2135 1609 2169 1643
rect 2227 1609 2261 1643
rect 2319 1609 2353 1643
rect 622 1544 656 1546
rect 622 1512 656 1544
rect 622 1442 656 1474
rect 622 1440 656 1442
rect 718 1544 752 1546
rect 718 1512 752 1544
rect 718 1442 752 1474
rect 718 1440 752 1442
rect 814 1544 848 1546
rect 814 1512 848 1544
rect 814 1442 848 1474
rect 814 1440 848 1442
rect 670 1356 704 1390
rect 590 1247 624 1281
rect 1020 1230 1054 1264
rect 69 1099 103 1133
rect 161 1099 195 1133
rect 253 1099 287 1133
rect 432 1109 466 1143
rect 1078 1109 1112 1143
rect 118 821 152 832
rect 118 798 120 821
rect 120 798 152 821
rect 679 1057 713 1091
rect 2106 1364 2140 1398
rect 2494 1909 2528 1911
rect 2494 1877 2528 1909
rect 2494 1807 2528 1839
rect 2494 1805 2528 1807
rect 2590 1909 2624 1911
rect 2590 1877 2624 1909
rect 2590 1807 2624 1839
rect 2590 1805 2624 1807
rect 4457 2113 4491 2147
rect 4526 2005 4560 2039
rect 2686 1909 2720 1911
rect 2686 1877 2720 1909
rect 2953 1875 2987 1882
rect 2953 1848 2957 1875
rect 2957 1848 2987 1875
rect 2686 1807 2720 1839
rect 2686 1805 2720 1807
rect 3127 1875 3161 1882
rect 3127 1848 3159 1875
rect 3159 1848 3161 1875
rect 4029 1875 4063 1884
rect 4029 1850 4031 1875
rect 4031 1850 4063 1875
rect 4202 1875 4236 1880
rect 4202 1846 4233 1875
rect 4233 1846 4236 1875
rect 2542 1677 2576 1711
rect 3041 1755 3073 1759
rect 3073 1755 3075 1759
rect 3041 1725 3075 1755
rect 4111 1755 4113 1764
rect 4113 1755 4145 1764
rect 4111 1730 4145 1755
rect 2654 1596 2688 1630
rect 2949 1609 2983 1643
rect 3041 1609 3075 1643
rect 3133 1609 3167 1643
rect 4023 1609 4057 1643
rect 4115 1609 4149 1643
rect 4207 1609 4241 1643
rect 2510 1544 2544 1546
rect 2510 1512 2544 1544
rect 2510 1442 2544 1474
rect 2510 1440 2544 1442
rect 2606 1544 2640 1546
rect 2606 1512 2640 1544
rect 2606 1442 2640 1474
rect 2606 1440 2640 1442
rect 2702 1544 2736 1546
rect 2702 1512 2736 1544
rect 2702 1442 2736 1474
rect 2702 1440 2736 1442
rect 2558 1356 2592 1390
rect 2478 1247 2512 1281
rect 2908 1230 2942 1264
rect 1265 1107 1299 1141
rect 1357 1107 1391 1141
rect 1449 1107 1483 1141
rect 388 1013 422 1015
rect 388 981 422 1013
rect 388 911 422 943
rect 388 909 422 911
rect 476 1013 510 1015
rect 476 981 510 1013
rect 1034 1013 1068 1015
rect 748 949 782 983
rect 1034 981 1068 1013
rect 476 911 510 943
rect 476 909 510 911
rect 1034 911 1068 943
rect 1034 909 1068 911
rect 604 853 638 855
rect 604 821 638 853
rect 432 781 466 815
rect 604 751 638 783
rect 604 749 638 751
rect 700 853 734 855
rect 700 821 734 853
rect 700 751 734 783
rect 700 749 734 751
rect 1611 1105 1645 1139
rect 1703 1105 1737 1139
rect 1795 1105 1829 1139
rect 1122 1013 1156 1015
rect 1122 981 1156 1013
rect 1122 911 1156 943
rect 1122 909 1156 911
rect 1957 1099 1991 1133
rect 2049 1099 2083 1133
rect 2141 1099 2175 1133
rect 2320 1109 2354 1143
rect 796 853 830 855
rect 796 821 830 853
rect 796 751 830 783
rect 1078 781 1112 815
rect 796 749 830 751
rect 1617 793 1619 826
rect 1619 793 1651 826
rect 1617 792 1651 793
rect 2966 1109 3000 1143
rect 1810 804 1844 838
rect 652 621 686 655
rect 69 555 103 589
rect 161 555 195 589
rect 253 555 287 589
rect 404 550 438 584
rect 1036 578 1070 612
rect 1396 711 1430 728
rect 1396 694 1430 711
rect 2006 821 2040 832
rect 2006 798 2008 821
rect 2008 798 2040 821
rect 764 540 798 574
rect 1265 563 1299 597
rect 1357 563 1391 597
rect 1449 563 1483 597
rect 2567 1057 2601 1091
rect 3994 1364 4028 1398
rect 4382 1909 4416 1911
rect 4382 1877 4416 1909
rect 4382 1807 4416 1839
rect 4382 1805 4416 1807
rect 4478 1909 4512 1911
rect 4478 1877 4512 1909
rect 4478 1807 4512 1839
rect 4478 1805 4512 1807
rect 6345 2113 6379 2147
rect 6414 2005 6448 2039
rect 4574 1909 4608 1911
rect 4574 1877 4608 1909
rect 4841 1875 4875 1882
rect 4841 1848 4845 1875
rect 4845 1848 4875 1875
rect 4574 1807 4608 1839
rect 4574 1805 4608 1807
rect 5015 1875 5049 1882
rect 5015 1848 5047 1875
rect 5047 1848 5049 1875
rect 5917 1875 5951 1884
rect 5917 1850 5919 1875
rect 5919 1850 5951 1875
rect 6090 1875 6124 1880
rect 6090 1846 6121 1875
rect 6121 1846 6124 1875
rect 4430 1677 4464 1711
rect 4929 1755 4961 1759
rect 4961 1755 4963 1759
rect 4929 1725 4963 1755
rect 5999 1755 6001 1764
rect 6001 1755 6033 1764
rect 5999 1730 6033 1755
rect 4542 1596 4576 1630
rect 4837 1609 4871 1643
rect 4929 1609 4963 1643
rect 5021 1609 5055 1643
rect 5911 1609 5945 1643
rect 6003 1609 6037 1643
rect 6095 1609 6129 1643
rect 4398 1544 4432 1546
rect 4398 1512 4432 1544
rect 4398 1442 4432 1474
rect 4398 1440 4432 1442
rect 4494 1544 4528 1546
rect 4494 1512 4528 1544
rect 4494 1442 4528 1474
rect 4494 1440 4528 1442
rect 4590 1544 4624 1546
rect 4590 1512 4624 1544
rect 4590 1442 4624 1474
rect 4590 1440 4624 1442
rect 4446 1356 4480 1390
rect 4366 1247 4400 1281
rect 4796 1230 4830 1264
rect 3153 1107 3187 1141
rect 3245 1107 3279 1141
rect 3337 1107 3371 1141
rect 2276 1013 2310 1015
rect 2276 981 2310 1013
rect 2276 911 2310 943
rect 2276 909 2310 911
rect 2364 1013 2398 1015
rect 2364 981 2398 1013
rect 2922 1013 2956 1015
rect 2636 949 2670 983
rect 2922 981 2956 1013
rect 2364 911 2398 943
rect 2364 909 2398 911
rect 2922 911 2956 943
rect 2922 909 2956 911
rect 2492 853 2526 855
rect 2492 821 2526 853
rect 2320 781 2354 815
rect 1611 561 1645 595
rect 1703 561 1737 595
rect 1795 561 1829 595
rect 2492 751 2526 783
rect 2492 749 2526 751
rect 2588 853 2622 855
rect 2588 821 2622 853
rect 2588 751 2622 783
rect 2588 749 2622 751
rect 3499 1105 3533 1139
rect 3591 1105 3625 1139
rect 3683 1105 3717 1139
rect 3010 1013 3044 1015
rect 3010 981 3044 1013
rect 3010 911 3044 943
rect 3010 909 3044 911
rect 3845 1099 3879 1133
rect 3937 1099 3971 1133
rect 4029 1099 4063 1133
rect 4208 1109 4242 1143
rect 2684 853 2718 855
rect 2684 821 2718 853
rect 2684 751 2718 783
rect 2966 781 3000 815
rect 2684 749 2718 751
rect 3505 793 3507 826
rect 3507 793 3539 826
rect 3505 792 3539 793
rect 4854 1109 4888 1143
rect 3698 804 3732 838
rect 2540 621 2574 655
rect 1957 555 1991 589
rect 2049 555 2083 589
rect 2141 555 2175 589
rect 2292 550 2326 584
rect 2924 578 2958 612
rect 3284 711 3318 728
rect 3284 694 3318 711
rect 3894 821 3928 832
rect 3894 798 3896 821
rect 3896 798 3928 821
rect 620 488 654 490
rect 620 456 654 488
rect 716 488 750 490
rect 716 456 750 488
rect 620 386 654 418
rect 620 384 654 386
rect 716 386 750 418
rect 716 384 750 386
rect 812 488 846 490
rect 812 456 846 488
rect 2652 540 2686 574
rect 3153 563 3187 597
rect 3245 563 3279 597
rect 3337 563 3371 597
rect 4455 1057 4489 1091
rect 5882 1364 5916 1398
rect 6270 1909 6304 1911
rect 6270 1877 6304 1909
rect 6270 1807 6304 1839
rect 6270 1805 6304 1807
rect 6366 1909 6400 1911
rect 6366 1877 6400 1909
rect 6366 1807 6400 1839
rect 6366 1805 6400 1807
rect 8233 2113 8267 2147
rect 8302 2005 8336 2039
rect 6462 1909 6496 1911
rect 6462 1877 6496 1909
rect 6729 1875 6763 1882
rect 6729 1848 6733 1875
rect 6733 1848 6763 1875
rect 6462 1807 6496 1839
rect 6462 1805 6496 1807
rect 6903 1875 6937 1882
rect 6903 1848 6935 1875
rect 6935 1848 6937 1875
rect 7805 1875 7839 1884
rect 7805 1850 7807 1875
rect 7807 1850 7839 1875
rect 7978 1875 8012 1880
rect 7978 1846 8009 1875
rect 8009 1846 8012 1875
rect 6318 1677 6352 1711
rect 6817 1755 6849 1759
rect 6849 1755 6851 1759
rect 6817 1725 6851 1755
rect 7887 1755 7889 1764
rect 7889 1755 7921 1764
rect 7887 1730 7921 1755
rect 6430 1596 6464 1630
rect 6725 1609 6759 1643
rect 6817 1609 6851 1643
rect 6909 1609 6943 1643
rect 7799 1609 7833 1643
rect 7891 1609 7925 1643
rect 7983 1609 8017 1643
rect 6286 1544 6320 1546
rect 6286 1512 6320 1544
rect 6286 1442 6320 1474
rect 6286 1440 6320 1442
rect 6382 1544 6416 1546
rect 6382 1512 6416 1544
rect 6382 1442 6416 1474
rect 6382 1440 6416 1442
rect 6478 1544 6512 1546
rect 6478 1512 6512 1544
rect 6478 1442 6512 1474
rect 6478 1440 6512 1442
rect 6334 1356 6368 1390
rect 6254 1247 6288 1281
rect 6684 1230 6718 1264
rect 5041 1107 5075 1141
rect 5133 1107 5167 1141
rect 5225 1107 5259 1141
rect 4164 1013 4198 1015
rect 4164 981 4198 1013
rect 4164 911 4198 943
rect 4164 909 4198 911
rect 4252 1013 4286 1015
rect 4252 981 4286 1013
rect 4810 1013 4844 1015
rect 4524 949 4558 983
rect 4810 981 4844 1013
rect 4252 911 4286 943
rect 4252 909 4286 911
rect 4810 911 4844 943
rect 4810 909 4844 911
rect 4380 853 4414 855
rect 4380 821 4414 853
rect 4208 781 4242 815
rect 3499 561 3533 595
rect 3591 561 3625 595
rect 3683 561 3717 595
rect 4380 751 4414 783
rect 4380 749 4414 751
rect 4476 853 4510 855
rect 4476 821 4510 853
rect 4476 751 4510 783
rect 4476 749 4510 751
rect 5387 1105 5421 1139
rect 5479 1105 5513 1139
rect 5571 1105 5605 1139
rect 4898 1013 4932 1015
rect 4898 981 4932 1013
rect 4898 911 4932 943
rect 4898 909 4932 911
rect 5733 1099 5767 1133
rect 5825 1099 5859 1133
rect 5917 1099 5951 1133
rect 6096 1109 6130 1143
rect 4572 853 4606 855
rect 4572 821 4606 853
rect 4572 751 4606 783
rect 4854 781 4888 815
rect 4572 749 4606 751
rect 5393 793 5395 826
rect 5395 793 5427 826
rect 5393 792 5427 793
rect 6742 1109 6776 1143
rect 5586 804 5620 838
rect 4428 621 4462 655
rect 3845 555 3879 589
rect 3937 555 3971 589
rect 4029 555 4063 589
rect 4180 550 4214 584
rect 4812 578 4846 612
rect 5172 711 5206 728
rect 5172 694 5206 711
rect 5782 821 5816 832
rect 5782 798 5784 821
rect 5784 798 5816 821
rect 812 386 846 418
rect 812 384 846 386
rect 2508 488 2542 490
rect 2508 456 2542 488
rect 2604 488 2638 490
rect 2604 456 2638 488
rect 2508 386 2542 418
rect 2508 384 2542 386
rect 2604 386 2638 418
rect 2604 384 2638 386
rect 2700 488 2734 490
rect 2700 456 2734 488
rect 4540 540 4574 574
rect 5041 563 5075 597
rect 5133 563 5167 597
rect 5225 563 5259 597
rect 6343 1057 6377 1091
rect 7770 1364 7804 1398
rect 8158 1909 8192 1911
rect 8158 1877 8192 1909
rect 8158 1807 8192 1839
rect 8158 1805 8192 1807
rect 8254 1909 8288 1911
rect 8254 1877 8288 1909
rect 8254 1807 8288 1839
rect 8254 1805 8288 1807
rect 10121 2113 10155 2147
rect 10190 2005 10224 2039
rect 8350 1909 8384 1911
rect 8350 1877 8384 1909
rect 8617 1875 8651 1882
rect 8617 1848 8621 1875
rect 8621 1848 8651 1875
rect 8350 1807 8384 1839
rect 8350 1805 8384 1807
rect 8791 1875 8825 1882
rect 8791 1848 8823 1875
rect 8823 1848 8825 1875
rect 9693 1875 9727 1884
rect 9693 1850 9695 1875
rect 9695 1850 9727 1875
rect 9866 1875 9900 1880
rect 9866 1846 9897 1875
rect 9897 1846 9900 1875
rect 8206 1677 8240 1711
rect 8705 1755 8737 1759
rect 8737 1755 8739 1759
rect 8705 1725 8739 1755
rect 9775 1755 9777 1764
rect 9777 1755 9809 1764
rect 9775 1730 9809 1755
rect 8318 1596 8352 1630
rect 8613 1609 8647 1643
rect 8705 1609 8739 1643
rect 8797 1609 8831 1643
rect 9687 1609 9721 1643
rect 9779 1609 9813 1643
rect 9871 1609 9905 1643
rect 8174 1544 8208 1546
rect 8174 1512 8208 1544
rect 8174 1442 8208 1474
rect 8174 1440 8208 1442
rect 8270 1544 8304 1546
rect 8270 1512 8304 1544
rect 8270 1442 8304 1474
rect 8270 1440 8304 1442
rect 8366 1544 8400 1546
rect 8366 1512 8400 1544
rect 8366 1442 8400 1474
rect 8366 1440 8400 1442
rect 8222 1356 8256 1390
rect 8142 1247 8176 1281
rect 8572 1230 8606 1264
rect 6929 1107 6963 1141
rect 7021 1107 7055 1141
rect 7113 1107 7147 1141
rect 6052 1013 6086 1015
rect 6052 981 6086 1013
rect 6052 911 6086 943
rect 6052 909 6086 911
rect 6140 1013 6174 1015
rect 6140 981 6174 1013
rect 6698 1013 6732 1015
rect 6412 949 6446 983
rect 6698 981 6732 1013
rect 6140 911 6174 943
rect 6140 909 6174 911
rect 6698 911 6732 943
rect 6698 909 6732 911
rect 6268 853 6302 855
rect 6268 821 6302 853
rect 6096 781 6130 815
rect 5387 561 5421 595
rect 5479 561 5513 595
rect 5571 561 5605 595
rect 6268 751 6302 783
rect 6268 749 6302 751
rect 6364 853 6398 855
rect 6364 821 6398 853
rect 6364 751 6398 783
rect 6364 749 6398 751
rect 7275 1105 7309 1139
rect 7367 1105 7401 1139
rect 7459 1105 7493 1139
rect 6786 1013 6820 1015
rect 6786 981 6820 1013
rect 6786 911 6820 943
rect 6786 909 6820 911
rect 7621 1099 7655 1133
rect 7713 1099 7747 1133
rect 7805 1099 7839 1133
rect 7984 1109 8018 1143
rect 6460 853 6494 855
rect 6460 821 6494 853
rect 6460 751 6494 783
rect 6742 781 6776 815
rect 6460 749 6494 751
rect 7281 793 7283 826
rect 7283 793 7315 826
rect 7281 792 7315 793
rect 8630 1109 8664 1143
rect 7474 804 7508 838
rect 6316 621 6350 655
rect 5733 555 5767 589
rect 5825 555 5859 589
rect 5917 555 5951 589
rect 6068 550 6102 584
rect 6700 578 6734 612
rect 7060 711 7094 728
rect 7060 694 7094 711
rect 7670 821 7704 832
rect 7670 798 7672 821
rect 7672 798 7704 821
rect 2700 386 2734 418
rect 2700 384 2734 386
rect 4396 488 4430 490
rect 4396 456 4430 488
rect 4492 488 4526 490
rect 4492 456 4526 488
rect 4396 386 4430 418
rect 4396 384 4430 386
rect 4492 386 4526 418
rect 4492 384 4526 386
rect 4588 488 4622 490
rect 4588 456 4622 488
rect 6428 540 6462 574
rect 6929 563 6963 597
rect 7021 563 7055 597
rect 7113 563 7147 597
rect 8231 1057 8265 1091
rect 9658 1364 9692 1398
rect 10046 1909 10080 1911
rect 10046 1877 10080 1909
rect 10046 1807 10080 1839
rect 10046 1805 10080 1807
rect 10142 1909 10176 1911
rect 10142 1877 10176 1909
rect 10142 1807 10176 1839
rect 10142 1805 10176 1807
rect 12009 2113 12043 2147
rect 12078 2005 12112 2039
rect 10238 1909 10272 1911
rect 10238 1877 10272 1909
rect 10505 1875 10539 1882
rect 10505 1848 10509 1875
rect 10509 1848 10539 1875
rect 10238 1807 10272 1839
rect 10238 1805 10272 1807
rect 10679 1875 10713 1882
rect 10679 1848 10711 1875
rect 10711 1848 10713 1875
rect 11581 1875 11615 1884
rect 11581 1850 11583 1875
rect 11583 1850 11615 1875
rect 11754 1875 11788 1880
rect 11754 1846 11785 1875
rect 11785 1846 11788 1875
rect 10094 1677 10128 1711
rect 10593 1755 10625 1759
rect 10625 1755 10627 1759
rect 10593 1725 10627 1755
rect 11663 1755 11665 1764
rect 11665 1755 11697 1764
rect 11663 1730 11697 1755
rect 10206 1596 10240 1630
rect 10501 1609 10535 1643
rect 10593 1609 10627 1643
rect 10685 1609 10719 1643
rect 11575 1609 11609 1643
rect 11667 1609 11701 1643
rect 11759 1609 11793 1643
rect 10062 1544 10096 1546
rect 10062 1512 10096 1544
rect 10062 1442 10096 1474
rect 10062 1440 10096 1442
rect 10158 1544 10192 1546
rect 10158 1512 10192 1544
rect 10158 1442 10192 1474
rect 10158 1440 10192 1442
rect 10254 1544 10288 1546
rect 10254 1512 10288 1544
rect 10254 1442 10288 1474
rect 10254 1440 10288 1442
rect 10110 1356 10144 1390
rect 10030 1247 10064 1281
rect 10460 1230 10494 1264
rect 8817 1107 8851 1141
rect 8909 1107 8943 1141
rect 9001 1107 9035 1141
rect 7940 1013 7974 1015
rect 7940 981 7974 1013
rect 7940 911 7974 943
rect 7940 909 7974 911
rect 8028 1013 8062 1015
rect 8028 981 8062 1013
rect 8586 1013 8620 1015
rect 8300 949 8334 983
rect 8586 981 8620 1013
rect 8028 911 8062 943
rect 8028 909 8062 911
rect 8586 911 8620 943
rect 8586 909 8620 911
rect 8156 853 8190 855
rect 8156 821 8190 853
rect 7984 781 8018 815
rect 7275 561 7309 595
rect 7367 561 7401 595
rect 7459 561 7493 595
rect 8156 751 8190 783
rect 8156 749 8190 751
rect 8252 853 8286 855
rect 8252 821 8286 853
rect 8252 751 8286 783
rect 8252 749 8286 751
rect 9163 1105 9197 1139
rect 9255 1105 9289 1139
rect 9347 1105 9381 1139
rect 8674 1013 8708 1015
rect 8674 981 8708 1013
rect 8674 911 8708 943
rect 8674 909 8708 911
rect 9509 1099 9543 1133
rect 9601 1099 9635 1133
rect 9693 1099 9727 1133
rect 9872 1109 9906 1143
rect 8348 853 8382 855
rect 8348 821 8382 853
rect 8348 751 8382 783
rect 8630 781 8664 815
rect 8348 749 8382 751
rect 9169 793 9171 826
rect 9171 793 9203 826
rect 9169 792 9203 793
rect 10518 1109 10552 1143
rect 9362 804 9396 838
rect 8204 621 8238 655
rect 7621 555 7655 589
rect 7713 555 7747 589
rect 7805 555 7839 589
rect 7956 550 7990 584
rect 8588 578 8622 612
rect 8948 711 8982 728
rect 8948 694 8982 711
rect 9558 821 9592 832
rect 9558 798 9560 821
rect 9560 798 9592 821
rect 4588 386 4622 418
rect 4588 384 4622 386
rect 6284 488 6318 490
rect 6284 456 6318 488
rect 6380 488 6414 490
rect 6380 456 6414 488
rect 6284 386 6318 418
rect 6284 384 6318 386
rect 6380 386 6414 418
rect 6380 384 6414 386
rect 6476 488 6510 490
rect 6476 456 6510 488
rect 8316 540 8350 574
rect 8817 563 8851 597
rect 8909 563 8943 597
rect 9001 563 9035 597
rect 10119 1057 10153 1091
rect 11546 1364 11580 1398
rect 11934 1909 11968 1911
rect 11934 1877 11968 1909
rect 11934 1807 11968 1839
rect 11934 1805 11968 1807
rect 12030 1909 12064 1911
rect 12030 1877 12064 1909
rect 12030 1807 12064 1839
rect 12030 1805 12064 1807
rect 13897 2113 13931 2147
rect 13966 2005 14000 2039
rect 12126 1909 12160 1911
rect 12126 1877 12160 1909
rect 12393 1875 12427 1882
rect 12393 1848 12397 1875
rect 12397 1848 12427 1875
rect 12126 1807 12160 1839
rect 12126 1805 12160 1807
rect 12567 1875 12601 1882
rect 12567 1848 12599 1875
rect 12599 1848 12601 1875
rect 13469 1875 13503 1884
rect 13469 1850 13471 1875
rect 13471 1850 13503 1875
rect 13642 1875 13676 1880
rect 13642 1846 13673 1875
rect 13673 1846 13676 1875
rect 11982 1677 12016 1711
rect 12481 1755 12513 1759
rect 12513 1755 12515 1759
rect 12481 1725 12515 1755
rect 13551 1755 13553 1764
rect 13553 1755 13585 1764
rect 13551 1730 13585 1755
rect 12094 1596 12128 1630
rect 12389 1609 12423 1643
rect 12481 1609 12515 1643
rect 12573 1609 12607 1643
rect 13463 1609 13497 1643
rect 13555 1609 13589 1643
rect 13647 1609 13681 1643
rect 11950 1544 11984 1546
rect 11950 1512 11984 1544
rect 11950 1442 11984 1474
rect 11950 1440 11984 1442
rect 12046 1544 12080 1546
rect 12046 1512 12080 1544
rect 12046 1442 12080 1474
rect 12046 1440 12080 1442
rect 12142 1544 12176 1546
rect 12142 1512 12176 1544
rect 12142 1442 12176 1474
rect 12142 1440 12176 1442
rect 11998 1356 12032 1390
rect 11918 1247 11952 1281
rect 12348 1230 12382 1264
rect 10705 1107 10739 1141
rect 10797 1107 10831 1141
rect 10889 1107 10923 1141
rect 9828 1013 9862 1015
rect 9828 981 9862 1013
rect 9828 911 9862 943
rect 9828 909 9862 911
rect 9916 1013 9950 1015
rect 9916 981 9950 1013
rect 10474 1013 10508 1015
rect 10188 949 10222 983
rect 10474 981 10508 1013
rect 9916 911 9950 943
rect 9916 909 9950 911
rect 10474 911 10508 943
rect 10474 909 10508 911
rect 10044 853 10078 855
rect 10044 821 10078 853
rect 9872 781 9906 815
rect 9163 561 9197 595
rect 9255 561 9289 595
rect 9347 561 9381 595
rect 10044 751 10078 783
rect 10044 749 10078 751
rect 10140 853 10174 855
rect 10140 821 10174 853
rect 10140 751 10174 783
rect 10140 749 10174 751
rect 11051 1105 11085 1139
rect 11143 1105 11177 1139
rect 11235 1105 11269 1139
rect 10562 1013 10596 1015
rect 10562 981 10596 1013
rect 10562 911 10596 943
rect 10562 909 10596 911
rect 11397 1099 11431 1133
rect 11489 1099 11523 1133
rect 11581 1099 11615 1133
rect 11760 1109 11794 1143
rect 10236 853 10270 855
rect 10236 821 10270 853
rect 10236 751 10270 783
rect 10518 781 10552 815
rect 10236 749 10270 751
rect 11057 793 11059 826
rect 11059 793 11091 826
rect 11057 792 11091 793
rect 12406 1109 12440 1143
rect 11250 804 11284 838
rect 10092 621 10126 655
rect 9509 555 9543 589
rect 9601 555 9635 589
rect 9693 555 9727 589
rect 9844 550 9878 584
rect 10476 578 10510 612
rect 10836 711 10870 728
rect 10836 694 10870 711
rect 11446 821 11480 832
rect 11446 798 11448 821
rect 11448 798 11480 821
rect 6476 386 6510 418
rect 6476 384 6510 386
rect 8172 488 8206 490
rect 8172 456 8206 488
rect 8268 488 8302 490
rect 8268 456 8302 488
rect 8172 386 8206 418
rect 8172 384 8206 386
rect 8268 386 8302 418
rect 8268 384 8302 386
rect 8364 488 8398 490
rect 8364 456 8398 488
rect 10204 540 10238 574
rect 10705 563 10739 597
rect 10797 563 10831 597
rect 10889 563 10923 597
rect 12007 1057 12041 1091
rect 13434 1364 13468 1398
rect 13822 1909 13856 1911
rect 13822 1877 13856 1909
rect 13822 1807 13856 1839
rect 13822 1805 13856 1807
rect 13918 1909 13952 1911
rect 13918 1877 13952 1909
rect 13918 1807 13952 1839
rect 13918 1805 13952 1807
rect 15779 2113 15813 2147
rect 15848 2005 15882 2039
rect 14014 1909 14048 1911
rect 14014 1877 14048 1909
rect 14281 1875 14315 1882
rect 14281 1848 14285 1875
rect 14285 1848 14315 1875
rect 14014 1807 14048 1839
rect 14014 1805 14048 1807
rect 14455 1875 14489 1882
rect 14455 1848 14487 1875
rect 14487 1848 14489 1875
rect 15351 1875 15385 1884
rect 15351 1850 15353 1875
rect 15353 1850 15385 1875
rect 15524 1875 15558 1880
rect 15524 1846 15555 1875
rect 15555 1846 15558 1875
rect 13870 1677 13904 1711
rect 14369 1755 14401 1759
rect 14401 1755 14403 1759
rect 14369 1725 14403 1755
rect 15433 1755 15435 1764
rect 15435 1755 15467 1764
rect 15433 1730 15467 1755
rect 13982 1596 14016 1630
rect 14277 1609 14311 1643
rect 14369 1609 14403 1643
rect 14461 1609 14495 1643
rect 15345 1609 15379 1643
rect 15437 1609 15471 1643
rect 15529 1609 15563 1643
rect 13838 1544 13872 1546
rect 13838 1512 13872 1544
rect 13838 1442 13872 1474
rect 13838 1440 13872 1442
rect 13934 1544 13968 1546
rect 13934 1512 13968 1544
rect 13934 1442 13968 1474
rect 13934 1440 13968 1442
rect 14030 1544 14064 1546
rect 14030 1512 14064 1544
rect 14030 1442 14064 1474
rect 14030 1440 14064 1442
rect 13886 1356 13920 1390
rect 13806 1247 13840 1281
rect 14236 1230 14270 1264
rect 12593 1107 12627 1141
rect 12685 1107 12719 1141
rect 12777 1107 12811 1141
rect 11716 1013 11750 1015
rect 11716 981 11750 1013
rect 11716 911 11750 943
rect 11716 909 11750 911
rect 11804 1013 11838 1015
rect 11804 981 11838 1013
rect 12362 1013 12396 1015
rect 12076 949 12110 983
rect 12362 981 12396 1013
rect 11804 911 11838 943
rect 11804 909 11838 911
rect 12362 911 12396 943
rect 12362 909 12396 911
rect 11932 853 11966 855
rect 11932 821 11966 853
rect 11760 781 11794 815
rect 11051 561 11085 595
rect 11143 561 11177 595
rect 11235 561 11269 595
rect 11932 751 11966 783
rect 11932 749 11966 751
rect 12028 853 12062 855
rect 12028 821 12062 853
rect 12028 751 12062 783
rect 12028 749 12062 751
rect 12939 1105 12973 1139
rect 13031 1105 13065 1139
rect 13123 1105 13157 1139
rect 12450 1013 12484 1015
rect 12450 981 12484 1013
rect 12450 911 12484 943
rect 12450 909 12484 911
rect 13285 1099 13319 1133
rect 13377 1099 13411 1133
rect 13469 1099 13503 1133
rect 13648 1109 13682 1143
rect 12124 853 12158 855
rect 12124 821 12158 853
rect 12124 751 12158 783
rect 12406 781 12440 815
rect 12124 749 12158 751
rect 12945 793 12947 826
rect 12947 793 12979 826
rect 12945 792 12979 793
rect 14294 1109 14328 1143
rect 13138 804 13172 838
rect 11980 621 12014 655
rect 11397 555 11431 589
rect 11489 555 11523 589
rect 11581 555 11615 589
rect 11732 550 11766 584
rect 12364 578 12398 612
rect 12724 711 12758 728
rect 12724 694 12758 711
rect 13334 821 13368 832
rect 13334 798 13336 821
rect 13336 798 13368 821
rect 8364 386 8398 418
rect 8364 384 8398 386
rect 10060 488 10094 490
rect 10060 456 10094 488
rect 10156 488 10190 490
rect 10156 456 10190 488
rect 10060 386 10094 418
rect 10060 384 10094 386
rect 10156 386 10190 418
rect 10156 384 10190 386
rect 10252 488 10286 490
rect 10252 456 10286 488
rect 12092 540 12126 574
rect 12593 563 12627 597
rect 12685 563 12719 597
rect 12777 563 12811 597
rect 13895 1057 13929 1091
rect 15316 1364 15350 1398
rect 15704 1909 15738 1911
rect 15704 1877 15738 1909
rect 15704 1807 15738 1839
rect 15704 1805 15738 1807
rect 15800 1909 15834 1911
rect 15800 1877 15834 1909
rect 15800 1807 15834 1839
rect 15800 1805 15834 1807
rect 17667 2113 17701 2147
rect 17736 2005 17770 2039
rect 15896 1909 15930 1911
rect 15896 1877 15930 1909
rect 16163 1875 16197 1882
rect 16163 1848 16167 1875
rect 16167 1848 16197 1875
rect 15896 1807 15930 1839
rect 15896 1805 15930 1807
rect 16337 1875 16371 1882
rect 16337 1848 16369 1875
rect 16369 1848 16371 1875
rect 17239 1875 17273 1884
rect 17239 1850 17241 1875
rect 17241 1850 17273 1875
rect 17412 1875 17446 1880
rect 17412 1846 17443 1875
rect 17443 1846 17446 1875
rect 15752 1677 15786 1711
rect 16251 1755 16283 1759
rect 16283 1755 16285 1759
rect 16251 1725 16285 1755
rect 17321 1755 17323 1764
rect 17323 1755 17355 1764
rect 17321 1730 17355 1755
rect 15864 1596 15898 1630
rect 16159 1609 16193 1643
rect 16251 1609 16285 1643
rect 16343 1609 16377 1643
rect 17233 1609 17267 1643
rect 17325 1609 17359 1643
rect 17417 1609 17451 1643
rect 15720 1544 15754 1546
rect 15720 1512 15754 1544
rect 15720 1442 15754 1474
rect 15720 1440 15754 1442
rect 15816 1544 15850 1546
rect 15816 1512 15850 1544
rect 15816 1442 15850 1474
rect 15816 1440 15850 1442
rect 15912 1544 15946 1546
rect 15912 1512 15946 1544
rect 15912 1442 15946 1474
rect 15912 1440 15946 1442
rect 15768 1356 15802 1390
rect 15688 1247 15722 1281
rect 16118 1230 16152 1264
rect 14481 1107 14515 1141
rect 14573 1107 14607 1141
rect 14665 1107 14699 1141
rect 13604 1013 13638 1015
rect 13604 981 13638 1013
rect 13604 911 13638 943
rect 13604 909 13638 911
rect 13692 1013 13726 1015
rect 13692 981 13726 1013
rect 14250 1013 14284 1015
rect 13964 949 13998 983
rect 14250 981 14284 1013
rect 13692 911 13726 943
rect 13692 909 13726 911
rect 14250 911 14284 943
rect 14250 909 14284 911
rect 13820 853 13854 855
rect 13820 821 13854 853
rect 13648 781 13682 815
rect 12939 561 12973 595
rect 13031 561 13065 595
rect 13123 561 13157 595
rect 13820 751 13854 783
rect 13820 749 13854 751
rect 13916 853 13950 855
rect 13916 821 13950 853
rect 13916 751 13950 783
rect 13916 749 13950 751
rect 14827 1105 14861 1139
rect 14919 1105 14953 1139
rect 15011 1105 15045 1139
rect 14338 1013 14372 1015
rect 14338 981 14372 1013
rect 14338 911 14372 943
rect 14338 909 14372 911
rect 15167 1099 15201 1133
rect 15259 1099 15293 1133
rect 15351 1099 15385 1133
rect 15530 1109 15564 1143
rect 14012 853 14046 855
rect 14012 821 14046 853
rect 14012 751 14046 783
rect 14294 781 14328 815
rect 14012 749 14046 751
rect 14833 793 14835 826
rect 14835 793 14867 826
rect 14833 792 14867 793
rect 16176 1109 16210 1143
rect 15026 804 15060 838
rect 13868 621 13902 655
rect 13285 555 13319 589
rect 13377 555 13411 589
rect 13469 555 13503 589
rect 13620 550 13654 584
rect 14252 578 14286 612
rect 14612 711 14646 728
rect 14612 694 14646 711
rect 15216 821 15250 832
rect 15216 798 15218 821
rect 15218 798 15250 821
rect 10252 386 10286 418
rect 10252 384 10286 386
rect 11948 488 11982 490
rect 11948 456 11982 488
rect 12044 488 12078 490
rect 12044 456 12078 488
rect 11948 386 11982 418
rect 11948 384 11982 386
rect 12044 386 12078 418
rect 12044 384 12078 386
rect 12140 488 12174 490
rect 12140 456 12174 488
rect 13980 540 14014 574
rect 14481 563 14515 597
rect 14573 563 14607 597
rect 14665 563 14699 597
rect 15777 1057 15811 1091
rect 17204 1364 17238 1398
rect 17592 1909 17626 1911
rect 17592 1877 17626 1909
rect 17592 1807 17626 1839
rect 17592 1805 17626 1807
rect 17688 1909 17722 1911
rect 17688 1877 17722 1909
rect 17688 1807 17722 1839
rect 17688 1805 17722 1807
rect 19555 2113 19589 2147
rect 19624 2005 19658 2039
rect 17784 1909 17818 1911
rect 17784 1877 17818 1909
rect 18051 1875 18085 1882
rect 18051 1848 18055 1875
rect 18055 1848 18085 1875
rect 17784 1807 17818 1839
rect 17784 1805 17818 1807
rect 18225 1875 18259 1882
rect 18225 1848 18257 1875
rect 18257 1848 18259 1875
rect 19127 1875 19161 1884
rect 19127 1850 19129 1875
rect 19129 1850 19161 1875
rect 19300 1875 19334 1880
rect 19300 1846 19331 1875
rect 19331 1846 19334 1875
rect 17640 1677 17674 1711
rect 18139 1755 18171 1759
rect 18171 1755 18173 1759
rect 18139 1725 18173 1755
rect 19209 1755 19211 1764
rect 19211 1755 19243 1764
rect 19209 1730 19243 1755
rect 17752 1596 17786 1630
rect 18047 1609 18081 1643
rect 18139 1609 18173 1643
rect 18231 1609 18265 1643
rect 19121 1609 19155 1643
rect 19213 1609 19247 1643
rect 19305 1609 19339 1643
rect 17608 1544 17642 1546
rect 17608 1512 17642 1544
rect 17608 1442 17642 1474
rect 17608 1440 17642 1442
rect 17704 1544 17738 1546
rect 17704 1512 17738 1544
rect 17704 1442 17738 1474
rect 17704 1440 17738 1442
rect 17800 1544 17834 1546
rect 17800 1512 17834 1544
rect 17800 1442 17834 1474
rect 17800 1440 17834 1442
rect 17656 1356 17690 1390
rect 17576 1247 17610 1281
rect 18006 1230 18040 1264
rect 16363 1107 16397 1141
rect 16455 1107 16489 1141
rect 16547 1107 16581 1141
rect 15486 1013 15520 1015
rect 15486 981 15520 1013
rect 15486 911 15520 943
rect 15486 909 15520 911
rect 15574 1013 15608 1015
rect 15574 981 15608 1013
rect 16132 1013 16166 1015
rect 15846 949 15880 983
rect 16132 981 16166 1013
rect 15574 911 15608 943
rect 15574 909 15608 911
rect 16132 911 16166 943
rect 16132 909 16166 911
rect 15702 853 15736 855
rect 15702 821 15736 853
rect 15530 781 15564 815
rect 14827 561 14861 595
rect 14919 561 14953 595
rect 15011 561 15045 595
rect 15702 751 15736 783
rect 15702 749 15736 751
rect 15798 853 15832 855
rect 15798 821 15832 853
rect 15798 751 15832 783
rect 15798 749 15832 751
rect 16709 1105 16743 1139
rect 16801 1105 16835 1139
rect 16893 1105 16927 1139
rect 16220 1013 16254 1015
rect 16220 981 16254 1013
rect 16220 911 16254 943
rect 16220 909 16254 911
rect 17055 1099 17089 1133
rect 17147 1099 17181 1133
rect 17239 1099 17273 1133
rect 17418 1109 17452 1143
rect 15894 853 15928 855
rect 15894 821 15928 853
rect 15894 751 15928 783
rect 16176 781 16210 815
rect 15894 749 15928 751
rect 16715 793 16717 826
rect 16717 793 16749 826
rect 16715 792 16749 793
rect 18064 1109 18098 1143
rect 16908 804 16942 838
rect 15750 621 15784 655
rect 15167 555 15201 589
rect 15259 555 15293 589
rect 15351 555 15385 589
rect 15502 550 15536 584
rect 16134 578 16168 612
rect 16494 711 16528 728
rect 16494 694 16528 711
rect 17104 821 17138 832
rect 17104 798 17106 821
rect 17106 798 17138 821
rect 12140 386 12174 418
rect 12140 384 12174 386
rect 13836 488 13870 490
rect 13836 456 13870 488
rect 13932 488 13966 490
rect 13932 456 13966 488
rect 13836 386 13870 418
rect 13836 384 13870 386
rect 13932 386 13966 418
rect 13932 384 13966 386
rect 14028 488 14062 490
rect 14028 456 14062 488
rect 15862 540 15896 574
rect 16363 563 16397 597
rect 16455 563 16489 597
rect 16547 563 16581 597
rect 17665 1057 17699 1091
rect 19092 1364 19126 1398
rect 19480 1909 19514 1911
rect 19480 1877 19514 1909
rect 19480 1807 19514 1839
rect 19480 1805 19514 1807
rect 19576 1909 19610 1911
rect 19576 1877 19610 1909
rect 19576 1807 19610 1839
rect 19576 1805 19610 1807
rect 21443 2113 21477 2147
rect 21512 2005 21546 2039
rect 19672 1909 19706 1911
rect 19672 1877 19706 1909
rect 19939 1875 19973 1882
rect 19939 1848 19943 1875
rect 19943 1848 19973 1875
rect 19672 1807 19706 1839
rect 19672 1805 19706 1807
rect 20113 1875 20147 1882
rect 20113 1848 20145 1875
rect 20145 1848 20147 1875
rect 21015 1875 21049 1884
rect 21015 1850 21017 1875
rect 21017 1850 21049 1875
rect 21188 1875 21222 1880
rect 21188 1846 21219 1875
rect 21219 1846 21222 1875
rect 19528 1677 19562 1711
rect 20027 1755 20059 1759
rect 20059 1755 20061 1759
rect 20027 1725 20061 1755
rect 21097 1755 21099 1764
rect 21099 1755 21131 1764
rect 21097 1730 21131 1755
rect 19640 1596 19674 1630
rect 19935 1609 19969 1643
rect 20027 1609 20061 1643
rect 20119 1609 20153 1643
rect 21009 1609 21043 1643
rect 21101 1609 21135 1643
rect 21193 1609 21227 1643
rect 19496 1544 19530 1546
rect 19496 1512 19530 1544
rect 19496 1442 19530 1474
rect 19496 1440 19530 1442
rect 19592 1544 19626 1546
rect 19592 1512 19626 1544
rect 19592 1442 19626 1474
rect 19592 1440 19626 1442
rect 19688 1544 19722 1546
rect 19688 1512 19722 1544
rect 19688 1442 19722 1474
rect 19688 1440 19722 1442
rect 19544 1356 19578 1390
rect 19464 1247 19498 1281
rect 19894 1230 19928 1264
rect 18251 1107 18285 1141
rect 18343 1107 18377 1141
rect 18435 1107 18469 1141
rect 17374 1013 17408 1015
rect 17374 981 17408 1013
rect 17374 911 17408 943
rect 17374 909 17408 911
rect 17462 1013 17496 1015
rect 17462 981 17496 1013
rect 18020 1013 18054 1015
rect 17734 949 17768 983
rect 18020 981 18054 1013
rect 17462 911 17496 943
rect 17462 909 17496 911
rect 18020 911 18054 943
rect 18020 909 18054 911
rect 17590 853 17624 855
rect 17590 821 17624 853
rect 17418 781 17452 815
rect 16709 561 16743 595
rect 16801 561 16835 595
rect 16893 561 16927 595
rect 17590 751 17624 783
rect 17590 749 17624 751
rect 17686 853 17720 855
rect 17686 821 17720 853
rect 17686 751 17720 783
rect 17686 749 17720 751
rect 18597 1105 18631 1139
rect 18689 1105 18723 1139
rect 18781 1105 18815 1139
rect 18108 1013 18142 1015
rect 18108 981 18142 1013
rect 18108 911 18142 943
rect 18108 909 18142 911
rect 18943 1099 18977 1133
rect 19035 1099 19069 1133
rect 19127 1099 19161 1133
rect 19306 1109 19340 1143
rect 17782 853 17816 855
rect 17782 821 17816 853
rect 17782 751 17816 783
rect 18064 781 18098 815
rect 17782 749 17816 751
rect 18603 793 18605 826
rect 18605 793 18637 826
rect 18603 792 18637 793
rect 19952 1109 19986 1143
rect 18796 804 18830 838
rect 17638 621 17672 655
rect 17055 555 17089 589
rect 17147 555 17181 589
rect 17239 555 17273 589
rect 17390 550 17424 584
rect 18022 578 18056 612
rect 18382 711 18416 728
rect 18382 694 18416 711
rect 18992 821 19026 832
rect 18992 798 18994 821
rect 18994 798 19026 821
rect 14028 386 14062 418
rect 14028 384 14062 386
rect 15718 488 15752 490
rect 15718 456 15752 488
rect 15814 488 15848 490
rect 15814 456 15848 488
rect 15718 386 15752 418
rect 15718 384 15752 386
rect 15814 386 15848 418
rect 15814 384 15848 386
rect 15910 488 15944 490
rect 15910 456 15944 488
rect 17750 540 17784 574
rect 18251 563 18285 597
rect 18343 563 18377 597
rect 18435 563 18469 597
rect 19553 1057 19587 1091
rect 20980 1364 21014 1398
rect 21368 1909 21402 1911
rect 21368 1877 21402 1909
rect 21368 1807 21402 1839
rect 21368 1805 21402 1807
rect 21464 1909 21498 1911
rect 21464 1877 21498 1909
rect 21464 1807 21498 1839
rect 21464 1805 21498 1807
rect 23331 2113 23365 2147
rect 23400 2005 23434 2039
rect 21560 1909 21594 1911
rect 21560 1877 21594 1909
rect 21827 1875 21861 1882
rect 21827 1848 21831 1875
rect 21831 1848 21861 1875
rect 21560 1807 21594 1839
rect 21560 1805 21594 1807
rect 22001 1875 22035 1882
rect 22001 1848 22033 1875
rect 22033 1848 22035 1875
rect 22903 1875 22937 1884
rect 22903 1850 22905 1875
rect 22905 1850 22937 1875
rect 23076 1875 23110 1880
rect 23076 1846 23107 1875
rect 23107 1846 23110 1875
rect 21416 1677 21450 1711
rect 21915 1755 21947 1759
rect 21947 1755 21949 1759
rect 21915 1725 21949 1755
rect 22985 1755 22987 1764
rect 22987 1755 23019 1764
rect 22985 1730 23019 1755
rect 21528 1596 21562 1630
rect 21823 1609 21857 1643
rect 21915 1609 21949 1643
rect 22007 1609 22041 1643
rect 22897 1609 22931 1643
rect 22989 1609 23023 1643
rect 23081 1609 23115 1643
rect 21384 1544 21418 1546
rect 21384 1512 21418 1544
rect 21384 1442 21418 1474
rect 21384 1440 21418 1442
rect 21480 1544 21514 1546
rect 21480 1512 21514 1544
rect 21480 1442 21514 1474
rect 21480 1440 21514 1442
rect 21576 1544 21610 1546
rect 21576 1512 21610 1544
rect 21576 1442 21610 1474
rect 21576 1440 21610 1442
rect 21432 1356 21466 1390
rect 21352 1247 21386 1281
rect 21782 1230 21816 1264
rect 20139 1107 20173 1141
rect 20231 1107 20265 1141
rect 20323 1107 20357 1141
rect 19262 1013 19296 1015
rect 19262 981 19296 1013
rect 19262 911 19296 943
rect 19262 909 19296 911
rect 19350 1013 19384 1015
rect 19350 981 19384 1013
rect 19908 1013 19942 1015
rect 19622 949 19656 983
rect 19908 981 19942 1013
rect 19350 911 19384 943
rect 19350 909 19384 911
rect 19908 911 19942 943
rect 19908 909 19942 911
rect 19478 853 19512 855
rect 19478 821 19512 853
rect 19306 781 19340 815
rect 18597 561 18631 595
rect 18689 561 18723 595
rect 18781 561 18815 595
rect 19478 751 19512 783
rect 19478 749 19512 751
rect 19574 853 19608 855
rect 19574 821 19608 853
rect 19574 751 19608 783
rect 19574 749 19608 751
rect 20485 1105 20519 1139
rect 20577 1105 20611 1139
rect 20669 1105 20703 1139
rect 19996 1013 20030 1015
rect 19996 981 20030 1013
rect 19996 911 20030 943
rect 19996 909 20030 911
rect 20831 1099 20865 1133
rect 20923 1099 20957 1133
rect 21015 1099 21049 1133
rect 21194 1109 21228 1143
rect 19670 853 19704 855
rect 19670 821 19704 853
rect 19670 751 19704 783
rect 19952 781 19986 815
rect 19670 749 19704 751
rect 20491 793 20493 826
rect 20493 793 20525 826
rect 20491 792 20525 793
rect 21840 1109 21874 1143
rect 20684 804 20718 838
rect 19526 621 19560 655
rect 18943 555 18977 589
rect 19035 555 19069 589
rect 19127 555 19161 589
rect 19278 550 19312 584
rect 19910 578 19944 612
rect 20270 711 20304 728
rect 20270 694 20304 711
rect 20880 821 20914 832
rect 20880 798 20882 821
rect 20882 798 20914 821
rect 15910 386 15944 418
rect 15910 384 15944 386
rect 17606 488 17640 490
rect 17606 456 17640 488
rect 17702 488 17736 490
rect 17702 456 17736 488
rect 17606 386 17640 418
rect 17606 384 17640 386
rect 17702 386 17736 418
rect 17702 384 17736 386
rect 17798 488 17832 490
rect 17798 456 17832 488
rect 19638 540 19672 574
rect 20139 563 20173 597
rect 20231 563 20265 597
rect 20323 563 20357 597
rect 21441 1057 21475 1091
rect 22868 1364 22902 1398
rect 23256 1909 23290 1911
rect 23256 1877 23290 1909
rect 23256 1807 23290 1839
rect 23256 1805 23290 1807
rect 23352 1909 23386 1911
rect 23352 1877 23386 1909
rect 23352 1807 23386 1839
rect 23352 1805 23386 1807
rect 25219 2113 25253 2147
rect 25288 2005 25322 2039
rect 23448 1909 23482 1911
rect 23448 1877 23482 1909
rect 23715 1875 23749 1882
rect 23715 1848 23719 1875
rect 23719 1848 23749 1875
rect 23448 1807 23482 1839
rect 23448 1805 23482 1807
rect 23889 1875 23923 1882
rect 23889 1848 23921 1875
rect 23921 1848 23923 1875
rect 24791 1875 24825 1884
rect 24791 1850 24793 1875
rect 24793 1850 24825 1875
rect 24964 1875 24998 1880
rect 24964 1846 24995 1875
rect 24995 1846 24998 1875
rect 23304 1677 23338 1711
rect 23803 1755 23835 1759
rect 23835 1755 23837 1759
rect 23803 1725 23837 1755
rect 24873 1755 24875 1764
rect 24875 1755 24907 1764
rect 24873 1730 24907 1755
rect 23416 1596 23450 1630
rect 23711 1609 23745 1643
rect 23803 1609 23837 1643
rect 23895 1609 23929 1643
rect 24785 1609 24819 1643
rect 24877 1609 24911 1643
rect 24969 1609 25003 1643
rect 23272 1544 23306 1546
rect 23272 1512 23306 1544
rect 23272 1442 23306 1474
rect 23272 1440 23306 1442
rect 23368 1544 23402 1546
rect 23368 1512 23402 1544
rect 23368 1442 23402 1474
rect 23368 1440 23402 1442
rect 23464 1544 23498 1546
rect 23464 1512 23498 1544
rect 23464 1442 23498 1474
rect 23464 1440 23498 1442
rect 23320 1356 23354 1390
rect 23240 1247 23274 1281
rect 23670 1230 23704 1264
rect 22027 1107 22061 1141
rect 22119 1107 22153 1141
rect 22211 1107 22245 1141
rect 21150 1013 21184 1015
rect 21150 981 21184 1013
rect 21150 911 21184 943
rect 21150 909 21184 911
rect 21238 1013 21272 1015
rect 21238 981 21272 1013
rect 21796 1013 21830 1015
rect 21510 949 21544 983
rect 21796 981 21830 1013
rect 21238 911 21272 943
rect 21238 909 21272 911
rect 21796 911 21830 943
rect 21796 909 21830 911
rect 21366 853 21400 855
rect 21366 821 21400 853
rect 21194 781 21228 815
rect 20485 561 20519 595
rect 20577 561 20611 595
rect 20669 561 20703 595
rect 21366 751 21400 783
rect 21366 749 21400 751
rect 21462 853 21496 855
rect 21462 821 21496 853
rect 21462 751 21496 783
rect 21462 749 21496 751
rect 22373 1105 22407 1139
rect 22465 1105 22499 1139
rect 22557 1105 22591 1139
rect 21884 1013 21918 1015
rect 21884 981 21918 1013
rect 21884 911 21918 943
rect 21884 909 21918 911
rect 22719 1099 22753 1133
rect 22811 1099 22845 1133
rect 22903 1099 22937 1133
rect 23082 1109 23116 1143
rect 21558 853 21592 855
rect 21558 821 21592 853
rect 21558 751 21592 783
rect 21840 781 21874 815
rect 21558 749 21592 751
rect 22379 793 22381 826
rect 22381 793 22413 826
rect 22379 792 22413 793
rect 23728 1109 23762 1143
rect 22572 804 22606 838
rect 21414 621 21448 655
rect 20831 555 20865 589
rect 20923 555 20957 589
rect 21015 555 21049 589
rect 21166 550 21200 584
rect 21798 578 21832 612
rect 22158 711 22192 728
rect 22158 694 22192 711
rect 22768 821 22802 832
rect 22768 798 22770 821
rect 22770 798 22802 821
rect 17798 386 17832 418
rect 17798 384 17832 386
rect 19494 488 19528 490
rect 19494 456 19528 488
rect 19590 488 19624 490
rect 19590 456 19624 488
rect 19494 386 19528 418
rect 19494 384 19528 386
rect 19590 386 19624 418
rect 19590 384 19624 386
rect 19686 488 19720 490
rect 19686 456 19720 488
rect 21526 540 21560 574
rect 22027 563 22061 597
rect 22119 563 22153 597
rect 22211 563 22245 597
rect 23329 1057 23363 1091
rect 24756 1364 24790 1398
rect 25144 1909 25178 1911
rect 25144 1877 25178 1909
rect 25144 1807 25178 1839
rect 25144 1805 25178 1807
rect 25240 1909 25274 1911
rect 25240 1877 25274 1909
rect 25240 1807 25274 1839
rect 25240 1805 25274 1807
rect 27107 2113 27141 2147
rect 27176 2005 27210 2039
rect 25336 1909 25370 1911
rect 25336 1877 25370 1909
rect 25603 1875 25637 1882
rect 25603 1848 25607 1875
rect 25607 1848 25637 1875
rect 25336 1807 25370 1839
rect 25336 1805 25370 1807
rect 25777 1875 25811 1882
rect 25777 1848 25809 1875
rect 25809 1848 25811 1875
rect 26679 1875 26713 1884
rect 26679 1850 26681 1875
rect 26681 1850 26713 1875
rect 26852 1875 26886 1880
rect 26852 1846 26883 1875
rect 26883 1846 26886 1875
rect 25192 1677 25226 1711
rect 25691 1755 25723 1759
rect 25723 1755 25725 1759
rect 25691 1725 25725 1755
rect 26761 1755 26763 1764
rect 26763 1755 26795 1764
rect 26761 1730 26795 1755
rect 25304 1596 25338 1630
rect 25599 1609 25633 1643
rect 25691 1609 25725 1643
rect 25783 1609 25817 1643
rect 26673 1609 26707 1643
rect 26765 1609 26799 1643
rect 26857 1609 26891 1643
rect 25160 1544 25194 1546
rect 25160 1512 25194 1544
rect 25160 1442 25194 1474
rect 25160 1440 25194 1442
rect 25256 1544 25290 1546
rect 25256 1512 25290 1544
rect 25256 1442 25290 1474
rect 25256 1440 25290 1442
rect 25352 1544 25386 1546
rect 25352 1512 25386 1544
rect 25352 1442 25386 1474
rect 25352 1440 25386 1442
rect 25208 1356 25242 1390
rect 25128 1247 25162 1281
rect 25558 1230 25592 1264
rect 23915 1107 23949 1141
rect 24007 1107 24041 1141
rect 24099 1107 24133 1141
rect 23038 1013 23072 1015
rect 23038 981 23072 1013
rect 23038 911 23072 943
rect 23038 909 23072 911
rect 23126 1013 23160 1015
rect 23126 981 23160 1013
rect 23684 1013 23718 1015
rect 23398 949 23432 983
rect 23684 981 23718 1013
rect 23126 911 23160 943
rect 23126 909 23160 911
rect 23684 911 23718 943
rect 23684 909 23718 911
rect 23254 853 23288 855
rect 23254 821 23288 853
rect 23082 781 23116 815
rect 22373 561 22407 595
rect 22465 561 22499 595
rect 22557 561 22591 595
rect 23254 751 23288 783
rect 23254 749 23288 751
rect 23350 853 23384 855
rect 23350 821 23384 853
rect 23350 751 23384 783
rect 23350 749 23384 751
rect 24261 1105 24295 1139
rect 24353 1105 24387 1139
rect 24445 1105 24479 1139
rect 23772 1013 23806 1015
rect 23772 981 23806 1013
rect 23772 911 23806 943
rect 23772 909 23806 911
rect 24607 1099 24641 1133
rect 24699 1099 24733 1133
rect 24791 1099 24825 1133
rect 24970 1109 25004 1143
rect 23446 853 23480 855
rect 23446 821 23480 853
rect 23446 751 23480 783
rect 23728 781 23762 815
rect 23446 749 23480 751
rect 24267 793 24269 826
rect 24269 793 24301 826
rect 24267 792 24301 793
rect 25616 1109 25650 1143
rect 24460 804 24494 838
rect 23302 621 23336 655
rect 22719 555 22753 589
rect 22811 555 22845 589
rect 22903 555 22937 589
rect 23054 550 23088 584
rect 23686 578 23720 612
rect 24046 711 24080 728
rect 24046 694 24080 711
rect 24656 821 24690 832
rect 24656 798 24658 821
rect 24658 798 24690 821
rect 19686 386 19720 418
rect 19686 384 19720 386
rect 21382 488 21416 490
rect 21382 456 21416 488
rect 21478 488 21512 490
rect 21478 456 21512 488
rect 21382 386 21416 418
rect 21382 384 21416 386
rect 21478 386 21512 418
rect 21478 384 21512 386
rect 21574 488 21608 490
rect 21574 456 21608 488
rect 23414 540 23448 574
rect 23915 563 23949 597
rect 24007 563 24041 597
rect 24099 563 24133 597
rect 25217 1057 25251 1091
rect 26644 1364 26678 1398
rect 27032 1909 27066 1911
rect 27032 1877 27066 1909
rect 27032 1807 27066 1839
rect 27032 1805 27066 1807
rect 27128 1909 27162 1911
rect 27128 1877 27162 1909
rect 27128 1807 27162 1839
rect 27128 1805 27162 1807
rect 28995 2113 29029 2147
rect 29064 2005 29098 2039
rect 27224 1909 27258 1911
rect 27224 1877 27258 1909
rect 27491 1875 27525 1882
rect 27491 1848 27495 1875
rect 27495 1848 27525 1875
rect 27224 1807 27258 1839
rect 27224 1805 27258 1807
rect 27665 1875 27699 1882
rect 27665 1848 27697 1875
rect 27697 1848 27699 1875
rect 28567 1875 28601 1884
rect 28567 1850 28569 1875
rect 28569 1850 28601 1875
rect 28740 1875 28774 1880
rect 28740 1846 28771 1875
rect 28771 1846 28774 1875
rect 27080 1677 27114 1711
rect 27579 1755 27611 1759
rect 27611 1755 27613 1759
rect 27579 1725 27613 1755
rect 28649 1755 28651 1764
rect 28651 1755 28683 1764
rect 28649 1730 28683 1755
rect 27192 1596 27226 1630
rect 27487 1609 27521 1643
rect 27579 1609 27613 1643
rect 27671 1609 27705 1643
rect 28561 1609 28595 1643
rect 28653 1609 28687 1643
rect 28745 1609 28779 1643
rect 27048 1544 27082 1546
rect 27048 1512 27082 1544
rect 27048 1442 27082 1474
rect 27048 1440 27082 1442
rect 27144 1544 27178 1546
rect 27144 1512 27178 1544
rect 27144 1442 27178 1474
rect 27144 1440 27178 1442
rect 27240 1544 27274 1546
rect 27240 1512 27274 1544
rect 27240 1442 27274 1474
rect 27240 1440 27274 1442
rect 27096 1356 27130 1390
rect 27016 1247 27050 1281
rect 27446 1230 27480 1264
rect 25803 1107 25837 1141
rect 25895 1107 25929 1141
rect 25987 1107 26021 1141
rect 24926 1013 24960 1015
rect 24926 981 24960 1013
rect 24926 911 24960 943
rect 24926 909 24960 911
rect 25014 1013 25048 1015
rect 25014 981 25048 1013
rect 25572 1013 25606 1015
rect 25286 949 25320 983
rect 25572 981 25606 1013
rect 25014 911 25048 943
rect 25014 909 25048 911
rect 25572 911 25606 943
rect 25572 909 25606 911
rect 25142 853 25176 855
rect 25142 821 25176 853
rect 24970 781 25004 815
rect 24261 561 24295 595
rect 24353 561 24387 595
rect 24445 561 24479 595
rect 25142 751 25176 783
rect 25142 749 25176 751
rect 25238 853 25272 855
rect 25238 821 25272 853
rect 25238 751 25272 783
rect 25238 749 25272 751
rect 26149 1105 26183 1139
rect 26241 1105 26275 1139
rect 26333 1105 26367 1139
rect 25660 1013 25694 1015
rect 25660 981 25694 1013
rect 25660 911 25694 943
rect 25660 909 25694 911
rect 26495 1099 26529 1133
rect 26587 1099 26621 1133
rect 26679 1099 26713 1133
rect 26858 1109 26892 1143
rect 25334 853 25368 855
rect 25334 821 25368 853
rect 25334 751 25368 783
rect 25616 781 25650 815
rect 25334 749 25368 751
rect 26155 793 26157 826
rect 26157 793 26189 826
rect 26155 792 26189 793
rect 27504 1109 27538 1143
rect 26348 804 26382 838
rect 25190 621 25224 655
rect 24607 555 24641 589
rect 24699 555 24733 589
rect 24791 555 24825 589
rect 24942 550 24976 584
rect 25574 578 25608 612
rect 25934 711 25968 728
rect 25934 694 25968 711
rect 26544 821 26578 832
rect 26544 798 26546 821
rect 26546 798 26578 821
rect 21574 386 21608 418
rect 21574 384 21608 386
rect 23270 488 23304 490
rect 23270 456 23304 488
rect 23366 488 23400 490
rect 23366 456 23400 488
rect 23270 386 23304 418
rect 23270 384 23304 386
rect 23366 386 23400 418
rect 23366 384 23400 386
rect 23462 488 23496 490
rect 23462 456 23496 488
rect 25302 540 25336 574
rect 25803 563 25837 597
rect 25895 563 25929 597
rect 25987 563 26021 597
rect 27105 1057 27139 1091
rect 28532 1364 28566 1398
rect 28920 1909 28954 1911
rect 28920 1877 28954 1909
rect 28920 1807 28954 1839
rect 28920 1805 28954 1807
rect 29016 1909 29050 1911
rect 29016 1877 29050 1909
rect 29016 1807 29050 1839
rect 29016 1805 29050 1807
rect 30883 2113 30917 2147
rect 30952 2005 30986 2039
rect 29112 1909 29146 1911
rect 29112 1877 29146 1909
rect 29379 1875 29413 1882
rect 29379 1848 29383 1875
rect 29383 1848 29413 1875
rect 29112 1807 29146 1839
rect 29112 1805 29146 1807
rect 29553 1875 29587 1882
rect 29553 1848 29585 1875
rect 29585 1848 29587 1875
rect 30455 1875 30489 1884
rect 30455 1850 30457 1875
rect 30457 1850 30489 1875
rect 30628 1875 30662 1880
rect 30628 1846 30659 1875
rect 30659 1846 30662 1875
rect 28968 1677 29002 1711
rect 29467 1755 29499 1759
rect 29499 1755 29501 1759
rect 29467 1725 29501 1755
rect 30537 1755 30539 1764
rect 30539 1755 30571 1764
rect 30537 1730 30571 1755
rect 29080 1596 29114 1630
rect 29375 1609 29409 1643
rect 29467 1609 29501 1643
rect 29559 1609 29593 1643
rect 30449 1609 30483 1643
rect 30541 1609 30575 1643
rect 30633 1609 30667 1643
rect 28936 1544 28970 1546
rect 28936 1512 28970 1544
rect 28936 1442 28970 1474
rect 28936 1440 28970 1442
rect 29032 1544 29066 1546
rect 29032 1512 29066 1544
rect 29032 1442 29066 1474
rect 29032 1440 29066 1442
rect 29128 1544 29162 1546
rect 29128 1512 29162 1544
rect 29128 1442 29162 1474
rect 29128 1440 29162 1442
rect 28984 1356 29018 1390
rect 28904 1247 28938 1281
rect 29334 1230 29368 1264
rect 27691 1107 27725 1141
rect 27783 1107 27817 1141
rect 27875 1107 27909 1141
rect 26814 1013 26848 1015
rect 26814 981 26848 1013
rect 26814 911 26848 943
rect 26814 909 26848 911
rect 26902 1013 26936 1015
rect 26902 981 26936 1013
rect 27460 1013 27494 1015
rect 27174 949 27208 983
rect 27460 981 27494 1013
rect 26902 911 26936 943
rect 26902 909 26936 911
rect 27460 911 27494 943
rect 27460 909 27494 911
rect 27030 853 27064 855
rect 27030 821 27064 853
rect 26858 781 26892 815
rect 26149 561 26183 595
rect 26241 561 26275 595
rect 26333 561 26367 595
rect 27030 751 27064 783
rect 27030 749 27064 751
rect 27126 853 27160 855
rect 27126 821 27160 853
rect 27126 751 27160 783
rect 27126 749 27160 751
rect 28037 1105 28071 1139
rect 28129 1105 28163 1139
rect 28221 1105 28255 1139
rect 27548 1013 27582 1015
rect 27548 981 27582 1013
rect 27548 911 27582 943
rect 27548 909 27582 911
rect 28383 1099 28417 1133
rect 28475 1099 28509 1133
rect 28567 1099 28601 1133
rect 28746 1109 28780 1143
rect 27222 853 27256 855
rect 27222 821 27256 853
rect 27222 751 27256 783
rect 27504 781 27538 815
rect 27222 749 27256 751
rect 28043 793 28045 826
rect 28045 793 28077 826
rect 28043 792 28077 793
rect 29392 1109 29426 1143
rect 28236 804 28270 838
rect 27078 621 27112 655
rect 26495 555 26529 589
rect 26587 555 26621 589
rect 26679 555 26713 589
rect 26830 550 26864 584
rect 27462 578 27496 612
rect 27822 711 27856 728
rect 27822 694 27856 711
rect 28432 821 28466 832
rect 28432 798 28434 821
rect 28434 798 28466 821
rect 23462 386 23496 418
rect 23462 384 23496 386
rect 25158 488 25192 490
rect 25158 456 25192 488
rect 25254 488 25288 490
rect 25254 456 25288 488
rect 25158 386 25192 418
rect 25158 384 25192 386
rect 25254 386 25288 418
rect 25254 384 25288 386
rect 25350 488 25384 490
rect 25350 456 25384 488
rect 27190 540 27224 574
rect 27691 563 27725 597
rect 27783 563 27817 597
rect 27875 563 27909 597
rect 28993 1057 29027 1091
rect 30420 1364 30454 1398
rect 30808 1909 30842 1911
rect 30808 1877 30842 1909
rect 30808 1807 30842 1839
rect 30808 1805 30842 1807
rect 30904 1909 30938 1911
rect 30904 1877 30938 1909
rect 30904 1807 30938 1839
rect 30904 1805 30938 1807
rect 32771 2113 32805 2147
rect 32840 2005 32874 2039
rect 31000 1909 31034 1911
rect 31000 1877 31034 1909
rect 31267 1875 31301 1882
rect 31267 1848 31271 1875
rect 31271 1848 31301 1875
rect 31000 1807 31034 1839
rect 31000 1805 31034 1807
rect 31441 1875 31475 1882
rect 31441 1848 31473 1875
rect 31473 1848 31475 1875
rect 32343 1875 32377 1884
rect 32343 1850 32345 1875
rect 32345 1850 32377 1875
rect 32516 1875 32550 1880
rect 32516 1846 32547 1875
rect 32547 1846 32550 1875
rect 30856 1677 30890 1711
rect 31355 1755 31387 1759
rect 31387 1755 31389 1759
rect 31355 1725 31389 1755
rect 32425 1755 32427 1764
rect 32427 1755 32459 1764
rect 32425 1730 32459 1755
rect 30968 1596 31002 1630
rect 31263 1609 31297 1643
rect 31355 1609 31389 1643
rect 31447 1609 31481 1643
rect 32337 1609 32371 1643
rect 32429 1609 32463 1643
rect 32521 1609 32555 1643
rect 30824 1544 30858 1546
rect 30824 1512 30858 1544
rect 30824 1442 30858 1474
rect 30824 1440 30858 1442
rect 30920 1544 30954 1546
rect 30920 1512 30954 1544
rect 30920 1442 30954 1474
rect 30920 1440 30954 1442
rect 31016 1544 31050 1546
rect 31016 1512 31050 1544
rect 31016 1442 31050 1474
rect 31016 1440 31050 1442
rect 30872 1356 30906 1390
rect 30792 1247 30826 1281
rect 31222 1230 31256 1264
rect 29579 1107 29613 1141
rect 29671 1107 29705 1141
rect 29763 1107 29797 1141
rect 28702 1013 28736 1015
rect 28702 981 28736 1013
rect 28702 911 28736 943
rect 28702 909 28736 911
rect 28790 1013 28824 1015
rect 28790 981 28824 1013
rect 29348 1013 29382 1015
rect 29062 949 29096 983
rect 29348 981 29382 1013
rect 28790 911 28824 943
rect 28790 909 28824 911
rect 29348 911 29382 943
rect 29348 909 29382 911
rect 28918 853 28952 855
rect 28918 821 28952 853
rect 28746 781 28780 815
rect 28037 561 28071 595
rect 28129 561 28163 595
rect 28221 561 28255 595
rect 28918 751 28952 783
rect 28918 749 28952 751
rect 29014 853 29048 855
rect 29014 821 29048 853
rect 29014 751 29048 783
rect 29014 749 29048 751
rect 29925 1105 29959 1139
rect 30017 1105 30051 1139
rect 30109 1105 30143 1139
rect 29436 1013 29470 1015
rect 29436 981 29470 1013
rect 29436 911 29470 943
rect 29436 909 29470 911
rect 30271 1099 30305 1133
rect 30363 1099 30397 1133
rect 30455 1099 30489 1133
rect 30634 1109 30668 1143
rect 29110 853 29144 855
rect 29110 821 29144 853
rect 29110 751 29144 783
rect 29392 781 29426 815
rect 29110 749 29144 751
rect 29931 793 29933 826
rect 29933 793 29965 826
rect 29931 792 29965 793
rect 31280 1109 31314 1143
rect 30124 804 30158 838
rect 28966 621 29000 655
rect 28383 555 28417 589
rect 28475 555 28509 589
rect 28567 555 28601 589
rect 28718 550 28752 584
rect 29350 578 29384 612
rect 29710 711 29744 728
rect 29710 694 29744 711
rect 30320 821 30354 832
rect 30320 798 30322 821
rect 30322 798 30354 821
rect 25350 386 25384 418
rect 25350 384 25384 386
rect 27046 488 27080 490
rect 27046 456 27080 488
rect 27142 488 27176 490
rect 27142 456 27176 488
rect 27046 386 27080 418
rect 27046 384 27080 386
rect 27142 386 27176 418
rect 27142 384 27176 386
rect 27238 488 27272 490
rect 27238 456 27272 488
rect 29078 540 29112 574
rect 29579 563 29613 597
rect 29671 563 29705 597
rect 29763 563 29797 597
rect 30881 1057 30915 1091
rect 32308 1364 32342 1398
rect 32696 1909 32730 1911
rect 32696 1877 32730 1909
rect 32696 1807 32730 1839
rect 32696 1805 32730 1807
rect 32792 1909 32826 1911
rect 32792 1877 32826 1909
rect 32792 1807 32826 1839
rect 32792 1805 32826 1807
rect 34659 2113 34693 2147
rect 34728 2005 34762 2039
rect 32888 1909 32922 1911
rect 32888 1877 32922 1909
rect 33155 1875 33189 1882
rect 33155 1848 33159 1875
rect 33159 1848 33189 1875
rect 32888 1807 32922 1839
rect 32888 1805 32922 1807
rect 33329 1875 33363 1882
rect 33329 1848 33361 1875
rect 33361 1848 33363 1875
rect 34231 1875 34265 1884
rect 34231 1850 34233 1875
rect 34233 1850 34265 1875
rect 34404 1875 34438 1880
rect 34404 1846 34435 1875
rect 34435 1846 34438 1875
rect 32744 1677 32778 1711
rect 33243 1755 33275 1759
rect 33275 1755 33277 1759
rect 33243 1725 33277 1755
rect 34313 1755 34315 1764
rect 34315 1755 34347 1764
rect 34313 1730 34347 1755
rect 32856 1596 32890 1630
rect 33151 1609 33185 1643
rect 33243 1609 33277 1643
rect 33335 1609 33369 1643
rect 34225 1609 34259 1643
rect 34317 1609 34351 1643
rect 34409 1609 34443 1643
rect 32712 1544 32746 1546
rect 32712 1512 32746 1544
rect 32712 1442 32746 1474
rect 32712 1440 32746 1442
rect 32808 1544 32842 1546
rect 32808 1512 32842 1544
rect 32808 1442 32842 1474
rect 32808 1440 32842 1442
rect 32904 1544 32938 1546
rect 32904 1512 32938 1544
rect 32904 1442 32938 1474
rect 32904 1440 32938 1442
rect 32760 1356 32794 1390
rect 32680 1247 32714 1281
rect 33110 1230 33144 1264
rect 31467 1107 31501 1141
rect 31559 1107 31593 1141
rect 31651 1107 31685 1141
rect 30590 1013 30624 1015
rect 30590 981 30624 1013
rect 30590 911 30624 943
rect 30590 909 30624 911
rect 30678 1013 30712 1015
rect 30678 981 30712 1013
rect 31236 1013 31270 1015
rect 30950 949 30984 983
rect 31236 981 31270 1013
rect 30678 911 30712 943
rect 30678 909 30712 911
rect 31236 911 31270 943
rect 31236 909 31270 911
rect 30806 853 30840 855
rect 30806 821 30840 853
rect 30634 781 30668 815
rect 29925 561 29959 595
rect 30017 561 30051 595
rect 30109 561 30143 595
rect 30806 751 30840 783
rect 30806 749 30840 751
rect 30902 853 30936 855
rect 30902 821 30936 853
rect 30902 751 30936 783
rect 30902 749 30936 751
rect 31813 1105 31847 1139
rect 31905 1105 31939 1139
rect 31997 1105 32031 1139
rect 31324 1013 31358 1015
rect 31324 981 31358 1013
rect 31324 911 31358 943
rect 31324 909 31358 911
rect 32159 1099 32193 1133
rect 32251 1099 32285 1133
rect 32343 1099 32377 1133
rect 32522 1109 32556 1143
rect 30998 853 31032 855
rect 30998 821 31032 853
rect 30998 751 31032 783
rect 31280 781 31314 815
rect 30998 749 31032 751
rect 31819 793 31821 826
rect 31821 793 31853 826
rect 31819 792 31853 793
rect 33168 1109 33202 1143
rect 32012 804 32046 838
rect 30854 621 30888 655
rect 30271 555 30305 589
rect 30363 555 30397 589
rect 30455 555 30489 589
rect 30606 550 30640 584
rect 31238 578 31272 612
rect 31598 711 31632 728
rect 31598 694 31632 711
rect 32208 821 32242 832
rect 32208 798 32210 821
rect 32210 798 32242 821
rect 27238 386 27272 418
rect 27238 384 27272 386
rect 28934 488 28968 490
rect 28934 456 28968 488
rect 29030 488 29064 490
rect 29030 456 29064 488
rect 28934 386 28968 418
rect 28934 384 28968 386
rect 29030 386 29064 418
rect 29030 384 29064 386
rect 29126 488 29160 490
rect 29126 456 29160 488
rect 30966 540 31000 574
rect 31467 563 31501 597
rect 31559 563 31593 597
rect 31651 563 31685 597
rect 32769 1057 32803 1091
rect 34196 1364 34230 1398
rect 34584 1909 34618 1911
rect 34584 1877 34618 1909
rect 34584 1807 34618 1839
rect 34584 1805 34618 1807
rect 34680 1909 34714 1911
rect 34680 1877 34714 1909
rect 34680 1807 34714 1839
rect 34680 1805 34714 1807
rect 36547 2113 36581 2147
rect 36616 2005 36650 2039
rect 34776 1909 34810 1911
rect 34776 1877 34810 1909
rect 35043 1875 35077 1882
rect 35043 1848 35047 1875
rect 35047 1848 35077 1875
rect 34776 1807 34810 1839
rect 34776 1805 34810 1807
rect 35217 1875 35251 1882
rect 35217 1848 35249 1875
rect 35249 1848 35251 1875
rect 36119 1875 36153 1884
rect 36119 1850 36121 1875
rect 36121 1850 36153 1875
rect 36292 1875 36326 1880
rect 36292 1846 36323 1875
rect 36323 1846 36326 1875
rect 34632 1677 34666 1711
rect 35131 1755 35163 1759
rect 35163 1755 35165 1759
rect 35131 1725 35165 1755
rect 36201 1755 36203 1764
rect 36203 1755 36235 1764
rect 36201 1730 36235 1755
rect 34744 1596 34778 1630
rect 35039 1609 35073 1643
rect 35131 1609 35165 1643
rect 35223 1609 35257 1643
rect 36113 1609 36147 1643
rect 36205 1609 36239 1643
rect 36297 1609 36331 1643
rect 34600 1544 34634 1546
rect 34600 1512 34634 1544
rect 34600 1442 34634 1474
rect 34600 1440 34634 1442
rect 34696 1544 34730 1546
rect 34696 1512 34730 1544
rect 34696 1442 34730 1474
rect 34696 1440 34730 1442
rect 34792 1544 34826 1546
rect 34792 1512 34826 1544
rect 34792 1442 34826 1474
rect 34792 1440 34826 1442
rect 34648 1356 34682 1390
rect 34568 1247 34602 1281
rect 34998 1230 35032 1264
rect 33355 1107 33389 1141
rect 33447 1107 33481 1141
rect 33539 1107 33573 1141
rect 32478 1013 32512 1015
rect 32478 981 32512 1013
rect 32478 911 32512 943
rect 32478 909 32512 911
rect 32566 1013 32600 1015
rect 32566 981 32600 1013
rect 33124 1013 33158 1015
rect 32838 949 32872 983
rect 33124 981 33158 1013
rect 32566 911 32600 943
rect 32566 909 32600 911
rect 33124 911 33158 943
rect 33124 909 33158 911
rect 32694 853 32728 855
rect 32694 821 32728 853
rect 32522 781 32556 815
rect 31813 561 31847 595
rect 31905 561 31939 595
rect 31997 561 32031 595
rect 32694 751 32728 783
rect 32694 749 32728 751
rect 32790 853 32824 855
rect 32790 821 32824 853
rect 32790 751 32824 783
rect 32790 749 32824 751
rect 33701 1105 33735 1139
rect 33793 1105 33827 1139
rect 33885 1105 33919 1139
rect 33212 1013 33246 1015
rect 33212 981 33246 1013
rect 33212 911 33246 943
rect 33212 909 33246 911
rect 34047 1099 34081 1133
rect 34139 1099 34173 1133
rect 34231 1099 34265 1133
rect 34410 1109 34444 1143
rect 32886 853 32920 855
rect 32886 821 32920 853
rect 32886 751 32920 783
rect 33168 781 33202 815
rect 32886 749 32920 751
rect 33707 793 33709 826
rect 33709 793 33741 826
rect 33707 792 33741 793
rect 35056 1109 35090 1143
rect 33900 804 33934 838
rect 32742 621 32776 655
rect 32159 555 32193 589
rect 32251 555 32285 589
rect 32343 555 32377 589
rect 32494 550 32528 584
rect 33126 578 33160 612
rect 33486 711 33520 728
rect 33486 694 33520 711
rect 34096 821 34130 832
rect 34096 798 34098 821
rect 34098 798 34130 821
rect 29126 386 29160 418
rect 29126 384 29160 386
rect 30822 488 30856 490
rect 30822 456 30856 488
rect 30918 488 30952 490
rect 30918 456 30952 488
rect 30822 386 30856 418
rect 30822 384 30856 386
rect 30918 386 30952 418
rect 30918 384 30952 386
rect 31014 488 31048 490
rect 31014 456 31048 488
rect 32854 540 32888 574
rect 33355 563 33389 597
rect 33447 563 33481 597
rect 33539 563 33573 597
rect 34657 1057 34691 1091
rect 36084 1364 36118 1398
rect 36472 1909 36506 1911
rect 36472 1877 36506 1909
rect 36472 1807 36506 1839
rect 36472 1805 36506 1807
rect 36568 1909 36602 1911
rect 36568 1877 36602 1909
rect 36568 1807 36602 1839
rect 36568 1805 36602 1807
rect 38435 2113 38469 2147
rect 38504 2005 38538 2039
rect 36664 1909 36698 1911
rect 36664 1877 36698 1909
rect 36931 1875 36965 1882
rect 36931 1848 36935 1875
rect 36935 1848 36965 1875
rect 36664 1807 36698 1839
rect 36664 1805 36698 1807
rect 37105 1875 37139 1882
rect 37105 1848 37137 1875
rect 37137 1848 37139 1875
rect 38007 1875 38041 1884
rect 38007 1850 38009 1875
rect 38009 1850 38041 1875
rect 38180 1875 38214 1880
rect 38180 1846 38211 1875
rect 38211 1846 38214 1875
rect 36520 1677 36554 1711
rect 37019 1755 37051 1759
rect 37051 1755 37053 1759
rect 37019 1725 37053 1755
rect 38089 1755 38091 1764
rect 38091 1755 38123 1764
rect 38089 1730 38123 1755
rect 36632 1596 36666 1630
rect 36927 1609 36961 1643
rect 37019 1609 37053 1643
rect 37111 1609 37145 1643
rect 38001 1609 38035 1643
rect 38093 1609 38127 1643
rect 38185 1609 38219 1643
rect 36488 1544 36522 1546
rect 36488 1512 36522 1544
rect 36488 1442 36522 1474
rect 36488 1440 36522 1442
rect 36584 1544 36618 1546
rect 36584 1512 36618 1544
rect 36584 1442 36618 1474
rect 36584 1440 36618 1442
rect 36680 1544 36714 1546
rect 36680 1512 36714 1544
rect 36680 1442 36714 1474
rect 36680 1440 36714 1442
rect 36536 1356 36570 1390
rect 36456 1247 36490 1281
rect 36886 1230 36920 1264
rect 35243 1107 35277 1141
rect 35335 1107 35369 1141
rect 35427 1107 35461 1141
rect 34366 1013 34400 1015
rect 34366 981 34400 1013
rect 34366 911 34400 943
rect 34366 909 34400 911
rect 34454 1013 34488 1015
rect 34454 981 34488 1013
rect 35012 1013 35046 1015
rect 34726 949 34760 983
rect 35012 981 35046 1013
rect 34454 911 34488 943
rect 34454 909 34488 911
rect 35012 911 35046 943
rect 35012 909 35046 911
rect 34582 853 34616 855
rect 34582 821 34616 853
rect 34410 781 34444 815
rect 33701 561 33735 595
rect 33793 561 33827 595
rect 33885 561 33919 595
rect 34582 751 34616 783
rect 34582 749 34616 751
rect 34678 853 34712 855
rect 34678 821 34712 853
rect 34678 751 34712 783
rect 34678 749 34712 751
rect 35589 1105 35623 1139
rect 35681 1105 35715 1139
rect 35773 1105 35807 1139
rect 35100 1013 35134 1015
rect 35100 981 35134 1013
rect 35100 911 35134 943
rect 35100 909 35134 911
rect 35935 1099 35969 1133
rect 36027 1099 36061 1133
rect 36119 1099 36153 1133
rect 36298 1109 36332 1143
rect 34774 853 34808 855
rect 34774 821 34808 853
rect 34774 751 34808 783
rect 35056 781 35090 815
rect 34774 749 34808 751
rect 35595 793 35597 826
rect 35597 793 35629 826
rect 35595 792 35629 793
rect 36944 1109 36978 1143
rect 35788 804 35822 838
rect 34630 621 34664 655
rect 34047 555 34081 589
rect 34139 555 34173 589
rect 34231 555 34265 589
rect 34382 550 34416 584
rect 35014 578 35048 612
rect 35374 711 35408 728
rect 35374 694 35408 711
rect 35984 821 36018 832
rect 35984 798 35986 821
rect 35986 798 36018 821
rect 31014 386 31048 418
rect 31014 384 31048 386
rect 32710 488 32744 490
rect 32710 456 32744 488
rect 32806 488 32840 490
rect 32806 456 32840 488
rect 32710 386 32744 418
rect 32710 384 32744 386
rect 32806 386 32840 418
rect 32806 384 32840 386
rect 32902 488 32936 490
rect 32902 456 32936 488
rect 34742 540 34776 574
rect 35243 563 35277 597
rect 35335 563 35369 597
rect 35427 563 35461 597
rect 36545 1057 36579 1091
rect 37972 1364 38006 1398
rect 38360 1909 38394 1911
rect 38360 1877 38394 1909
rect 38360 1807 38394 1839
rect 38360 1805 38394 1807
rect 38456 1909 38490 1911
rect 38456 1877 38490 1909
rect 38456 1807 38490 1839
rect 38456 1805 38490 1807
rect 40323 2113 40357 2147
rect 40392 2005 40426 2039
rect 38552 1909 38586 1911
rect 38552 1877 38586 1909
rect 38819 1875 38853 1882
rect 38819 1848 38823 1875
rect 38823 1848 38853 1875
rect 38552 1807 38586 1839
rect 38552 1805 38586 1807
rect 38993 1875 39027 1882
rect 38993 1848 39025 1875
rect 39025 1848 39027 1875
rect 39895 1875 39929 1884
rect 39895 1850 39897 1875
rect 39897 1850 39929 1875
rect 40068 1875 40102 1880
rect 40068 1846 40099 1875
rect 40099 1846 40102 1875
rect 38408 1677 38442 1711
rect 38907 1755 38939 1759
rect 38939 1755 38941 1759
rect 38907 1725 38941 1755
rect 39977 1755 39979 1764
rect 39979 1755 40011 1764
rect 39977 1730 40011 1755
rect 38520 1596 38554 1630
rect 38815 1609 38849 1643
rect 38907 1609 38941 1643
rect 38999 1609 39033 1643
rect 39889 1609 39923 1643
rect 39981 1609 40015 1643
rect 40073 1609 40107 1643
rect 38376 1544 38410 1546
rect 38376 1512 38410 1544
rect 38376 1442 38410 1474
rect 38376 1440 38410 1442
rect 38472 1544 38506 1546
rect 38472 1512 38506 1544
rect 38472 1442 38506 1474
rect 38472 1440 38506 1442
rect 38568 1544 38602 1546
rect 38568 1512 38602 1544
rect 38568 1442 38602 1474
rect 38568 1440 38602 1442
rect 38424 1356 38458 1390
rect 38344 1247 38378 1281
rect 38774 1230 38808 1264
rect 37131 1107 37165 1141
rect 37223 1107 37257 1141
rect 37315 1107 37349 1141
rect 36254 1013 36288 1015
rect 36254 981 36288 1013
rect 36254 911 36288 943
rect 36254 909 36288 911
rect 36342 1013 36376 1015
rect 36342 981 36376 1013
rect 36900 1013 36934 1015
rect 36614 949 36648 983
rect 36900 981 36934 1013
rect 36342 911 36376 943
rect 36342 909 36376 911
rect 36900 911 36934 943
rect 36900 909 36934 911
rect 36470 853 36504 855
rect 36470 821 36504 853
rect 36298 781 36332 815
rect 35589 561 35623 595
rect 35681 561 35715 595
rect 35773 561 35807 595
rect 36470 751 36504 783
rect 36470 749 36504 751
rect 36566 853 36600 855
rect 36566 821 36600 853
rect 36566 751 36600 783
rect 36566 749 36600 751
rect 37477 1105 37511 1139
rect 37569 1105 37603 1139
rect 37661 1105 37695 1139
rect 36988 1013 37022 1015
rect 36988 981 37022 1013
rect 36988 911 37022 943
rect 36988 909 37022 911
rect 37823 1099 37857 1133
rect 37915 1099 37949 1133
rect 38007 1099 38041 1133
rect 38186 1109 38220 1143
rect 36662 853 36696 855
rect 36662 821 36696 853
rect 36662 751 36696 783
rect 36944 781 36978 815
rect 36662 749 36696 751
rect 37483 793 37485 826
rect 37485 793 37517 826
rect 37483 792 37517 793
rect 38832 1109 38866 1143
rect 37676 804 37710 838
rect 36518 621 36552 655
rect 35935 555 35969 589
rect 36027 555 36061 589
rect 36119 555 36153 589
rect 36270 550 36304 584
rect 36902 578 36936 612
rect 37262 711 37296 728
rect 37262 694 37296 711
rect 37872 821 37906 832
rect 37872 798 37874 821
rect 37874 798 37906 821
rect 32902 386 32936 418
rect 32902 384 32936 386
rect 34598 488 34632 490
rect 34598 456 34632 488
rect 34694 488 34728 490
rect 34694 456 34728 488
rect 34598 386 34632 418
rect 34598 384 34632 386
rect 34694 386 34728 418
rect 34694 384 34728 386
rect 34790 488 34824 490
rect 34790 456 34824 488
rect 36630 540 36664 574
rect 37131 563 37165 597
rect 37223 563 37257 597
rect 37315 563 37349 597
rect 38433 1057 38467 1091
rect 39860 1364 39894 1398
rect 40248 1909 40282 1911
rect 40248 1877 40282 1909
rect 40248 1807 40282 1839
rect 40248 1805 40282 1807
rect 40344 1909 40378 1911
rect 40344 1877 40378 1909
rect 40344 1807 40378 1839
rect 40344 1805 40378 1807
rect 42211 2113 42245 2147
rect 42280 2005 42314 2039
rect 40440 1909 40474 1911
rect 40440 1877 40474 1909
rect 40707 1875 40741 1882
rect 40707 1848 40711 1875
rect 40711 1848 40741 1875
rect 40440 1807 40474 1839
rect 40440 1805 40474 1807
rect 40881 1875 40915 1882
rect 40881 1848 40913 1875
rect 40913 1848 40915 1875
rect 41783 1875 41817 1884
rect 41783 1850 41785 1875
rect 41785 1850 41817 1875
rect 41956 1875 41990 1880
rect 41956 1846 41987 1875
rect 41987 1846 41990 1875
rect 40296 1677 40330 1711
rect 40795 1755 40827 1759
rect 40827 1755 40829 1759
rect 40795 1725 40829 1755
rect 41865 1755 41867 1764
rect 41867 1755 41899 1764
rect 41865 1730 41899 1755
rect 40408 1596 40442 1630
rect 40703 1609 40737 1643
rect 40795 1609 40829 1643
rect 40887 1609 40921 1643
rect 41777 1609 41811 1643
rect 41869 1609 41903 1643
rect 41961 1609 41995 1643
rect 40264 1544 40298 1546
rect 40264 1512 40298 1544
rect 40264 1442 40298 1474
rect 40264 1440 40298 1442
rect 40360 1544 40394 1546
rect 40360 1512 40394 1544
rect 40360 1442 40394 1474
rect 40360 1440 40394 1442
rect 40456 1544 40490 1546
rect 40456 1512 40490 1544
rect 40456 1442 40490 1474
rect 40456 1440 40490 1442
rect 40312 1356 40346 1390
rect 40232 1247 40266 1281
rect 40662 1230 40696 1264
rect 39019 1107 39053 1141
rect 39111 1107 39145 1141
rect 39203 1107 39237 1141
rect 38142 1013 38176 1015
rect 38142 981 38176 1013
rect 38142 911 38176 943
rect 38142 909 38176 911
rect 38230 1013 38264 1015
rect 38230 981 38264 1013
rect 38788 1013 38822 1015
rect 38502 949 38536 983
rect 38788 981 38822 1013
rect 38230 911 38264 943
rect 38230 909 38264 911
rect 38788 911 38822 943
rect 38788 909 38822 911
rect 38358 853 38392 855
rect 38358 821 38392 853
rect 38186 781 38220 815
rect 37477 561 37511 595
rect 37569 561 37603 595
rect 37661 561 37695 595
rect 38358 751 38392 783
rect 38358 749 38392 751
rect 38454 853 38488 855
rect 38454 821 38488 853
rect 38454 751 38488 783
rect 38454 749 38488 751
rect 39365 1105 39399 1139
rect 39457 1105 39491 1139
rect 39549 1105 39583 1139
rect 38876 1013 38910 1015
rect 38876 981 38910 1013
rect 38876 911 38910 943
rect 38876 909 38910 911
rect 39711 1099 39745 1133
rect 39803 1099 39837 1133
rect 39895 1099 39929 1133
rect 40074 1109 40108 1143
rect 38550 853 38584 855
rect 38550 821 38584 853
rect 38550 751 38584 783
rect 38832 781 38866 815
rect 38550 749 38584 751
rect 39371 793 39373 826
rect 39373 793 39405 826
rect 39371 792 39405 793
rect 40720 1109 40754 1143
rect 39564 804 39598 838
rect 38406 621 38440 655
rect 37823 555 37857 589
rect 37915 555 37949 589
rect 38007 555 38041 589
rect 38158 550 38192 584
rect 38790 578 38824 612
rect 39150 711 39184 728
rect 39150 694 39184 711
rect 39760 821 39794 832
rect 39760 798 39762 821
rect 39762 798 39794 821
rect 34790 386 34824 418
rect 34790 384 34824 386
rect 36486 488 36520 490
rect 36486 456 36520 488
rect 36582 488 36616 490
rect 36582 456 36616 488
rect 36486 386 36520 418
rect 36486 384 36520 386
rect 36582 386 36616 418
rect 36582 384 36616 386
rect 36678 488 36712 490
rect 36678 456 36712 488
rect 38518 540 38552 574
rect 39019 563 39053 597
rect 39111 563 39145 597
rect 39203 563 39237 597
rect 40321 1057 40355 1091
rect 41748 1364 41782 1398
rect 42136 1909 42170 1911
rect 42136 1877 42170 1909
rect 42136 1807 42170 1839
rect 42136 1805 42170 1807
rect 42232 1909 42266 1911
rect 42232 1877 42266 1909
rect 42232 1807 42266 1839
rect 42232 1805 42266 1807
rect 44099 2113 44133 2147
rect 44168 2005 44202 2039
rect 42328 1909 42362 1911
rect 42328 1877 42362 1909
rect 42595 1875 42629 1882
rect 42595 1848 42599 1875
rect 42599 1848 42629 1875
rect 42328 1807 42362 1839
rect 42328 1805 42362 1807
rect 42769 1875 42803 1882
rect 42769 1848 42801 1875
rect 42801 1848 42803 1875
rect 43671 1875 43705 1884
rect 43671 1850 43673 1875
rect 43673 1850 43705 1875
rect 43844 1875 43878 1880
rect 43844 1846 43875 1875
rect 43875 1846 43878 1875
rect 42184 1677 42218 1711
rect 42683 1755 42715 1759
rect 42715 1755 42717 1759
rect 42683 1725 42717 1755
rect 43753 1755 43755 1764
rect 43755 1755 43787 1764
rect 43753 1730 43787 1755
rect 42296 1596 42330 1630
rect 42591 1609 42625 1643
rect 42683 1609 42717 1643
rect 42775 1609 42809 1643
rect 43665 1609 43699 1643
rect 43757 1609 43791 1643
rect 43849 1609 43883 1643
rect 42152 1544 42186 1546
rect 42152 1512 42186 1544
rect 42152 1442 42186 1474
rect 42152 1440 42186 1442
rect 42248 1544 42282 1546
rect 42248 1512 42282 1544
rect 42248 1442 42282 1474
rect 42248 1440 42282 1442
rect 42344 1544 42378 1546
rect 42344 1512 42378 1544
rect 42344 1442 42378 1474
rect 42344 1440 42378 1442
rect 42200 1356 42234 1390
rect 42120 1247 42154 1281
rect 42550 1230 42584 1264
rect 40907 1107 40941 1141
rect 40999 1107 41033 1141
rect 41091 1107 41125 1141
rect 40030 1013 40064 1015
rect 40030 981 40064 1013
rect 40030 911 40064 943
rect 40030 909 40064 911
rect 40118 1013 40152 1015
rect 40118 981 40152 1013
rect 40676 1013 40710 1015
rect 40390 949 40424 983
rect 40676 981 40710 1013
rect 40118 911 40152 943
rect 40118 909 40152 911
rect 40676 911 40710 943
rect 40676 909 40710 911
rect 40246 853 40280 855
rect 40246 821 40280 853
rect 40074 781 40108 815
rect 39365 561 39399 595
rect 39457 561 39491 595
rect 39549 561 39583 595
rect 40246 751 40280 783
rect 40246 749 40280 751
rect 40342 853 40376 855
rect 40342 821 40376 853
rect 40342 751 40376 783
rect 40342 749 40376 751
rect 41253 1105 41287 1139
rect 41345 1105 41379 1139
rect 41437 1105 41471 1139
rect 40764 1013 40798 1015
rect 40764 981 40798 1013
rect 40764 911 40798 943
rect 40764 909 40798 911
rect 41599 1099 41633 1133
rect 41691 1099 41725 1133
rect 41783 1099 41817 1133
rect 41962 1109 41996 1143
rect 40438 853 40472 855
rect 40438 821 40472 853
rect 40438 751 40472 783
rect 40720 781 40754 815
rect 40438 749 40472 751
rect 41259 793 41261 826
rect 41261 793 41293 826
rect 41259 792 41293 793
rect 42608 1109 42642 1143
rect 41452 804 41486 838
rect 40294 621 40328 655
rect 39711 555 39745 589
rect 39803 555 39837 589
rect 39895 555 39929 589
rect 40046 550 40080 584
rect 40678 578 40712 612
rect 41038 711 41072 728
rect 41038 694 41072 711
rect 41648 821 41682 832
rect 41648 798 41650 821
rect 41650 798 41682 821
rect 36678 386 36712 418
rect 36678 384 36712 386
rect 38374 488 38408 490
rect 38374 456 38408 488
rect 38470 488 38504 490
rect 38470 456 38504 488
rect 38374 386 38408 418
rect 38374 384 38408 386
rect 38470 386 38504 418
rect 38470 384 38504 386
rect 38566 488 38600 490
rect 38566 456 38600 488
rect 40406 540 40440 574
rect 40907 563 40941 597
rect 40999 563 41033 597
rect 41091 563 41125 597
rect 42209 1057 42243 1091
rect 43636 1364 43670 1398
rect 44024 1909 44058 1911
rect 44024 1877 44058 1909
rect 44024 1807 44058 1839
rect 44024 1805 44058 1807
rect 44120 1909 44154 1911
rect 44120 1877 44154 1909
rect 44120 1807 44154 1839
rect 44120 1805 44154 1807
rect 45981 2113 46015 2147
rect 46050 2005 46084 2039
rect 44216 1909 44250 1911
rect 44216 1877 44250 1909
rect 44483 1875 44517 1882
rect 44483 1848 44487 1875
rect 44487 1848 44517 1875
rect 44216 1807 44250 1839
rect 44216 1805 44250 1807
rect 44657 1875 44691 1882
rect 44657 1848 44689 1875
rect 44689 1848 44691 1875
rect 45553 1875 45587 1884
rect 45553 1850 45555 1875
rect 45555 1850 45587 1875
rect 45726 1875 45760 1880
rect 45726 1846 45757 1875
rect 45757 1846 45760 1875
rect 44072 1677 44106 1711
rect 44571 1755 44603 1759
rect 44603 1755 44605 1759
rect 44571 1725 44605 1755
rect 45635 1755 45637 1764
rect 45637 1755 45669 1764
rect 45635 1730 45669 1755
rect 44184 1596 44218 1630
rect 44479 1609 44513 1643
rect 44571 1609 44605 1643
rect 44663 1609 44697 1643
rect 45547 1609 45581 1643
rect 45639 1609 45673 1643
rect 45731 1609 45765 1643
rect 44040 1544 44074 1546
rect 44040 1512 44074 1544
rect 44040 1442 44074 1474
rect 44040 1440 44074 1442
rect 44136 1544 44170 1546
rect 44136 1512 44170 1544
rect 44136 1442 44170 1474
rect 44136 1440 44170 1442
rect 44232 1544 44266 1546
rect 44232 1512 44266 1544
rect 44232 1442 44266 1474
rect 44232 1440 44266 1442
rect 44088 1356 44122 1390
rect 44008 1247 44042 1281
rect 44438 1230 44472 1264
rect 42795 1107 42829 1141
rect 42887 1107 42921 1141
rect 42979 1107 43013 1141
rect 41918 1013 41952 1015
rect 41918 981 41952 1013
rect 41918 911 41952 943
rect 41918 909 41952 911
rect 42006 1013 42040 1015
rect 42006 981 42040 1013
rect 42564 1013 42598 1015
rect 42278 949 42312 983
rect 42564 981 42598 1013
rect 42006 911 42040 943
rect 42006 909 42040 911
rect 42564 911 42598 943
rect 42564 909 42598 911
rect 42134 853 42168 855
rect 42134 821 42168 853
rect 41962 781 41996 815
rect 41253 561 41287 595
rect 41345 561 41379 595
rect 41437 561 41471 595
rect 42134 751 42168 783
rect 42134 749 42168 751
rect 42230 853 42264 855
rect 42230 821 42264 853
rect 42230 751 42264 783
rect 42230 749 42264 751
rect 43141 1105 43175 1139
rect 43233 1105 43267 1139
rect 43325 1105 43359 1139
rect 42652 1013 42686 1015
rect 42652 981 42686 1013
rect 42652 911 42686 943
rect 42652 909 42686 911
rect 43487 1099 43521 1133
rect 43579 1099 43613 1133
rect 43671 1099 43705 1133
rect 43850 1109 43884 1143
rect 42326 853 42360 855
rect 42326 821 42360 853
rect 42326 751 42360 783
rect 42608 781 42642 815
rect 42326 749 42360 751
rect 43147 793 43149 826
rect 43149 793 43181 826
rect 43147 792 43181 793
rect 44496 1109 44530 1143
rect 43340 804 43374 838
rect 42182 621 42216 655
rect 41599 555 41633 589
rect 41691 555 41725 589
rect 41783 555 41817 589
rect 41934 550 41968 584
rect 42566 578 42600 612
rect 42926 711 42960 728
rect 42926 694 42960 711
rect 43536 821 43570 832
rect 43536 798 43538 821
rect 43538 798 43570 821
rect 38566 386 38600 418
rect 38566 384 38600 386
rect 40262 488 40296 490
rect 40262 456 40296 488
rect 40358 488 40392 490
rect 40358 456 40392 488
rect 40262 386 40296 418
rect 40262 384 40296 386
rect 40358 386 40392 418
rect 40358 384 40392 386
rect 40454 488 40488 490
rect 40454 456 40488 488
rect 42294 540 42328 574
rect 42795 563 42829 597
rect 42887 563 42921 597
rect 42979 563 43013 597
rect 44097 1057 44131 1091
rect 45518 1364 45552 1398
rect 45906 1909 45940 1911
rect 45906 1877 45940 1909
rect 45906 1807 45940 1839
rect 45906 1805 45940 1807
rect 46002 1909 46036 1911
rect 46002 1877 46036 1909
rect 46002 1807 46036 1839
rect 46002 1805 46036 1807
rect 47869 2113 47903 2147
rect 47938 2005 47972 2039
rect 46098 1909 46132 1911
rect 46098 1877 46132 1909
rect 46365 1875 46399 1882
rect 46365 1848 46369 1875
rect 46369 1848 46399 1875
rect 46098 1807 46132 1839
rect 46098 1805 46132 1807
rect 46539 1875 46573 1882
rect 46539 1848 46571 1875
rect 46571 1848 46573 1875
rect 47441 1875 47475 1884
rect 47441 1850 47443 1875
rect 47443 1850 47475 1875
rect 47614 1875 47648 1880
rect 47614 1846 47645 1875
rect 47645 1846 47648 1875
rect 45954 1677 45988 1711
rect 46453 1755 46485 1759
rect 46485 1755 46487 1759
rect 46453 1725 46487 1755
rect 47523 1755 47525 1764
rect 47525 1755 47557 1764
rect 47523 1730 47557 1755
rect 46066 1596 46100 1630
rect 46361 1609 46395 1643
rect 46453 1609 46487 1643
rect 46545 1609 46579 1643
rect 47435 1609 47469 1643
rect 47527 1609 47561 1643
rect 47619 1609 47653 1643
rect 45922 1544 45956 1546
rect 45922 1512 45956 1544
rect 45922 1442 45956 1474
rect 45922 1440 45956 1442
rect 46018 1544 46052 1546
rect 46018 1512 46052 1544
rect 46018 1442 46052 1474
rect 46018 1440 46052 1442
rect 46114 1544 46148 1546
rect 46114 1512 46148 1544
rect 46114 1442 46148 1474
rect 46114 1440 46148 1442
rect 45970 1356 46004 1390
rect 45890 1247 45924 1281
rect 46320 1230 46354 1264
rect 44683 1107 44717 1141
rect 44775 1107 44809 1141
rect 44867 1107 44901 1141
rect 43806 1013 43840 1015
rect 43806 981 43840 1013
rect 43806 911 43840 943
rect 43806 909 43840 911
rect 43894 1013 43928 1015
rect 43894 981 43928 1013
rect 44452 1013 44486 1015
rect 44166 949 44200 983
rect 44452 981 44486 1013
rect 43894 911 43928 943
rect 43894 909 43928 911
rect 44452 911 44486 943
rect 44452 909 44486 911
rect 44022 853 44056 855
rect 44022 821 44056 853
rect 43850 781 43884 815
rect 43141 561 43175 595
rect 43233 561 43267 595
rect 43325 561 43359 595
rect 44022 751 44056 783
rect 44022 749 44056 751
rect 44118 853 44152 855
rect 44118 821 44152 853
rect 44118 751 44152 783
rect 44118 749 44152 751
rect 45029 1105 45063 1139
rect 45121 1105 45155 1139
rect 45213 1105 45247 1139
rect 44540 1013 44574 1015
rect 44540 981 44574 1013
rect 44540 911 44574 943
rect 44540 909 44574 911
rect 45369 1099 45403 1133
rect 45461 1099 45495 1133
rect 45553 1099 45587 1133
rect 45732 1109 45766 1143
rect 44214 853 44248 855
rect 44214 821 44248 853
rect 44214 751 44248 783
rect 44496 781 44530 815
rect 44214 749 44248 751
rect 45035 793 45037 826
rect 45037 793 45069 826
rect 45035 792 45069 793
rect 46378 1109 46412 1143
rect 45228 804 45262 838
rect 44070 621 44104 655
rect 43487 555 43521 589
rect 43579 555 43613 589
rect 43671 555 43705 589
rect 43822 550 43856 584
rect 44454 578 44488 612
rect 44814 711 44848 728
rect 44814 694 44848 711
rect 45418 821 45452 832
rect 45418 798 45420 821
rect 45420 798 45452 821
rect 40454 386 40488 418
rect 40454 384 40488 386
rect 42150 488 42184 490
rect 42150 456 42184 488
rect 42246 488 42280 490
rect 42246 456 42280 488
rect 42150 386 42184 418
rect 42150 384 42184 386
rect 42246 386 42280 418
rect 42246 384 42280 386
rect 42342 488 42376 490
rect 42342 456 42376 488
rect 44182 540 44216 574
rect 44683 563 44717 597
rect 44775 563 44809 597
rect 44867 563 44901 597
rect 45979 1057 46013 1091
rect 47406 1364 47440 1398
rect 47794 1909 47828 1911
rect 47794 1877 47828 1909
rect 47794 1807 47828 1839
rect 47794 1805 47828 1807
rect 47890 1909 47924 1911
rect 47890 1877 47924 1909
rect 47890 1807 47924 1839
rect 47890 1805 47924 1807
rect 49757 2113 49791 2147
rect 49826 2005 49860 2039
rect 47986 1909 48020 1911
rect 47986 1877 48020 1909
rect 48253 1875 48287 1882
rect 48253 1848 48257 1875
rect 48257 1848 48287 1875
rect 47986 1807 48020 1839
rect 47986 1805 48020 1807
rect 48427 1875 48461 1882
rect 48427 1848 48459 1875
rect 48459 1848 48461 1875
rect 49329 1875 49363 1884
rect 49329 1850 49331 1875
rect 49331 1850 49363 1875
rect 49502 1875 49536 1880
rect 49502 1846 49533 1875
rect 49533 1846 49536 1875
rect 47842 1677 47876 1711
rect 48341 1755 48373 1759
rect 48373 1755 48375 1759
rect 48341 1725 48375 1755
rect 49411 1755 49413 1764
rect 49413 1755 49445 1764
rect 49411 1730 49445 1755
rect 47954 1596 47988 1630
rect 48249 1609 48283 1643
rect 48341 1609 48375 1643
rect 48433 1609 48467 1643
rect 49323 1609 49357 1643
rect 49415 1609 49449 1643
rect 49507 1609 49541 1643
rect 47810 1544 47844 1546
rect 47810 1512 47844 1544
rect 47810 1442 47844 1474
rect 47810 1440 47844 1442
rect 47906 1544 47940 1546
rect 47906 1512 47940 1544
rect 47906 1442 47940 1474
rect 47906 1440 47940 1442
rect 48002 1544 48036 1546
rect 48002 1512 48036 1544
rect 48002 1442 48036 1474
rect 48002 1440 48036 1442
rect 47858 1356 47892 1390
rect 47778 1247 47812 1281
rect 48208 1230 48242 1264
rect 46565 1107 46599 1141
rect 46657 1107 46691 1141
rect 46749 1107 46783 1141
rect 45688 1013 45722 1015
rect 45688 981 45722 1013
rect 45688 911 45722 943
rect 45688 909 45722 911
rect 45776 1013 45810 1015
rect 45776 981 45810 1013
rect 46334 1013 46368 1015
rect 46048 949 46082 983
rect 46334 981 46368 1013
rect 45776 911 45810 943
rect 45776 909 45810 911
rect 46334 911 46368 943
rect 46334 909 46368 911
rect 45904 853 45938 855
rect 45904 821 45938 853
rect 45732 781 45766 815
rect 45029 561 45063 595
rect 45121 561 45155 595
rect 45213 561 45247 595
rect 45904 751 45938 783
rect 45904 749 45938 751
rect 46000 853 46034 855
rect 46000 821 46034 853
rect 46000 751 46034 783
rect 46000 749 46034 751
rect 46911 1105 46945 1139
rect 47003 1105 47037 1139
rect 47095 1105 47129 1139
rect 46422 1013 46456 1015
rect 46422 981 46456 1013
rect 46422 911 46456 943
rect 46422 909 46456 911
rect 47257 1099 47291 1133
rect 47349 1099 47383 1133
rect 47441 1099 47475 1133
rect 47620 1109 47654 1143
rect 46096 853 46130 855
rect 46096 821 46130 853
rect 46096 751 46130 783
rect 46378 781 46412 815
rect 46096 749 46130 751
rect 46917 793 46919 826
rect 46919 793 46951 826
rect 46917 792 46951 793
rect 48266 1109 48300 1143
rect 47110 804 47144 838
rect 45952 621 45986 655
rect 45369 555 45403 589
rect 45461 555 45495 589
rect 45553 555 45587 589
rect 45704 550 45738 584
rect 46336 578 46370 612
rect 46696 711 46730 728
rect 46696 694 46730 711
rect 47306 821 47340 832
rect 47306 798 47308 821
rect 47308 798 47340 821
rect 42342 386 42376 418
rect 42342 384 42376 386
rect 44038 488 44072 490
rect 44038 456 44072 488
rect 44134 488 44168 490
rect 44134 456 44168 488
rect 44038 386 44072 418
rect 44038 384 44072 386
rect 44134 386 44168 418
rect 44134 384 44168 386
rect 44230 488 44264 490
rect 44230 456 44264 488
rect 46064 540 46098 574
rect 46565 563 46599 597
rect 46657 563 46691 597
rect 46749 563 46783 597
rect 47867 1057 47901 1091
rect 49294 1364 49328 1398
rect 49682 1909 49716 1911
rect 49682 1877 49716 1909
rect 49682 1807 49716 1839
rect 49682 1805 49716 1807
rect 49778 1909 49812 1911
rect 49778 1877 49812 1909
rect 49778 1807 49812 1839
rect 49778 1805 49812 1807
rect 51645 2113 51679 2147
rect 51714 2005 51748 2039
rect 49874 1909 49908 1911
rect 49874 1877 49908 1909
rect 50141 1875 50175 1882
rect 50141 1848 50145 1875
rect 50145 1848 50175 1875
rect 49874 1807 49908 1839
rect 49874 1805 49908 1807
rect 50315 1875 50349 1882
rect 50315 1848 50347 1875
rect 50347 1848 50349 1875
rect 51217 1875 51251 1884
rect 51217 1850 51219 1875
rect 51219 1850 51251 1875
rect 51390 1875 51424 1880
rect 51390 1846 51421 1875
rect 51421 1846 51424 1875
rect 49730 1677 49764 1711
rect 50229 1755 50261 1759
rect 50261 1755 50263 1759
rect 50229 1725 50263 1755
rect 51299 1755 51301 1764
rect 51301 1755 51333 1764
rect 51299 1730 51333 1755
rect 49842 1596 49876 1630
rect 50137 1609 50171 1643
rect 50229 1609 50263 1643
rect 50321 1609 50355 1643
rect 51211 1609 51245 1643
rect 51303 1609 51337 1643
rect 51395 1609 51429 1643
rect 49698 1544 49732 1546
rect 49698 1512 49732 1544
rect 49698 1442 49732 1474
rect 49698 1440 49732 1442
rect 49794 1544 49828 1546
rect 49794 1512 49828 1544
rect 49794 1442 49828 1474
rect 49794 1440 49828 1442
rect 49890 1544 49924 1546
rect 49890 1512 49924 1544
rect 49890 1442 49924 1474
rect 49890 1440 49924 1442
rect 49746 1356 49780 1390
rect 49666 1247 49700 1281
rect 50096 1230 50130 1264
rect 48453 1107 48487 1141
rect 48545 1107 48579 1141
rect 48637 1107 48671 1141
rect 47576 1013 47610 1015
rect 47576 981 47610 1013
rect 47576 911 47610 943
rect 47576 909 47610 911
rect 47664 1013 47698 1015
rect 47664 981 47698 1013
rect 48222 1013 48256 1015
rect 47936 949 47970 983
rect 48222 981 48256 1013
rect 47664 911 47698 943
rect 47664 909 47698 911
rect 48222 911 48256 943
rect 48222 909 48256 911
rect 47792 853 47826 855
rect 47792 821 47826 853
rect 47620 781 47654 815
rect 46911 561 46945 595
rect 47003 561 47037 595
rect 47095 561 47129 595
rect 47792 751 47826 783
rect 47792 749 47826 751
rect 47888 853 47922 855
rect 47888 821 47922 853
rect 47888 751 47922 783
rect 47888 749 47922 751
rect 48799 1105 48833 1139
rect 48891 1105 48925 1139
rect 48983 1105 49017 1139
rect 48310 1013 48344 1015
rect 48310 981 48344 1013
rect 48310 911 48344 943
rect 48310 909 48344 911
rect 49145 1099 49179 1133
rect 49237 1099 49271 1133
rect 49329 1099 49363 1133
rect 49508 1109 49542 1143
rect 47984 853 48018 855
rect 47984 821 48018 853
rect 47984 751 48018 783
rect 48266 781 48300 815
rect 47984 749 48018 751
rect 48805 793 48807 826
rect 48807 793 48839 826
rect 48805 792 48839 793
rect 50154 1109 50188 1143
rect 48998 804 49032 838
rect 47840 621 47874 655
rect 47257 555 47291 589
rect 47349 555 47383 589
rect 47441 555 47475 589
rect 47592 550 47626 584
rect 48224 578 48258 612
rect 48584 711 48618 728
rect 48584 694 48618 711
rect 49194 821 49228 832
rect 49194 798 49196 821
rect 49196 798 49228 821
rect 44230 386 44264 418
rect 44230 384 44264 386
rect 45920 488 45954 490
rect 45920 456 45954 488
rect 46016 488 46050 490
rect 46016 456 46050 488
rect 45920 386 45954 418
rect 45920 384 45954 386
rect 46016 386 46050 418
rect 46016 384 46050 386
rect 46112 488 46146 490
rect 46112 456 46146 488
rect 47952 540 47986 574
rect 48453 563 48487 597
rect 48545 563 48579 597
rect 48637 563 48671 597
rect 49755 1057 49789 1091
rect 51182 1364 51216 1398
rect 51570 1909 51604 1911
rect 51570 1877 51604 1909
rect 51570 1807 51604 1839
rect 51570 1805 51604 1807
rect 51666 1909 51700 1911
rect 51666 1877 51700 1909
rect 51666 1807 51700 1839
rect 51666 1805 51700 1807
rect 53533 2113 53567 2147
rect 53602 2005 53636 2039
rect 51762 1909 51796 1911
rect 51762 1877 51796 1909
rect 52029 1875 52063 1882
rect 52029 1848 52033 1875
rect 52033 1848 52063 1875
rect 51762 1807 51796 1839
rect 51762 1805 51796 1807
rect 52203 1875 52237 1882
rect 52203 1848 52235 1875
rect 52235 1848 52237 1875
rect 53105 1875 53139 1884
rect 53105 1850 53107 1875
rect 53107 1850 53139 1875
rect 53278 1875 53312 1880
rect 53278 1846 53309 1875
rect 53309 1846 53312 1875
rect 51618 1677 51652 1711
rect 52117 1755 52149 1759
rect 52149 1755 52151 1759
rect 52117 1725 52151 1755
rect 53187 1755 53189 1764
rect 53189 1755 53221 1764
rect 53187 1730 53221 1755
rect 51730 1596 51764 1630
rect 52025 1609 52059 1643
rect 52117 1609 52151 1643
rect 52209 1609 52243 1643
rect 53099 1609 53133 1643
rect 53191 1609 53225 1643
rect 53283 1609 53317 1643
rect 51586 1544 51620 1546
rect 51586 1512 51620 1544
rect 51586 1442 51620 1474
rect 51586 1440 51620 1442
rect 51682 1544 51716 1546
rect 51682 1512 51716 1544
rect 51682 1442 51716 1474
rect 51682 1440 51716 1442
rect 51778 1544 51812 1546
rect 51778 1512 51812 1544
rect 51778 1442 51812 1474
rect 51778 1440 51812 1442
rect 51634 1356 51668 1390
rect 51554 1247 51588 1281
rect 51984 1230 52018 1264
rect 50341 1107 50375 1141
rect 50433 1107 50467 1141
rect 50525 1107 50559 1141
rect 49464 1013 49498 1015
rect 49464 981 49498 1013
rect 49464 911 49498 943
rect 49464 909 49498 911
rect 49552 1013 49586 1015
rect 49552 981 49586 1013
rect 50110 1013 50144 1015
rect 49824 949 49858 983
rect 50110 981 50144 1013
rect 49552 911 49586 943
rect 49552 909 49586 911
rect 50110 911 50144 943
rect 50110 909 50144 911
rect 49680 853 49714 855
rect 49680 821 49714 853
rect 49508 781 49542 815
rect 48799 561 48833 595
rect 48891 561 48925 595
rect 48983 561 49017 595
rect 49680 751 49714 783
rect 49680 749 49714 751
rect 49776 853 49810 855
rect 49776 821 49810 853
rect 49776 751 49810 783
rect 49776 749 49810 751
rect 50687 1105 50721 1139
rect 50779 1105 50813 1139
rect 50871 1105 50905 1139
rect 50198 1013 50232 1015
rect 50198 981 50232 1013
rect 50198 911 50232 943
rect 50198 909 50232 911
rect 51033 1099 51067 1133
rect 51125 1099 51159 1133
rect 51217 1099 51251 1133
rect 51396 1109 51430 1143
rect 49872 853 49906 855
rect 49872 821 49906 853
rect 49872 751 49906 783
rect 50154 781 50188 815
rect 49872 749 49906 751
rect 50693 793 50695 826
rect 50695 793 50727 826
rect 50693 792 50727 793
rect 52042 1109 52076 1143
rect 50886 804 50920 838
rect 49728 621 49762 655
rect 49145 555 49179 589
rect 49237 555 49271 589
rect 49329 555 49363 589
rect 49480 550 49514 584
rect 50112 578 50146 612
rect 50472 711 50506 728
rect 50472 694 50506 711
rect 51082 821 51116 832
rect 51082 798 51084 821
rect 51084 798 51116 821
rect 46112 386 46146 418
rect 46112 384 46146 386
rect 47808 488 47842 490
rect 47808 456 47842 488
rect 47904 488 47938 490
rect 47904 456 47938 488
rect 47808 386 47842 418
rect 47808 384 47842 386
rect 47904 386 47938 418
rect 47904 384 47938 386
rect 48000 488 48034 490
rect 48000 456 48034 488
rect 49840 540 49874 574
rect 50341 563 50375 597
rect 50433 563 50467 597
rect 50525 563 50559 597
rect 51643 1057 51677 1091
rect 53070 1364 53104 1398
rect 53458 1909 53492 1911
rect 53458 1877 53492 1909
rect 53458 1807 53492 1839
rect 53458 1805 53492 1807
rect 53554 1909 53588 1911
rect 53554 1877 53588 1909
rect 53554 1807 53588 1839
rect 53554 1805 53588 1807
rect 55421 2113 55455 2147
rect 55490 2005 55524 2039
rect 53650 1909 53684 1911
rect 53650 1877 53684 1909
rect 53917 1875 53951 1882
rect 53917 1848 53921 1875
rect 53921 1848 53951 1875
rect 53650 1807 53684 1839
rect 53650 1805 53684 1807
rect 54091 1875 54125 1882
rect 54091 1848 54123 1875
rect 54123 1848 54125 1875
rect 54993 1875 55027 1884
rect 54993 1850 54995 1875
rect 54995 1850 55027 1875
rect 55166 1875 55200 1880
rect 55166 1846 55197 1875
rect 55197 1846 55200 1875
rect 53506 1677 53540 1711
rect 54005 1755 54037 1759
rect 54037 1755 54039 1759
rect 54005 1725 54039 1755
rect 55075 1755 55077 1764
rect 55077 1755 55109 1764
rect 55075 1730 55109 1755
rect 53618 1596 53652 1630
rect 53913 1609 53947 1643
rect 54005 1609 54039 1643
rect 54097 1609 54131 1643
rect 54987 1609 55021 1643
rect 55079 1609 55113 1643
rect 55171 1609 55205 1643
rect 53474 1544 53508 1546
rect 53474 1512 53508 1544
rect 53474 1442 53508 1474
rect 53474 1440 53508 1442
rect 53570 1544 53604 1546
rect 53570 1512 53604 1544
rect 53570 1442 53604 1474
rect 53570 1440 53604 1442
rect 53666 1544 53700 1546
rect 53666 1512 53700 1544
rect 53666 1442 53700 1474
rect 53666 1440 53700 1442
rect 53522 1356 53556 1390
rect 53442 1247 53476 1281
rect 53872 1230 53906 1264
rect 52229 1107 52263 1141
rect 52321 1107 52355 1141
rect 52413 1107 52447 1141
rect 51352 1013 51386 1015
rect 51352 981 51386 1013
rect 51352 911 51386 943
rect 51352 909 51386 911
rect 51440 1013 51474 1015
rect 51440 981 51474 1013
rect 51998 1013 52032 1015
rect 51712 949 51746 983
rect 51998 981 52032 1013
rect 51440 911 51474 943
rect 51440 909 51474 911
rect 51998 911 52032 943
rect 51998 909 52032 911
rect 51568 853 51602 855
rect 51568 821 51602 853
rect 51396 781 51430 815
rect 50687 561 50721 595
rect 50779 561 50813 595
rect 50871 561 50905 595
rect 51568 751 51602 783
rect 51568 749 51602 751
rect 51664 853 51698 855
rect 51664 821 51698 853
rect 51664 751 51698 783
rect 51664 749 51698 751
rect 52575 1105 52609 1139
rect 52667 1105 52701 1139
rect 52759 1105 52793 1139
rect 52086 1013 52120 1015
rect 52086 981 52120 1013
rect 52086 911 52120 943
rect 52086 909 52120 911
rect 52921 1099 52955 1133
rect 53013 1099 53047 1133
rect 53105 1099 53139 1133
rect 53284 1109 53318 1143
rect 51760 853 51794 855
rect 51760 821 51794 853
rect 51760 751 51794 783
rect 52042 781 52076 815
rect 51760 749 51794 751
rect 52581 793 52583 826
rect 52583 793 52615 826
rect 52581 792 52615 793
rect 53930 1109 53964 1143
rect 52774 804 52808 838
rect 51616 621 51650 655
rect 51033 555 51067 589
rect 51125 555 51159 589
rect 51217 555 51251 589
rect 51368 550 51402 584
rect 52000 578 52034 612
rect 52360 711 52394 728
rect 52360 694 52394 711
rect 52970 821 53004 832
rect 52970 798 52972 821
rect 52972 798 53004 821
rect 48000 386 48034 418
rect 48000 384 48034 386
rect 49696 488 49730 490
rect 49696 456 49730 488
rect 49792 488 49826 490
rect 49792 456 49826 488
rect 49696 386 49730 418
rect 49696 384 49730 386
rect 49792 386 49826 418
rect 49792 384 49826 386
rect 49888 488 49922 490
rect 49888 456 49922 488
rect 51728 540 51762 574
rect 52229 563 52263 597
rect 52321 563 52355 597
rect 52413 563 52447 597
rect 53531 1057 53565 1091
rect 54958 1364 54992 1398
rect 55346 1909 55380 1911
rect 55346 1877 55380 1909
rect 55346 1807 55380 1839
rect 55346 1805 55380 1807
rect 55442 1909 55476 1911
rect 55442 1877 55476 1909
rect 55442 1807 55476 1839
rect 55442 1805 55476 1807
rect 57309 2113 57343 2147
rect 57378 2005 57412 2039
rect 55538 1909 55572 1911
rect 55538 1877 55572 1909
rect 55805 1875 55839 1882
rect 55805 1848 55809 1875
rect 55809 1848 55839 1875
rect 55538 1807 55572 1839
rect 55538 1805 55572 1807
rect 55979 1875 56013 1882
rect 55979 1848 56011 1875
rect 56011 1848 56013 1875
rect 56881 1875 56915 1884
rect 56881 1850 56883 1875
rect 56883 1850 56915 1875
rect 57054 1875 57088 1880
rect 57054 1846 57085 1875
rect 57085 1846 57088 1875
rect 55394 1677 55428 1711
rect 55893 1755 55925 1759
rect 55925 1755 55927 1759
rect 55893 1725 55927 1755
rect 56963 1755 56965 1764
rect 56965 1755 56997 1764
rect 56963 1730 56997 1755
rect 55506 1596 55540 1630
rect 55801 1609 55835 1643
rect 55893 1609 55927 1643
rect 55985 1609 56019 1643
rect 56875 1609 56909 1643
rect 56967 1609 57001 1643
rect 57059 1609 57093 1643
rect 55362 1544 55396 1546
rect 55362 1512 55396 1544
rect 55362 1442 55396 1474
rect 55362 1440 55396 1442
rect 55458 1544 55492 1546
rect 55458 1512 55492 1544
rect 55458 1442 55492 1474
rect 55458 1440 55492 1442
rect 55554 1544 55588 1546
rect 55554 1512 55588 1544
rect 55554 1442 55588 1474
rect 55554 1440 55588 1442
rect 55410 1356 55444 1390
rect 55330 1247 55364 1281
rect 55760 1230 55794 1264
rect 54117 1107 54151 1141
rect 54209 1107 54243 1141
rect 54301 1107 54335 1141
rect 53240 1013 53274 1015
rect 53240 981 53274 1013
rect 53240 911 53274 943
rect 53240 909 53274 911
rect 53328 1013 53362 1015
rect 53328 981 53362 1013
rect 53886 1013 53920 1015
rect 53600 949 53634 983
rect 53886 981 53920 1013
rect 53328 911 53362 943
rect 53328 909 53362 911
rect 53886 911 53920 943
rect 53886 909 53920 911
rect 53456 853 53490 855
rect 53456 821 53490 853
rect 53284 781 53318 815
rect 52575 561 52609 595
rect 52667 561 52701 595
rect 52759 561 52793 595
rect 53456 751 53490 783
rect 53456 749 53490 751
rect 53552 853 53586 855
rect 53552 821 53586 853
rect 53552 751 53586 783
rect 53552 749 53586 751
rect 54463 1105 54497 1139
rect 54555 1105 54589 1139
rect 54647 1105 54681 1139
rect 53974 1013 54008 1015
rect 53974 981 54008 1013
rect 53974 911 54008 943
rect 53974 909 54008 911
rect 54809 1099 54843 1133
rect 54901 1099 54935 1133
rect 54993 1099 55027 1133
rect 55172 1109 55206 1143
rect 53648 853 53682 855
rect 53648 821 53682 853
rect 53648 751 53682 783
rect 53930 781 53964 815
rect 53648 749 53682 751
rect 54469 793 54471 826
rect 54471 793 54503 826
rect 54469 792 54503 793
rect 55818 1109 55852 1143
rect 54662 804 54696 838
rect 53504 621 53538 655
rect 52921 555 52955 589
rect 53013 555 53047 589
rect 53105 555 53139 589
rect 53256 550 53290 584
rect 53888 578 53922 612
rect 54248 711 54282 728
rect 54248 694 54282 711
rect 54858 821 54892 832
rect 54858 798 54860 821
rect 54860 798 54892 821
rect 49888 386 49922 418
rect 49888 384 49922 386
rect 51584 488 51618 490
rect 51584 456 51618 488
rect 51680 488 51714 490
rect 51680 456 51714 488
rect 51584 386 51618 418
rect 51584 384 51618 386
rect 51680 386 51714 418
rect 51680 384 51714 386
rect 51776 488 51810 490
rect 51776 456 51810 488
rect 53616 540 53650 574
rect 54117 563 54151 597
rect 54209 563 54243 597
rect 54301 563 54335 597
rect 55419 1057 55453 1091
rect 56846 1364 56880 1398
rect 57234 1909 57268 1911
rect 57234 1877 57268 1909
rect 57234 1807 57268 1839
rect 57234 1805 57268 1807
rect 57330 1909 57364 1911
rect 57330 1877 57364 1909
rect 57330 1807 57364 1839
rect 57330 1805 57364 1807
rect 59197 2113 59231 2147
rect 59266 2005 59300 2039
rect 57426 1909 57460 1911
rect 57426 1877 57460 1909
rect 57693 1875 57727 1882
rect 57693 1848 57697 1875
rect 57697 1848 57727 1875
rect 57426 1807 57460 1839
rect 57426 1805 57460 1807
rect 57867 1875 57901 1882
rect 57867 1848 57899 1875
rect 57899 1848 57901 1875
rect 58769 1875 58803 1884
rect 58769 1850 58771 1875
rect 58771 1850 58803 1875
rect 58942 1875 58976 1880
rect 58942 1846 58973 1875
rect 58973 1846 58976 1875
rect 57282 1677 57316 1711
rect 57781 1755 57813 1759
rect 57813 1755 57815 1759
rect 57781 1725 57815 1755
rect 58851 1755 58853 1764
rect 58853 1755 58885 1764
rect 58851 1730 58885 1755
rect 57394 1596 57428 1630
rect 57689 1609 57723 1643
rect 57781 1609 57815 1643
rect 57873 1609 57907 1643
rect 58763 1609 58797 1643
rect 58855 1609 58889 1643
rect 58947 1609 58981 1643
rect 57250 1544 57284 1546
rect 57250 1512 57284 1544
rect 57250 1442 57284 1474
rect 57250 1440 57284 1442
rect 57346 1544 57380 1546
rect 57346 1512 57380 1544
rect 57346 1442 57380 1474
rect 57346 1440 57380 1442
rect 57442 1544 57476 1546
rect 57442 1512 57476 1544
rect 57442 1442 57476 1474
rect 57442 1440 57476 1442
rect 57298 1356 57332 1390
rect 57218 1247 57252 1281
rect 57648 1230 57682 1264
rect 56005 1107 56039 1141
rect 56097 1107 56131 1141
rect 56189 1107 56223 1141
rect 55128 1013 55162 1015
rect 55128 981 55162 1013
rect 55128 911 55162 943
rect 55128 909 55162 911
rect 55216 1013 55250 1015
rect 55216 981 55250 1013
rect 55774 1013 55808 1015
rect 55488 949 55522 983
rect 55774 981 55808 1013
rect 55216 911 55250 943
rect 55216 909 55250 911
rect 55774 911 55808 943
rect 55774 909 55808 911
rect 55344 853 55378 855
rect 55344 821 55378 853
rect 55172 781 55206 815
rect 54463 561 54497 595
rect 54555 561 54589 595
rect 54647 561 54681 595
rect 55344 751 55378 783
rect 55344 749 55378 751
rect 55440 853 55474 855
rect 55440 821 55474 853
rect 55440 751 55474 783
rect 55440 749 55474 751
rect 56351 1105 56385 1139
rect 56443 1105 56477 1139
rect 56535 1105 56569 1139
rect 55862 1013 55896 1015
rect 55862 981 55896 1013
rect 55862 911 55896 943
rect 55862 909 55896 911
rect 56697 1099 56731 1133
rect 56789 1099 56823 1133
rect 56881 1099 56915 1133
rect 57060 1109 57094 1143
rect 55536 853 55570 855
rect 55536 821 55570 853
rect 55536 751 55570 783
rect 55818 781 55852 815
rect 55536 749 55570 751
rect 56357 793 56359 826
rect 56359 793 56391 826
rect 56357 792 56391 793
rect 57706 1109 57740 1143
rect 56550 804 56584 838
rect 55392 621 55426 655
rect 54809 555 54843 589
rect 54901 555 54935 589
rect 54993 555 55027 589
rect 55144 550 55178 584
rect 55776 578 55810 612
rect 56136 711 56170 728
rect 56136 694 56170 711
rect 56746 821 56780 832
rect 56746 798 56748 821
rect 56748 798 56780 821
rect 51776 386 51810 418
rect 51776 384 51810 386
rect 53472 488 53506 490
rect 53472 456 53506 488
rect 53568 488 53602 490
rect 53568 456 53602 488
rect 53472 386 53506 418
rect 53472 384 53506 386
rect 53568 386 53602 418
rect 53568 384 53602 386
rect 53664 488 53698 490
rect 53664 456 53698 488
rect 55504 540 55538 574
rect 56005 563 56039 597
rect 56097 563 56131 597
rect 56189 563 56223 597
rect 57307 1057 57341 1091
rect 58734 1364 58768 1398
rect 59122 1909 59156 1911
rect 59122 1877 59156 1909
rect 59122 1807 59156 1839
rect 59122 1805 59156 1807
rect 59218 1909 59252 1911
rect 59218 1877 59252 1909
rect 59218 1807 59252 1839
rect 59218 1805 59252 1807
rect 59314 1909 59348 1911
rect 59314 1877 59348 1909
rect 59581 1875 59615 1882
rect 59581 1848 59585 1875
rect 59585 1848 59615 1875
rect 59314 1807 59348 1839
rect 59314 1805 59348 1807
rect 59755 1875 59789 1882
rect 59755 1848 59787 1875
rect 59787 1848 59789 1875
rect 59170 1677 59204 1711
rect 59669 1755 59701 1759
rect 59701 1755 59703 1759
rect 59669 1725 59703 1755
rect 59282 1596 59316 1630
rect 59577 1609 59611 1643
rect 59669 1609 59703 1643
rect 59761 1609 59795 1643
rect 59138 1544 59172 1546
rect 59138 1512 59172 1544
rect 59138 1442 59172 1474
rect 59138 1440 59172 1442
rect 59234 1544 59268 1546
rect 59234 1512 59268 1544
rect 59234 1442 59268 1474
rect 59234 1440 59268 1442
rect 59330 1544 59364 1546
rect 59330 1512 59364 1544
rect 59330 1442 59364 1474
rect 59330 1440 59364 1442
rect 59186 1356 59220 1390
rect 59106 1247 59140 1281
rect 59536 1230 59570 1264
rect 57893 1107 57927 1141
rect 57985 1107 58019 1141
rect 58077 1107 58111 1141
rect 57016 1013 57050 1015
rect 57016 981 57050 1013
rect 57016 911 57050 943
rect 57016 909 57050 911
rect 57104 1013 57138 1015
rect 57104 981 57138 1013
rect 57662 1013 57696 1015
rect 57376 949 57410 983
rect 57662 981 57696 1013
rect 57104 911 57138 943
rect 57104 909 57138 911
rect 57662 911 57696 943
rect 57662 909 57696 911
rect 57232 853 57266 855
rect 57232 821 57266 853
rect 57060 781 57094 815
rect 56351 561 56385 595
rect 56443 561 56477 595
rect 56535 561 56569 595
rect 57232 751 57266 783
rect 57232 749 57266 751
rect 57328 853 57362 855
rect 57328 821 57362 853
rect 57328 751 57362 783
rect 57328 749 57362 751
rect 58239 1105 58273 1139
rect 58331 1105 58365 1139
rect 58423 1105 58457 1139
rect 57750 1013 57784 1015
rect 57750 981 57784 1013
rect 57750 911 57784 943
rect 57750 909 57784 911
rect 58585 1099 58619 1133
rect 58677 1099 58711 1133
rect 58769 1099 58803 1133
rect 58948 1109 58982 1143
rect 57424 853 57458 855
rect 57424 821 57458 853
rect 57424 751 57458 783
rect 57706 781 57740 815
rect 57424 749 57458 751
rect 58245 793 58247 826
rect 58247 793 58279 826
rect 58245 792 58279 793
rect 59594 1109 59628 1143
rect 58438 804 58472 838
rect 57280 621 57314 655
rect 56697 555 56731 589
rect 56789 555 56823 589
rect 56881 555 56915 589
rect 57032 550 57066 584
rect 57664 578 57698 612
rect 58024 711 58058 728
rect 58024 694 58058 711
rect 58634 821 58668 832
rect 58634 798 58636 821
rect 58636 798 58668 821
rect 53664 386 53698 418
rect 53664 384 53698 386
rect 55360 488 55394 490
rect 55360 456 55394 488
rect 55456 488 55490 490
rect 55456 456 55490 488
rect 55360 386 55394 418
rect 55360 384 55394 386
rect 55456 386 55490 418
rect 55456 384 55490 386
rect 55552 488 55586 490
rect 55552 456 55586 488
rect 57392 540 57426 574
rect 57893 563 57927 597
rect 57985 563 58019 597
rect 58077 563 58111 597
rect 59195 1057 59229 1091
rect 59781 1107 59815 1141
rect 59873 1107 59907 1141
rect 59965 1107 59999 1141
rect 58904 1013 58938 1015
rect 58904 981 58938 1013
rect 58904 911 58938 943
rect 58904 909 58938 911
rect 58992 1013 59026 1015
rect 58992 981 59026 1013
rect 59550 1013 59584 1015
rect 59264 949 59298 983
rect 59550 981 59584 1013
rect 58992 911 59026 943
rect 58992 909 59026 911
rect 59550 911 59584 943
rect 59550 909 59584 911
rect 59120 853 59154 855
rect 59120 821 59154 853
rect 58948 781 58982 815
rect 58239 561 58273 595
rect 58331 561 58365 595
rect 58423 561 58457 595
rect 59120 751 59154 783
rect 59120 749 59154 751
rect 59216 853 59250 855
rect 59216 821 59250 853
rect 59216 751 59250 783
rect 59216 749 59250 751
rect 60127 1105 60161 1139
rect 60219 1105 60253 1139
rect 60311 1105 60345 1139
rect 59638 1013 59672 1015
rect 59638 981 59672 1013
rect 59638 911 59672 943
rect 59638 909 59672 911
rect 59312 853 59346 855
rect 59312 821 59346 853
rect 59312 751 59346 783
rect 59594 781 59628 815
rect 59312 749 59346 751
rect 60133 793 60135 826
rect 60135 793 60167 826
rect 60133 792 60167 793
rect 60326 804 60360 838
rect 59168 621 59202 655
rect 58585 555 58619 589
rect 58677 555 58711 589
rect 58769 555 58803 589
rect 58920 550 58954 584
rect 59552 578 59586 612
rect 59912 711 59946 728
rect 59912 694 59946 711
rect 55552 386 55586 418
rect 55552 384 55586 386
rect 57248 488 57282 490
rect 57248 456 57282 488
rect 57344 488 57378 490
rect 57344 456 57378 488
rect 57248 386 57282 418
rect 57248 384 57282 386
rect 57344 386 57378 418
rect 57344 384 57378 386
rect 57440 488 57474 490
rect 57440 456 57474 488
rect 59280 540 59314 574
rect 59781 563 59815 597
rect 59873 563 59907 597
rect 59965 563 59999 597
rect 60127 561 60161 595
rect 60219 561 60253 595
rect 60311 561 60345 595
rect 57440 386 57474 418
rect 57440 384 57474 386
rect 59136 488 59170 490
rect 59136 456 59170 488
rect 59232 488 59266 490
rect 59232 456 59266 488
rect 59136 386 59170 418
rect 59136 384 59170 386
rect 59232 386 59266 418
rect 59232 384 59266 386
rect 59328 488 59362 490
rect 59328 456 59362 488
rect 59328 386 59362 418
rect 59328 384 59362 386
rect 668 300 702 334
rect 2556 300 2590 334
rect 4444 300 4478 334
rect 6332 300 6366 334
rect 8220 300 8254 334
rect 10108 300 10142 334
rect 11996 300 12030 334
rect 13884 300 13918 334
rect 15766 300 15800 334
rect 17654 300 17688 334
rect 19542 300 19576 334
rect 21430 300 21464 334
rect 23318 300 23352 334
rect 25206 300 25240 334
rect 27094 300 27128 334
rect 28982 300 29016 334
rect 30870 300 30904 334
rect 32758 300 32792 334
rect 34646 300 34680 334
rect 36534 300 36568 334
rect 38422 300 38456 334
rect 40310 300 40344 334
rect 42198 300 42232 334
rect 44086 300 44120 334
rect 45968 300 46002 334
rect 47856 300 47890 334
rect 49744 300 49778 334
rect 51632 300 51666 334
rect 53520 300 53554 334
rect 55408 300 55442 334
rect 57296 300 57330 334
rect 59184 300 59218 334
rect 588 191 622 225
rect 2476 191 2510 225
rect 4364 191 4398 225
rect 6252 191 6286 225
rect 8140 191 8174 225
rect 10028 191 10062 225
rect 11916 191 11950 225
rect 13804 191 13838 225
rect 15686 191 15720 225
rect 17574 191 17608 225
rect 19462 191 19496 225
rect 21350 191 21384 225
rect 23238 191 23272 225
rect 25126 191 25160 225
rect 27014 191 27048 225
rect 28902 191 28936 225
rect 30790 191 30824 225
rect 32678 191 32712 225
rect 34566 191 34600 225
rect 36454 191 36488 225
rect 38342 191 38376 225
rect 40230 191 40264 225
rect 42118 191 42152 225
rect 44006 191 44040 225
rect 45888 191 45922 225
rect 47776 191 47810 225
rect 49664 191 49698 225
rect 51552 191 51586 225
rect 53440 191 53474 225
rect 55328 191 55362 225
rect 57216 191 57250 225
rect 59104 191 59138 225
<< metal1 >>
rect -430 7376 59974 7440
rect -430 7260 -377 7376
rect -69 7260 1511 7376
rect 1819 7260 3399 7376
rect 3707 7260 5287 7376
rect 5595 7260 7175 7376
rect 7483 7260 9063 7376
rect 9371 7260 10951 7376
rect 11259 7260 12839 7376
rect 13147 7260 14721 7376
rect 15029 7260 16609 7376
rect 16917 7260 18497 7376
rect 18805 7260 20385 7376
rect 20693 7260 22273 7376
rect 22581 7260 24161 7376
rect 24469 7260 26049 7376
rect 26357 7260 27937 7376
rect 28245 7260 29825 7376
rect 30133 7260 31713 7376
rect 32021 7260 33601 7376
rect 33909 7260 35489 7376
rect 35797 7260 37377 7376
rect 37685 7260 39265 7376
rect 39573 7260 41153 7376
rect 41461 7260 43041 7376
rect 43349 7260 44923 7376
rect 45231 7260 46811 7376
rect 47119 7260 48699 7376
rect 49007 7260 50587 7376
rect 50895 7260 52475 7376
rect 52783 7260 54363 7376
rect 54671 7260 56251 7376
rect 56559 7260 58139 7376
rect 58447 7260 59974 7376
rect -430 7249 59974 7260
rect -430 7215 844 7249
rect 878 7215 2732 7249
rect 2766 7215 4620 7249
rect 4654 7215 6508 7249
rect 6542 7215 8396 7249
rect 8430 7215 10284 7249
rect 10318 7215 12172 7249
rect 12206 7215 14060 7249
rect 14094 7215 15942 7249
rect 15976 7215 17830 7249
rect 17864 7215 19718 7249
rect 19752 7215 21606 7249
rect 21640 7215 23494 7249
rect 23528 7215 25382 7249
rect 25416 7215 27270 7249
rect 27304 7215 29158 7249
rect 29192 7215 31046 7249
rect 31080 7215 32934 7249
rect 32968 7215 34822 7249
rect 34856 7215 36710 7249
rect 36744 7215 38598 7249
rect 38632 7215 40486 7249
rect 40520 7215 42374 7249
rect 42408 7215 44262 7249
rect 44296 7215 46144 7249
rect 46178 7215 48032 7249
rect 48066 7215 49920 7249
rect 49954 7215 51808 7249
rect 51842 7215 53696 7249
rect 53730 7215 55584 7249
rect 55618 7215 57472 7249
rect 57506 7215 59360 7249
rect 59394 7215 59974 7249
rect -430 7186 59974 7215
rect 132 6910 230 7186
rect -392 6879 230 6910
rect -392 6845 -363 6879
rect -329 6845 -271 6879
rect -237 6845 -179 6879
rect -145 6877 230 6879
rect -145 6845 -17 6877
rect -392 6843 -17 6845
rect 17 6843 75 6877
rect 109 6843 167 6877
rect 201 6843 230 6877
rect 492 7140 812 7158
rect 492 7106 764 7140
rect 798 7106 812 7140
rect 492 7096 812 7106
rect -392 6812 230 6843
rect 370 6868 446 6874
rect 370 6816 386 6868
rect 438 6816 446 6868
rect 370 6810 446 6816
rect 492 6766 552 7096
rect 614 7056 660 7068
rect 24 6746 552 6766
rect 24 6712 36 6746
rect 70 6732 552 6746
rect 70 6712 82 6732
rect 24 6698 82 6712
rect -406 6636 -332 6660
rect -406 6602 -378 6636
rect -344 6602 -332 6636
rect -406 6582 -332 6602
rect -208 6652 -136 6664
rect -208 6600 -197 6652
rect -145 6600 -136 6652
rect 338 6659 404 6668
rect 338 6625 354 6659
rect 388 6625 404 6659
rect 338 6612 404 6625
rect -208 6596 -136 6600
rect 304 6531 350 6578
rect 304 6497 310 6531
rect 344 6497 350 6531
rect 304 6459 350 6497
rect 304 6425 310 6459
rect 344 6425 350 6459
rect 392 6531 438 6578
rect 392 6497 398 6531
rect 432 6497 438 6531
rect 392 6459 438 6497
rect 492 6500 552 6732
rect 580 7022 620 7056
rect 654 7022 660 7056
rect 580 6984 660 7022
rect 700 7062 766 7068
rect 700 7010 706 7062
rect 758 7010 766 7062
rect 700 7004 766 7010
rect 806 7056 908 7068
rect 806 7022 812 7056
rect 846 7022 908 7056
rect 580 6950 620 6984
rect 654 6950 660 6984
rect 580 6938 660 6950
rect 710 6984 756 7004
rect 710 6950 716 6984
rect 750 6950 756 6984
rect 710 6938 756 6950
rect 806 6984 908 7022
rect 806 6950 812 6984
rect 846 6950 908 6984
rect 806 6938 908 6950
rect 580 6738 626 6938
rect 656 6900 714 6910
rect 656 6866 668 6900
rect 702 6866 714 6900
rect 656 6848 714 6866
rect 858 6858 908 6938
rect 1274 6916 1358 7186
rect 1016 6906 1074 6912
rect 1008 6900 1082 6906
rect 768 6819 826 6836
rect 768 6785 780 6819
rect 814 6785 826 6819
rect 768 6770 826 6785
rect 858 6792 928 6858
rect 1008 6848 1019 6900
rect 1071 6848 1082 6900
rect 1008 6842 1082 6848
rect 1150 6890 1426 6916
rect 2020 6910 2118 7186
rect 1150 6885 1251 6890
rect 1303 6885 1426 6890
rect 1150 6851 1179 6885
rect 1213 6851 1251 6885
rect 1305 6851 1363 6885
rect 1397 6851 1426 6885
rect 1016 6834 1074 6842
rect 1150 6838 1251 6851
rect 1303 6838 1426 6851
rect 1150 6820 1426 6838
rect 1496 6879 2118 6910
rect 1496 6845 1525 6879
rect 1559 6845 1617 6879
rect 1651 6845 1709 6879
rect 1743 6877 2118 6879
rect 1743 6845 1871 6877
rect 1496 6843 1871 6845
rect 1905 6843 1963 6877
rect 1997 6843 2055 6877
rect 2089 6843 2118 6877
rect 2380 7140 2700 7158
rect 2380 7106 2652 7140
rect 2686 7106 2700 7140
rect 2380 7096 2700 7106
rect 1496 6812 2118 6843
rect 2258 6868 2334 6874
rect 2258 6816 2274 6868
rect 2326 6816 2334 6868
rect 2258 6810 2334 6816
rect 858 6738 908 6792
rect 2380 6766 2440 7096
rect 2502 7056 2548 7068
rect 580 6691 676 6738
rect 580 6657 636 6691
rect 670 6657 676 6691
rect 580 6619 676 6657
rect 580 6585 636 6619
rect 670 6585 676 6619
rect 726 6691 772 6738
rect 726 6657 732 6691
rect 766 6657 772 6691
rect 726 6619 772 6657
rect 726 6598 732 6619
rect 580 6538 676 6585
rect 716 6590 732 6598
rect 766 6598 772 6619
rect 822 6691 908 6738
rect 1912 6746 2440 6766
rect 1912 6712 1924 6746
rect 1958 6732 2440 6746
rect 1958 6712 1970 6732
rect 1912 6698 1970 6712
rect 822 6657 828 6691
rect 862 6657 908 6691
rect 822 6619 908 6657
rect 766 6590 782 6598
rect 716 6538 724 6590
rect 776 6538 782 6590
rect 822 6585 828 6619
rect 862 6585 908 6619
rect 984 6659 1050 6672
rect 984 6625 1000 6659
rect 1034 6625 1050 6659
rect 1378 6652 1446 6654
rect 984 6614 1050 6625
rect 1294 6648 1446 6652
rect 1294 6642 1387 6648
rect 1294 6608 1314 6642
rect 1348 6608 1387 6642
rect 1294 6602 1387 6608
rect 1378 6596 1387 6602
rect 1439 6596 1446 6648
rect 1378 6590 1446 6596
rect 1482 6636 1556 6660
rect 1482 6602 1510 6636
rect 1544 6602 1556 6636
rect 822 6542 908 6585
rect 1482 6582 1556 6602
rect 1680 6652 1752 6664
rect 1680 6600 1691 6652
rect 1743 6600 1752 6652
rect 2226 6659 2292 6668
rect 2226 6625 2242 6659
rect 2276 6625 2292 6659
rect 2226 6612 2292 6625
rect 1680 6596 1752 6600
rect 822 6538 868 6542
rect 716 6530 782 6538
rect 950 6531 996 6578
rect 492 6491 730 6500
rect 492 6468 684 6491
rect 392 6442 398 6459
rect 304 6378 350 6425
rect 380 6436 398 6442
rect 432 6442 438 6459
rect 490 6457 684 6468
rect 718 6457 730 6491
rect 950 6497 956 6531
rect 990 6497 996 6531
rect 950 6464 996 6497
rect 432 6436 446 6442
rect 380 6384 386 6436
rect 438 6384 446 6436
rect 380 6378 446 6384
rect 490 6440 730 6457
rect -394 6348 230 6366
rect -394 6335 148 6348
rect -394 6301 -363 6335
rect -329 6301 -271 6335
rect -237 6301 -179 6335
rect -145 6333 148 6335
rect 200 6333 230 6348
rect -145 6301 -17 6333
rect -394 6299 -17 6301
rect 17 6299 75 6333
rect 109 6299 148 6333
rect 201 6299 230 6333
rect -394 6296 148 6299
rect 200 6296 230 6299
rect -394 6264 230 6296
rect 338 6331 404 6342
rect 338 6297 354 6331
rect 388 6297 404 6331
rect 338 6286 404 6297
rect 490 6294 524 6440
rect 672 6438 730 6440
rect 928 6459 996 6464
rect 928 6456 956 6459
rect 928 6404 936 6456
rect 990 6425 996 6459
rect 988 6404 996 6425
rect 726 6383 816 6404
rect 928 6398 996 6404
rect 726 6349 753 6383
rect 787 6349 816 6383
rect 950 6378 996 6398
rect 1038 6531 1084 6578
rect 1038 6497 1044 6531
rect 1078 6497 1084 6531
rect 1038 6459 1084 6497
rect 1038 6425 1044 6459
rect 1078 6425 1084 6459
rect 1038 6404 1084 6425
rect 2192 6531 2238 6578
rect 2192 6497 2198 6531
rect 2232 6497 2238 6531
rect 2192 6459 2238 6497
rect 2192 6425 2198 6459
rect 2232 6425 2238 6459
rect 2280 6531 2326 6578
rect 2280 6497 2286 6531
rect 2320 6497 2326 6531
rect 2280 6459 2326 6497
rect 2380 6500 2440 6732
rect 2468 7022 2508 7056
rect 2542 7022 2548 7056
rect 2468 6984 2548 7022
rect 2588 7062 2654 7068
rect 2588 7010 2594 7062
rect 2646 7010 2654 7062
rect 2588 7004 2654 7010
rect 2694 7056 2796 7068
rect 2694 7022 2700 7056
rect 2734 7022 2796 7056
rect 2468 6950 2508 6984
rect 2542 6950 2548 6984
rect 2468 6938 2548 6950
rect 2598 6984 2644 7004
rect 2598 6950 2604 6984
rect 2638 6950 2644 6984
rect 2598 6938 2644 6950
rect 2694 6984 2796 7022
rect 2694 6950 2700 6984
rect 2734 6950 2796 6984
rect 2694 6938 2796 6950
rect 2468 6738 2514 6938
rect 2544 6900 2602 6910
rect 2544 6866 2556 6900
rect 2590 6866 2602 6900
rect 2544 6848 2602 6866
rect 2746 6858 2796 6938
rect 3162 6916 3246 7186
rect 2904 6906 2962 6912
rect 2896 6900 2970 6906
rect 2656 6819 2714 6836
rect 2656 6785 2668 6819
rect 2702 6785 2714 6819
rect 2656 6770 2714 6785
rect 2746 6792 2816 6858
rect 2896 6848 2907 6900
rect 2959 6848 2970 6900
rect 2896 6842 2970 6848
rect 3038 6890 3314 6916
rect 3908 6910 4006 7186
rect 3038 6885 3139 6890
rect 3191 6885 3314 6890
rect 3038 6851 3067 6885
rect 3101 6851 3139 6885
rect 3193 6851 3251 6885
rect 3285 6851 3314 6885
rect 2904 6834 2962 6842
rect 3038 6838 3139 6851
rect 3191 6838 3314 6851
rect 3038 6820 3314 6838
rect 3384 6879 4006 6910
rect 3384 6845 3413 6879
rect 3447 6845 3505 6879
rect 3539 6845 3597 6879
rect 3631 6877 4006 6879
rect 3631 6845 3759 6877
rect 3384 6843 3759 6845
rect 3793 6843 3851 6877
rect 3885 6843 3943 6877
rect 3977 6843 4006 6877
rect 4268 7140 4588 7158
rect 4268 7106 4540 7140
rect 4574 7106 4588 7140
rect 4268 7096 4588 7106
rect 3384 6812 4006 6843
rect 4146 6868 4222 6874
rect 4146 6816 4162 6868
rect 4214 6816 4222 6868
rect 4146 6810 4222 6816
rect 2746 6738 2796 6792
rect 4268 6766 4328 7096
rect 4390 7056 4436 7068
rect 2468 6691 2564 6738
rect 2468 6657 2524 6691
rect 2558 6657 2564 6691
rect 2468 6619 2564 6657
rect 2468 6585 2524 6619
rect 2558 6585 2564 6619
rect 2614 6691 2660 6738
rect 2614 6657 2620 6691
rect 2654 6657 2660 6691
rect 2614 6619 2660 6657
rect 2614 6598 2620 6619
rect 2468 6538 2564 6585
rect 2604 6590 2620 6598
rect 2654 6598 2660 6619
rect 2710 6691 2796 6738
rect 3800 6746 4328 6766
rect 3800 6712 3812 6746
rect 3846 6732 4328 6746
rect 3846 6712 3858 6732
rect 3800 6698 3858 6712
rect 2710 6657 2716 6691
rect 2750 6657 2796 6691
rect 2710 6619 2796 6657
rect 2654 6590 2670 6598
rect 2604 6538 2612 6590
rect 2664 6538 2670 6590
rect 2710 6585 2716 6619
rect 2750 6585 2796 6619
rect 2872 6659 2938 6672
rect 2872 6625 2888 6659
rect 2922 6625 2938 6659
rect 3266 6652 3334 6654
rect 2872 6614 2938 6625
rect 3182 6648 3334 6652
rect 3182 6642 3275 6648
rect 3182 6608 3202 6642
rect 3236 6608 3275 6642
rect 3182 6602 3275 6608
rect 3266 6596 3275 6602
rect 3327 6596 3334 6648
rect 3266 6590 3334 6596
rect 3370 6636 3444 6660
rect 3370 6602 3398 6636
rect 3432 6602 3444 6636
rect 2710 6542 2796 6585
rect 3370 6582 3444 6602
rect 3568 6652 3640 6664
rect 3568 6600 3579 6652
rect 3631 6600 3640 6652
rect 4114 6659 4180 6668
rect 4114 6625 4130 6659
rect 4164 6625 4180 6659
rect 4114 6612 4180 6625
rect 3568 6596 3640 6600
rect 2710 6538 2756 6542
rect 2604 6530 2670 6538
rect 2838 6531 2884 6578
rect 2380 6491 2618 6500
rect 2380 6468 2572 6491
rect 2280 6442 2286 6459
rect 1038 6376 1110 6404
rect 2192 6378 2238 6425
rect 2268 6436 2286 6442
rect 2320 6442 2326 6459
rect 2378 6457 2572 6468
rect 2606 6457 2618 6491
rect 2838 6497 2844 6531
rect 2878 6497 2884 6531
rect 2838 6464 2884 6497
rect 2320 6436 2334 6442
rect 2268 6384 2274 6436
rect 2326 6384 2334 6436
rect 2268 6378 2334 6384
rect 2378 6440 2618 6457
rect 726 6328 816 6349
rect 984 6331 1050 6340
rect 984 6297 1000 6331
rect 1034 6297 1050 6331
rect 984 6294 1050 6297
rect 490 6266 1050 6294
rect 394 6210 462 6224
rect 394 6176 412 6210
rect 446 6176 462 6210
rect 394 6166 462 6176
rect 434 5862 462 6166
rect 490 6084 524 6266
rect 822 6200 894 6212
rect 822 6148 832 6200
rect 884 6148 894 6200
rect 822 6136 894 6148
rect 746 6084 810 6102
rect 490 6050 762 6084
rect 796 6050 810 6084
rect 746 6040 810 6050
rect 1082 6026 1110 6376
rect 1150 6342 1426 6372
rect 1150 6341 1182 6342
rect 1234 6341 1426 6342
rect 1150 6307 1179 6341
rect 1234 6307 1271 6341
rect 1305 6307 1363 6341
rect 1397 6307 1426 6341
rect 1150 6290 1182 6307
rect 1234 6290 1426 6307
rect 1150 6276 1426 6290
rect 1494 6348 2118 6366
rect 1494 6335 2036 6348
rect 1494 6301 1525 6335
rect 1559 6301 1617 6335
rect 1651 6301 1709 6335
rect 1743 6333 2036 6335
rect 2088 6333 2118 6348
rect 1743 6301 1871 6333
rect 1494 6299 1871 6301
rect 1905 6299 1963 6333
rect 1997 6299 2036 6333
rect 2089 6299 2118 6333
rect 1494 6296 2036 6299
rect 2088 6296 2118 6299
rect 1200 6084 1266 6090
rect 1200 6032 1206 6084
rect 1258 6032 1266 6084
rect 1200 6026 1266 6032
rect 856 6012 1110 6026
rect 612 6000 658 6012
rect 158 5834 462 5862
rect 578 5966 618 6000
rect 652 5966 658 6000
rect 578 5928 658 5966
rect 698 6006 764 6012
rect 698 5954 704 6006
rect 756 5954 764 6006
rect 698 5948 764 5954
rect 804 6000 1110 6012
rect 804 5966 810 6000
rect 844 5998 1110 6000
rect 844 5966 906 5998
rect 578 5894 618 5928
rect 652 5894 658 5928
rect 578 5882 658 5894
rect 708 5928 754 5948
rect 708 5894 714 5928
rect 748 5894 754 5928
rect 708 5882 754 5894
rect 804 5928 906 5966
rect 804 5894 810 5928
rect 844 5894 906 5928
rect 804 5882 906 5894
rect 1026 5951 1260 5960
rect 1026 5899 1032 5951
rect 1084 5932 1208 5951
rect 1084 5899 1090 5932
rect 1026 5892 1090 5899
rect 1202 5899 1208 5932
rect 1260 5899 1266 5932
rect 1202 5892 1266 5899
rect 158 5831 434 5834
rect 158 5797 187 5831
rect 221 5797 279 5831
rect 313 5797 371 5831
rect 405 5797 434 5831
rect 158 5766 434 5797
rect 264 5718 328 5724
rect 264 5666 270 5718
rect 322 5666 328 5718
rect 264 5660 328 5666
rect 578 5682 624 5882
rect 654 5844 712 5854
rect 654 5810 666 5844
rect 700 5810 712 5844
rect 654 5792 712 5810
rect 766 5763 824 5780
rect 766 5729 778 5763
rect 812 5729 824 5763
rect 766 5714 824 5729
rect 856 5682 906 5882
rect 972 5831 1248 5862
rect 972 5797 1001 5831
rect 1035 5797 1093 5831
rect 1127 5797 1185 5831
rect 1219 5797 1248 5831
rect 972 5766 1248 5797
rect 578 5635 674 5682
rect 176 5602 240 5608
rect 176 5550 182 5602
rect 234 5550 240 5602
rect 176 5544 240 5550
rect 346 5592 416 5610
rect 346 5558 367 5592
rect 401 5558 416 5592
rect 346 5550 416 5558
rect 578 5601 634 5635
rect 668 5601 674 5635
rect 578 5563 674 5601
rect 346 5514 374 5550
rect 578 5529 634 5563
rect 668 5529 674 5563
rect 724 5635 770 5682
rect 724 5601 730 5635
rect 764 5601 770 5635
rect 724 5563 770 5601
rect 724 5542 730 5563
rect 578 5514 674 5529
rect 346 5482 674 5514
rect 714 5534 730 5542
rect 764 5542 770 5563
rect 820 5635 906 5682
rect 1078 5716 1146 5726
rect 1078 5664 1086 5716
rect 1138 5664 1146 5716
rect 1078 5658 1146 5664
rect 820 5601 826 5635
rect 860 5601 906 5635
rect 820 5563 906 5601
rect 764 5534 780 5542
rect 714 5482 722 5534
rect 774 5482 780 5534
rect 820 5529 826 5563
rect 860 5529 906 5563
rect 988 5604 1056 5610
rect 988 5552 994 5604
rect 1046 5552 1056 5604
rect 988 5546 1056 5552
rect 1162 5590 1228 5602
rect 1162 5556 1179 5590
rect 1213 5556 1228 5590
rect 1162 5548 1228 5556
rect 820 5510 906 5529
rect 1200 5510 1228 5548
rect 820 5482 1228 5510
rect 714 5474 780 5482
rect 862 5478 1228 5482
rect 666 5435 728 5444
rect 666 5401 682 5435
rect 716 5401 728 5435
rect 666 5384 728 5401
rect 670 5382 728 5384
rect 724 5327 814 5348
rect 724 5318 751 5327
rect -430 5293 751 5318
rect 785 5318 814 5327
rect 1328 5318 1406 6276
rect 1494 6264 2118 6296
rect 2226 6331 2292 6342
rect 2226 6297 2242 6331
rect 2276 6297 2292 6331
rect 2226 6286 2292 6297
rect 2378 6294 2412 6440
rect 2560 6438 2618 6440
rect 2816 6459 2884 6464
rect 2816 6456 2844 6459
rect 2816 6404 2824 6456
rect 2878 6425 2884 6459
rect 2876 6404 2884 6425
rect 2614 6383 2704 6404
rect 2816 6398 2884 6404
rect 2614 6349 2641 6383
rect 2675 6349 2704 6383
rect 2838 6378 2884 6398
rect 2926 6531 2972 6578
rect 2926 6497 2932 6531
rect 2966 6497 2972 6531
rect 2926 6459 2972 6497
rect 2926 6425 2932 6459
rect 2966 6425 2972 6459
rect 2926 6404 2972 6425
rect 4080 6531 4126 6578
rect 4080 6497 4086 6531
rect 4120 6497 4126 6531
rect 4080 6459 4126 6497
rect 4080 6425 4086 6459
rect 4120 6425 4126 6459
rect 4168 6531 4214 6578
rect 4168 6497 4174 6531
rect 4208 6497 4214 6531
rect 4168 6459 4214 6497
rect 4268 6500 4328 6732
rect 4356 7022 4396 7056
rect 4430 7022 4436 7056
rect 4356 6984 4436 7022
rect 4476 7062 4542 7068
rect 4476 7010 4482 7062
rect 4534 7010 4542 7062
rect 4476 7004 4542 7010
rect 4582 7056 4684 7068
rect 4582 7022 4588 7056
rect 4622 7022 4684 7056
rect 4356 6950 4396 6984
rect 4430 6950 4436 6984
rect 4356 6938 4436 6950
rect 4486 6984 4532 7004
rect 4486 6950 4492 6984
rect 4526 6950 4532 6984
rect 4486 6938 4532 6950
rect 4582 6984 4684 7022
rect 4582 6950 4588 6984
rect 4622 6950 4684 6984
rect 4582 6938 4684 6950
rect 4356 6738 4402 6938
rect 4432 6900 4490 6910
rect 4432 6866 4444 6900
rect 4478 6866 4490 6900
rect 4432 6848 4490 6866
rect 4634 6858 4684 6938
rect 5050 6916 5134 7186
rect 4792 6906 4850 6912
rect 4784 6900 4858 6906
rect 4544 6819 4602 6836
rect 4544 6785 4556 6819
rect 4590 6785 4602 6819
rect 4544 6770 4602 6785
rect 4634 6792 4704 6858
rect 4784 6848 4795 6900
rect 4847 6848 4858 6900
rect 4784 6842 4858 6848
rect 4926 6890 5202 6916
rect 5796 6910 5894 7186
rect 4926 6885 5027 6890
rect 5079 6885 5202 6890
rect 4926 6851 4955 6885
rect 4989 6851 5027 6885
rect 5081 6851 5139 6885
rect 5173 6851 5202 6885
rect 4792 6834 4850 6842
rect 4926 6838 5027 6851
rect 5079 6838 5202 6851
rect 4926 6820 5202 6838
rect 5272 6879 5894 6910
rect 5272 6845 5301 6879
rect 5335 6845 5393 6879
rect 5427 6845 5485 6879
rect 5519 6877 5894 6879
rect 5519 6845 5647 6877
rect 5272 6843 5647 6845
rect 5681 6843 5739 6877
rect 5773 6843 5831 6877
rect 5865 6843 5894 6877
rect 6156 7140 6476 7158
rect 6156 7106 6428 7140
rect 6462 7106 6476 7140
rect 6156 7096 6476 7106
rect 5272 6812 5894 6843
rect 6034 6868 6110 6874
rect 6034 6816 6050 6868
rect 6102 6816 6110 6868
rect 6034 6810 6110 6816
rect 4634 6738 4684 6792
rect 6156 6766 6216 7096
rect 6278 7056 6324 7068
rect 4356 6691 4452 6738
rect 4356 6657 4412 6691
rect 4446 6657 4452 6691
rect 4356 6619 4452 6657
rect 4356 6585 4412 6619
rect 4446 6585 4452 6619
rect 4502 6691 4548 6738
rect 4502 6657 4508 6691
rect 4542 6657 4548 6691
rect 4502 6619 4548 6657
rect 4502 6598 4508 6619
rect 4356 6538 4452 6585
rect 4492 6590 4508 6598
rect 4542 6598 4548 6619
rect 4598 6691 4684 6738
rect 5688 6746 6216 6766
rect 5688 6712 5700 6746
rect 5734 6732 6216 6746
rect 5734 6712 5746 6732
rect 5688 6698 5746 6712
rect 4598 6657 4604 6691
rect 4638 6657 4684 6691
rect 4598 6619 4684 6657
rect 4542 6590 4558 6598
rect 4492 6538 4500 6590
rect 4552 6538 4558 6590
rect 4598 6585 4604 6619
rect 4638 6585 4684 6619
rect 4760 6659 4826 6672
rect 4760 6625 4776 6659
rect 4810 6625 4826 6659
rect 5154 6652 5222 6654
rect 4760 6614 4826 6625
rect 5070 6648 5222 6652
rect 5070 6642 5163 6648
rect 5070 6608 5090 6642
rect 5124 6608 5163 6642
rect 5070 6602 5163 6608
rect 5154 6596 5163 6602
rect 5215 6596 5222 6648
rect 5154 6590 5222 6596
rect 5258 6636 5332 6660
rect 5258 6602 5286 6636
rect 5320 6602 5332 6636
rect 4598 6542 4684 6585
rect 5258 6582 5332 6602
rect 5456 6652 5528 6664
rect 5456 6600 5467 6652
rect 5519 6600 5528 6652
rect 6002 6659 6068 6668
rect 6002 6625 6018 6659
rect 6052 6625 6068 6659
rect 6002 6612 6068 6625
rect 5456 6596 5528 6600
rect 4598 6538 4644 6542
rect 4492 6530 4558 6538
rect 4726 6531 4772 6578
rect 4268 6491 4506 6500
rect 4268 6468 4460 6491
rect 4168 6442 4174 6459
rect 2926 6376 2998 6404
rect 4080 6378 4126 6425
rect 4156 6436 4174 6442
rect 4208 6442 4214 6459
rect 4266 6457 4460 6468
rect 4494 6457 4506 6491
rect 4726 6497 4732 6531
rect 4766 6497 4772 6531
rect 4726 6464 4772 6497
rect 4208 6436 4222 6442
rect 4156 6384 4162 6436
rect 4214 6384 4222 6436
rect 4156 6378 4222 6384
rect 4266 6440 4506 6457
rect 2614 6328 2704 6349
rect 2872 6331 2938 6340
rect 2872 6297 2888 6331
rect 2922 6297 2938 6331
rect 2872 6294 2938 6297
rect 2378 6266 2938 6294
rect 2282 6210 2350 6224
rect 2282 6176 2300 6210
rect 2334 6176 2350 6210
rect 2282 6166 2350 6176
rect 2322 5862 2350 6166
rect 2378 6084 2412 6266
rect 2710 6200 2782 6212
rect 2710 6148 2720 6200
rect 2772 6148 2782 6200
rect 2710 6136 2782 6148
rect 2634 6084 2698 6102
rect 2378 6050 2650 6084
rect 2684 6050 2698 6084
rect 2634 6040 2698 6050
rect 2970 6026 2998 6376
rect 3038 6342 3314 6372
rect 3038 6341 3070 6342
rect 3122 6341 3314 6342
rect 3038 6307 3067 6341
rect 3122 6307 3159 6341
rect 3193 6307 3251 6341
rect 3285 6307 3314 6341
rect 3038 6290 3070 6307
rect 3122 6290 3314 6307
rect 3038 6276 3314 6290
rect 3382 6348 4006 6366
rect 3382 6335 3924 6348
rect 3382 6301 3413 6335
rect 3447 6301 3505 6335
rect 3539 6301 3597 6335
rect 3631 6333 3924 6335
rect 3976 6333 4006 6348
rect 3631 6301 3759 6333
rect 3382 6299 3759 6301
rect 3793 6299 3851 6333
rect 3885 6299 3924 6333
rect 3977 6299 4006 6333
rect 3382 6296 3924 6299
rect 3976 6296 4006 6299
rect 3088 6084 3154 6090
rect 3088 6032 3094 6084
rect 3146 6032 3154 6084
rect 3088 6026 3154 6032
rect 2744 6012 2998 6026
rect 2500 6000 2546 6012
rect 2046 5834 2350 5862
rect 2466 5966 2506 6000
rect 2540 5966 2546 6000
rect 2466 5928 2546 5966
rect 2586 6006 2652 6012
rect 2586 5954 2592 6006
rect 2644 5954 2652 6006
rect 2586 5948 2652 5954
rect 2692 6000 2998 6012
rect 2692 5966 2698 6000
rect 2732 5998 2998 6000
rect 2732 5966 2794 5998
rect 2466 5894 2506 5928
rect 2540 5894 2546 5928
rect 2466 5882 2546 5894
rect 2596 5928 2642 5948
rect 2596 5894 2602 5928
rect 2636 5894 2642 5928
rect 2596 5882 2642 5894
rect 2692 5928 2794 5966
rect 2692 5894 2698 5928
rect 2732 5894 2794 5928
rect 2692 5882 2794 5894
rect 2914 5951 3148 5960
rect 2914 5899 2920 5951
rect 2972 5932 3096 5951
rect 2972 5899 2978 5932
rect 2914 5892 2978 5899
rect 3090 5899 3096 5932
rect 3148 5899 3154 5932
rect 3090 5892 3154 5899
rect 2046 5831 2322 5834
rect 2046 5797 2075 5831
rect 2109 5797 2167 5831
rect 2201 5797 2259 5831
rect 2293 5797 2322 5831
rect 2046 5766 2322 5797
rect 2152 5718 2216 5724
rect 2152 5666 2158 5718
rect 2210 5666 2216 5718
rect 2152 5660 2216 5666
rect 2466 5682 2512 5882
rect 2542 5844 2600 5854
rect 2542 5810 2554 5844
rect 2588 5810 2600 5844
rect 2542 5792 2600 5810
rect 2654 5763 2712 5780
rect 2654 5729 2666 5763
rect 2700 5729 2712 5763
rect 2654 5714 2712 5729
rect 2744 5682 2794 5882
rect 2860 5831 3136 5862
rect 2860 5797 2889 5831
rect 2923 5797 2981 5831
rect 3015 5797 3073 5831
rect 3107 5797 3136 5831
rect 2860 5766 3136 5797
rect 2466 5635 2562 5682
rect 2064 5602 2128 5608
rect 2064 5550 2070 5602
rect 2122 5550 2128 5602
rect 2064 5544 2128 5550
rect 2234 5592 2304 5610
rect 2234 5558 2255 5592
rect 2289 5558 2304 5592
rect 2234 5550 2304 5558
rect 2466 5601 2522 5635
rect 2556 5601 2562 5635
rect 2466 5563 2562 5601
rect 2234 5514 2262 5550
rect 2466 5529 2522 5563
rect 2556 5529 2562 5563
rect 2612 5635 2658 5682
rect 2612 5601 2618 5635
rect 2652 5601 2658 5635
rect 2612 5563 2658 5601
rect 2612 5542 2618 5563
rect 2466 5514 2562 5529
rect 2234 5482 2562 5514
rect 2602 5534 2618 5542
rect 2652 5542 2658 5563
rect 2708 5635 2794 5682
rect 2966 5716 3034 5726
rect 2966 5664 2974 5716
rect 3026 5664 3034 5716
rect 2966 5658 3034 5664
rect 2708 5601 2714 5635
rect 2748 5601 2794 5635
rect 2708 5563 2794 5601
rect 2652 5534 2668 5542
rect 2602 5482 2610 5534
rect 2662 5482 2668 5534
rect 2708 5529 2714 5563
rect 2748 5529 2794 5563
rect 2876 5604 2944 5610
rect 2876 5552 2882 5604
rect 2934 5552 2944 5604
rect 2876 5546 2944 5552
rect 3050 5590 3116 5602
rect 3050 5556 3067 5590
rect 3101 5556 3116 5590
rect 3050 5548 3116 5556
rect 2708 5510 2794 5529
rect 3088 5510 3116 5548
rect 2708 5482 3116 5510
rect 2602 5474 2668 5482
rect 2750 5478 3116 5482
rect 2554 5435 2616 5444
rect 2554 5401 2570 5435
rect 2604 5401 2616 5435
rect 2554 5384 2616 5401
rect 2558 5382 2616 5384
rect 2612 5327 2702 5348
rect 2612 5318 2639 5327
rect 785 5293 2639 5318
rect 2673 5318 2702 5327
rect 3216 5318 3294 6276
rect 3382 6264 4006 6296
rect 4114 6331 4180 6342
rect 4114 6297 4130 6331
rect 4164 6297 4180 6331
rect 4114 6286 4180 6297
rect 4266 6294 4300 6440
rect 4448 6438 4506 6440
rect 4704 6459 4772 6464
rect 4704 6456 4732 6459
rect 4704 6404 4712 6456
rect 4766 6425 4772 6459
rect 4764 6404 4772 6425
rect 4502 6383 4592 6404
rect 4704 6398 4772 6404
rect 4502 6349 4529 6383
rect 4563 6349 4592 6383
rect 4726 6378 4772 6398
rect 4814 6531 4860 6578
rect 4814 6497 4820 6531
rect 4854 6497 4860 6531
rect 4814 6459 4860 6497
rect 4814 6425 4820 6459
rect 4854 6425 4860 6459
rect 4814 6404 4860 6425
rect 5968 6531 6014 6578
rect 5968 6497 5974 6531
rect 6008 6497 6014 6531
rect 5968 6459 6014 6497
rect 5968 6425 5974 6459
rect 6008 6425 6014 6459
rect 6056 6531 6102 6578
rect 6056 6497 6062 6531
rect 6096 6497 6102 6531
rect 6056 6459 6102 6497
rect 6156 6500 6216 6732
rect 6244 7022 6284 7056
rect 6318 7022 6324 7056
rect 6244 6984 6324 7022
rect 6364 7062 6430 7068
rect 6364 7010 6370 7062
rect 6422 7010 6430 7062
rect 6364 7004 6430 7010
rect 6470 7056 6572 7068
rect 6470 7022 6476 7056
rect 6510 7022 6572 7056
rect 6244 6950 6284 6984
rect 6318 6950 6324 6984
rect 6244 6938 6324 6950
rect 6374 6984 6420 7004
rect 6374 6950 6380 6984
rect 6414 6950 6420 6984
rect 6374 6938 6420 6950
rect 6470 6984 6572 7022
rect 6470 6950 6476 6984
rect 6510 6950 6572 6984
rect 6470 6938 6572 6950
rect 6244 6738 6290 6938
rect 6320 6900 6378 6910
rect 6320 6866 6332 6900
rect 6366 6866 6378 6900
rect 6320 6848 6378 6866
rect 6522 6858 6572 6938
rect 6938 6916 7022 7186
rect 6680 6906 6738 6912
rect 6672 6900 6746 6906
rect 6432 6819 6490 6836
rect 6432 6785 6444 6819
rect 6478 6785 6490 6819
rect 6432 6770 6490 6785
rect 6522 6792 6592 6858
rect 6672 6848 6683 6900
rect 6735 6848 6746 6900
rect 6672 6842 6746 6848
rect 6814 6890 7090 6916
rect 7684 6910 7782 7186
rect 6814 6885 6915 6890
rect 6967 6885 7090 6890
rect 6814 6851 6843 6885
rect 6877 6851 6915 6885
rect 6969 6851 7027 6885
rect 7061 6851 7090 6885
rect 6680 6834 6738 6842
rect 6814 6838 6915 6851
rect 6967 6838 7090 6851
rect 6814 6820 7090 6838
rect 7160 6879 7782 6910
rect 7160 6845 7189 6879
rect 7223 6845 7281 6879
rect 7315 6845 7373 6879
rect 7407 6877 7782 6879
rect 7407 6845 7535 6877
rect 7160 6843 7535 6845
rect 7569 6843 7627 6877
rect 7661 6843 7719 6877
rect 7753 6843 7782 6877
rect 8044 7140 8364 7158
rect 8044 7106 8316 7140
rect 8350 7106 8364 7140
rect 8044 7096 8364 7106
rect 7160 6812 7782 6843
rect 7922 6868 7998 6874
rect 7922 6816 7938 6868
rect 7990 6816 7998 6868
rect 7922 6810 7998 6816
rect 6522 6738 6572 6792
rect 8044 6766 8104 7096
rect 8166 7056 8212 7068
rect 6244 6691 6340 6738
rect 6244 6657 6300 6691
rect 6334 6657 6340 6691
rect 6244 6619 6340 6657
rect 6244 6585 6300 6619
rect 6334 6585 6340 6619
rect 6390 6691 6436 6738
rect 6390 6657 6396 6691
rect 6430 6657 6436 6691
rect 6390 6619 6436 6657
rect 6390 6598 6396 6619
rect 6244 6538 6340 6585
rect 6380 6590 6396 6598
rect 6430 6598 6436 6619
rect 6486 6691 6572 6738
rect 7576 6746 8104 6766
rect 7576 6712 7588 6746
rect 7622 6732 8104 6746
rect 7622 6712 7634 6732
rect 7576 6698 7634 6712
rect 6486 6657 6492 6691
rect 6526 6657 6572 6691
rect 6486 6619 6572 6657
rect 6430 6590 6446 6598
rect 6380 6538 6388 6590
rect 6440 6538 6446 6590
rect 6486 6585 6492 6619
rect 6526 6585 6572 6619
rect 6648 6659 6714 6672
rect 6648 6625 6664 6659
rect 6698 6625 6714 6659
rect 7042 6652 7110 6654
rect 6648 6614 6714 6625
rect 6958 6648 7110 6652
rect 6958 6642 7051 6648
rect 6958 6608 6978 6642
rect 7012 6608 7051 6642
rect 6958 6602 7051 6608
rect 7042 6596 7051 6602
rect 7103 6596 7110 6648
rect 7042 6590 7110 6596
rect 7146 6636 7220 6660
rect 7146 6602 7174 6636
rect 7208 6602 7220 6636
rect 6486 6542 6572 6585
rect 7146 6582 7220 6602
rect 7344 6652 7416 6664
rect 7344 6600 7355 6652
rect 7407 6600 7416 6652
rect 7890 6659 7956 6668
rect 7890 6625 7906 6659
rect 7940 6625 7956 6659
rect 7890 6612 7956 6625
rect 7344 6596 7416 6600
rect 6486 6538 6532 6542
rect 6380 6530 6446 6538
rect 6614 6531 6660 6578
rect 6156 6491 6394 6500
rect 6156 6468 6348 6491
rect 6056 6442 6062 6459
rect 4814 6376 4886 6404
rect 5968 6378 6014 6425
rect 6044 6436 6062 6442
rect 6096 6442 6102 6459
rect 6154 6457 6348 6468
rect 6382 6457 6394 6491
rect 6614 6497 6620 6531
rect 6654 6497 6660 6531
rect 6614 6464 6660 6497
rect 6096 6436 6110 6442
rect 6044 6384 6050 6436
rect 6102 6384 6110 6436
rect 6044 6378 6110 6384
rect 6154 6440 6394 6457
rect 4502 6328 4592 6349
rect 4760 6331 4826 6340
rect 4760 6297 4776 6331
rect 4810 6297 4826 6331
rect 4760 6294 4826 6297
rect 4266 6266 4826 6294
rect 4170 6210 4238 6224
rect 4170 6176 4188 6210
rect 4222 6176 4238 6210
rect 4170 6166 4238 6176
rect 4210 5862 4238 6166
rect 4266 6084 4300 6266
rect 4598 6200 4670 6212
rect 4598 6148 4608 6200
rect 4660 6148 4670 6200
rect 4598 6136 4670 6148
rect 4522 6084 4586 6102
rect 4266 6050 4538 6084
rect 4572 6050 4586 6084
rect 4522 6040 4586 6050
rect 4858 6026 4886 6376
rect 4926 6342 5202 6372
rect 4926 6341 4958 6342
rect 5010 6341 5202 6342
rect 4926 6307 4955 6341
rect 5010 6307 5047 6341
rect 5081 6307 5139 6341
rect 5173 6307 5202 6341
rect 4926 6290 4958 6307
rect 5010 6290 5202 6307
rect 4926 6276 5202 6290
rect 5270 6348 5894 6366
rect 5270 6335 5812 6348
rect 5270 6301 5301 6335
rect 5335 6301 5393 6335
rect 5427 6301 5485 6335
rect 5519 6333 5812 6335
rect 5864 6333 5894 6348
rect 5519 6301 5647 6333
rect 5270 6299 5647 6301
rect 5681 6299 5739 6333
rect 5773 6299 5812 6333
rect 5865 6299 5894 6333
rect 5270 6296 5812 6299
rect 5864 6296 5894 6299
rect 4976 6084 5042 6090
rect 4976 6032 4982 6084
rect 5034 6032 5042 6084
rect 4976 6026 5042 6032
rect 4632 6012 4886 6026
rect 4388 6000 4434 6012
rect 3934 5834 4238 5862
rect 4354 5966 4394 6000
rect 4428 5966 4434 6000
rect 4354 5928 4434 5966
rect 4474 6006 4540 6012
rect 4474 5954 4480 6006
rect 4532 5954 4540 6006
rect 4474 5948 4540 5954
rect 4580 6000 4886 6012
rect 4580 5966 4586 6000
rect 4620 5998 4886 6000
rect 4620 5966 4682 5998
rect 4354 5894 4394 5928
rect 4428 5894 4434 5928
rect 4354 5882 4434 5894
rect 4484 5928 4530 5948
rect 4484 5894 4490 5928
rect 4524 5894 4530 5928
rect 4484 5882 4530 5894
rect 4580 5928 4682 5966
rect 4580 5894 4586 5928
rect 4620 5894 4682 5928
rect 4580 5882 4682 5894
rect 4802 5951 5036 5960
rect 4802 5899 4808 5951
rect 4860 5932 4984 5951
rect 4860 5899 4866 5932
rect 4802 5892 4866 5899
rect 4978 5899 4984 5932
rect 5036 5899 5042 5932
rect 4978 5892 5042 5899
rect 3934 5831 4210 5834
rect 3934 5797 3963 5831
rect 3997 5797 4055 5831
rect 4089 5797 4147 5831
rect 4181 5797 4210 5831
rect 3934 5766 4210 5797
rect 4040 5718 4104 5724
rect 4040 5666 4046 5718
rect 4098 5666 4104 5718
rect 4040 5660 4104 5666
rect 4354 5682 4400 5882
rect 4430 5844 4488 5854
rect 4430 5810 4442 5844
rect 4476 5810 4488 5844
rect 4430 5792 4488 5810
rect 4542 5763 4600 5780
rect 4542 5729 4554 5763
rect 4588 5729 4600 5763
rect 4542 5714 4600 5729
rect 4632 5682 4682 5882
rect 4748 5831 5024 5862
rect 4748 5797 4777 5831
rect 4811 5797 4869 5831
rect 4903 5797 4961 5831
rect 4995 5797 5024 5831
rect 4748 5766 5024 5797
rect 4354 5635 4450 5682
rect 3952 5602 4016 5608
rect 3952 5550 3958 5602
rect 4010 5550 4016 5602
rect 3952 5544 4016 5550
rect 4122 5592 4192 5610
rect 4122 5558 4143 5592
rect 4177 5558 4192 5592
rect 4122 5550 4192 5558
rect 4354 5601 4410 5635
rect 4444 5601 4450 5635
rect 4354 5563 4450 5601
rect 4122 5514 4150 5550
rect 4354 5529 4410 5563
rect 4444 5529 4450 5563
rect 4500 5635 4546 5682
rect 4500 5601 4506 5635
rect 4540 5601 4546 5635
rect 4500 5563 4546 5601
rect 4500 5542 4506 5563
rect 4354 5514 4450 5529
rect 4122 5482 4450 5514
rect 4490 5534 4506 5542
rect 4540 5542 4546 5563
rect 4596 5635 4682 5682
rect 4854 5716 4922 5726
rect 4854 5664 4862 5716
rect 4914 5664 4922 5716
rect 4854 5658 4922 5664
rect 4596 5601 4602 5635
rect 4636 5601 4682 5635
rect 4596 5563 4682 5601
rect 4540 5534 4556 5542
rect 4490 5482 4498 5534
rect 4550 5482 4556 5534
rect 4596 5529 4602 5563
rect 4636 5529 4682 5563
rect 4764 5604 4832 5610
rect 4764 5552 4770 5604
rect 4822 5552 4832 5604
rect 4764 5546 4832 5552
rect 4938 5590 5004 5602
rect 4938 5556 4955 5590
rect 4989 5556 5004 5590
rect 4938 5548 5004 5556
rect 4596 5510 4682 5529
rect 4976 5510 5004 5548
rect 4596 5482 5004 5510
rect 4490 5474 4556 5482
rect 4638 5478 5004 5482
rect 4442 5435 4504 5444
rect 4442 5401 4458 5435
rect 4492 5401 4504 5435
rect 4442 5384 4504 5401
rect 4446 5382 4504 5384
rect 4500 5327 4590 5348
rect 4500 5318 4527 5327
rect 2673 5293 4527 5318
rect 4561 5318 4590 5327
rect 5104 5318 5182 6276
rect 5270 6264 5894 6296
rect 6002 6331 6068 6342
rect 6002 6297 6018 6331
rect 6052 6297 6068 6331
rect 6002 6286 6068 6297
rect 6154 6294 6188 6440
rect 6336 6438 6394 6440
rect 6592 6459 6660 6464
rect 6592 6456 6620 6459
rect 6592 6404 6600 6456
rect 6654 6425 6660 6459
rect 6652 6404 6660 6425
rect 6390 6383 6480 6404
rect 6592 6398 6660 6404
rect 6390 6349 6417 6383
rect 6451 6349 6480 6383
rect 6614 6378 6660 6398
rect 6702 6531 6748 6578
rect 6702 6497 6708 6531
rect 6742 6497 6748 6531
rect 6702 6459 6748 6497
rect 6702 6425 6708 6459
rect 6742 6425 6748 6459
rect 6702 6404 6748 6425
rect 7856 6531 7902 6578
rect 7856 6497 7862 6531
rect 7896 6497 7902 6531
rect 7856 6459 7902 6497
rect 7856 6425 7862 6459
rect 7896 6425 7902 6459
rect 7944 6531 7990 6578
rect 7944 6497 7950 6531
rect 7984 6497 7990 6531
rect 7944 6459 7990 6497
rect 8044 6500 8104 6732
rect 8132 7022 8172 7056
rect 8206 7022 8212 7056
rect 8132 6984 8212 7022
rect 8252 7062 8318 7068
rect 8252 7010 8258 7062
rect 8310 7010 8318 7062
rect 8252 7004 8318 7010
rect 8358 7056 8460 7068
rect 8358 7022 8364 7056
rect 8398 7022 8460 7056
rect 8132 6950 8172 6984
rect 8206 6950 8212 6984
rect 8132 6938 8212 6950
rect 8262 6984 8308 7004
rect 8262 6950 8268 6984
rect 8302 6950 8308 6984
rect 8262 6938 8308 6950
rect 8358 6984 8460 7022
rect 8358 6950 8364 6984
rect 8398 6950 8460 6984
rect 8358 6938 8460 6950
rect 8132 6738 8178 6938
rect 8208 6900 8266 6910
rect 8208 6866 8220 6900
rect 8254 6866 8266 6900
rect 8208 6848 8266 6866
rect 8410 6858 8460 6938
rect 8826 6916 8910 7186
rect 8568 6906 8626 6912
rect 8560 6900 8634 6906
rect 8320 6819 8378 6836
rect 8320 6785 8332 6819
rect 8366 6785 8378 6819
rect 8320 6770 8378 6785
rect 8410 6792 8480 6858
rect 8560 6848 8571 6900
rect 8623 6848 8634 6900
rect 8560 6842 8634 6848
rect 8702 6890 8978 6916
rect 9572 6910 9670 7186
rect 8702 6885 8803 6890
rect 8855 6885 8978 6890
rect 8702 6851 8731 6885
rect 8765 6851 8803 6885
rect 8857 6851 8915 6885
rect 8949 6851 8978 6885
rect 8568 6834 8626 6842
rect 8702 6838 8803 6851
rect 8855 6838 8978 6851
rect 8702 6820 8978 6838
rect 9048 6879 9670 6910
rect 9048 6845 9077 6879
rect 9111 6845 9169 6879
rect 9203 6845 9261 6879
rect 9295 6877 9670 6879
rect 9295 6845 9423 6877
rect 9048 6843 9423 6845
rect 9457 6843 9515 6877
rect 9549 6843 9607 6877
rect 9641 6843 9670 6877
rect 9932 7140 10252 7158
rect 9932 7106 10204 7140
rect 10238 7106 10252 7140
rect 9932 7096 10252 7106
rect 9048 6812 9670 6843
rect 9810 6868 9886 6874
rect 9810 6816 9826 6868
rect 9878 6816 9886 6868
rect 9810 6810 9886 6816
rect 8410 6738 8460 6792
rect 9932 6766 9992 7096
rect 10054 7056 10100 7068
rect 8132 6691 8228 6738
rect 8132 6657 8188 6691
rect 8222 6657 8228 6691
rect 8132 6619 8228 6657
rect 8132 6585 8188 6619
rect 8222 6585 8228 6619
rect 8278 6691 8324 6738
rect 8278 6657 8284 6691
rect 8318 6657 8324 6691
rect 8278 6619 8324 6657
rect 8278 6598 8284 6619
rect 8132 6538 8228 6585
rect 8268 6590 8284 6598
rect 8318 6598 8324 6619
rect 8374 6691 8460 6738
rect 9464 6746 9992 6766
rect 9464 6712 9476 6746
rect 9510 6732 9992 6746
rect 9510 6712 9522 6732
rect 9464 6698 9522 6712
rect 8374 6657 8380 6691
rect 8414 6657 8460 6691
rect 8374 6619 8460 6657
rect 8318 6590 8334 6598
rect 8268 6538 8276 6590
rect 8328 6538 8334 6590
rect 8374 6585 8380 6619
rect 8414 6585 8460 6619
rect 8536 6659 8602 6672
rect 8536 6625 8552 6659
rect 8586 6625 8602 6659
rect 8930 6652 8998 6654
rect 8536 6614 8602 6625
rect 8846 6648 8998 6652
rect 8846 6642 8939 6648
rect 8846 6608 8866 6642
rect 8900 6608 8939 6642
rect 8846 6602 8939 6608
rect 8930 6596 8939 6602
rect 8991 6596 8998 6648
rect 8930 6590 8998 6596
rect 9034 6636 9108 6660
rect 9034 6602 9062 6636
rect 9096 6602 9108 6636
rect 8374 6542 8460 6585
rect 9034 6582 9108 6602
rect 9232 6652 9304 6664
rect 9232 6600 9243 6652
rect 9295 6600 9304 6652
rect 9778 6659 9844 6668
rect 9778 6625 9794 6659
rect 9828 6625 9844 6659
rect 9778 6612 9844 6625
rect 9232 6596 9304 6600
rect 8374 6538 8420 6542
rect 8268 6530 8334 6538
rect 8502 6531 8548 6578
rect 8044 6491 8282 6500
rect 8044 6468 8236 6491
rect 7944 6442 7950 6459
rect 6702 6376 6774 6404
rect 7856 6378 7902 6425
rect 7932 6436 7950 6442
rect 7984 6442 7990 6459
rect 8042 6457 8236 6468
rect 8270 6457 8282 6491
rect 8502 6497 8508 6531
rect 8542 6497 8548 6531
rect 8502 6464 8548 6497
rect 7984 6436 7998 6442
rect 7932 6384 7938 6436
rect 7990 6384 7998 6436
rect 7932 6378 7998 6384
rect 8042 6440 8282 6457
rect 6390 6328 6480 6349
rect 6648 6331 6714 6340
rect 6648 6297 6664 6331
rect 6698 6297 6714 6331
rect 6648 6294 6714 6297
rect 6154 6266 6714 6294
rect 6058 6210 6126 6224
rect 6058 6176 6076 6210
rect 6110 6176 6126 6210
rect 6058 6166 6126 6176
rect 6098 5862 6126 6166
rect 6154 6084 6188 6266
rect 6486 6200 6558 6212
rect 6486 6148 6496 6200
rect 6548 6148 6558 6200
rect 6486 6136 6558 6148
rect 6410 6084 6474 6102
rect 6154 6050 6426 6084
rect 6460 6050 6474 6084
rect 6410 6040 6474 6050
rect 6746 6026 6774 6376
rect 6814 6342 7090 6372
rect 6814 6341 6846 6342
rect 6898 6341 7090 6342
rect 6814 6307 6843 6341
rect 6898 6307 6935 6341
rect 6969 6307 7027 6341
rect 7061 6307 7090 6341
rect 6814 6290 6846 6307
rect 6898 6290 7090 6307
rect 6814 6276 7090 6290
rect 7158 6348 7782 6366
rect 7158 6335 7700 6348
rect 7158 6301 7189 6335
rect 7223 6301 7281 6335
rect 7315 6301 7373 6335
rect 7407 6333 7700 6335
rect 7752 6333 7782 6348
rect 7407 6301 7535 6333
rect 7158 6299 7535 6301
rect 7569 6299 7627 6333
rect 7661 6299 7700 6333
rect 7753 6299 7782 6333
rect 7158 6296 7700 6299
rect 7752 6296 7782 6299
rect 6864 6084 6930 6090
rect 6864 6032 6870 6084
rect 6922 6032 6930 6084
rect 6864 6026 6930 6032
rect 6520 6012 6774 6026
rect 6276 6000 6322 6012
rect 5822 5834 6126 5862
rect 6242 5966 6282 6000
rect 6316 5966 6322 6000
rect 6242 5928 6322 5966
rect 6362 6006 6428 6012
rect 6362 5954 6368 6006
rect 6420 5954 6428 6006
rect 6362 5948 6428 5954
rect 6468 6000 6774 6012
rect 6468 5966 6474 6000
rect 6508 5998 6774 6000
rect 6508 5966 6570 5998
rect 6242 5894 6282 5928
rect 6316 5894 6322 5928
rect 6242 5882 6322 5894
rect 6372 5928 6418 5948
rect 6372 5894 6378 5928
rect 6412 5894 6418 5928
rect 6372 5882 6418 5894
rect 6468 5928 6570 5966
rect 6468 5894 6474 5928
rect 6508 5894 6570 5928
rect 6468 5882 6570 5894
rect 6690 5951 6924 5960
rect 6690 5899 6696 5951
rect 6748 5932 6872 5951
rect 6748 5899 6754 5932
rect 6690 5892 6754 5899
rect 6866 5899 6872 5932
rect 6924 5899 6930 5932
rect 6866 5892 6930 5899
rect 5822 5831 6098 5834
rect 5822 5797 5851 5831
rect 5885 5797 5943 5831
rect 5977 5797 6035 5831
rect 6069 5797 6098 5831
rect 5822 5766 6098 5797
rect 5928 5718 5992 5724
rect 5928 5666 5934 5718
rect 5986 5666 5992 5718
rect 5928 5660 5992 5666
rect 6242 5682 6288 5882
rect 6318 5844 6376 5854
rect 6318 5810 6330 5844
rect 6364 5810 6376 5844
rect 6318 5792 6376 5810
rect 6430 5763 6488 5780
rect 6430 5729 6442 5763
rect 6476 5729 6488 5763
rect 6430 5714 6488 5729
rect 6520 5682 6570 5882
rect 6636 5831 6912 5862
rect 6636 5797 6665 5831
rect 6699 5797 6757 5831
rect 6791 5797 6849 5831
rect 6883 5797 6912 5831
rect 6636 5766 6912 5797
rect 6242 5635 6338 5682
rect 5840 5602 5904 5608
rect 5840 5550 5846 5602
rect 5898 5550 5904 5602
rect 5840 5544 5904 5550
rect 6010 5592 6080 5610
rect 6010 5558 6031 5592
rect 6065 5558 6080 5592
rect 6010 5550 6080 5558
rect 6242 5601 6298 5635
rect 6332 5601 6338 5635
rect 6242 5563 6338 5601
rect 6010 5514 6038 5550
rect 6242 5529 6298 5563
rect 6332 5529 6338 5563
rect 6388 5635 6434 5682
rect 6388 5601 6394 5635
rect 6428 5601 6434 5635
rect 6388 5563 6434 5601
rect 6388 5542 6394 5563
rect 6242 5514 6338 5529
rect 6010 5482 6338 5514
rect 6378 5534 6394 5542
rect 6428 5542 6434 5563
rect 6484 5635 6570 5682
rect 6742 5716 6810 5726
rect 6742 5664 6750 5716
rect 6802 5664 6810 5716
rect 6742 5658 6810 5664
rect 6484 5601 6490 5635
rect 6524 5601 6570 5635
rect 6484 5563 6570 5601
rect 6428 5534 6444 5542
rect 6378 5482 6386 5534
rect 6438 5482 6444 5534
rect 6484 5529 6490 5563
rect 6524 5529 6570 5563
rect 6652 5604 6720 5610
rect 6652 5552 6658 5604
rect 6710 5552 6720 5604
rect 6652 5546 6720 5552
rect 6826 5590 6892 5602
rect 6826 5556 6843 5590
rect 6877 5556 6892 5590
rect 6826 5548 6892 5556
rect 6484 5510 6570 5529
rect 6864 5510 6892 5548
rect 6484 5482 6892 5510
rect 6378 5474 6444 5482
rect 6526 5478 6892 5482
rect 6330 5435 6392 5444
rect 6330 5401 6346 5435
rect 6380 5401 6392 5435
rect 6330 5384 6392 5401
rect 6334 5382 6392 5384
rect 6388 5327 6478 5348
rect 6388 5318 6415 5327
rect 4561 5293 6415 5318
rect 6449 5318 6478 5327
rect 6992 5318 7070 6276
rect 7158 6264 7782 6296
rect 7890 6331 7956 6342
rect 7890 6297 7906 6331
rect 7940 6297 7956 6331
rect 7890 6286 7956 6297
rect 8042 6294 8076 6440
rect 8224 6438 8282 6440
rect 8480 6459 8548 6464
rect 8480 6456 8508 6459
rect 8480 6404 8488 6456
rect 8542 6425 8548 6459
rect 8540 6404 8548 6425
rect 8278 6383 8368 6404
rect 8480 6398 8548 6404
rect 8278 6349 8305 6383
rect 8339 6349 8368 6383
rect 8502 6378 8548 6398
rect 8590 6531 8636 6578
rect 8590 6497 8596 6531
rect 8630 6497 8636 6531
rect 8590 6459 8636 6497
rect 8590 6425 8596 6459
rect 8630 6425 8636 6459
rect 8590 6404 8636 6425
rect 9744 6531 9790 6578
rect 9744 6497 9750 6531
rect 9784 6497 9790 6531
rect 9744 6459 9790 6497
rect 9744 6425 9750 6459
rect 9784 6425 9790 6459
rect 9832 6531 9878 6578
rect 9832 6497 9838 6531
rect 9872 6497 9878 6531
rect 9832 6459 9878 6497
rect 9932 6500 9992 6732
rect 10020 7022 10060 7056
rect 10094 7022 10100 7056
rect 10020 6984 10100 7022
rect 10140 7062 10206 7068
rect 10140 7010 10146 7062
rect 10198 7010 10206 7062
rect 10140 7004 10206 7010
rect 10246 7056 10348 7068
rect 10246 7022 10252 7056
rect 10286 7022 10348 7056
rect 10020 6950 10060 6984
rect 10094 6950 10100 6984
rect 10020 6938 10100 6950
rect 10150 6984 10196 7004
rect 10150 6950 10156 6984
rect 10190 6950 10196 6984
rect 10150 6938 10196 6950
rect 10246 6984 10348 7022
rect 10246 6950 10252 6984
rect 10286 6950 10348 6984
rect 10246 6938 10348 6950
rect 10020 6738 10066 6938
rect 10096 6900 10154 6910
rect 10096 6866 10108 6900
rect 10142 6866 10154 6900
rect 10096 6848 10154 6866
rect 10298 6858 10348 6938
rect 10714 6916 10798 7186
rect 10456 6906 10514 6912
rect 10448 6900 10522 6906
rect 10208 6819 10266 6836
rect 10208 6785 10220 6819
rect 10254 6785 10266 6819
rect 10208 6770 10266 6785
rect 10298 6792 10368 6858
rect 10448 6848 10459 6900
rect 10511 6848 10522 6900
rect 10448 6842 10522 6848
rect 10590 6890 10866 6916
rect 11460 6910 11558 7186
rect 10590 6885 10691 6890
rect 10743 6885 10866 6890
rect 10590 6851 10619 6885
rect 10653 6851 10691 6885
rect 10745 6851 10803 6885
rect 10837 6851 10866 6885
rect 10456 6834 10514 6842
rect 10590 6838 10691 6851
rect 10743 6838 10866 6851
rect 10590 6820 10866 6838
rect 10936 6879 11558 6910
rect 10936 6845 10965 6879
rect 10999 6845 11057 6879
rect 11091 6845 11149 6879
rect 11183 6877 11558 6879
rect 11183 6845 11311 6877
rect 10936 6843 11311 6845
rect 11345 6843 11403 6877
rect 11437 6843 11495 6877
rect 11529 6843 11558 6877
rect 11820 7140 12140 7158
rect 11820 7106 12092 7140
rect 12126 7106 12140 7140
rect 11820 7096 12140 7106
rect 10936 6812 11558 6843
rect 11698 6868 11774 6874
rect 11698 6816 11714 6868
rect 11766 6816 11774 6868
rect 11698 6810 11774 6816
rect 10298 6738 10348 6792
rect 11820 6766 11880 7096
rect 11942 7056 11988 7068
rect 10020 6691 10116 6738
rect 10020 6657 10076 6691
rect 10110 6657 10116 6691
rect 10020 6619 10116 6657
rect 10020 6585 10076 6619
rect 10110 6585 10116 6619
rect 10166 6691 10212 6738
rect 10166 6657 10172 6691
rect 10206 6657 10212 6691
rect 10166 6619 10212 6657
rect 10166 6598 10172 6619
rect 10020 6538 10116 6585
rect 10156 6590 10172 6598
rect 10206 6598 10212 6619
rect 10262 6691 10348 6738
rect 11352 6746 11880 6766
rect 11352 6712 11364 6746
rect 11398 6732 11880 6746
rect 11398 6712 11410 6732
rect 11352 6698 11410 6712
rect 10262 6657 10268 6691
rect 10302 6657 10348 6691
rect 10262 6619 10348 6657
rect 10206 6590 10222 6598
rect 10156 6538 10164 6590
rect 10216 6538 10222 6590
rect 10262 6585 10268 6619
rect 10302 6585 10348 6619
rect 10424 6659 10490 6672
rect 10424 6625 10440 6659
rect 10474 6625 10490 6659
rect 10818 6652 10886 6654
rect 10424 6614 10490 6625
rect 10734 6648 10886 6652
rect 10734 6642 10827 6648
rect 10734 6608 10754 6642
rect 10788 6608 10827 6642
rect 10734 6602 10827 6608
rect 10818 6596 10827 6602
rect 10879 6596 10886 6648
rect 10818 6590 10886 6596
rect 10922 6636 10996 6660
rect 10922 6602 10950 6636
rect 10984 6602 10996 6636
rect 10262 6542 10348 6585
rect 10922 6582 10996 6602
rect 11120 6652 11192 6664
rect 11120 6600 11131 6652
rect 11183 6600 11192 6652
rect 11666 6659 11732 6668
rect 11666 6625 11682 6659
rect 11716 6625 11732 6659
rect 11666 6612 11732 6625
rect 11120 6596 11192 6600
rect 10262 6538 10308 6542
rect 10156 6530 10222 6538
rect 10390 6531 10436 6578
rect 9932 6491 10170 6500
rect 9932 6468 10124 6491
rect 9832 6442 9838 6459
rect 8590 6376 8662 6404
rect 9744 6378 9790 6425
rect 9820 6436 9838 6442
rect 9872 6442 9878 6459
rect 9930 6457 10124 6468
rect 10158 6457 10170 6491
rect 10390 6497 10396 6531
rect 10430 6497 10436 6531
rect 10390 6464 10436 6497
rect 9872 6436 9886 6442
rect 9820 6384 9826 6436
rect 9878 6384 9886 6436
rect 9820 6378 9886 6384
rect 9930 6440 10170 6457
rect 8278 6328 8368 6349
rect 8536 6331 8602 6340
rect 8536 6297 8552 6331
rect 8586 6297 8602 6331
rect 8536 6294 8602 6297
rect 8042 6266 8602 6294
rect 7946 6210 8014 6224
rect 7946 6176 7964 6210
rect 7998 6176 8014 6210
rect 7946 6166 8014 6176
rect 7986 5862 8014 6166
rect 8042 6084 8076 6266
rect 8374 6200 8446 6212
rect 8374 6148 8384 6200
rect 8436 6148 8446 6200
rect 8374 6136 8446 6148
rect 8298 6084 8362 6102
rect 8042 6050 8314 6084
rect 8348 6050 8362 6084
rect 8298 6040 8362 6050
rect 8634 6026 8662 6376
rect 8702 6342 8978 6372
rect 8702 6341 8734 6342
rect 8786 6341 8978 6342
rect 8702 6307 8731 6341
rect 8786 6307 8823 6341
rect 8857 6307 8915 6341
rect 8949 6307 8978 6341
rect 8702 6290 8734 6307
rect 8786 6290 8978 6307
rect 8702 6276 8978 6290
rect 9046 6348 9670 6366
rect 9046 6335 9588 6348
rect 9046 6301 9077 6335
rect 9111 6301 9169 6335
rect 9203 6301 9261 6335
rect 9295 6333 9588 6335
rect 9640 6333 9670 6348
rect 9295 6301 9423 6333
rect 9046 6299 9423 6301
rect 9457 6299 9515 6333
rect 9549 6299 9588 6333
rect 9641 6299 9670 6333
rect 9046 6296 9588 6299
rect 9640 6296 9670 6299
rect 8752 6084 8818 6090
rect 8752 6032 8758 6084
rect 8810 6032 8818 6084
rect 8752 6026 8818 6032
rect 8408 6012 8662 6026
rect 8164 6000 8210 6012
rect 7710 5834 8014 5862
rect 8130 5966 8170 6000
rect 8204 5966 8210 6000
rect 8130 5928 8210 5966
rect 8250 6006 8316 6012
rect 8250 5954 8256 6006
rect 8308 5954 8316 6006
rect 8250 5948 8316 5954
rect 8356 6000 8662 6012
rect 8356 5966 8362 6000
rect 8396 5998 8662 6000
rect 8396 5966 8458 5998
rect 8130 5894 8170 5928
rect 8204 5894 8210 5928
rect 8130 5882 8210 5894
rect 8260 5928 8306 5948
rect 8260 5894 8266 5928
rect 8300 5894 8306 5928
rect 8260 5882 8306 5894
rect 8356 5928 8458 5966
rect 8356 5894 8362 5928
rect 8396 5894 8458 5928
rect 8356 5882 8458 5894
rect 8578 5951 8812 5960
rect 8578 5899 8584 5951
rect 8636 5932 8760 5951
rect 8636 5899 8642 5932
rect 8578 5892 8642 5899
rect 8754 5899 8760 5932
rect 8812 5899 8818 5932
rect 8754 5892 8818 5899
rect 7710 5831 7986 5834
rect 7710 5797 7739 5831
rect 7773 5797 7831 5831
rect 7865 5797 7923 5831
rect 7957 5797 7986 5831
rect 7710 5766 7986 5797
rect 7816 5718 7880 5724
rect 7816 5666 7822 5718
rect 7874 5666 7880 5718
rect 7816 5660 7880 5666
rect 8130 5682 8176 5882
rect 8206 5844 8264 5854
rect 8206 5810 8218 5844
rect 8252 5810 8264 5844
rect 8206 5792 8264 5810
rect 8318 5763 8376 5780
rect 8318 5729 8330 5763
rect 8364 5729 8376 5763
rect 8318 5714 8376 5729
rect 8408 5682 8458 5882
rect 8524 5831 8800 5862
rect 8524 5797 8553 5831
rect 8587 5797 8645 5831
rect 8679 5797 8737 5831
rect 8771 5797 8800 5831
rect 8524 5766 8800 5797
rect 8130 5635 8226 5682
rect 7728 5602 7792 5608
rect 7728 5550 7734 5602
rect 7786 5550 7792 5602
rect 7728 5544 7792 5550
rect 7898 5592 7968 5610
rect 7898 5558 7919 5592
rect 7953 5558 7968 5592
rect 7898 5550 7968 5558
rect 8130 5601 8186 5635
rect 8220 5601 8226 5635
rect 8130 5563 8226 5601
rect 7898 5514 7926 5550
rect 8130 5529 8186 5563
rect 8220 5529 8226 5563
rect 8276 5635 8322 5682
rect 8276 5601 8282 5635
rect 8316 5601 8322 5635
rect 8276 5563 8322 5601
rect 8276 5542 8282 5563
rect 8130 5514 8226 5529
rect 7898 5482 8226 5514
rect 8266 5534 8282 5542
rect 8316 5542 8322 5563
rect 8372 5635 8458 5682
rect 8630 5716 8698 5726
rect 8630 5664 8638 5716
rect 8690 5664 8698 5716
rect 8630 5658 8698 5664
rect 8372 5601 8378 5635
rect 8412 5601 8458 5635
rect 8372 5563 8458 5601
rect 8316 5534 8332 5542
rect 8266 5482 8274 5534
rect 8326 5482 8332 5534
rect 8372 5529 8378 5563
rect 8412 5529 8458 5563
rect 8540 5604 8608 5610
rect 8540 5552 8546 5604
rect 8598 5552 8608 5604
rect 8540 5546 8608 5552
rect 8714 5590 8780 5602
rect 8714 5556 8731 5590
rect 8765 5556 8780 5590
rect 8714 5548 8780 5556
rect 8372 5510 8458 5529
rect 8752 5510 8780 5548
rect 8372 5482 8780 5510
rect 8266 5474 8332 5482
rect 8414 5478 8780 5482
rect 8218 5435 8280 5444
rect 8218 5401 8234 5435
rect 8268 5401 8280 5435
rect 8218 5384 8280 5401
rect 8222 5382 8280 5384
rect 8276 5327 8366 5348
rect 8276 5318 8303 5327
rect 6449 5293 8303 5318
rect 8337 5318 8366 5327
rect 8880 5318 8958 6276
rect 9046 6264 9670 6296
rect 9778 6331 9844 6342
rect 9778 6297 9794 6331
rect 9828 6297 9844 6331
rect 9778 6286 9844 6297
rect 9930 6294 9964 6440
rect 10112 6438 10170 6440
rect 10368 6459 10436 6464
rect 10368 6456 10396 6459
rect 10368 6404 10376 6456
rect 10430 6425 10436 6459
rect 10428 6404 10436 6425
rect 10166 6383 10256 6404
rect 10368 6398 10436 6404
rect 10166 6349 10193 6383
rect 10227 6349 10256 6383
rect 10390 6378 10436 6398
rect 10478 6531 10524 6578
rect 10478 6497 10484 6531
rect 10518 6497 10524 6531
rect 10478 6459 10524 6497
rect 10478 6425 10484 6459
rect 10518 6425 10524 6459
rect 10478 6404 10524 6425
rect 11632 6531 11678 6578
rect 11632 6497 11638 6531
rect 11672 6497 11678 6531
rect 11632 6459 11678 6497
rect 11632 6425 11638 6459
rect 11672 6425 11678 6459
rect 11720 6531 11766 6578
rect 11720 6497 11726 6531
rect 11760 6497 11766 6531
rect 11720 6459 11766 6497
rect 11820 6500 11880 6732
rect 11908 7022 11948 7056
rect 11982 7022 11988 7056
rect 11908 6984 11988 7022
rect 12028 7062 12094 7068
rect 12028 7010 12034 7062
rect 12086 7010 12094 7062
rect 12028 7004 12094 7010
rect 12134 7056 12236 7068
rect 12134 7022 12140 7056
rect 12174 7022 12236 7056
rect 11908 6950 11948 6984
rect 11982 6950 11988 6984
rect 11908 6938 11988 6950
rect 12038 6984 12084 7004
rect 12038 6950 12044 6984
rect 12078 6950 12084 6984
rect 12038 6938 12084 6950
rect 12134 6984 12236 7022
rect 12134 6950 12140 6984
rect 12174 6950 12236 6984
rect 12134 6938 12236 6950
rect 11908 6738 11954 6938
rect 11984 6900 12042 6910
rect 11984 6866 11996 6900
rect 12030 6866 12042 6900
rect 11984 6848 12042 6866
rect 12186 6858 12236 6938
rect 12602 6916 12686 7186
rect 12344 6906 12402 6912
rect 12336 6900 12410 6906
rect 12096 6819 12154 6836
rect 12096 6785 12108 6819
rect 12142 6785 12154 6819
rect 12096 6770 12154 6785
rect 12186 6792 12256 6858
rect 12336 6848 12347 6900
rect 12399 6848 12410 6900
rect 12336 6842 12410 6848
rect 12478 6890 12754 6916
rect 13348 6910 13446 7186
rect 12478 6885 12579 6890
rect 12631 6885 12754 6890
rect 12478 6851 12507 6885
rect 12541 6851 12579 6885
rect 12633 6851 12691 6885
rect 12725 6851 12754 6885
rect 12344 6834 12402 6842
rect 12478 6838 12579 6851
rect 12631 6838 12754 6851
rect 12478 6820 12754 6838
rect 12824 6879 13446 6910
rect 12824 6845 12853 6879
rect 12887 6845 12945 6879
rect 12979 6845 13037 6879
rect 13071 6877 13446 6879
rect 13071 6845 13199 6877
rect 12824 6843 13199 6845
rect 13233 6843 13291 6877
rect 13325 6843 13383 6877
rect 13417 6843 13446 6877
rect 13708 7140 14028 7158
rect 13708 7106 13980 7140
rect 14014 7106 14028 7140
rect 13708 7096 14028 7106
rect 12824 6812 13446 6843
rect 13586 6868 13662 6874
rect 13586 6816 13602 6868
rect 13654 6816 13662 6868
rect 13586 6810 13662 6816
rect 12186 6738 12236 6792
rect 13708 6766 13768 7096
rect 13830 7056 13876 7068
rect 11908 6691 12004 6738
rect 11908 6657 11964 6691
rect 11998 6657 12004 6691
rect 11908 6619 12004 6657
rect 11908 6585 11964 6619
rect 11998 6585 12004 6619
rect 12054 6691 12100 6738
rect 12054 6657 12060 6691
rect 12094 6657 12100 6691
rect 12054 6619 12100 6657
rect 12054 6598 12060 6619
rect 11908 6538 12004 6585
rect 12044 6590 12060 6598
rect 12094 6598 12100 6619
rect 12150 6691 12236 6738
rect 13240 6746 13768 6766
rect 13240 6712 13252 6746
rect 13286 6732 13768 6746
rect 13286 6712 13298 6732
rect 13240 6698 13298 6712
rect 12150 6657 12156 6691
rect 12190 6657 12236 6691
rect 12150 6619 12236 6657
rect 12094 6590 12110 6598
rect 12044 6538 12052 6590
rect 12104 6538 12110 6590
rect 12150 6585 12156 6619
rect 12190 6585 12236 6619
rect 12312 6659 12378 6672
rect 12312 6625 12328 6659
rect 12362 6625 12378 6659
rect 12706 6652 12774 6654
rect 12312 6614 12378 6625
rect 12622 6648 12774 6652
rect 12622 6642 12715 6648
rect 12622 6608 12642 6642
rect 12676 6608 12715 6642
rect 12622 6602 12715 6608
rect 12706 6596 12715 6602
rect 12767 6596 12774 6648
rect 12706 6590 12774 6596
rect 12810 6636 12884 6660
rect 12810 6602 12838 6636
rect 12872 6602 12884 6636
rect 12150 6542 12236 6585
rect 12810 6582 12884 6602
rect 13008 6652 13080 6664
rect 13008 6600 13019 6652
rect 13071 6600 13080 6652
rect 13554 6659 13620 6668
rect 13554 6625 13570 6659
rect 13604 6625 13620 6659
rect 13554 6612 13620 6625
rect 13008 6596 13080 6600
rect 12150 6538 12196 6542
rect 12044 6530 12110 6538
rect 12278 6531 12324 6578
rect 11820 6491 12058 6500
rect 11820 6468 12012 6491
rect 11720 6442 11726 6459
rect 10478 6376 10550 6404
rect 11632 6378 11678 6425
rect 11708 6436 11726 6442
rect 11760 6442 11766 6459
rect 11818 6457 12012 6468
rect 12046 6457 12058 6491
rect 12278 6497 12284 6531
rect 12318 6497 12324 6531
rect 12278 6464 12324 6497
rect 11760 6436 11774 6442
rect 11708 6384 11714 6436
rect 11766 6384 11774 6436
rect 11708 6378 11774 6384
rect 11818 6440 12058 6457
rect 10166 6328 10256 6349
rect 10424 6331 10490 6340
rect 10424 6297 10440 6331
rect 10474 6297 10490 6331
rect 10424 6294 10490 6297
rect 9930 6266 10490 6294
rect 9834 6210 9902 6224
rect 9834 6176 9852 6210
rect 9886 6176 9902 6210
rect 9834 6166 9902 6176
rect 9874 5862 9902 6166
rect 9930 6084 9964 6266
rect 10262 6200 10334 6212
rect 10262 6148 10272 6200
rect 10324 6148 10334 6200
rect 10262 6136 10334 6148
rect 10186 6084 10250 6102
rect 9930 6050 10202 6084
rect 10236 6050 10250 6084
rect 10186 6040 10250 6050
rect 10522 6026 10550 6376
rect 10590 6342 10866 6372
rect 10590 6341 10622 6342
rect 10674 6341 10866 6342
rect 10590 6307 10619 6341
rect 10674 6307 10711 6341
rect 10745 6307 10803 6341
rect 10837 6307 10866 6341
rect 10590 6290 10622 6307
rect 10674 6290 10866 6307
rect 10590 6276 10866 6290
rect 10934 6348 11558 6366
rect 10934 6335 11476 6348
rect 10934 6301 10965 6335
rect 10999 6301 11057 6335
rect 11091 6301 11149 6335
rect 11183 6333 11476 6335
rect 11528 6333 11558 6348
rect 11183 6301 11311 6333
rect 10934 6299 11311 6301
rect 11345 6299 11403 6333
rect 11437 6299 11476 6333
rect 11529 6299 11558 6333
rect 10934 6296 11476 6299
rect 11528 6296 11558 6299
rect 10640 6084 10706 6090
rect 10640 6032 10646 6084
rect 10698 6032 10706 6084
rect 10640 6026 10706 6032
rect 10296 6012 10550 6026
rect 10052 6000 10098 6012
rect 9598 5834 9902 5862
rect 10018 5966 10058 6000
rect 10092 5966 10098 6000
rect 10018 5928 10098 5966
rect 10138 6006 10204 6012
rect 10138 5954 10144 6006
rect 10196 5954 10204 6006
rect 10138 5948 10204 5954
rect 10244 6000 10550 6012
rect 10244 5966 10250 6000
rect 10284 5998 10550 6000
rect 10284 5966 10346 5998
rect 10018 5894 10058 5928
rect 10092 5894 10098 5928
rect 10018 5882 10098 5894
rect 10148 5928 10194 5948
rect 10148 5894 10154 5928
rect 10188 5894 10194 5928
rect 10148 5882 10194 5894
rect 10244 5928 10346 5966
rect 10244 5894 10250 5928
rect 10284 5894 10346 5928
rect 10244 5882 10346 5894
rect 10466 5951 10700 5960
rect 10466 5899 10472 5951
rect 10524 5932 10648 5951
rect 10524 5899 10530 5932
rect 10466 5892 10530 5899
rect 10642 5899 10648 5932
rect 10700 5899 10706 5932
rect 10642 5892 10706 5899
rect 9598 5831 9874 5834
rect 9598 5797 9627 5831
rect 9661 5797 9719 5831
rect 9753 5797 9811 5831
rect 9845 5797 9874 5831
rect 9598 5766 9874 5797
rect 9704 5718 9768 5724
rect 9704 5666 9710 5718
rect 9762 5666 9768 5718
rect 9704 5660 9768 5666
rect 10018 5682 10064 5882
rect 10094 5844 10152 5854
rect 10094 5810 10106 5844
rect 10140 5810 10152 5844
rect 10094 5792 10152 5810
rect 10206 5763 10264 5780
rect 10206 5729 10218 5763
rect 10252 5729 10264 5763
rect 10206 5714 10264 5729
rect 10296 5682 10346 5882
rect 10412 5831 10688 5862
rect 10412 5797 10441 5831
rect 10475 5797 10533 5831
rect 10567 5797 10625 5831
rect 10659 5797 10688 5831
rect 10412 5766 10688 5797
rect 10018 5635 10114 5682
rect 9616 5602 9680 5608
rect 9616 5550 9622 5602
rect 9674 5550 9680 5602
rect 9616 5544 9680 5550
rect 9786 5592 9856 5610
rect 9786 5558 9807 5592
rect 9841 5558 9856 5592
rect 9786 5550 9856 5558
rect 10018 5601 10074 5635
rect 10108 5601 10114 5635
rect 10018 5563 10114 5601
rect 9786 5514 9814 5550
rect 10018 5529 10074 5563
rect 10108 5529 10114 5563
rect 10164 5635 10210 5682
rect 10164 5601 10170 5635
rect 10204 5601 10210 5635
rect 10164 5563 10210 5601
rect 10164 5542 10170 5563
rect 10018 5514 10114 5529
rect 9786 5482 10114 5514
rect 10154 5534 10170 5542
rect 10204 5542 10210 5563
rect 10260 5635 10346 5682
rect 10518 5716 10586 5726
rect 10518 5664 10526 5716
rect 10578 5664 10586 5716
rect 10518 5658 10586 5664
rect 10260 5601 10266 5635
rect 10300 5601 10346 5635
rect 10260 5563 10346 5601
rect 10204 5534 10220 5542
rect 10154 5482 10162 5534
rect 10214 5482 10220 5534
rect 10260 5529 10266 5563
rect 10300 5529 10346 5563
rect 10428 5604 10496 5610
rect 10428 5552 10434 5604
rect 10486 5552 10496 5604
rect 10428 5546 10496 5552
rect 10602 5590 10668 5602
rect 10602 5556 10619 5590
rect 10653 5556 10668 5590
rect 10602 5548 10668 5556
rect 10260 5510 10346 5529
rect 10640 5510 10668 5548
rect 10260 5482 10668 5510
rect 10154 5474 10220 5482
rect 10302 5478 10668 5482
rect 10106 5435 10168 5444
rect 10106 5401 10122 5435
rect 10156 5401 10168 5435
rect 10106 5384 10168 5401
rect 10110 5382 10168 5384
rect 10164 5327 10254 5348
rect 10164 5318 10191 5327
rect 8337 5293 10191 5318
rect 10225 5318 10254 5327
rect 10768 5318 10846 6276
rect 10934 6264 11558 6296
rect 11666 6331 11732 6342
rect 11666 6297 11682 6331
rect 11716 6297 11732 6331
rect 11666 6286 11732 6297
rect 11818 6294 11852 6440
rect 12000 6438 12058 6440
rect 12256 6459 12324 6464
rect 12256 6456 12284 6459
rect 12256 6404 12264 6456
rect 12318 6425 12324 6459
rect 12316 6404 12324 6425
rect 12054 6383 12144 6404
rect 12256 6398 12324 6404
rect 12054 6349 12081 6383
rect 12115 6349 12144 6383
rect 12278 6378 12324 6398
rect 12366 6531 12412 6578
rect 12366 6497 12372 6531
rect 12406 6497 12412 6531
rect 12366 6459 12412 6497
rect 12366 6425 12372 6459
rect 12406 6425 12412 6459
rect 12366 6404 12412 6425
rect 13520 6531 13566 6578
rect 13520 6497 13526 6531
rect 13560 6497 13566 6531
rect 13520 6459 13566 6497
rect 13520 6425 13526 6459
rect 13560 6425 13566 6459
rect 13608 6531 13654 6578
rect 13608 6497 13614 6531
rect 13648 6497 13654 6531
rect 13608 6459 13654 6497
rect 13708 6500 13768 6732
rect 13796 7022 13836 7056
rect 13870 7022 13876 7056
rect 13796 6984 13876 7022
rect 13916 7062 13982 7068
rect 13916 7010 13922 7062
rect 13974 7010 13982 7062
rect 13916 7004 13982 7010
rect 14022 7056 14124 7068
rect 14022 7022 14028 7056
rect 14062 7022 14124 7056
rect 13796 6950 13836 6984
rect 13870 6950 13876 6984
rect 13796 6938 13876 6950
rect 13926 6984 13972 7004
rect 13926 6950 13932 6984
rect 13966 6950 13972 6984
rect 13926 6938 13972 6950
rect 14022 6984 14124 7022
rect 14022 6950 14028 6984
rect 14062 6950 14124 6984
rect 14022 6938 14124 6950
rect 13796 6738 13842 6938
rect 13872 6900 13930 6910
rect 13872 6866 13884 6900
rect 13918 6866 13930 6900
rect 13872 6848 13930 6866
rect 14074 6858 14124 6938
rect 14490 6916 14574 7186
rect 14232 6906 14290 6912
rect 14224 6900 14298 6906
rect 13984 6819 14042 6836
rect 13984 6785 13996 6819
rect 14030 6785 14042 6819
rect 13984 6770 14042 6785
rect 14074 6792 14144 6858
rect 14224 6848 14235 6900
rect 14287 6848 14298 6900
rect 14224 6842 14298 6848
rect 14366 6890 14642 6916
rect 15230 6910 15328 7186
rect 14366 6885 14467 6890
rect 14519 6885 14642 6890
rect 14366 6851 14395 6885
rect 14429 6851 14467 6885
rect 14521 6851 14579 6885
rect 14613 6851 14642 6885
rect 14232 6834 14290 6842
rect 14366 6838 14467 6851
rect 14519 6838 14642 6851
rect 14366 6820 14642 6838
rect 14706 6879 15328 6910
rect 14706 6845 14735 6879
rect 14769 6845 14827 6879
rect 14861 6845 14919 6879
rect 14953 6877 15328 6879
rect 14953 6845 15081 6877
rect 14706 6843 15081 6845
rect 15115 6843 15173 6877
rect 15207 6843 15265 6877
rect 15299 6843 15328 6877
rect 15590 7140 15910 7158
rect 15590 7106 15862 7140
rect 15896 7106 15910 7140
rect 15590 7096 15910 7106
rect 14706 6812 15328 6843
rect 15468 6868 15544 6874
rect 15468 6816 15484 6868
rect 15536 6816 15544 6868
rect 15468 6810 15544 6816
rect 14074 6738 14124 6792
rect 15590 6766 15650 7096
rect 15712 7056 15758 7068
rect 13796 6691 13892 6738
rect 13796 6657 13852 6691
rect 13886 6657 13892 6691
rect 13796 6619 13892 6657
rect 13796 6585 13852 6619
rect 13886 6585 13892 6619
rect 13942 6691 13988 6738
rect 13942 6657 13948 6691
rect 13982 6657 13988 6691
rect 13942 6619 13988 6657
rect 13942 6598 13948 6619
rect 13796 6538 13892 6585
rect 13932 6590 13948 6598
rect 13982 6598 13988 6619
rect 14038 6691 14124 6738
rect 15122 6746 15650 6766
rect 15122 6712 15134 6746
rect 15168 6732 15650 6746
rect 15168 6712 15180 6732
rect 15122 6698 15180 6712
rect 14038 6657 14044 6691
rect 14078 6657 14124 6691
rect 14038 6619 14124 6657
rect 13982 6590 13998 6598
rect 13932 6538 13940 6590
rect 13992 6538 13998 6590
rect 14038 6585 14044 6619
rect 14078 6585 14124 6619
rect 14200 6659 14266 6672
rect 14200 6625 14216 6659
rect 14250 6625 14266 6659
rect 14594 6652 14662 6654
rect 14200 6614 14266 6625
rect 14510 6648 14662 6652
rect 14510 6642 14603 6648
rect 14510 6608 14530 6642
rect 14564 6608 14603 6642
rect 14510 6602 14603 6608
rect 14594 6596 14603 6602
rect 14655 6596 14662 6648
rect 14594 6590 14662 6596
rect 14692 6636 14766 6660
rect 14692 6602 14720 6636
rect 14754 6602 14766 6636
rect 14038 6542 14124 6585
rect 14692 6582 14766 6602
rect 14890 6652 14962 6664
rect 14890 6600 14901 6652
rect 14953 6600 14962 6652
rect 15436 6659 15502 6668
rect 15436 6625 15452 6659
rect 15486 6625 15502 6659
rect 15436 6612 15502 6625
rect 14890 6596 14962 6600
rect 14038 6538 14084 6542
rect 13932 6530 13998 6538
rect 14166 6531 14212 6578
rect 13708 6491 13946 6500
rect 13708 6468 13900 6491
rect 13608 6442 13614 6459
rect 12366 6376 12438 6404
rect 13520 6378 13566 6425
rect 13596 6436 13614 6442
rect 13648 6442 13654 6459
rect 13706 6457 13900 6468
rect 13934 6457 13946 6491
rect 14166 6497 14172 6531
rect 14206 6497 14212 6531
rect 14166 6464 14212 6497
rect 13648 6436 13662 6442
rect 13596 6384 13602 6436
rect 13654 6384 13662 6436
rect 13596 6378 13662 6384
rect 13706 6440 13946 6457
rect 12054 6328 12144 6349
rect 12312 6331 12378 6340
rect 12312 6297 12328 6331
rect 12362 6297 12378 6331
rect 12312 6294 12378 6297
rect 11818 6266 12378 6294
rect 11722 6210 11790 6224
rect 11722 6176 11740 6210
rect 11774 6176 11790 6210
rect 11722 6166 11790 6176
rect 11762 5862 11790 6166
rect 11818 6084 11852 6266
rect 12150 6200 12222 6212
rect 12150 6148 12160 6200
rect 12212 6148 12222 6200
rect 12150 6136 12222 6148
rect 12074 6084 12138 6102
rect 11818 6050 12090 6084
rect 12124 6050 12138 6084
rect 12074 6040 12138 6050
rect 12410 6026 12438 6376
rect 12478 6342 12754 6372
rect 12478 6341 12510 6342
rect 12562 6341 12754 6342
rect 12478 6307 12507 6341
rect 12562 6307 12599 6341
rect 12633 6307 12691 6341
rect 12725 6307 12754 6341
rect 12478 6290 12510 6307
rect 12562 6290 12754 6307
rect 12478 6276 12754 6290
rect 12822 6348 13446 6366
rect 12822 6335 13364 6348
rect 12822 6301 12853 6335
rect 12887 6301 12945 6335
rect 12979 6301 13037 6335
rect 13071 6333 13364 6335
rect 13416 6333 13446 6348
rect 13071 6301 13199 6333
rect 12822 6299 13199 6301
rect 13233 6299 13291 6333
rect 13325 6299 13364 6333
rect 13417 6299 13446 6333
rect 12822 6296 13364 6299
rect 13416 6296 13446 6299
rect 12528 6084 12594 6090
rect 12528 6032 12534 6084
rect 12586 6032 12594 6084
rect 12528 6026 12594 6032
rect 12184 6012 12438 6026
rect 11940 6000 11986 6012
rect 11486 5834 11790 5862
rect 11906 5966 11946 6000
rect 11980 5966 11986 6000
rect 11906 5928 11986 5966
rect 12026 6006 12092 6012
rect 12026 5954 12032 6006
rect 12084 5954 12092 6006
rect 12026 5948 12092 5954
rect 12132 6000 12438 6012
rect 12132 5966 12138 6000
rect 12172 5998 12438 6000
rect 12172 5966 12234 5998
rect 11906 5894 11946 5928
rect 11980 5894 11986 5928
rect 11906 5882 11986 5894
rect 12036 5928 12082 5948
rect 12036 5894 12042 5928
rect 12076 5894 12082 5928
rect 12036 5882 12082 5894
rect 12132 5928 12234 5966
rect 12132 5894 12138 5928
rect 12172 5894 12234 5928
rect 12132 5882 12234 5894
rect 12354 5951 12588 5960
rect 12354 5899 12360 5951
rect 12412 5932 12536 5951
rect 12412 5899 12418 5932
rect 12354 5892 12418 5899
rect 12530 5899 12536 5932
rect 12588 5899 12594 5932
rect 12530 5892 12594 5899
rect 11486 5831 11762 5834
rect 11486 5797 11515 5831
rect 11549 5797 11607 5831
rect 11641 5797 11699 5831
rect 11733 5797 11762 5831
rect 11486 5766 11762 5797
rect 11592 5718 11656 5724
rect 11592 5666 11598 5718
rect 11650 5666 11656 5718
rect 11592 5660 11656 5666
rect 11906 5682 11952 5882
rect 11982 5844 12040 5854
rect 11982 5810 11994 5844
rect 12028 5810 12040 5844
rect 11982 5792 12040 5810
rect 12094 5763 12152 5780
rect 12094 5729 12106 5763
rect 12140 5729 12152 5763
rect 12094 5714 12152 5729
rect 12184 5682 12234 5882
rect 12300 5831 12576 5862
rect 12300 5797 12329 5831
rect 12363 5797 12421 5831
rect 12455 5797 12513 5831
rect 12547 5797 12576 5831
rect 12300 5766 12576 5797
rect 11906 5635 12002 5682
rect 11504 5602 11568 5608
rect 11504 5550 11510 5602
rect 11562 5550 11568 5602
rect 11504 5544 11568 5550
rect 11674 5592 11744 5610
rect 11674 5558 11695 5592
rect 11729 5558 11744 5592
rect 11674 5550 11744 5558
rect 11906 5601 11962 5635
rect 11996 5601 12002 5635
rect 11906 5563 12002 5601
rect 11674 5514 11702 5550
rect 11906 5529 11962 5563
rect 11996 5529 12002 5563
rect 12052 5635 12098 5682
rect 12052 5601 12058 5635
rect 12092 5601 12098 5635
rect 12052 5563 12098 5601
rect 12052 5542 12058 5563
rect 11906 5514 12002 5529
rect 11674 5482 12002 5514
rect 12042 5534 12058 5542
rect 12092 5542 12098 5563
rect 12148 5635 12234 5682
rect 12406 5716 12474 5726
rect 12406 5664 12414 5716
rect 12466 5664 12474 5716
rect 12406 5658 12474 5664
rect 12148 5601 12154 5635
rect 12188 5601 12234 5635
rect 12148 5563 12234 5601
rect 12092 5534 12108 5542
rect 12042 5482 12050 5534
rect 12102 5482 12108 5534
rect 12148 5529 12154 5563
rect 12188 5529 12234 5563
rect 12316 5604 12384 5610
rect 12316 5552 12322 5604
rect 12374 5552 12384 5604
rect 12316 5546 12384 5552
rect 12490 5590 12556 5602
rect 12490 5556 12507 5590
rect 12541 5556 12556 5590
rect 12490 5548 12556 5556
rect 12148 5510 12234 5529
rect 12528 5510 12556 5548
rect 12148 5482 12556 5510
rect 12042 5474 12108 5482
rect 12190 5478 12556 5482
rect 11994 5435 12056 5444
rect 11994 5401 12010 5435
rect 12044 5401 12056 5435
rect 11994 5384 12056 5401
rect 11998 5382 12056 5384
rect 12052 5327 12142 5348
rect 12052 5318 12079 5327
rect 10225 5293 12079 5318
rect 12113 5318 12142 5327
rect 12656 5318 12734 6276
rect 12822 6264 13446 6296
rect 13554 6331 13620 6342
rect 13554 6297 13570 6331
rect 13604 6297 13620 6331
rect 13554 6286 13620 6297
rect 13706 6294 13740 6440
rect 13888 6438 13946 6440
rect 14144 6459 14212 6464
rect 14144 6456 14172 6459
rect 14144 6404 14152 6456
rect 14206 6425 14212 6459
rect 14204 6404 14212 6425
rect 13942 6383 14032 6404
rect 14144 6398 14212 6404
rect 13942 6349 13969 6383
rect 14003 6349 14032 6383
rect 14166 6378 14212 6398
rect 14254 6531 14300 6578
rect 14254 6497 14260 6531
rect 14294 6497 14300 6531
rect 14254 6459 14300 6497
rect 14254 6425 14260 6459
rect 14294 6425 14300 6459
rect 14254 6404 14300 6425
rect 15402 6531 15448 6578
rect 15402 6497 15408 6531
rect 15442 6497 15448 6531
rect 15402 6459 15448 6497
rect 15402 6425 15408 6459
rect 15442 6425 15448 6459
rect 15490 6531 15536 6578
rect 15490 6497 15496 6531
rect 15530 6497 15536 6531
rect 15490 6459 15536 6497
rect 15590 6500 15650 6732
rect 15678 7022 15718 7056
rect 15752 7022 15758 7056
rect 15678 6984 15758 7022
rect 15798 7062 15864 7068
rect 15798 7010 15804 7062
rect 15856 7010 15864 7062
rect 15798 7004 15864 7010
rect 15904 7056 16006 7068
rect 15904 7022 15910 7056
rect 15944 7022 16006 7056
rect 15678 6950 15718 6984
rect 15752 6950 15758 6984
rect 15678 6938 15758 6950
rect 15808 6984 15854 7004
rect 15808 6950 15814 6984
rect 15848 6950 15854 6984
rect 15808 6938 15854 6950
rect 15904 6984 16006 7022
rect 15904 6950 15910 6984
rect 15944 6950 16006 6984
rect 15904 6938 16006 6950
rect 15678 6738 15724 6938
rect 15754 6900 15812 6910
rect 15754 6866 15766 6900
rect 15800 6866 15812 6900
rect 15754 6848 15812 6866
rect 15956 6858 16006 6938
rect 16372 6916 16456 7186
rect 16114 6906 16172 6912
rect 16106 6900 16180 6906
rect 15866 6819 15924 6836
rect 15866 6785 15878 6819
rect 15912 6785 15924 6819
rect 15866 6770 15924 6785
rect 15956 6792 16026 6858
rect 16106 6848 16117 6900
rect 16169 6848 16180 6900
rect 16106 6842 16180 6848
rect 16248 6890 16524 6916
rect 17118 6910 17216 7186
rect 16248 6885 16349 6890
rect 16401 6885 16524 6890
rect 16248 6851 16277 6885
rect 16311 6851 16349 6885
rect 16403 6851 16461 6885
rect 16495 6851 16524 6885
rect 16114 6834 16172 6842
rect 16248 6838 16349 6851
rect 16401 6838 16524 6851
rect 16248 6820 16524 6838
rect 16594 6879 17216 6910
rect 16594 6845 16623 6879
rect 16657 6845 16715 6879
rect 16749 6845 16807 6879
rect 16841 6877 17216 6879
rect 16841 6845 16969 6877
rect 16594 6843 16969 6845
rect 17003 6843 17061 6877
rect 17095 6843 17153 6877
rect 17187 6843 17216 6877
rect 17478 7140 17798 7158
rect 17478 7106 17750 7140
rect 17784 7106 17798 7140
rect 17478 7096 17798 7106
rect 16594 6812 17216 6843
rect 17356 6868 17432 6874
rect 17356 6816 17372 6868
rect 17424 6816 17432 6868
rect 17356 6810 17432 6816
rect 15956 6738 16006 6792
rect 17478 6766 17538 7096
rect 17600 7056 17646 7068
rect 15678 6691 15774 6738
rect 15678 6657 15734 6691
rect 15768 6657 15774 6691
rect 15678 6619 15774 6657
rect 15678 6585 15734 6619
rect 15768 6585 15774 6619
rect 15824 6691 15870 6738
rect 15824 6657 15830 6691
rect 15864 6657 15870 6691
rect 15824 6619 15870 6657
rect 15824 6598 15830 6619
rect 15678 6538 15774 6585
rect 15814 6590 15830 6598
rect 15864 6598 15870 6619
rect 15920 6691 16006 6738
rect 17010 6746 17538 6766
rect 17010 6712 17022 6746
rect 17056 6732 17538 6746
rect 17056 6712 17068 6732
rect 17010 6698 17068 6712
rect 15920 6657 15926 6691
rect 15960 6657 16006 6691
rect 15920 6619 16006 6657
rect 15864 6590 15880 6598
rect 15814 6538 15822 6590
rect 15874 6538 15880 6590
rect 15920 6585 15926 6619
rect 15960 6585 16006 6619
rect 16082 6659 16148 6672
rect 16082 6625 16098 6659
rect 16132 6625 16148 6659
rect 16476 6652 16544 6654
rect 16082 6614 16148 6625
rect 16392 6648 16544 6652
rect 16392 6642 16485 6648
rect 16392 6608 16412 6642
rect 16446 6608 16485 6642
rect 16392 6602 16485 6608
rect 16476 6596 16485 6602
rect 16537 6596 16544 6648
rect 16476 6590 16544 6596
rect 16580 6636 16654 6660
rect 16580 6602 16608 6636
rect 16642 6602 16654 6636
rect 15920 6542 16006 6585
rect 16580 6582 16654 6602
rect 16778 6652 16850 6664
rect 16778 6600 16789 6652
rect 16841 6600 16850 6652
rect 17324 6659 17390 6668
rect 17324 6625 17340 6659
rect 17374 6625 17390 6659
rect 17324 6612 17390 6625
rect 16778 6596 16850 6600
rect 15920 6538 15966 6542
rect 15814 6530 15880 6538
rect 16048 6531 16094 6578
rect 15590 6491 15828 6500
rect 15590 6468 15782 6491
rect 15490 6442 15496 6459
rect 14254 6376 14326 6404
rect 15402 6378 15448 6425
rect 15478 6436 15496 6442
rect 15530 6442 15536 6459
rect 15588 6457 15782 6468
rect 15816 6457 15828 6491
rect 16048 6497 16054 6531
rect 16088 6497 16094 6531
rect 16048 6464 16094 6497
rect 15530 6436 15544 6442
rect 15478 6384 15484 6436
rect 15536 6384 15544 6436
rect 15478 6378 15544 6384
rect 15588 6440 15828 6457
rect 13942 6328 14032 6349
rect 14200 6331 14266 6340
rect 14200 6297 14216 6331
rect 14250 6297 14266 6331
rect 14200 6294 14266 6297
rect 13706 6266 14266 6294
rect 13610 6210 13678 6224
rect 13610 6176 13628 6210
rect 13662 6176 13678 6210
rect 13610 6166 13678 6176
rect 13650 5862 13678 6166
rect 13706 6084 13740 6266
rect 14038 6200 14110 6212
rect 14038 6148 14048 6200
rect 14100 6148 14110 6200
rect 14038 6136 14110 6148
rect 13962 6084 14026 6102
rect 13706 6050 13978 6084
rect 14012 6050 14026 6084
rect 13962 6040 14026 6050
rect 14298 6026 14326 6376
rect 14366 6342 14642 6372
rect 14366 6341 14398 6342
rect 14450 6341 14642 6342
rect 14366 6307 14395 6341
rect 14450 6307 14487 6341
rect 14521 6307 14579 6341
rect 14613 6307 14642 6341
rect 14366 6290 14398 6307
rect 14450 6290 14642 6307
rect 14366 6276 14642 6290
rect 14704 6348 15328 6366
rect 14704 6335 15246 6348
rect 14704 6301 14735 6335
rect 14769 6301 14827 6335
rect 14861 6301 14919 6335
rect 14953 6333 15246 6335
rect 15298 6333 15328 6348
rect 14953 6301 15081 6333
rect 14704 6299 15081 6301
rect 15115 6299 15173 6333
rect 15207 6299 15246 6333
rect 15299 6299 15328 6333
rect 14704 6296 15246 6299
rect 15298 6296 15328 6299
rect 14416 6084 14482 6090
rect 14416 6032 14422 6084
rect 14474 6032 14482 6084
rect 14416 6026 14482 6032
rect 14072 6012 14326 6026
rect 13828 6000 13874 6012
rect 13374 5834 13678 5862
rect 13794 5966 13834 6000
rect 13868 5966 13874 6000
rect 13794 5928 13874 5966
rect 13914 6006 13980 6012
rect 13914 5954 13920 6006
rect 13972 5954 13980 6006
rect 13914 5948 13980 5954
rect 14020 6000 14326 6012
rect 14020 5966 14026 6000
rect 14060 5998 14326 6000
rect 14060 5966 14122 5998
rect 13794 5894 13834 5928
rect 13868 5894 13874 5928
rect 13794 5882 13874 5894
rect 13924 5928 13970 5948
rect 13924 5894 13930 5928
rect 13964 5894 13970 5928
rect 13924 5882 13970 5894
rect 14020 5928 14122 5966
rect 14020 5894 14026 5928
rect 14060 5894 14122 5928
rect 14020 5882 14122 5894
rect 14242 5951 14476 5960
rect 14242 5899 14248 5951
rect 14300 5932 14424 5951
rect 14300 5899 14306 5932
rect 14242 5892 14306 5899
rect 14418 5899 14424 5932
rect 14476 5899 14482 5932
rect 14418 5892 14482 5899
rect 13374 5831 13650 5834
rect 13374 5797 13403 5831
rect 13437 5797 13495 5831
rect 13529 5797 13587 5831
rect 13621 5797 13650 5831
rect 13374 5766 13650 5797
rect 13480 5718 13544 5724
rect 13480 5666 13486 5718
rect 13538 5666 13544 5718
rect 13480 5660 13544 5666
rect 13794 5682 13840 5882
rect 13870 5844 13928 5854
rect 13870 5810 13882 5844
rect 13916 5810 13928 5844
rect 13870 5792 13928 5810
rect 13982 5763 14040 5780
rect 13982 5729 13994 5763
rect 14028 5729 14040 5763
rect 13982 5714 14040 5729
rect 14072 5682 14122 5882
rect 14188 5831 14464 5862
rect 14188 5797 14217 5831
rect 14251 5797 14309 5831
rect 14343 5797 14401 5831
rect 14435 5797 14464 5831
rect 14188 5766 14464 5797
rect 13794 5635 13890 5682
rect 13392 5602 13456 5608
rect 13392 5550 13398 5602
rect 13450 5550 13456 5602
rect 13392 5544 13456 5550
rect 13562 5592 13632 5610
rect 13562 5558 13583 5592
rect 13617 5558 13632 5592
rect 13562 5550 13632 5558
rect 13794 5601 13850 5635
rect 13884 5601 13890 5635
rect 13794 5563 13890 5601
rect 13562 5514 13590 5550
rect 13794 5529 13850 5563
rect 13884 5529 13890 5563
rect 13940 5635 13986 5682
rect 13940 5601 13946 5635
rect 13980 5601 13986 5635
rect 13940 5563 13986 5601
rect 13940 5542 13946 5563
rect 13794 5514 13890 5529
rect 13562 5482 13890 5514
rect 13930 5534 13946 5542
rect 13980 5542 13986 5563
rect 14036 5635 14122 5682
rect 14294 5716 14362 5726
rect 14294 5664 14302 5716
rect 14354 5664 14362 5716
rect 14294 5658 14362 5664
rect 14036 5601 14042 5635
rect 14076 5601 14122 5635
rect 14036 5563 14122 5601
rect 13980 5534 13996 5542
rect 13930 5482 13938 5534
rect 13990 5482 13996 5534
rect 14036 5529 14042 5563
rect 14076 5529 14122 5563
rect 14204 5604 14272 5610
rect 14204 5552 14210 5604
rect 14262 5552 14272 5604
rect 14204 5546 14272 5552
rect 14378 5590 14444 5602
rect 14378 5556 14395 5590
rect 14429 5556 14444 5590
rect 14378 5548 14444 5556
rect 14036 5510 14122 5529
rect 14416 5510 14444 5548
rect 14036 5482 14444 5510
rect 13930 5474 13996 5482
rect 14078 5478 14444 5482
rect 13882 5435 13944 5444
rect 13882 5401 13898 5435
rect 13932 5401 13944 5435
rect 13882 5384 13944 5401
rect 13886 5382 13944 5384
rect 13940 5327 14030 5348
rect 13940 5318 13967 5327
rect 12113 5293 13967 5318
rect 14001 5318 14030 5327
rect 14544 5318 14622 6276
rect 14704 6264 15328 6296
rect 15436 6331 15502 6342
rect 15436 6297 15452 6331
rect 15486 6297 15502 6331
rect 15436 6286 15502 6297
rect 15588 6294 15622 6440
rect 15770 6438 15828 6440
rect 16026 6459 16094 6464
rect 16026 6456 16054 6459
rect 16026 6404 16034 6456
rect 16088 6425 16094 6459
rect 16086 6404 16094 6425
rect 15824 6383 15914 6404
rect 16026 6398 16094 6404
rect 15824 6349 15851 6383
rect 15885 6349 15914 6383
rect 16048 6378 16094 6398
rect 16136 6531 16182 6578
rect 16136 6497 16142 6531
rect 16176 6497 16182 6531
rect 16136 6459 16182 6497
rect 16136 6425 16142 6459
rect 16176 6425 16182 6459
rect 16136 6404 16182 6425
rect 17290 6531 17336 6578
rect 17290 6497 17296 6531
rect 17330 6497 17336 6531
rect 17290 6459 17336 6497
rect 17290 6425 17296 6459
rect 17330 6425 17336 6459
rect 17378 6531 17424 6578
rect 17378 6497 17384 6531
rect 17418 6497 17424 6531
rect 17378 6459 17424 6497
rect 17478 6500 17538 6732
rect 17566 7022 17606 7056
rect 17640 7022 17646 7056
rect 17566 6984 17646 7022
rect 17686 7062 17752 7068
rect 17686 7010 17692 7062
rect 17744 7010 17752 7062
rect 17686 7004 17752 7010
rect 17792 7056 17894 7068
rect 17792 7022 17798 7056
rect 17832 7022 17894 7056
rect 17566 6950 17606 6984
rect 17640 6950 17646 6984
rect 17566 6938 17646 6950
rect 17696 6984 17742 7004
rect 17696 6950 17702 6984
rect 17736 6950 17742 6984
rect 17696 6938 17742 6950
rect 17792 6984 17894 7022
rect 17792 6950 17798 6984
rect 17832 6950 17894 6984
rect 17792 6938 17894 6950
rect 17566 6738 17612 6938
rect 17642 6900 17700 6910
rect 17642 6866 17654 6900
rect 17688 6866 17700 6900
rect 17642 6848 17700 6866
rect 17844 6858 17894 6938
rect 18260 6916 18344 7186
rect 18002 6906 18060 6912
rect 17994 6900 18068 6906
rect 17754 6819 17812 6836
rect 17754 6785 17766 6819
rect 17800 6785 17812 6819
rect 17754 6770 17812 6785
rect 17844 6792 17914 6858
rect 17994 6848 18005 6900
rect 18057 6848 18068 6900
rect 17994 6842 18068 6848
rect 18136 6890 18412 6916
rect 19006 6910 19104 7186
rect 18136 6885 18237 6890
rect 18289 6885 18412 6890
rect 18136 6851 18165 6885
rect 18199 6851 18237 6885
rect 18291 6851 18349 6885
rect 18383 6851 18412 6885
rect 18002 6834 18060 6842
rect 18136 6838 18237 6851
rect 18289 6838 18412 6851
rect 18136 6820 18412 6838
rect 18482 6879 19104 6910
rect 18482 6845 18511 6879
rect 18545 6845 18603 6879
rect 18637 6845 18695 6879
rect 18729 6877 19104 6879
rect 18729 6845 18857 6877
rect 18482 6843 18857 6845
rect 18891 6843 18949 6877
rect 18983 6843 19041 6877
rect 19075 6843 19104 6877
rect 19366 7140 19686 7158
rect 19366 7106 19638 7140
rect 19672 7106 19686 7140
rect 19366 7096 19686 7106
rect 18482 6812 19104 6843
rect 19244 6868 19320 6874
rect 19244 6816 19260 6868
rect 19312 6816 19320 6868
rect 19244 6810 19320 6816
rect 17844 6738 17894 6792
rect 19366 6766 19426 7096
rect 19488 7056 19534 7068
rect 17566 6691 17662 6738
rect 17566 6657 17622 6691
rect 17656 6657 17662 6691
rect 17566 6619 17662 6657
rect 17566 6585 17622 6619
rect 17656 6585 17662 6619
rect 17712 6691 17758 6738
rect 17712 6657 17718 6691
rect 17752 6657 17758 6691
rect 17712 6619 17758 6657
rect 17712 6598 17718 6619
rect 17566 6538 17662 6585
rect 17702 6590 17718 6598
rect 17752 6598 17758 6619
rect 17808 6691 17894 6738
rect 18898 6746 19426 6766
rect 18898 6712 18910 6746
rect 18944 6732 19426 6746
rect 18944 6712 18956 6732
rect 18898 6698 18956 6712
rect 17808 6657 17814 6691
rect 17848 6657 17894 6691
rect 17808 6619 17894 6657
rect 17752 6590 17768 6598
rect 17702 6538 17710 6590
rect 17762 6538 17768 6590
rect 17808 6585 17814 6619
rect 17848 6585 17894 6619
rect 17970 6659 18036 6672
rect 17970 6625 17986 6659
rect 18020 6625 18036 6659
rect 18364 6652 18432 6654
rect 17970 6614 18036 6625
rect 18280 6648 18432 6652
rect 18280 6642 18373 6648
rect 18280 6608 18300 6642
rect 18334 6608 18373 6642
rect 18280 6602 18373 6608
rect 18364 6596 18373 6602
rect 18425 6596 18432 6648
rect 18364 6590 18432 6596
rect 18468 6636 18542 6660
rect 18468 6602 18496 6636
rect 18530 6602 18542 6636
rect 17808 6542 17894 6585
rect 18468 6582 18542 6602
rect 18666 6652 18738 6664
rect 18666 6600 18677 6652
rect 18729 6600 18738 6652
rect 19212 6659 19278 6668
rect 19212 6625 19228 6659
rect 19262 6625 19278 6659
rect 19212 6612 19278 6625
rect 18666 6596 18738 6600
rect 17808 6538 17854 6542
rect 17702 6530 17768 6538
rect 17936 6531 17982 6578
rect 17478 6491 17716 6500
rect 17478 6468 17670 6491
rect 17378 6442 17384 6459
rect 16136 6376 16208 6404
rect 17290 6378 17336 6425
rect 17366 6436 17384 6442
rect 17418 6442 17424 6459
rect 17476 6457 17670 6468
rect 17704 6457 17716 6491
rect 17936 6497 17942 6531
rect 17976 6497 17982 6531
rect 17936 6464 17982 6497
rect 17418 6436 17432 6442
rect 17366 6384 17372 6436
rect 17424 6384 17432 6436
rect 17366 6378 17432 6384
rect 17476 6440 17716 6457
rect 15824 6328 15914 6349
rect 16082 6331 16148 6340
rect 16082 6297 16098 6331
rect 16132 6297 16148 6331
rect 16082 6294 16148 6297
rect 15588 6266 16148 6294
rect 15492 6210 15560 6224
rect 15492 6176 15510 6210
rect 15544 6176 15560 6210
rect 15492 6166 15560 6176
rect 15532 5862 15560 6166
rect 15588 6084 15622 6266
rect 15920 6200 15992 6212
rect 15920 6148 15930 6200
rect 15982 6148 15992 6200
rect 15920 6136 15992 6148
rect 15844 6084 15908 6102
rect 15588 6050 15860 6084
rect 15894 6050 15908 6084
rect 15844 6040 15908 6050
rect 16180 6026 16208 6376
rect 16248 6342 16524 6372
rect 16248 6341 16280 6342
rect 16332 6341 16524 6342
rect 16248 6307 16277 6341
rect 16332 6307 16369 6341
rect 16403 6307 16461 6341
rect 16495 6307 16524 6341
rect 16248 6290 16280 6307
rect 16332 6290 16524 6307
rect 16248 6276 16524 6290
rect 16592 6348 17216 6366
rect 16592 6335 17134 6348
rect 16592 6301 16623 6335
rect 16657 6301 16715 6335
rect 16749 6301 16807 6335
rect 16841 6333 17134 6335
rect 17186 6333 17216 6348
rect 16841 6301 16969 6333
rect 16592 6299 16969 6301
rect 17003 6299 17061 6333
rect 17095 6299 17134 6333
rect 17187 6299 17216 6333
rect 16592 6296 17134 6299
rect 17186 6296 17216 6299
rect 16298 6084 16364 6090
rect 16298 6032 16304 6084
rect 16356 6032 16364 6084
rect 16298 6026 16364 6032
rect 15954 6012 16208 6026
rect 15710 6000 15756 6012
rect 15256 5834 15560 5862
rect 15676 5966 15716 6000
rect 15750 5966 15756 6000
rect 15676 5928 15756 5966
rect 15796 6006 15862 6012
rect 15796 5954 15802 6006
rect 15854 5954 15862 6006
rect 15796 5948 15862 5954
rect 15902 6000 16208 6012
rect 15902 5966 15908 6000
rect 15942 5998 16208 6000
rect 15942 5966 16004 5998
rect 15676 5894 15716 5928
rect 15750 5894 15756 5928
rect 15676 5882 15756 5894
rect 15806 5928 15852 5948
rect 15806 5894 15812 5928
rect 15846 5894 15852 5928
rect 15806 5882 15852 5894
rect 15902 5928 16004 5966
rect 15902 5894 15908 5928
rect 15942 5894 16004 5928
rect 15902 5882 16004 5894
rect 16124 5951 16358 5960
rect 16124 5899 16130 5951
rect 16182 5932 16306 5951
rect 16182 5899 16188 5932
rect 16124 5892 16188 5899
rect 16300 5899 16306 5932
rect 16358 5899 16364 5932
rect 16300 5892 16364 5899
rect 15256 5831 15532 5834
rect 15256 5797 15285 5831
rect 15319 5797 15377 5831
rect 15411 5797 15469 5831
rect 15503 5797 15532 5831
rect 15256 5766 15532 5797
rect 15362 5718 15426 5724
rect 15362 5666 15368 5718
rect 15420 5666 15426 5718
rect 15362 5660 15426 5666
rect 15676 5682 15722 5882
rect 15752 5844 15810 5854
rect 15752 5810 15764 5844
rect 15798 5810 15810 5844
rect 15752 5792 15810 5810
rect 15864 5763 15922 5780
rect 15864 5729 15876 5763
rect 15910 5729 15922 5763
rect 15864 5714 15922 5729
rect 15954 5682 16004 5882
rect 16070 5831 16346 5862
rect 16070 5797 16099 5831
rect 16133 5797 16191 5831
rect 16225 5797 16283 5831
rect 16317 5797 16346 5831
rect 16070 5766 16346 5797
rect 15676 5635 15772 5682
rect 15274 5602 15338 5608
rect 15274 5550 15280 5602
rect 15332 5550 15338 5602
rect 15274 5544 15338 5550
rect 15444 5592 15514 5610
rect 15444 5558 15465 5592
rect 15499 5558 15514 5592
rect 15444 5550 15514 5558
rect 15676 5601 15732 5635
rect 15766 5601 15772 5635
rect 15676 5563 15772 5601
rect 15444 5514 15472 5550
rect 15676 5529 15732 5563
rect 15766 5529 15772 5563
rect 15822 5635 15868 5682
rect 15822 5601 15828 5635
rect 15862 5601 15868 5635
rect 15822 5563 15868 5601
rect 15822 5542 15828 5563
rect 15676 5514 15772 5529
rect 15444 5482 15772 5514
rect 15812 5534 15828 5542
rect 15862 5542 15868 5563
rect 15918 5635 16004 5682
rect 16176 5716 16244 5726
rect 16176 5664 16184 5716
rect 16236 5664 16244 5716
rect 16176 5658 16244 5664
rect 15918 5601 15924 5635
rect 15958 5601 16004 5635
rect 15918 5563 16004 5601
rect 15862 5534 15878 5542
rect 15812 5482 15820 5534
rect 15872 5482 15878 5534
rect 15918 5529 15924 5563
rect 15958 5529 16004 5563
rect 16086 5604 16154 5610
rect 16086 5552 16092 5604
rect 16144 5552 16154 5604
rect 16086 5546 16154 5552
rect 16260 5590 16326 5602
rect 16260 5556 16277 5590
rect 16311 5556 16326 5590
rect 16260 5548 16326 5556
rect 15918 5510 16004 5529
rect 16298 5510 16326 5548
rect 15918 5482 16326 5510
rect 15812 5474 15878 5482
rect 15960 5478 16326 5482
rect 15764 5435 15826 5444
rect 15764 5401 15780 5435
rect 15814 5401 15826 5435
rect 15764 5384 15826 5401
rect 15768 5382 15826 5384
rect 15822 5327 15912 5348
rect 15822 5318 15849 5327
rect 14001 5293 15849 5318
rect 15883 5318 15912 5327
rect 16426 5318 16504 6276
rect 16592 6264 17216 6296
rect 17324 6331 17390 6342
rect 17324 6297 17340 6331
rect 17374 6297 17390 6331
rect 17324 6286 17390 6297
rect 17476 6294 17510 6440
rect 17658 6438 17716 6440
rect 17914 6459 17982 6464
rect 17914 6456 17942 6459
rect 17914 6404 17922 6456
rect 17976 6425 17982 6459
rect 17974 6404 17982 6425
rect 17712 6383 17802 6404
rect 17914 6398 17982 6404
rect 17712 6349 17739 6383
rect 17773 6349 17802 6383
rect 17936 6378 17982 6398
rect 18024 6531 18070 6578
rect 18024 6497 18030 6531
rect 18064 6497 18070 6531
rect 18024 6459 18070 6497
rect 18024 6425 18030 6459
rect 18064 6425 18070 6459
rect 18024 6404 18070 6425
rect 19178 6531 19224 6578
rect 19178 6497 19184 6531
rect 19218 6497 19224 6531
rect 19178 6459 19224 6497
rect 19178 6425 19184 6459
rect 19218 6425 19224 6459
rect 19266 6531 19312 6578
rect 19266 6497 19272 6531
rect 19306 6497 19312 6531
rect 19266 6459 19312 6497
rect 19366 6500 19426 6732
rect 19454 7022 19494 7056
rect 19528 7022 19534 7056
rect 19454 6984 19534 7022
rect 19574 7062 19640 7068
rect 19574 7010 19580 7062
rect 19632 7010 19640 7062
rect 19574 7004 19640 7010
rect 19680 7056 19782 7068
rect 19680 7022 19686 7056
rect 19720 7022 19782 7056
rect 19454 6950 19494 6984
rect 19528 6950 19534 6984
rect 19454 6938 19534 6950
rect 19584 6984 19630 7004
rect 19584 6950 19590 6984
rect 19624 6950 19630 6984
rect 19584 6938 19630 6950
rect 19680 6984 19782 7022
rect 19680 6950 19686 6984
rect 19720 6950 19782 6984
rect 19680 6938 19782 6950
rect 19454 6738 19500 6938
rect 19530 6900 19588 6910
rect 19530 6866 19542 6900
rect 19576 6866 19588 6900
rect 19530 6848 19588 6866
rect 19732 6858 19782 6938
rect 20148 6916 20232 7186
rect 19890 6906 19948 6912
rect 19882 6900 19956 6906
rect 19642 6819 19700 6836
rect 19642 6785 19654 6819
rect 19688 6785 19700 6819
rect 19642 6770 19700 6785
rect 19732 6792 19802 6858
rect 19882 6848 19893 6900
rect 19945 6848 19956 6900
rect 19882 6842 19956 6848
rect 20024 6890 20300 6916
rect 20894 6910 20992 7186
rect 20024 6885 20125 6890
rect 20177 6885 20300 6890
rect 20024 6851 20053 6885
rect 20087 6851 20125 6885
rect 20179 6851 20237 6885
rect 20271 6851 20300 6885
rect 19890 6834 19948 6842
rect 20024 6838 20125 6851
rect 20177 6838 20300 6851
rect 20024 6820 20300 6838
rect 20370 6879 20992 6910
rect 20370 6845 20399 6879
rect 20433 6845 20491 6879
rect 20525 6845 20583 6879
rect 20617 6877 20992 6879
rect 20617 6845 20745 6877
rect 20370 6843 20745 6845
rect 20779 6843 20837 6877
rect 20871 6843 20929 6877
rect 20963 6843 20992 6877
rect 21254 7140 21574 7158
rect 21254 7106 21526 7140
rect 21560 7106 21574 7140
rect 21254 7096 21574 7106
rect 20370 6812 20992 6843
rect 21132 6868 21208 6874
rect 21132 6816 21148 6868
rect 21200 6816 21208 6868
rect 21132 6810 21208 6816
rect 19732 6738 19782 6792
rect 21254 6766 21314 7096
rect 21376 7056 21422 7068
rect 19454 6691 19550 6738
rect 19454 6657 19510 6691
rect 19544 6657 19550 6691
rect 19454 6619 19550 6657
rect 19454 6585 19510 6619
rect 19544 6585 19550 6619
rect 19600 6691 19646 6738
rect 19600 6657 19606 6691
rect 19640 6657 19646 6691
rect 19600 6619 19646 6657
rect 19600 6598 19606 6619
rect 19454 6538 19550 6585
rect 19590 6590 19606 6598
rect 19640 6598 19646 6619
rect 19696 6691 19782 6738
rect 20786 6746 21314 6766
rect 20786 6712 20798 6746
rect 20832 6732 21314 6746
rect 20832 6712 20844 6732
rect 20786 6698 20844 6712
rect 19696 6657 19702 6691
rect 19736 6657 19782 6691
rect 19696 6619 19782 6657
rect 19640 6590 19656 6598
rect 19590 6538 19598 6590
rect 19650 6538 19656 6590
rect 19696 6585 19702 6619
rect 19736 6585 19782 6619
rect 19858 6659 19924 6672
rect 19858 6625 19874 6659
rect 19908 6625 19924 6659
rect 20252 6652 20320 6654
rect 19858 6614 19924 6625
rect 20168 6648 20320 6652
rect 20168 6642 20261 6648
rect 20168 6608 20188 6642
rect 20222 6608 20261 6642
rect 20168 6602 20261 6608
rect 20252 6596 20261 6602
rect 20313 6596 20320 6648
rect 20252 6590 20320 6596
rect 20356 6636 20430 6660
rect 20356 6602 20384 6636
rect 20418 6602 20430 6636
rect 19696 6542 19782 6585
rect 20356 6582 20430 6602
rect 20554 6652 20626 6664
rect 20554 6600 20565 6652
rect 20617 6600 20626 6652
rect 21100 6659 21166 6668
rect 21100 6625 21116 6659
rect 21150 6625 21166 6659
rect 21100 6612 21166 6625
rect 20554 6596 20626 6600
rect 19696 6538 19742 6542
rect 19590 6530 19656 6538
rect 19824 6531 19870 6578
rect 19366 6491 19604 6500
rect 19366 6468 19558 6491
rect 19266 6442 19272 6459
rect 18024 6376 18096 6404
rect 19178 6378 19224 6425
rect 19254 6436 19272 6442
rect 19306 6442 19312 6459
rect 19364 6457 19558 6468
rect 19592 6457 19604 6491
rect 19824 6497 19830 6531
rect 19864 6497 19870 6531
rect 19824 6464 19870 6497
rect 19306 6436 19320 6442
rect 19254 6384 19260 6436
rect 19312 6384 19320 6436
rect 19254 6378 19320 6384
rect 19364 6440 19604 6457
rect 17712 6328 17802 6349
rect 17970 6331 18036 6340
rect 17970 6297 17986 6331
rect 18020 6297 18036 6331
rect 17970 6294 18036 6297
rect 17476 6266 18036 6294
rect 17380 6210 17448 6224
rect 17380 6176 17398 6210
rect 17432 6176 17448 6210
rect 17380 6166 17448 6176
rect 17420 5862 17448 6166
rect 17476 6084 17510 6266
rect 17808 6200 17880 6212
rect 17808 6148 17818 6200
rect 17870 6148 17880 6200
rect 17808 6136 17880 6148
rect 17732 6084 17796 6102
rect 17476 6050 17748 6084
rect 17782 6050 17796 6084
rect 17732 6040 17796 6050
rect 18068 6026 18096 6376
rect 18136 6342 18412 6372
rect 18136 6341 18168 6342
rect 18220 6341 18412 6342
rect 18136 6307 18165 6341
rect 18220 6307 18257 6341
rect 18291 6307 18349 6341
rect 18383 6307 18412 6341
rect 18136 6290 18168 6307
rect 18220 6290 18412 6307
rect 18136 6276 18412 6290
rect 18480 6348 19104 6366
rect 18480 6335 19022 6348
rect 18480 6301 18511 6335
rect 18545 6301 18603 6335
rect 18637 6301 18695 6335
rect 18729 6333 19022 6335
rect 19074 6333 19104 6348
rect 18729 6301 18857 6333
rect 18480 6299 18857 6301
rect 18891 6299 18949 6333
rect 18983 6299 19022 6333
rect 19075 6299 19104 6333
rect 18480 6296 19022 6299
rect 19074 6296 19104 6299
rect 18186 6084 18252 6090
rect 18186 6032 18192 6084
rect 18244 6032 18252 6084
rect 18186 6026 18252 6032
rect 17842 6012 18096 6026
rect 17598 6000 17644 6012
rect 17144 5834 17448 5862
rect 17564 5966 17604 6000
rect 17638 5966 17644 6000
rect 17564 5928 17644 5966
rect 17684 6006 17750 6012
rect 17684 5954 17690 6006
rect 17742 5954 17750 6006
rect 17684 5948 17750 5954
rect 17790 6000 18096 6012
rect 17790 5966 17796 6000
rect 17830 5998 18096 6000
rect 17830 5966 17892 5998
rect 17564 5894 17604 5928
rect 17638 5894 17644 5928
rect 17564 5882 17644 5894
rect 17694 5928 17740 5948
rect 17694 5894 17700 5928
rect 17734 5894 17740 5928
rect 17694 5882 17740 5894
rect 17790 5928 17892 5966
rect 17790 5894 17796 5928
rect 17830 5894 17892 5928
rect 17790 5882 17892 5894
rect 18012 5951 18246 5960
rect 18012 5899 18018 5951
rect 18070 5932 18194 5951
rect 18070 5899 18076 5932
rect 18012 5892 18076 5899
rect 18188 5899 18194 5932
rect 18246 5899 18252 5932
rect 18188 5892 18252 5899
rect 17144 5831 17420 5834
rect 17144 5797 17173 5831
rect 17207 5797 17265 5831
rect 17299 5797 17357 5831
rect 17391 5797 17420 5831
rect 17144 5766 17420 5797
rect 17250 5718 17314 5724
rect 17250 5666 17256 5718
rect 17308 5666 17314 5718
rect 17250 5660 17314 5666
rect 17564 5682 17610 5882
rect 17640 5844 17698 5854
rect 17640 5810 17652 5844
rect 17686 5810 17698 5844
rect 17640 5792 17698 5810
rect 17752 5763 17810 5780
rect 17752 5729 17764 5763
rect 17798 5729 17810 5763
rect 17752 5714 17810 5729
rect 17842 5682 17892 5882
rect 17958 5831 18234 5862
rect 17958 5797 17987 5831
rect 18021 5797 18079 5831
rect 18113 5797 18171 5831
rect 18205 5797 18234 5831
rect 17958 5766 18234 5797
rect 17564 5635 17660 5682
rect 17162 5602 17226 5608
rect 17162 5550 17168 5602
rect 17220 5550 17226 5602
rect 17162 5544 17226 5550
rect 17332 5592 17402 5610
rect 17332 5558 17353 5592
rect 17387 5558 17402 5592
rect 17332 5550 17402 5558
rect 17564 5601 17620 5635
rect 17654 5601 17660 5635
rect 17564 5563 17660 5601
rect 17332 5514 17360 5550
rect 17564 5529 17620 5563
rect 17654 5529 17660 5563
rect 17710 5635 17756 5682
rect 17710 5601 17716 5635
rect 17750 5601 17756 5635
rect 17710 5563 17756 5601
rect 17710 5542 17716 5563
rect 17564 5514 17660 5529
rect 17332 5482 17660 5514
rect 17700 5534 17716 5542
rect 17750 5542 17756 5563
rect 17806 5635 17892 5682
rect 18064 5716 18132 5726
rect 18064 5664 18072 5716
rect 18124 5664 18132 5716
rect 18064 5658 18132 5664
rect 17806 5601 17812 5635
rect 17846 5601 17892 5635
rect 17806 5563 17892 5601
rect 17750 5534 17766 5542
rect 17700 5482 17708 5534
rect 17760 5482 17766 5534
rect 17806 5529 17812 5563
rect 17846 5529 17892 5563
rect 17974 5604 18042 5610
rect 17974 5552 17980 5604
rect 18032 5552 18042 5604
rect 17974 5546 18042 5552
rect 18148 5590 18214 5602
rect 18148 5556 18165 5590
rect 18199 5556 18214 5590
rect 18148 5548 18214 5556
rect 17806 5510 17892 5529
rect 18186 5510 18214 5548
rect 17806 5482 18214 5510
rect 17700 5474 17766 5482
rect 17848 5478 18214 5482
rect 17652 5435 17714 5444
rect 17652 5401 17668 5435
rect 17702 5401 17714 5435
rect 17652 5384 17714 5401
rect 17656 5382 17714 5384
rect 17710 5327 17800 5348
rect 17710 5318 17737 5327
rect 15883 5293 17737 5318
rect 17771 5318 17800 5327
rect 18314 5318 18392 6276
rect 18480 6264 19104 6296
rect 19212 6331 19278 6342
rect 19212 6297 19228 6331
rect 19262 6297 19278 6331
rect 19212 6286 19278 6297
rect 19364 6294 19398 6440
rect 19546 6438 19604 6440
rect 19802 6459 19870 6464
rect 19802 6456 19830 6459
rect 19802 6404 19810 6456
rect 19864 6425 19870 6459
rect 19862 6404 19870 6425
rect 19600 6383 19690 6404
rect 19802 6398 19870 6404
rect 19600 6349 19627 6383
rect 19661 6349 19690 6383
rect 19824 6378 19870 6398
rect 19912 6531 19958 6578
rect 19912 6497 19918 6531
rect 19952 6497 19958 6531
rect 19912 6459 19958 6497
rect 19912 6425 19918 6459
rect 19952 6425 19958 6459
rect 19912 6404 19958 6425
rect 21066 6531 21112 6578
rect 21066 6497 21072 6531
rect 21106 6497 21112 6531
rect 21066 6459 21112 6497
rect 21066 6425 21072 6459
rect 21106 6425 21112 6459
rect 21154 6531 21200 6578
rect 21154 6497 21160 6531
rect 21194 6497 21200 6531
rect 21154 6459 21200 6497
rect 21254 6500 21314 6732
rect 21342 7022 21382 7056
rect 21416 7022 21422 7056
rect 21342 6984 21422 7022
rect 21462 7062 21528 7068
rect 21462 7010 21468 7062
rect 21520 7010 21528 7062
rect 21462 7004 21528 7010
rect 21568 7056 21670 7068
rect 21568 7022 21574 7056
rect 21608 7022 21670 7056
rect 21342 6950 21382 6984
rect 21416 6950 21422 6984
rect 21342 6938 21422 6950
rect 21472 6984 21518 7004
rect 21472 6950 21478 6984
rect 21512 6950 21518 6984
rect 21472 6938 21518 6950
rect 21568 6984 21670 7022
rect 21568 6950 21574 6984
rect 21608 6950 21670 6984
rect 21568 6938 21670 6950
rect 21342 6738 21388 6938
rect 21418 6900 21476 6910
rect 21418 6866 21430 6900
rect 21464 6866 21476 6900
rect 21418 6848 21476 6866
rect 21620 6858 21670 6938
rect 22036 6916 22120 7186
rect 21778 6906 21836 6912
rect 21770 6900 21844 6906
rect 21530 6819 21588 6836
rect 21530 6785 21542 6819
rect 21576 6785 21588 6819
rect 21530 6770 21588 6785
rect 21620 6792 21690 6858
rect 21770 6848 21781 6900
rect 21833 6848 21844 6900
rect 21770 6842 21844 6848
rect 21912 6890 22188 6916
rect 22782 6910 22880 7186
rect 21912 6885 22013 6890
rect 22065 6885 22188 6890
rect 21912 6851 21941 6885
rect 21975 6851 22013 6885
rect 22067 6851 22125 6885
rect 22159 6851 22188 6885
rect 21778 6834 21836 6842
rect 21912 6838 22013 6851
rect 22065 6838 22188 6851
rect 21912 6820 22188 6838
rect 22258 6879 22880 6910
rect 22258 6845 22287 6879
rect 22321 6845 22379 6879
rect 22413 6845 22471 6879
rect 22505 6877 22880 6879
rect 22505 6845 22633 6877
rect 22258 6843 22633 6845
rect 22667 6843 22725 6877
rect 22759 6843 22817 6877
rect 22851 6843 22880 6877
rect 23142 7140 23462 7158
rect 23142 7106 23414 7140
rect 23448 7106 23462 7140
rect 23142 7096 23462 7106
rect 22258 6812 22880 6843
rect 23020 6868 23096 6874
rect 23020 6816 23036 6868
rect 23088 6816 23096 6868
rect 23020 6810 23096 6816
rect 21620 6738 21670 6792
rect 23142 6766 23202 7096
rect 23264 7056 23310 7068
rect 21342 6691 21438 6738
rect 21342 6657 21398 6691
rect 21432 6657 21438 6691
rect 21342 6619 21438 6657
rect 21342 6585 21398 6619
rect 21432 6585 21438 6619
rect 21488 6691 21534 6738
rect 21488 6657 21494 6691
rect 21528 6657 21534 6691
rect 21488 6619 21534 6657
rect 21488 6598 21494 6619
rect 21342 6538 21438 6585
rect 21478 6590 21494 6598
rect 21528 6598 21534 6619
rect 21584 6691 21670 6738
rect 22674 6746 23202 6766
rect 22674 6712 22686 6746
rect 22720 6732 23202 6746
rect 22720 6712 22732 6732
rect 22674 6698 22732 6712
rect 21584 6657 21590 6691
rect 21624 6657 21670 6691
rect 21584 6619 21670 6657
rect 21528 6590 21544 6598
rect 21478 6538 21486 6590
rect 21538 6538 21544 6590
rect 21584 6585 21590 6619
rect 21624 6585 21670 6619
rect 21746 6659 21812 6672
rect 21746 6625 21762 6659
rect 21796 6625 21812 6659
rect 22140 6652 22208 6654
rect 21746 6614 21812 6625
rect 22056 6648 22208 6652
rect 22056 6642 22149 6648
rect 22056 6608 22076 6642
rect 22110 6608 22149 6642
rect 22056 6602 22149 6608
rect 22140 6596 22149 6602
rect 22201 6596 22208 6648
rect 22140 6590 22208 6596
rect 22244 6636 22318 6660
rect 22244 6602 22272 6636
rect 22306 6602 22318 6636
rect 21584 6542 21670 6585
rect 22244 6582 22318 6602
rect 22442 6652 22514 6664
rect 22442 6600 22453 6652
rect 22505 6600 22514 6652
rect 22988 6659 23054 6668
rect 22988 6625 23004 6659
rect 23038 6625 23054 6659
rect 22988 6612 23054 6625
rect 22442 6596 22514 6600
rect 21584 6538 21630 6542
rect 21478 6530 21544 6538
rect 21712 6531 21758 6578
rect 21254 6491 21492 6500
rect 21254 6468 21446 6491
rect 21154 6442 21160 6459
rect 19912 6376 19984 6404
rect 21066 6378 21112 6425
rect 21142 6436 21160 6442
rect 21194 6442 21200 6459
rect 21252 6457 21446 6468
rect 21480 6457 21492 6491
rect 21712 6497 21718 6531
rect 21752 6497 21758 6531
rect 21712 6464 21758 6497
rect 21194 6436 21208 6442
rect 21142 6384 21148 6436
rect 21200 6384 21208 6436
rect 21142 6378 21208 6384
rect 21252 6440 21492 6457
rect 19600 6328 19690 6349
rect 19858 6331 19924 6340
rect 19858 6297 19874 6331
rect 19908 6297 19924 6331
rect 19858 6294 19924 6297
rect 19364 6266 19924 6294
rect 19268 6210 19336 6224
rect 19268 6176 19286 6210
rect 19320 6176 19336 6210
rect 19268 6166 19336 6176
rect 19308 5862 19336 6166
rect 19364 6084 19398 6266
rect 19696 6200 19768 6212
rect 19696 6148 19706 6200
rect 19758 6148 19768 6200
rect 19696 6136 19768 6148
rect 19620 6084 19684 6102
rect 19364 6050 19636 6084
rect 19670 6050 19684 6084
rect 19620 6040 19684 6050
rect 19956 6026 19984 6376
rect 20024 6342 20300 6372
rect 20024 6341 20056 6342
rect 20108 6341 20300 6342
rect 20024 6307 20053 6341
rect 20108 6307 20145 6341
rect 20179 6307 20237 6341
rect 20271 6307 20300 6341
rect 20024 6290 20056 6307
rect 20108 6290 20300 6307
rect 20024 6276 20300 6290
rect 20368 6348 20992 6366
rect 20368 6335 20910 6348
rect 20368 6301 20399 6335
rect 20433 6301 20491 6335
rect 20525 6301 20583 6335
rect 20617 6333 20910 6335
rect 20962 6333 20992 6348
rect 20617 6301 20745 6333
rect 20368 6299 20745 6301
rect 20779 6299 20837 6333
rect 20871 6299 20910 6333
rect 20963 6299 20992 6333
rect 20368 6296 20910 6299
rect 20962 6296 20992 6299
rect 20074 6084 20140 6090
rect 20074 6032 20080 6084
rect 20132 6032 20140 6084
rect 20074 6026 20140 6032
rect 19730 6012 19984 6026
rect 19486 6000 19532 6012
rect 19032 5834 19336 5862
rect 19452 5966 19492 6000
rect 19526 5966 19532 6000
rect 19452 5928 19532 5966
rect 19572 6006 19638 6012
rect 19572 5954 19578 6006
rect 19630 5954 19638 6006
rect 19572 5948 19638 5954
rect 19678 6000 19984 6012
rect 19678 5966 19684 6000
rect 19718 5998 19984 6000
rect 19718 5966 19780 5998
rect 19452 5894 19492 5928
rect 19526 5894 19532 5928
rect 19452 5882 19532 5894
rect 19582 5928 19628 5948
rect 19582 5894 19588 5928
rect 19622 5894 19628 5928
rect 19582 5882 19628 5894
rect 19678 5928 19780 5966
rect 19678 5894 19684 5928
rect 19718 5894 19780 5928
rect 19678 5882 19780 5894
rect 19900 5951 20134 5960
rect 19900 5899 19906 5951
rect 19958 5932 20082 5951
rect 19958 5899 19964 5932
rect 19900 5892 19964 5899
rect 20076 5899 20082 5932
rect 20134 5899 20140 5932
rect 20076 5892 20140 5899
rect 19032 5831 19308 5834
rect 19032 5797 19061 5831
rect 19095 5797 19153 5831
rect 19187 5797 19245 5831
rect 19279 5797 19308 5831
rect 19032 5766 19308 5797
rect 19138 5718 19202 5724
rect 19138 5666 19144 5718
rect 19196 5666 19202 5718
rect 19138 5660 19202 5666
rect 19452 5682 19498 5882
rect 19528 5844 19586 5854
rect 19528 5810 19540 5844
rect 19574 5810 19586 5844
rect 19528 5792 19586 5810
rect 19640 5763 19698 5780
rect 19640 5729 19652 5763
rect 19686 5729 19698 5763
rect 19640 5714 19698 5729
rect 19730 5682 19780 5882
rect 19846 5831 20122 5862
rect 19846 5797 19875 5831
rect 19909 5797 19967 5831
rect 20001 5797 20059 5831
rect 20093 5797 20122 5831
rect 19846 5766 20122 5797
rect 19452 5635 19548 5682
rect 19050 5602 19114 5608
rect 19050 5550 19056 5602
rect 19108 5550 19114 5602
rect 19050 5544 19114 5550
rect 19220 5592 19290 5610
rect 19220 5558 19241 5592
rect 19275 5558 19290 5592
rect 19220 5550 19290 5558
rect 19452 5601 19508 5635
rect 19542 5601 19548 5635
rect 19452 5563 19548 5601
rect 19220 5514 19248 5550
rect 19452 5529 19508 5563
rect 19542 5529 19548 5563
rect 19598 5635 19644 5682
rect 19598 5601 19604 5635
rect 19638 5601 19644 5635
rect 19598 5563 19644 5601
rect 19598 5542 19604 5563
rect 19452 5514 19548 5529
rect 19220 5482 19548 5514
rect 19588 5534 19604 5542
rect 19638 5542 19644 5563
rect 19694 5635 19780 5682
rect 19952 5716 20020 5726
rect 19952 5664 19960 5716
rect 20012 5664 20020 5716
rect 19952 5658 20020 5664
rect 19694 5601 19700 5635
rect 19734 5601 19780 5635
rect 19694 5563 19780 5601
rect 19638 5534 19654 5542
rect 19588 5482 19596 5534
rect 19648 5482 19654 5534
rect 19694 5529 19700 5563
rect 19734 5529 19780 5563
rect 19862 5604 19930 5610
rect 19862 5552 19868 5604
rect 19920 5552 19930 5604
rect 19862 5546 19930 5552
rect 20036 5590 20102 5602
rect 20036 5556 20053 5590
rect 20087 5556 20102 5590
rect 20036 5548 20102 5556
rect 19694 5510 19780 5529
rect 20074 5510 20102 5548
rect 19694 5482 20102 5510
rect 19588 5474 19654 5482
rect 19736 5478 20102 5482
rect 19540 5435 19602 5444
rect 19540 5401 19556 5435
rect 19590 5401 19602 5435
rect 19540 5384 19602 5401
rect 19544 5382 19602 5384
rect 19598 5327 19688 5348
rect 19598 5318 19625 5327
rect 17771 5293 19625 5318
rect 19659 5318 19688 5327
rect 20202 5318 20280 6276
rect 20368 6264 20992 6296
rect 21100 6331 21166 6342
rect 21100 6297 21116 6331
rect 21150 6297 21166 6331
rect 21100 6286 21166 6297
rect 21252 6294 21286 6440
rect 21434 6438 21492 6440
rect 21690 6459 21758 6464
rect 21690 6456 21718 6459
rect 21690 6404 21698 6456
rect 21752 6425 21758 6459
rect 21750 6404 21758 6425
rect 21488 6383 21578 6404
rect 21690 6398 21758 6404
rect 21488 6349 21515 6383
rect 21549 6349 21578 6383
rect 21712 6378 21758 6398
rect 21800 6531 21846 6578
rect 21800 6497 21806 6531
rect 21840 6497 21846 6531
rect 21800 6459 21846 6497
rect 21800 6425 21806 6459
rect 21840 6425 21846 6459
rect 21800 6404 21846 6425
rect 22954 6531 23000 6578
rect 22954 6497 22960 6531
rect 22994 6497 23000 6531
rect 22954 6459 23000 6497
rect 22954 6425 22960 6459
rect 22994 6425 23000 6459
rect 23042 6531 23088 6578
rect 23042 6497 23048 6531
rect 23082 6497 23088 6531
rect 23042 6459 23088 6497
rect 23142 6500 23202 6732
rect 23230 7022 23270 7056
rect 23304 7022 23310 7056
rect 23230 6984 23310 7022
rect 23350 7062 23416 7068
rect 23350 7010 23356 7062
rect 23408 7010 23416 7062
rect 23350 7004 23416 7010
rect 23456 7056 23558 7068
rect 23456 7022 23462 7056
rect 23496 7022 23558 7056
rect 23230 6950 23270 6984
rect 23304 6950 23310 6984
rect 23230 6938 23310 6950
rect 23360 6984 23406 7004
rect 23360 6950 23366 6984
rect 23400 6950 23406 6984
rect 23360 6938 23406 6950
rect 23456 6984 23558 7022
rect 23456 6950 23462 6984
rect 23496 6950 23558 6984
rect 23456 6938 23558 6950
rect 23230 6738 23276 6938
rect 23306 6900 23364 6910
rect 23306 6866 23318 6900
rect 23352 6866 23364 6900
rect 23306 6848 23364 6866
rect 23508 6858 23558 6938
rect 23924 6916 24008 7186
rect 23666 6906 23724 6912
rect 23658 6900 23732 6906
rect 23418 6819 23476 6836
rect 23418 6785 23430 6819
rect 23464 6785 23476 6819
rect 23418 6770 23476 6785
rect 23508 6792 23578 6858
rect 23658 6848 23669 6900
rect 23721 6848 23732 6900
rect 23658 6842 23732 6848
rect 23800 6890 24076 6916
rect 24670 6910 24768 7186
rect 23800 6885 23901 6890
rect 23953 6885 24076 6890
rect 23800 6851 23829 6885
rect 23863 6851 23901 6885
rect 23955 6851 24013 6885
rect 24047 6851 24076 6885
rect 23666 6834 23724 6842
rect 23800 6838 23901 6851
rect 23953 6838 24076 6851
rect 23800 6820 24076 6838
rect 24146 6879 24768 6910
rect 24146 6845 24175 6879
rect 24209 6845 24267 6879
rect 24301 6845 24359 6879
rect 24393 6877 24768 6879
rect 24393 6845 24521 6877
rect 24146 6843 24521 6845
rect 24555 6843 24613 6877
rect 24647 6843 24705 6877
rect 24739 6843 24768 6877
rect 25030 7140 25350 7158
rect 25030 7106 25302 7140
rect 25336 7106 25350 7140
rect 25030 7096 25350 7106
rect 24146 6812 24768 6843
rect 24908 6868 24984 6874
rect 24908 6816 24924 6868
rect 24976 6816 24984 6868
rect 24908 6810 24984 6816
rect 23508 6738 23558 6792
rect 25030 6766 25090 7096
rect 25152 7056 25198 7068
rect 23230 6691 23326 6738
rect 23230 6657 23286 6691
rect 23320 6657 23326 6691
rect 23230 6619 23326 6657
rect 23230 6585 23286 6619
rect 23320 6585 23326 6619
rect 23376 6691 23422 6738
rect 23376 6657 23382 6691
rect 23416 6657 23422 6691
rect 23376 6619 23422 6657
rect 23376 6598 23382 6619
rect 23230 6538 23326 6585
rect 23366 6590 23382 6598
rect 23416 6598 23422 6619
rect 23472 6691 23558 6738
rect 24562 6746 25090 6766
rect 24562 6712 24574 6746
rect 24608 6732 25090 6746
rect 24608 6712 24620 6732
rect 24562 6698 24620 6712
rect 23472 6657 23478 6691
rect 23512 6657 23558 6691
rect 23472 6619 23558 6657
rect 23416 6590 23432 6598
rect 23366 6538 23374 6590
rect 23426 6538 23432 6590
rect 23472 6585 23478 6619
rect 23512 6585 23558 6619
rect 23634 6659 23700 6672
rect 23634 6625 23650 6659
rect 23684 6625 23700 6659
rect 24028 6652 24096 6654
rect 23634 6614 23700 6625
rect 23944 6648 24096 6652
rect 23944 6642 24037 6648
rect 23944 6608 23964 6642
rect 23998 6608 24037 6642
rect 23944 6602 24037 6608
rect 24028 6596 24037 6602
rect 24089 6596 24096 6648
rect 24028 6590 24096 6596
rect 24132 6636 24206 6660
rect 24132 6602 24160 6636
rect 24194 6602 24206 6636
rect 23472 6542 23558 6585
rect 24132 6582 24206 6602
rect 24330 6652 24402 6664
rect 24330 6600 24341 6652
rect 24393 6600 24402 6652
rect 24876 6659 24942 6668
rect 24876 6625 24892 6659
rect 24926 6625 24942 6659
rect 24876 6612 24942 6625
rect 24330 6596 24402 6600
rect 23472 6538 23518 6542
rect 23366 6530 23432 6538
rect 23600 6531 23646 6578
rect 23142 6491 23380 6500
rect 23142 6468 23334 6491
rect 23042 6442 23048 6459
rect 21800 6376 21872 6404
rect 22954 6378 23000 6425
rect 23030 6436 23048 6442
rect 23082 6442 23088 6459
rect 23140 6457 23334 6468
rect 23368 6457 23380 6491
rect 23600 6497 23606 6531
rect 23640 6497 23646 6531
rect 23600 6464 23646 6497
rect 23082 6436 23096 6442
rect 23030 6384 23036 6436
rect 23088 6384 23096 6436
rect 23030 6378 23096 6384
rect 23140 6440 23380 6457
rect 21488 6328 21578 6349
rect 21746 6331 21812 6340
rect 21746 6297 21762 6331
rect 21796 6297 21812 6331
rect 21746 6294 21812 6297
rect 21252 6266 21812 6294
rect 21156 6210 21224 6224
rect 21156 6176 21174 6210
rect 21208 6176 21224 6210
rect 21156 6166 21224 6176
rect 21196 5862 21224 6166
rect 21252 6084 21286 6266
rect 21584 6200 21656 6212
rect 21584 6148 21594 6200
rect 21646 6148 21656 6200
rect 21584 6136 21656 6148
rect 21508 6084 21572 6102
rect 21252 6050 21524 6084
rect 21558 6050 21572 6084
rect 21508 6040 21572 6050
rect 21844 6026 21872 6376
rect 21912 6342 22188 6372
rect 21912 6341 21944 6342
rect 21996 6341 22188 6342
rect 21912 6307 21941 6341
rect 21996 6307 22033 6341
rect 22067 6307 22125 6341
rect 22159 6307 22188 6341
rect 21912 6290 21944 6307
rect 21996 6290 22188 6307
rect 21912 6276 22188 6290
rect 22256 6348 22880 6366
rect 22256 6335 22798 6348
rect 22256 6301 22287 6335
rect 22321 6301 22379 6335
rect 22413 6301 22471 6335
rect 22505 6333 22798 6335
rect 22850 6333 22880 6348
rect 22505 6301 22633 6333
rect 22256 6299 22633 6301
rect 22667 6299 22725 6333
rect 22759 6299 22798 6333
rect 22851 6299 22880 6333
rect 22256 6296 22798 6299
rect 22850 6296 22880 6299
rect 21962 6084 22028 6090
rect 21962 6032 21968 6084
rect 22020 6032 22028 6084
rect 21962 6026 22028 6032
rect 21618 6012 21872 6026
rect 21374 6000 21420 6012
rect 20920 5834 21224 5862
rect 21340 5966 21380 6000
rect 21414 5966 21420 6000
rect 21340 5928 21420 5966
rect 21460 6006 21526 6012
rect 21460 5954 21466 6006
rect 21518 5954 21526 6006
rect 21460 5948 21526 5954
rect 21566 6000 21872 6012
rect 21566 5966 21572 6000
rect 21606 5998 21872 6000
rect 21606 5966 21668 5998
rect 21340 5894 21380 5928
rect 21414 5894 21420 5928
rect 21340 5882 21420 5894
rect 21470 5928 21516 5948
rect 21470 5894 21476 5928
rect 21510 5894 21516 5928
rect 21470 5882 21516 5894
rect 21566 5928 21668 5966
rect 21566 5894 21572 5928
rect 21606 5894 21668 5928
rect 21566 5882 21668 5894
rect 21788 5951 22022 5960
rect 21788 5899 21794 5951
rect 21846 5932 21970 5951
rect 21846 5899 21852 5932
rect 21788 5892 21852 5899
rect 21964 5899 21970 5932
rect 22022 5899 22028 5932
rect 21964 5892 22028 5899
rect 20920 5831 21196 5834
rect 20920 5797 20949 5831
rect 20983 5797 21041 5831
rect 21075 5797 21133 5831
rect 21167 5797 21196 5831
rect 20920 5766 21196 5797
rect 21026 5718 21090 5724
rect 21026 5666 21032 5718
rect 21084 5666 21090 5718
rect 21026 5660 21090 5666
rect 21340 5682 21386 5882
rect 21416 5844 21474 5854
rect 21416 5810 21428 5844
rect 21462 5810 21474 5844
rect 21416 5792 21474 5810
rect 21528 5763 21586 5780
rect 21528 5729 21540 5763
rect 21574 5729 21586 5763
rect 21528 5714 21586 5729
rect 21618 5682 21668 5882
rect 21734 5831 22010 5862
rect 21734 5797 21763 5831
rect 21797 5797 21855 5831
rect 21889 5797 21947 5831
rect 21981 5797 22010 5831
rect 21734 5766 22010 5797
rect 21340 5635 21436 5682
rect 20938 5602 21002 5608
rect 20938 5550 20944 5602
rect 20996 5550 21002 5602
rect 20938 5544 21002 5550
rect 21108 5592 21178 5610
rect 21108 5558 21129 5592
rect 21163 5558 21178 5592
rect 21108 5550 21178 5558
rect 21340 5601 21396 5635
rect 21430 5601 21436 5635
rect 21340 5563 21436 5601
rect 21108 5514 21136 5550
rect 21340 5529 21396 5563
rect 21430 5529 21436 5563
rect 21486 5635 21532 5682
rect 21486 5601 21492 5635
rect 21526 5601 21532 5635
rect 21486 5563 21532 5601
rect 21486 5542 21492 5563
rect 21340 5514 21436 5529
rect 21108 5482 21436 5514
rect 21476 5534 21492 5542
rect 21526 5542 21532 5563
rect 21582 5635 21668 5682
rect 21840 5716 21908 5726
rect 21840 5664 21848 5716
rect 21900 5664 21908 5716
rect 21840 5658 21908 5664
rect 21582 5601 21588 5635
rect 21622 5601 21668 5635
rect 21582 5563 21668 5601
rect 21526 5534 21542 5542
rect 21476 5482 21484 5534
rect 21536 5482 21542 5534
rect 21582 5529 21588 5563
rect 21622 5529 21668 5563
rect 21750 5604 21818 5610
rect 21750 5552 21756 5604
rect 21808 5552 21818 5604
rect 21750 5546 21818 5552
rect 21924 5590 21990 5602
rect 21924 5556 21941 5590
rect 21975 5556 21990 5590
rect 21924 5548 21990 5556
rect 21582 5510 21668 5529
rect 21962 5510 21990 5548
rect 21582 5482 21990 5510
rect 21476 5474 21542 5482
rect 21624 5478 21990 5482
rect 21428 5435 21490 5444
rect 21428 5401 21444 5435
rect 21478 5401 21490 5435
rect 21428 5384 21490 5401
rect 21432 5382 21490 5384
rect 21486 5327 21576 5348
rect 21486 5318 21513 5327
rect 19659 5293 21513 5318
rect 21547 5318 21576 5327
rect 22090 5318 22168 6276
rect 22256 6264 22880 6296
rect 22988 6331 23054 6342
rect 22988 6297 23004 6331
rect 23038 6297 23054 6331
rect 22988 6286 23054 6297
rect 23140 6294 23174 6440
rect 23322 6438 23380 6440
rect 23578 6459 23646 6464
rect 23578 6456 23606 6459
rect 23578 6404 23586 6456
rect 23640 6425 23646 6459
rect 23638 6404 23646 6425
rect 23376 6383 23466 6404
rect 23578 6398 23646 6404
rect 23376 6349 23403 6383
rect 23437 6349 23466 6383
rect 23600 6378 23646 6398
rect 23688 6531 23734 6578
rect 23688 6497 23694 6531
rect 23728 6497 23734 6531
rect 23688 6459 23734 6497
rect 23688 6425 23694 6459
rect 23728 6425 23734 6459
rect 23688 6404 23734 6425
rect 24842 6531 24888 6578
rect 24842 6497 24848 6531
rect 24882 6497 24888 6531
rect 24842 6459 24888 6497
rect 24842 6425 24848 6459
rect 24882 6425 24888 6459
rect 24930 6531 24976 6578
rect 24930 6497 24936 6531
rect 24970 6497 24976 6531
rect 24930 6459 24976 6497
rect 25030 6500 25090 6732
rect 25118 7022 25158 7056
rect 25192 7022 25198 7056
rect 25118 6984 25198 7022
rect 25238 7062 25304 7068
rect 25238 7010 25244 7062
rect 25296 7010 25304 7062
rect 25238 7004 25304 7010
rect 25344 7056 25446 7068
rect 25344 7022 25350 7056
rect 25384 7022 25446 7056
rect 25118 6950 25158 6984
rect 25192 6950 25198 6984
rect 25118 6938 25198 6950
rect 25248 6984 25294 7004
rect 25248 6950 25254 6984
rect 25288 6950 25294 6984
rect 25248 6938 25294 6950
rect 25344 6984 25446 7022
rect 25344 6950 25350 6984
rect 25384 6950 25446 6984
rect 25344 6938 25446 6950
rect 25118 6738 25164 6938
rect 25194 6900 25252 6910
rect 25194 6866 25206 6900
rect 25240 6866 25252 6900
rect 25194 6848 25252 6866
rect 25396 6858 25446 6938
rect 25812 6916 25896 7186
rect 25554 6906 25612 6912
rect 25546 6900 25620 6906
rect 25306 6819 25364 6836
rect 25306 6785 25318 6819
rect 25352 6785 25364 6819
rect 25306 6770 25364 6785
rect 25396 6792 25466 6858
rect 25546 6848 25557 6900
rect 25609 6848 25620 6900
rect 25546 6842 25620 6848
rect 25688 6890 25964 6916
rect 26558 6910 26656 7186
rect 25688 6885 25789 6890
rect 25841 6885 25964 6890
rect 25688 6851 25717 6885
rect 25751 6851 25789 6885
rect 25843 6851 25901 6885
rect 25935 6851 25964 6885
rect 25554 6834 25612 6842
rect 25688 6838 25789 6851
rect 25841 6838 25964 6851
rect 25688 6820 25964 6838
rect 26034 6879 26656 6910
rect 26034 6845 26063 6879
rect 26097 6845 26155 6879
rect 26189 6845 26247 6879
rect 26281 6877 26656 6879
rect 26281 6845 26409 6877
rect 26034 6843 26409 6845
rect 26443 6843 26501 6877
rect 26535 6843 26593 6877
rect 26627 6843 26656 6877
rect 26918 7140 27238 7158
rect 26918 7106 27190 7140
rect 27224 7106 27238 7140
rect 26918 7096 27238 7106
rect 26034 6812 26656 6843
rect 26796 6868 26872 6874
rect 26796 6816 26812 6868
rect 26864 6816 26872 6868
rect 26796 6810 26872 6816
rect 25396 6738 25446 6792
rect 26918 6766 26978 7096
rect 27040 7056 27086 7068
rect 25118 6691 25214 6738
rect 25118 6657 25174 6691
rect 25208 6657 25214 6691
rect 25118 6619 25214 6657
rect 25118 6585 25174 6619
rect 25208 6585 25214 6619
rect 25264 6691 25310 6738
rect 25264 6657 25270 6691
rect 25304 6657 25310 6691
rect 25264 6619 25310 6657
rect 25264 6598 25270 6619
rect 25118 6538 25214 6585
rect 25254 6590 25270 6598
rect 25304 6598 25310 6619
rect 25360 6691 25446 6738
rect 26450 6746 26978 6766
rect 26450 6712 26462 6746
rect 26496 6732 26978 6746
rect 26496 6712 26508 6732
rect 26450 6698 26508 6712
rect 25360 6657 25366 6691
rect 25400 6657 25446 6691
rect 25360 6619 25446 6657
rect 25304 6590 25320 6598
rect 25254 6538 25262 6590
rect 25314 6538 25320 6590
rect 25360 6585 25366 6619
rect 25400 6585 25446 6619
rect 25522 6659 25588 6672
rect 25522 6625 25538 6659
rect 25572 6625 25588 6659
rect 25916 6652 25984 6654
rect 25522 6614 25588 6625
rect 25832 6648 25984 6652
rect 25832 6642 25925 6648
rect 25832 6608 25852 6642
rect 25886 6608 25925 6642
rect 25832 6602 25925 6608
rect 25916 6596 25925 6602
rect 25977 6596 25984 6648
rect 25916 6590 25984 6596
rect 26020 6636 26094 6660
rect 26020 6602 26048 6636
rect 26082 6602 26094 6636
rect 25360 6542 25446 6585
rect 26020 6582 26094 6602
rect 26218 6652 26290 6664
rect 26218 6600 26229 6652
rect 26281 6600 26290 6652
rect 26764 6659 26830 6668
rect 26764 6625 26780 6659
rect 26814 6625 26830 6659
rect 26764 6612 26830 6625
rect 26218 6596 26290 6600
rect 25360 6538 25406 6542
rect 25254 6530 25320 6538
rect 25488 6531 25534 6578
rect 25030 6491 25268 6500
rect 25030 6468 25222 6491
rect 24930 6442 24936 6459
rect 23688 6376 23760 6404
rect 24842 6378 24888 6425
rect 24918 6436 24936 6442
rect 24970 6442 24976 6459
rect 25028 6457 25222 6468
rect 25256 6457 25268 6491
rect 25488 6497 25494 6531
rect 25528 6497 25534 6531
rect 25488 6464 25534 6497
rect 24970 6436 24984 6442
rect 24918 6384 24924 6436
rect 24976 6384 24984 6436
rect 24918 6378 24984 6384
rect 25028 6440 25268 6457
rect 23376 6328 23466 6349
rect 23634 6331 23700 6340
rect 23634 6297 23650 6331
rect 23684 6297 23700 6331
rect 23634 6294 23700 6297
rect 23140 6266 23700 6294
rect 23044 6210 23112 6224
rect 23044 6176 23062 6210
rect 23096 6176 23112 6210
rect 23044 6166 23112 6176
rect 23084 5862 23112 6166
rect 23140 6084 23174 6266
rect 23472 6200 23544 6212
rect 23472 6148 23482 6200
rect 23534 6148 23544 6200
rect 23472 6136 23544 6148
rect 23396 6084 23460 6102
rect 23140 6050 23412 6084
rect 23446 6050 23460 6084
rect 23396 6040 23460 6050
rect 23732 6026 23760 6376
rect 23800 6342 24076 6372
rect 23800 6341 23832 6342
rect 23884 6341 24076 6342
rect 23800 6307 23829 6341
rect 23884 6307 23921 6341
rect 23955 6307 24013 6341
rect 24047 6307 24076 6341
rect 23800 6290 23832 6307
rect 23884 6290 24076 6307
rect 23800 6276 24076 6290
rect 24144 6348 24768 6366
rect 24144 6335 24686 6348
rect 24144 6301 24175 6335
rect 24209 6301 24267 6335
rect 24301 6301 24359 6335
rect 24393 6333 24686 6335
rect 24738 6333 24768 6348
rect 24393 6301 24521 6333
rect 24144 6299 24521 6301
rect 24555 6299 24613 6333
rect 24647 6299 24686 6333
rect 24739 6299 24768 6333
rect 24144 6296 24686 6299
rect 24738 6296 24768 6299
rect 23850 6084 23916 6090
rect 23850 6032 23856 6084
rect 23908 6032 23916 6084
rect 23850 6026 23916 6032
rect 23506 6012 23760 6026
rect 23262 6000 23308 6012
rect 22808 5834 23112 5862
rect 23228 5966 23268 6000
rect 23302 5966 23308 6000
rect 23228 5928 23308 5966
rect 23348 6006 23414 6012
rect 23348 5954 23354 6006
rect 23406 5954 23414 6006
rect 23348 5948 23414 5954
rect 23454 6000 23760 6012
rect 23454 5966 23460 6000
rect 23494 5998 23760 6000
rect 23494 5966 23556 5998
rect 23228 5894 23268 5928
rect 23302 5894 23308 5928
rect 23228 5882 23308 5894
rect 23358 5928 23404 5948
rect 23358 5894 23364 5928
rect 23398 5894 23404 5928
rect 23358 5882 23404 5894
rect 23454 5928 23556 5966
rect 23454 5894 23460 5928
rect 23494 5894 23556 5928
rect 23454 5882 23556 5894
rect 23676 5951 23910 5960
rect 23676 5899 23682 5951
rect 23734 5932 23858 5951
rect 23734 5899 23740 5932
rect 23676 5892 23740 5899
rect 23852 5899 23858 5932
rect 23910 5899 23916 5932
rect 23852 5892 23916 5899
rect 22808 5831 23084 5834
rect 22808 5797 22837 5831
rect 22871 5797 22929 5831
rect 22963 5797 23021 5831
rect 23055 5797 23084 5831
rect 22808 5766 23084 5797
rect 22914 5718 22978 5724
rect 22914 5666 22920 5718
rect 22972 5666 22978 5718
rect 22914 5660 22978 5666
rect 23228 5682 23274 5882
rect 23304 5844 23362 5854
rect 23304 5810 23316 5844
rect 23350 5810 23362 5844
rect 23304 5792 23362 5810
rect 23416 5763 23474 5780
rect 23416 5729 23428 5763
rect 23462 5729 23474 5763
rect 23416 5714 23474 5729
rect 23506 5682 23556 5882
rect 23622 5831 23898 5862
rect 23622 5797 23651 5831
rect 23685 5797 23743 5831
rect 23777 5797 23835 5831
rect 23869 5797 23898 5831
rect 23622 5766 23898 5797
rect 23228 5635 23324 5682
rect 22826 5602 22890 5608
rect 22826 5550 22832 5602
rect 22884 5550 22890 5602
rect 22826 5544 22890 5550
rect 22996 5592 23066 5610
rect 22996 5558 23017 5592
rect 23051 5558 23066 5592
rect 22996 5550 23066 5558
rect 23228 5601 23284 5635
rect 23318 5601 23324 5635
rect 23228 5563 23324 5601
rect 22996 5514 23024 5550
rect 23228 5529 23284 5563
rect 23318 5529 23324 5563
rect 23374 5635 23420 5682
rect 23374 5601 23380 5635
rect 23414 5601 23420 5635
rect 23374 5563 23420 5601
rect 23374 5542 23380 5563
rect 23228 5514 23324 5529
rect 22996 5482 23324 5514
rect 23364 5534 23380 5542
rect 23414 5542 23420 5563
rect 23470 5635 23556 5682
rect 23728 5716 23796 5726
rect 23728 5664 23736 5716
rect 23788 5664 23796 5716
rect 23728 5658 23796 5664
rect 23470 5601 23476 5635
rect 23510 5601 23556 5635
rect 23470 5563 23556 5601
rect 23414 5534 23430 5542
rect 23364 5482 23372 5534
rect 23424 5482 23430 5534
rect 23470 5529 23476 5563
rect 23510 5529 23556 5563
rect 23638 5604 23706 5610
rect 23638 5552 23644 5604
rect 23696 5552 23706 5604
rect 23638 5546 23706 5552
rect 23812 5590 23878 5602
rect 23812 5556 23829 5590
rect 23863 5556 23878 5590
rect 23812 5548 23878 5556
rect 23470 5510 23556 5529
rect 23850 5510 23878 5548
rect 23470 5482 23878 5510
rect 23364 5474 23430 5482
rect 23512 5478 23878 5482
rect 23316 5435 23378 5444
rect 23316 5401 23332 5435
rect 23366 5401 23378 5435
rect 23316 5384 23378 5401
rect 23320 5382 23378 5384
rect 23374 5327 23464 5348
rect 23374 5318 23401 5327
rect 21547 5293 23401 5318
rect 23435 5318 23464 5327
rect 23978 5318 24056 6276
rect 24144 6264 24768 6296
rect 24876 6331 24942 6342
rect 24876 6297 24892 6331
rect 24926 6297 24942 6331
rect 24876 6286 24942 6297
rect 25028 6294 25062 6440
rect 25210 6438 25268 6440
rect 25466 6459 25534 6464
rect 25466 6456 25494 6459
rect 25466 6404 25474 6456
rect 25528 6425 25534 6459
rect 25526 6404 25534 6425
rect 25264 6383 25354 6404
rect 25466 6398 25534 6404
rect 25264 6349 25291 6383
rect 25325 6349 25354 6383
rect 25488 6378 25534 6398
rect 25576 6531 25622 6578
rect 25576 6497 25582 6531
rect 25616 6497 25622 6531
rect 25576 6459 25622 6497
rect 25576 6425 25582 6459
rect 25616 6425 25622 6459
rect 25576 6404 25622 6425
rect 26730 6531 26776 6578
rect 26730 6497 26736 6531
rect 26770 6497 26776 6531
rect 26730 6459 26776 6497
rect 26730 6425 26736 6459
rect 26770 6425 26776 6459
rect 26818 6531 26864 6578
rect 26818 6497 26824 6531
rect 26858 6497 26864 6531
rect 26818 6459 26864 6497
rect 26918 6500 26978 6732
rect 27006 7022 27046 7056
rect 27080 7022 27086 7056
rect 27006 6984 27086 7022
rect 27126 7062 27192 7068
rect 27126 7010 27132 7062
rect 27184 7010 27192 7062
rect 27126 7004 27192 7010
rect 27232 7056 27334 7068
rect 27232 7022 27238 7056
rect 27272 7022 27334 7056
rect 27006 6950 27046 6984
rect 27080 6950 27086 6984
rect 27006 6938 27086 6950
rect 27136 6984 27182 7004
rect 27136 6950 27142 6984
rect 27176 6950 27182 6984
rect 27136 6938 27182 6950
rect 27232 6984 27334 7022
rect 27232 6950 27238 6984
rect 27272 6950 27334 6984
rect 27232 6938 27334 6950
rect 27006 6738 27052 6938
rect 27082 6900 27140 6910
rect 27082 6866 27094 6900
rect 27128 6866 27140 6900
rect 27082 6848 27140 6866
rect 27284 6858 27334 6938
rect 27700 6916 27784 7186
rect 27442 6906 27500 6912
rect 27434 6900 27508 6906
rect 27194 6819 27252 6836
rect 27194 6785 27206 6819
rect 27240 6785 27252 6819
rect 27194 6770 27252 6785
rect 27284 6792 27354 6858
rect 27434 6848 27445 6900
rect 27497 6848 27508 6900
rect 27434 6842 27508 6848
rect 27576 6890 27852 6916
rect 28446 6910 28544 7186
rect 27576 6885 27677 6890
rect 27729 6885 27852 6890
rect 27576 6851 27605 6885
rect 27639 6851 27677 6885
rect 27731 6851 27789 6885
rect 27823 6851 27852 6885
rect 27442 6834 27500 6842
rect 27576 6838 27677 6851
rect 27729 6838 27852 6851
rect 27576 6820 27852 6838
rect 27922 6879 28544 6910
rect 27922 6845 27951 6879
rect 27985 6845 28043 6879
rect 28077 6845 28135 6879
rect 28169 6877 28544 6879
rect 28169 6845 28297 6877
rect 27922 6843 28297 6845
rect 28331 6843 28389 6877
rect 28423 6843 28481 6877
rect 28515 6843 28544 6877
rect 28806 7140 29126 7158
rect 28806 7106 29078 7140
rect 29112 7106 29126 7140
rect 28806 7096 29126 7106
rect 27922 6812 28544 6843
rect 28684 6868 28760 6874
rect 28684 6816 28700 6868
rect 28752 6816 28760 6868
rect 28684 6810 28760 6816
rect 27284 6738 27334 6792
rect 28806 6766 28866 7096
rect 28928 7056 28974 7068
rect 27006 6691 27102 6738
rect 27006 6657 27062 6691
rect 27096 6657 27102 6691
rect 27006 6619 27102 6657
rect 27006 6585 27062 6619
rect 27096 6585 27102 6619
rect 27152 6691 27198 6738
rect 27152 6657 27158 6691
rect 27192 6657 27198 6691
rect 27152 6619 27198 6657
rect 27152 6598 27158 6619
rect 27006 6538 27102 6585
rect 27142 6590 27158 6598
rect 27192 6598 27198 6619
rect 27248 6691 27334 6738
rect 28338 6746 28866 6766
rect 28338 6712 28350 6746
rect 28384 6732 28866 6746
rect 28384 6712 28396 6732
rect 28338 6698 28396 6712
rect 27248 6657 27254 6691
rect 27288 6657 27334 6691
rect 27248 6619 27334 6657
rect 27192 6590 27208 6598
rect 27142 6538 27150 6590
rect 27202 6538 27208 6590
rect 27248 6585 27254 6619
rect 27288 6585 27334 6619
rect 27410 6659 27476 6672
rect 27410 6625 27426 6659
rect 27460 6625 27476 6659
rect 27804 6652 27872 6654
rect 27410 6614 27476 6625
rect 27720 6648 27872 6652
rect 27720 6642 27813 6648
rect 27720 6608 27740 6642
rect 27774 6608 27813 6642
rect 27720 6602 27813 6608
rect 27804 6596 27813 6602
rect 27865 6596 27872 6648
rect 27804 6590 27872 6596
rect 27908 6636 27982 6660
rect 27908 6602 27936 6636
rect 27970 6602 27982 6636
rect 27248 6542 27334 6585
rect 27908 6582 27982 6602
rect 28106 6652 28178 6664
rect 28106 6600 28117 6652
rect 28169 6600 28178 6652
rect 28652 6659 28718 6668
rect 28652 6625 28668 6659
rect 28702 6625 28718 6659
rect 28652 6612 28718 6625
rect 28106 6596 28178 6600
rect 27248 6538 27294 6542
rect 27142 6530 27208 6538
rect 27376 6531 27422 6578
rect 26918 6491 27156 6500
rect 26918 6468 27110 6491
rect 26818 6442 26824 6459
rect 25576 6376 25648 6404
rect 26730 6378 26776 6425
rect 26806 6436 26824 6442
rect 26858 6442 26864 6459
rect 26916 6457 27110 6468
rect 27144 6457 27156 6491
rect 27376 6497 27382 6531
rect 27416 6497 27422 6531
rect 27376 6464 27422 6497
rect 26858 6436 26872 6442
rect 26806 6384 26812 6436
rect 26864 6384 26872 6436
rect 26806 6378 26872 6384
rect 26916 6440 27156 6457
rect 25264 6328 25354 6349
rect 25522 6331 25588 6340
rect 25522 6297 25538 6331
rect 25572 6297 25588 6331
rect 25522 6294 25588 6297
rect 25028 6266 25588 6294
rect 24932 6210 25000 6224
rect 24932 6176 24950 6210
rect 24984 6176 25000 6210
rect 24932 6166 25000 6176
rect 24972 5862 25000 6166
rect 25028 6084 25062 6266
rect 25360 6200 25432 6212
rect 25360 6148 25370 6200
rect 25422 6148 25432 6200
rect 25360 6136 25432 6148
rect 25284 6084 25348 6102
rect 25028 6050 25300 6084
rect 25334 6050 25348 6084
rect 25284 6040 25348 6050
rect 25620 6026 25648 6376
rect 25688 6342 25964 6372
rect 25688 6341 25720 6342
rect 25772 6341 25964 6342
rect 25688 6307 25717 6341
rect 25772 6307 25809 6341
rect 25843 6307 25901 6341
rect 25935 6307 25964 6341
rect 25688 6290 25720 6307
rect 25772 6290 25964 6307
rect 25688 6276 25964 6290
rect 26032 6348 26656 6366
rect 26032 6335 26574 6348
rect 26032 6301 26063 6335
rect 26097 6301 26155 6335
rect 26189 6301 26247 6335
rect 26281 6333 26574 6335
rect 26626 6333 26656 6348
rect 26281 6301 26409 6333
rect 26032 6299 26409 6301
rect 26443 6299 26501 6333
rect 26535 6299 26574 6333
rect 26627 6299 26656 6333
rect 26032 6296 26574 6299
rect 26626 6296 26656 6299
rect 25738 6084 25804 6090
rect 25738 6032 25744 6084
rect 25796 6032 25804 6084
rect 25738 6026 25804 6032
rect 25394 6012 25648 6026
rect 25150 6000 25196 6012
rect 24696 5834 25000 5862
rect 25116 5966 25156 6000
rect 25190 5966 25196 6000
rect 25116 5928 25196 5966
rect 25236 6006 25302 6012
rect 25236 5954 25242 6006
rect 25294 5954 25302 6006
rect 25236 5948 25302 5954
rect 25342 6000 25648 6012
rect 25342 5966 25348 6000
rect 25382 5998 25648 6000
rect 25382 5966 25444 5998
rect 25116 5894 25156 5928
rect 25190 5894 25196 5928
rect 25116 5882 25196 5894
rect 25246 5928 25292 5948
rect 25246 5894 25252 5928
rect 25286 5894 25292 5928
rect 25246 5882 25292 5894
rect 25342 5928 25444 5966
rect 25342 5894 25348 5928
rect 25382 5894 25444 5928
rect 25342 5882 25444 5894
rect 25564 5951 25798 5960
rect 25564 5899 25570 5951
rect 25622 5932 25746 5951
rect 25622 5899 25628 5932
rect 25564 5892 25628 5899
rect 25740 5899 25746 5932
rect 25798 5899 25804 5932
rect 25740 5892 25804 5899
rect 24696 5831 24972 5834
rect 24696 5797 24725 5831
rect 24759 5797 24817 5831
rect 24851 5797 24909 5831
rect 24943 5797 24972 5831
rect 24696 5766 24972 5797
rect 24802 5718 24866 5724
rect 24802 5666 24808 5718
rect 24860 5666 24866 5718
rect 24802 5660 24866 5666
rect 25116 5682 25162 5882
rect 25192 5844 25250 5854
rect 25192 5810 25204 5844
rect 25238 5810 25250 5844
rect 25192 5792 25250 5810
rect 25304 5763 25362 5780
rect 25304 5729 25316 5763
rect 25350 5729 25362 5763
rect 25304 5714 25362 5729
rect 25394 5682 25444 5882
rect 25510 5831 25786 5862
rect 25510 5797 25539 5831
rect 25573 5797 25631 5831
rect 25665 5797 25723 5831
rect 25757 5797 25786 5831
rect 25510 5766 25786 5797
rect 25116 5635 25212 5682
rect 24714 5602 24778 5608
rect 24714 5550 24720 5602
rect 24772 5550 24778 5602
rect 24714 5544 24778 5550
rect 24884 5592 24954 5610
rect 24884 5558 24905 5592
rect 24939 5558 24954 5592
rect 24884 5550 24954 5558
rect 25116 5601 25172 5635
rect 25206 5601 25212 5635
rect 25116 5563 25212 5601
rect 24884 5514 24912 5550
rect 25116 5529 25172 5563
rect 25206 5529 25212 5563
rect 25262 5635 25308 5682
rect 25262 5601 25268 5635
rect 25302 5601 25308 5635
rect 25262 5563 25308 5601
rect 25262 5542 25268 5563
rect 25116 5514 25212 5529
rect 24884 5482 25212 5514
rect 25252 5534 25268 5542
rect 25302 5542 25308 5563
rect 25358 5635 25444 5682
rect 25616 5716 25684 5726
rect 25616 5664 25624 5716
rect 25676 5664 25684 5716
rect 25616 5658 25684 5664
rect 25358 5601 25364 5635
rect 25398 5601 25444 5635
rect 25358 5563 25444 5601
rect 25302 5534 25318 5542
rect 25252 5482 25260 5534
rect 25312 5482 25318 5534
rect 25358 5529 25364 5563
rect 25398 5529 25444 5563
rect 25526 5604 25594 5610
rect 25526 5552 25532 5604
rect 25584 5552 25594 5604
rect 25526 5546 25594 5552
rect 25700 5590 25766 5602
rect 25700 5556 25717 5590
rect 25751 5556 25766 5590
rect 25700 5548 25766 5556
rect 25358 5510 25444 5529
rect 25738 5510 25766 5548
rect 25358 5482 25766 5510
rect 25252 5474 25318 5482
rect 25400 5478 25766 5482
rect 25204 5435 25266 5444
rect 25204 5401 25220 5435
rect 25254 5401 25266 5435
rect 25204 5384 25266 5401
rect 25208 5382 25266 5384
rect 25262 5327 25352 5348
rect 25262 5318 25289 5327
rect 23435 5293 25289 5318
rect 25323 5318 25352 5327
rect 25866 5318 25944 6276
rect 26032 6264 26656 6296
rect 26764 6331 26830 6342
rect 26764 6297 26780 6331
rect 26814 6297 26830 6331
rect 26764 6286 26830 6297
rect 26916 6294 26950 6440
rect 27098 6438 27156 6440
rect 27354 6459 27422 6464
rect 27354 6456 27382 6459
rect 27354 6404 27362 6456
rect 27416 6425 27422 6459
rect 27414 6404 27422 6425
rect 27152 6383 27242 6404
rect 27354 6398 27422 6404
rect 27152 6349 27179 6383
rect 27213 6349 27242 6383
rect 27376 6378 27422 6398
rect 27464 6531 27510 6578
rect 27464 6497 27470 6531
rect 27504 6497 27510 6531
rect 27464 6459 27510 6497
rect 27464 6425 27470 6459
rect 27504 6425 27510 6459
rect 27464 6404 27510 6425
rect 28618 6531 28664 6578
rect 28618 6497 28624 6531
rect 28658 6497 28664 6531
rect 28618 6459 28664 6497
rect 28618 6425 28624 6459
rect 28658 6425 28664 6459
rect 28706 6531 28752 6578
rect 28706 6497 28712 6531
rect 28746 6497 28752 6531
rect 28706 6459 28752 6497
rect 28806 6500 28866 6732
rect 28894 7022 28934 7056
rect 28968 7022 28974 7056
rect 28894 6984 28974 7022
rect 29014 7062 29080 7068
rect 29014 7010 29020 7062
rect 29072 7010 29080 7062
rect 29014 7004 29080 7010
rect 29120 7056 29222 7068
rect 29120 7022 29126 7056
rect 29160 7022 29222 7056
rect 28894 6950 28934 6984
rect 28968 6950 28974 6984
rect 28894 6938 28974 6950
rect 29024 6984 29070 7004
rect 29024 6950 29030 6984
rect 29064 6950 29070 6984
rect 29024 6938 29070 6950
rect 29120 6984 29222 7022
rect 29120 6950 29126 6984
rect 29160 6950 29222 6984
rect 29120 6938 29222 6950
rect 28894 6738 28940 6938
rect 28970 6900 29028 6910
rect 28970 6866 28982 6900
rect 29016 6866 29028 6900
rect 28970 6848 29028 6866
rect 29172 6858 29222 6938
rect 29588 6916 29672 7186
rect 29330 6906 29388 6912
rect 29322 6900 29396 6906
rect 29082 6819 29140 6836
rect 29082 6785 29094 6819
rect 29128 6785 29140 6819
rect 29082 6770 29140 6785
rect 29172 6792 29242 6858
rect 29322 6848 29333 6900
rect 29385 6848 29396 6900
rect 29322 6842 29396 6848
rect 29464 6890 29740 6916
rect 30334 6910 30432 7186
rect 29464 6885 29565 6890
rect 29617 6885 29740 6890
rect 29464 6851 29493 6885
rect 29527 6851 29565 6885
rect 29619 6851 29677 6885
rect 29711 6851 29740 6885
rect 29330 6834 29388 6842
rect 29464 6838 29565 6851
rect 29617 6838 29740 6851
rect 29464 6820 29740 6838
rect 29810 6879 30432 6910
rect 29810 6845 29839 6879
rect 29873 6845 29931 6879
rect 29965 6845 30023 6879
rect 30057 6877 30432 6879
rect 30057 6845 30185 6877
rect 29810 6843 30185 6845
rect 30219 6843 30277 6877
rect 30311 6843 30369 6877
rect 30403 6843 30432 6877
rect 30694 7140 31014 7158
rect 30694 7106 30966 7140
rect 31000 7106 31014 7140
rect 30694 7096 31014 7106
rect 29810 6812 30432 6843
rect 30572 6868 30648 6874
rect 30572 6816 30588 6868
rect 30640 6816 30648 6868
rect 30572 6810 30648 6816
rect 29172 6738 29222 6792
rect 30694 6766 30754 7096
rect 30816 7056 30862 7068
rect 28894 6691 28990 6738
rect 28894 6657 28950 6691
rect 28984 6657 28990 6691
rect 28894 6619 28990 6657
rect 28894 6585 28950 6619
rect 28984 6585 28990 6619
rect 29040 6691 29086 6738
rect 29040 6657 29046 6691
rect 29080 6657 29086 6691
rect 29040 6619 29086 6657
rect 29040 6598 29046 6619
rect 28894 6538 28990 6585
rect 29030 6590 29046 6598
rect 29080 6598 29086 6619
rect 29136 6691 29222 6738
rect 30226 6746 30754 6766
rect 30226 6712 30238 6746
rect 30272 6732 30754 6746
rect 30272 6712 30284 6732
rect 30226 6698 30284 6712
rect 29136 6657 29142 6691
rect 29176 6657 29222 6691
rect 29136 6619 29222 6657
rect 29080 6590 29096 6598
rect 29030 6538 29038 6590
rect 29090 6538 29096 6590
rect 29136 6585 29142 6619
rect 29176 6585 29222 6619
rect 29298 6659 29364 6672
rect 29298 6625 29314 6659
rect 29348 6625 29364 6659
rect 29692 6652 29760 6654
rect 29298 6614 29364 6625
rect 29608 6648 29760 6652
rect 29608 6642 29701 6648
rect 29608 6608 29628 6642
rect 29662 6608 29701 6642
rect 29608 6602 29701 6608
rect 29692 6596 29701 6602
rect 29753 6596 29760 6648
rect 29692 6590 29760 6596
rect 29796 6636 29870 6660
rect 29796 6602 29824 6636
rect 29858 6602 29870 6636
rect 29136 6542 29222 6585
rect 29796 6582 29870 6602
rect 29994 6652 30066 6664
rect 29994 6600 30005 6652
rect 30057 6600 30066 6652
rect 30540 6659 30606 6668
rect 30540 6625 30556 6659
rect 30590 6625 30606 6659
rect 30540 6612 30606 6625
rect 29994 6596 30066 6600
rect 29136 6538 29182 6542
rect 29030 6530 29096 6538
rect 29264 6531 29310 6578
rect 28806 6491 29044 6500
rect 28806 6468 28998 6491
rect 28706 6442 28712 6459
rect 27464 6376 27536 6404
rect 28618 6378 28664 6425
rect 28694 6436 28712 6442
rect 28746 6442 28752 6459
rect 28804 6457 28998 6468
rect 29032 6457 29044 6491
rect 29264 6497 29270 6531
rect 29304 6497 29310 6531
rect 29264 6464 29310 6497
rect 28746 6436 28760 6442
rect 28694 6384 28700 6436
rect 28752 6384 28760 6436
rect 28694 6378 28760 6384
rect 28804 6440 29044 6457
rect 27152 6328 27242 6349
rect 27410 6331 27476 6340
rect 27410 6297 27426 6331
rect 27460 6297 27476 6331
rect 27410 6294 27476 6297
rect 26916 6266 27476 6294
rect 26820 6210 26888 6224
rect 26820 6176 26838 6210
rect 26872 6176 26888 6210
rect 26820 6166 26888 6176
rect 26860 5862 26888 6166
rect 26916 6084 26950 6266
rect 27248 6200 27320 6212
rect 27248 6148 27258 6200
rect 27310 6148 27320 6200
rect 27248 6136 27320 6148
rect 27172 6084 27236 6102
rect 26916 6050 27188 6084
rect 27222 6050 27236 6084
rect 27172 6040 27236 6050
rect 27508 6026 27536 6376
rect 27576 6342 27852 6372
rect 27576 6341 27608 6342
rect 27660 6341 27852 6342
rect 27576 6307 27605 6341
rect 27660 6307 27697 6341
rect 27731 6307 27789 6341
rect 27823 6307 27852 6341
rect 27576 6290 27608 6307
rect 27660 6290 27852 6307
rect 27576 6276 27852 6290
rect 27920 6348 28544 6366
rect 27920 6335 28462 6348
rect 27920 6301 27951 6335
rect 27985 6301 28043 6335
rect 28077 6301 28135 6335
rect 28169 6333 28462 6335
rect 28514 6333 28544 6348
rect 28169 6301 28297 6333
rect 27920 6299 28297 6301
rect 28331 6299 28389 6333
rect 28423 6299 28462 6333
rect 28515 6299 28544 6333
rect 27920 6296 28462 6299
rect 28514 6296 28544 6299
rect 27626 6084 27692 6090
rect 27626 6032 27632 6084
rect 27684 6032 27692 6084
rect 27626 6026 27692 6032
rect 27282 6012 27536 6026
rect 27038 6000 27084 6012
rect 26584 5834 26888 5862
rect 27004 5966 27044 6000
rect 27078 5966 27084 6000
rect 27004 5928 27084 5966
rect 27124 6006 27190 6012
rect 27124 5954 27130 6006
rect 27182 5954 27190 6006
rect 27124 5948 27190 5954
rect 27230 6000 27536 6012
rect 27230 5966 27236 6000
rect 27270 5998 27536 6000
rect 27270 5966 27332 5998
rect 27004 5894 27044 5928
rect 27078 5894 27084 5928
rect 27004 5882 27084 5894
rect 27134 5928 27180 5948
rect 27134 5894 27140 5928
rect 27174 5894 27180 5928
rect 27134 5882 27180 5894
rect 27230 5928 27332 5966
rect 27230 5894 27236 5928
rect 27270 5894 27332 5928
rect 27230 5882 27332 5894
rect 27452 5951 27686 5960
rect 27452 5899 27458 5951
rect 27510 5932 27634 5951
rect 27510 5899 27516 5932
rect 27452 5892 27516 5899
rect 27628 5899 27634 5932
rect 27686 5899 27692 5932
rect 27628 5892 27692 5899
rect 26584 5831 26860 5834
rect 26584 5797 26613 5831
rect 26647 5797 26705 5831
rect 26739 5797 26797 5831
rect 26831 5797 26860 5831
rect 26584 5766 26860 5797
rect 26690 5718 26754 5724
rect 26690 5666 26696 5718
rect 26748 5666 26754 5718
rect 26690 5660 26754 5666
rect 27004 5682 27050 5882
rect 27080 5844 27138 5854
rect 27080 5810 27092 5844
rect 27126 5810 27138 5844
rect 27080 5792 27138 5810
rect 27192 5763 27250 5780
rect 27192 5729 27204 5763
rect 27238 5729 27250 5763
rect 27192 5714 27250 5729
rect 27282 5682 27332 5882
rect 27398 5831 27674 5862
rect 27398 5797 27427 5831
rect 27461 5797 27519 5831
rect 27553 5797 27611 5831
rect 27645 5797 27674 5831
rect 27398 5766 27674 5797
rect 27004 5635 27100 5682
rect 26602 5602 26666 5608
rect 26602 5550 26608 5602
rect 26660 5550 26666 5602
rect 26602 5544 26666 5550
rect 26772 5592 26842 5610
rect 26772 5558 26793 5592
rect 26827 5558 26842 5592
rect 26772 5550 26842 5558
rect 27004 5601 27060 5635
rect 27094 5601 27100 5635
rect 27004 5563 27100 5601
rect 26772 5514 26800 5550
rect 27004 5529 27060 5563
rect 27094 5529 27100 5563
rect 27150 5635 27196 5682
rect 27150 5601 27156 5635
rect 27190 5601 27196 5635
rect 27150 5563 27196 5601
rect 27150 5542 27156 5563
rect 27004 5514 27100 5529
rect 26772 5482 27100 5514
rect 27140 5534 27156 5542
rect 27190 5542 27196 5563
rect 27246 5635 27332 5682
rect 27504 5716 27572 5726
rect 27504 5664 27512 5716
rect 27564 5664 27572 5716
rect 27504 5658 27572 5664
rect 27246 5601 27252 5635
rect 27286 5601 27332 5635
rect 27246 5563 27332 5601
rect 27190 5534 27206 5542
rect 27140 5482 27148 5534
rect 27200 5482 27206 5534
rect 27246 5529 27252 5563
rect 27286 5529 27332 5563
rect 27414 5604 27482 5610
rect 27414 5552 27420 5604
rect 27472 5552 27482 5604
rect 27414 5546 27482 5552
rect 27588 5590 27654 5602
rect 27588 5556 27605 5590
rect 27639 5556 27654 5590
rect 27588 5548 27654 5556
rect 27246 5510 27332 5529
rect 27626 5510 27654 5548
rect 27246 5482 27654 5510
rect 27140 5474 27206 5482
rect 27288 5478 27654 5482
rect 27092 5435 27154 5444
rect 27092 5401 27108 5435
rect 27142 5401 27154 5435
rect 27092 5384 27154 5401
rect 27096 5382 27154 5384
rect 27150 5327 27240 5348
rect 27150 5318 27177 5327
rect 25323 5293 27177 5318
rect 27211 5318 27240 5327
rect 27754 5318 27832 6276
rect 27920 6264 28544 6296
rect 28652 6331 28718 6342
rect 28652 6297 28668 6331
rect 28702 6297 28718 6331
rect 28652 6286 28718 6297
rect 28804 6294 28838 6440
rect 28986 6438 29044 6440
rect 29242 6459 29310 6464
rect 29242 6456 29270 6459
rect 29242 6404 29250 6456
rect 29304 6425 29310 6459
rect 29302 6404 29310 6425
rect 29040 6383 29130 6404
rect 29242 6398 29310 6404
rect 29040 6349 29067 6383
rect 29101 6349 29130 6383
rect 29264 6378 29310 6398
rect 29352 6531 29398 6578
rect 29352 6497 29358 6531
rect 29392 6497 29398 6531
rect 29352 6459 29398 6497
rect 29352 6425 29358 6459
rect 29392 6425 29398 6459
rect 29352 6404 29398 6425
rect 30506 6531 30552 6578
rect 30506 6497 30512 6531
rect 30546 6497 30552 6531
rect 30506 6459 30552 6497
rect 30506 6425 30512 6459
rect 30546 6425 30552 6459
rect 30594 6531 30640 6578
rect 30594 6497 30600 6531
rect 30634 6497 30640 6531
rect 30594 6459 30640 6497
rect 30694 6500 30754 6732
rect 30782 7022 30822 7056
rect 30856 7022 30862 7056
rect 30782 6984 30862 7022
rect 30902 7062 30968 7068
rect 30902 7010 30908 7062
rect 30960 7010 30968 7062
rect 30902 7004 30968 7010
rect 31008 7056 31110 7068
rect 31008 7022 31014 7056
rect 31048 7022 31110 7056
rect 30782 6950 30822 6984
rect 30856 6950 30862 6984
rect 30782 6938 30862 6950
rect 30912 6984 30958 7004
rect 30912 6950 30918 6984
rect 30952 6950 30958 6984
rect 30912 6938 30958 6950
rect 31008 6984 31110 7022
rect 31008 6950 31014 6984
rect 31048 6950 31110 6984
rect 31008 6938 31110 6950
rect 30782 6738 30828 6938
rect 30858 6900 30916 6910
rect 30858 6866 30870 6900
rect 30904 6866 30916 6900
rect 30858 6848 30916 6866
rect 31060 6858 31110 6938
rect 31476 6916 31560 7186
rect 31218 6906 31276 6912
rect 31210 6900 31284 6906
rect 30970 6819 31028 6836
rect 30970 6785 30982 6819
rect 31016 6785 31028 6819
rect 30970 6770 31028 6785
rect 31060 6792 31130 6858
rect 31210 6848 31221 6900
rect 31273 6848 31284 6900
rect 31210 6842 31284 6848
rect 31352 6890 31628 6916
rect 32222 6910 32320 7186
rect 31352 6885 31453 6890
rect 31505 6885 31628 6890
rect 31352 6851 31381 6885
rect 31415 6851 31453 6885
rect 31507 6851 31565 6885
rect 31599 6851 31628 6885
rect 31218 6834 31276 6842
rect 31352 6838 31453 6851
rect 31505 6838 31628 6851
rect 31352 6820 31628 6838
rect 31698 6879 32320 6910
rect 31698 6845 31727 6879
rect 31761 6845 31819 6879
rect 31853 6845 31911 6879
rect 31945 6877 32320 6879
rect 31945 6845 32073 6877
rect 31698 6843 32073 6845
rect 32107 6843 32165 6877
rect 32199 6843 32257 6877
rect 32291 6843 32320 6877
rect 32582 7140 32902 7158
rect 32582 7106 32854 7140
rect 32888 7106 32902 7140
rect 32582 7096 32902 7106
rect 31698 6812 32320 6843
rect 32460 6868 32536 6874
rect 32460 6816 32476 6868
rect 32528 6816 32536 6868
rect 32460 6810 32536 6816
rect 31060 6738 31110 6792
rect 32582 6766 32642 7096
rect 32704 7056 32750 7068
rect 30782 6691 30878 6738
rect 30782 6657 30838 6691
rect 30872 6657 30878 6691
rect 30782 6619 30878 6657
rect 30782 6585 30838 6619
rect 30872 6585 30878 6619
rect 30928 6691 30974 6738
rect 30928 6657 30934 6691
rect 30968 6657 30974 6691
rect 30928 6619 30974 6657
rect 30928 6598 30934 6619
rect 30782 6538 30878 6585
rect 30918 6590 30934 6598
rect 30968 6598 30974 6619
rect 31024 6691 31110 6738
rect 32114 6746 32642 6766
rect 32114 6712 32126 6746
rect 32160 6732 32642 6746
rect 32160 6712 32172 6732
rect 32114 6698 32172 6712
rect 31024 6657 31030 6691
rect 31064 6657 31110 6691
rect 31024 6619 31110 6657
rect 30968 6590 30984 6598
rect 30918 6538 30926 6590
rect 30978 6538 30984 6590
rect 31024 6585 31030 6619
rect 31064 6585 31110 6619
rect 31186 6659 31252 6672
rect 31186 6625 31202 6659
rect 31236 6625 31252 6659
rect 31580 6652 31648 6654
rect 31186 6614 31252 6625
rect 31496 6648 31648 6652
rect 31496 6642 31589 6648
rect 31496 6608 31516 6642
rect 31550 6608 31589 6642
rect 31496 6602 31589 6608
rect 31580 6596 31589 6602
rect 31641 6596 31648 6648
rect 31580 6590 31648 6596
rect 31684 6636 31758 6660
rect 31684 6602 31712 6636
rect 31746 6602 31758 6636
rect 31024 6542 31110 6585
rect 31684 6582 31758 6602
rect 31882 6652 31954 6664
rect 31882 6600 31893 6652
rect 31945 6600 31954 6652
rect 32428 6659 32494 6668
rect 32428 6625 32444 6659
rect 32478 6625 32494 6659
rect 32428 6612 32494 6625
rect 31882 6596 31954 6600
rect 31024 6538 31070 6542
rect 30918 6530 30984 6538
rect 31152 6531 31198 6578
rect 30694 6491 30932 6500
rect 30694 6468 30886 6491
rect 30594 6442 30600 6459
rect 29352 6376 29424 6404
rect 30506 6378 30552 6425
rect 30582 6436 30600 6442
rect 30634 6442 30640 6459
rect 30692 6457 30886 6468
rect 30920 6457 30932 6491
rect 31152 6497 31158 6531
rect 31192 6497 31198 6531
rect 31152 6464 31198 6497
rect 30634 6436 30648 6442
rect 30582 6384 30588 6436
rect 30640 6384 30648 6436
rect 30582 6378 30648 6384
rect 30692 6440 30932 6457
rect 29040 6328 29130 6349
rect 29298 6331 29364 6340
rect 29298 6297 29314 6331
rect 29348 6297 29364 6331
rect 29298 6294 29364 6297
rect 28804 6266 29364 6294
rect 28708 6210 28776 6224
rect 28708 6176 28726 6210
rect 28760 6176 28776 6210
rect 28708 6166 28776 6176
rect 28748 5862 28776 6166
rect 28804 6084 28838 6266
rect 29136 6200 29208 6212
rect 29136 6148 29146 6200
rect 29198 6148 29208 6200
rect 29136 6136 29208 6148
rect 29060 6084 29124 6102
rect 28804 6050 29076 6084
rect 29110 6050 29124 6084
rect 29060 6040 29124 6050
rect 29396 6026 29424 6376
rect 29464 6342 29740 6372
rect 29464 6341 29496 6342
rect 29548 6341 29740 6342
rect 29464 6307 29493 6341
rect 29548 6307 29585 6341
rect 29619 6307 29677 6341
rect 29711 6307 29740 6341
rect 29464 6290 29496 6307
rect 29548 6290 29740 6307
rect 29464 6276 29740 6290
rect 29808 6348 30432 6366
rect 29808 6335 30350 6348
rect 29808 6301 29839 6335
rect 29873 6301 29931 6335
rect 29965 6301 30023 6335
rect 30057 6333 30350 6335
rect 30402 6333 30432 6348
rect 30057 6301 30185 6333
rect 29808 6299 30185 6301
rect 30219 6299 30277 6333
rect 30311 6299 30350 6333
rect 30403 6299 30432 6333
rect 29808 6296 30350 6299
rect 30402 6296 30432 6299
rect 29514 6084 29580 6090
rect 29514 6032 29520 6084
rect 29572 6032 29580 6084
rect 29514 6026 29580 6032
rect 29170 6012 29424 6026
rect 28926 6000 28972 6012
rect 28472 5834 28776 5862
rect 28892 5966 28932 6000
rect 28966 5966 28972 6000
rect 28892 5928 28972 5966
rect 29012 6006 29078 6012
rect 29012 5954 29018 6006
rect 29070 5954 29078 6006
rect 29012 5948 29078 5954
rect 29118 6000 29424 6012
rect 29118 5966 29124 6000
rect 29158 5998 29424 6000
rect 29158 5966 29220 5998
rect 28892 5894 28932 5928
rect 28966 5894 28972 5928
rect 28892 5882 28972 5894
rect 29022 5928 29068 5948
rect 29022 5894 29028 5928
rect 29062 5894 29068 5928
rect 29022 5882 29068 5894
rect 29118 5928 29220 5966
rect 29118 5894 29124 5928
rect 29158 5894 29220 5928
rect 29118 5882 29220 5894
rect 29340 5951 29574 5960
rect 29340 5899 29346 5951
rect 29398 5932 29522 5951
rect 29398 5899 29404 5932
rect 29340 5892 29404 5899
rect 29516 5899 29522 5932
rect 29574 5899 29580 5932
rect 29516 5892 29580 5899
rect 28472 5831 28748 5834
rect 28472 5797 28501 5831
rect 28535 5797 28593 5831
rect 28627 5797 28685 5831
rect 28719 5797 28748 5831
rect 28472 5766 28748 5797
rect 28578 5718 28642 5724
rect 28578 5666 28584 5718
rect 28636 5666 28642 5718
rect 28578 5660 28642 5666
rect 28892 5682 28938 5882
rect 28968 5844 29026 5854
rect 28968 5810 28980 5844
rect 29014 5810 29026 5844
rect 28968 5792 29026 5810
rect 29080 5763 29138 5780
rect 29080 5729 29092 5763
rect 29126 5729 29138 5763
rect 29080 5714 29138 5729
rect 29170 5682 29220 5882
rect 29286 5831 29562 5862
rect 29286 5797 29315 5831
rect 29349 5797 29407 5831
rect 29441 5797 29499 5831
rect 29533 5797 29562 5831
rect 29286 5766 29562 5797
rect 28892 5635 28988 5682
rect 28490 5602 28554 5608
rect 28490 5550 28496 5602
rect 28548 5550 28554 5602
rect 28490 5544 28554 5550
rect 28660 5592 28730 5610
rect 28660 5558 28681 5592
rect 28715 5558 28730 5592
rect 28660 5550 28730 5558
rect 28892 5601 28948 5635
rect 28982 5601 28988 5635
rect 28892 5563 28988 5601
rect 28660 5514 28688 5550
rect 28892 5529 28948 5563
rect 28982 5529 28988 5563
rect 29038 5635 29084 5682
rect 29038 5601 29044 5635
rect 29078 5601 29084 5635
rect 29038 5563 29084 5601
rect 29038 5542 29044 5563
rect 28892 5514 28988 5529
rect 28660 5482 28988 5514
rect 29028 5534 29044 5542
rect 29078 5542 29084 5563
rect 29134 5635 29220 5682
rect 29392 5716 29460 5726
rect 29392 5664 29400 5716
rect 29452 5664 29460 5716
rect 29392 5658 29460 5664
rect 29134 5601 29140 5635
rect 29174 5601 29220 5635
rect 29134 5563 29220 5601
rect 29078 5534 29094 5542
rect 29028 5482 29036 5534
rect 29088 5482 29094 5534
rect 29134 5529 29140 5563
rect 29174 5529 29220 5563
rect 29302 5604 29370 5610
rect 29302 5552 29308 5604
rect 29360 5552 29370 5604
rect 29302 5546 29370 5552
rect 29476 5590 29542 5602
rect 29476 5556 29493 5590
rect 29527 5556 29542 5590
rect 29476 5548 29542 5556
rect 29134 5510 29220 5529
rect 29514 5510 29542 5548
rect 29134 5482 29542 5510
rect 29028 5474 29094 5482
rect 29176 5478 29542 5482
rect 28980 5435 29042 5444
rect 28980 5401 28996 5435
rect 29030 5401 29042 5435
rect 28980 5384 29042 5401
rect 28984 5382 29042 5384
rect 29038 5327 29128 5348
rect 29038 5318 29065 5327
rect 27211 5293 29065 5318
rect 29099 5318 29128 5327
rect 29642 5318 29720 6276
rect 29808 6264 30432 6296
rect 30540 6331 30606 6342
rect 30540 6297 30556 6331
rect 30590 6297 30606 6331
rect 30540 6286 30606 6297
rect 30692 6294 30726 6440
rect 30874 6438 30932 6440
rect 31130 6459 31198 6464
rect 31130 6456 31158 6459
rect 31130 6404 31138 6456
rect 31192 6425 31198 6459
rect 31190 6404 31198 6425
rect 30928 6383 31018 6404
rect 31130 6398 31198 6404
rect 30928 6349 30955 6383
rect 30989 6349 31018 6383
rect 31152 6378 31198 6398
rect 31240 6531 31286 6578
rect 31240 6497 31246 6531
rect 31280 6497 31286 6531
rect 31240 6459 31286 6497
rect 31240 6425 31246 6459
rect 31280 6425 31286 6459
rect 31240 6404 31286 6425
rect 32394 6531 32440 6578
rect 32394 6497 32400 6531
rect 32434 6497 32440 6531
rect 32394 6459 32440 6497
rect 32394 6425 32400 6459
rect 32434 6425 32440 6459
rect 32482 6531 32528 6578
rect 32482 6497 32488 6531
rect 32522 6497 32528 6531
rect 32482 6459 32528 6497
rect 32582 6500 32642 6732
rect 32670 7022 32710 7056
rect 32744 7022 32750 7056
rect 32670 6984 32750 7022
rect 32790 7062 32856 7068
rect 32790 7010 32796 7062
rect 32848 7010 32856 7062
rect 32790 7004 32856 7010
rect 32896 7056 32998 7068
rect 32896 7022 32902 7056
rect 32936 7022 32998 7056
rect 32670 6950 32710 6984
rect 32744 6950 32750 6984
rect 32670 6938 32750 6950
rect 32800 6984 32846 7004
rect 32800 6950 32806 6984
rect 32840 6950 32846 6984
rect 32800 6938 32846 6950
rect 32896 6984 32998 7022
rect 32896 6950 32902 6984
rect 32936 6950 32998 6984
rect 32896 6938 32998 6950
rect 32670 6738 32716 6938
rect 32746 6900 32804 6910
rect 32746 6866 32758 6900
rect 32792 6866 32804 6900
rect 32746 6848 32804 6866
rect 32948 6858 32998 6938
rect 33364 6916 33448 7186
rect 33106 6906 33164 6912
rect 33098 6900 33172 6906
rect 32858 6819 32916 6836
rect 32858 6785 32870 6819
rect 32904 6785 32916 6819
rect 32858 6770 32916 6785
rect 32948 6792 33018 6858
rect 33098 6848 33109 6900
rect 33161 6848 33172 6900
rect 33098 6842 33172 6848
rect 33240 6890 33516 6916
rect 34110 6910 34208 7186
rect 33240 6885 33341 6890
rect 33393 6885 33516 6890
rect 33240 6851 33269 6885
rect 33303 6851 33341 6885
rect 33395 6851 33453 6885
rect 33487 6851 33516 6885
rect 33106 6834 33164 6842
rect 33240 6838 33341 6851
rect 33393 6838 33516 6851
rect 33240 6820 33516 6838
rect 33586 6879 34208 6910
rect 33586 6845 33615 6879
rect 33649 6845 33707 6879
rect 33741 6845 33799 6879
rect 33833 6877 34208 6879
rect 33833 6845 33961 6877
rect 33586 6843 33961 6845
rect 33995 6843 34053 6877
rect 34087 6843 34145 6877
rect 34179 6843 34208 6877
rect 34470 7140 34790 7158
rect 34470 7106 34742 7140
rect 34776 7106 34790 7140
rect 34470 7096 34790 7106
rect 33586 6812 34208 6843
rect 34348 6868 34424 6874
rect 34348 6816 34364 6868
rect 34416 6816 34424 6868
rect 34348 6810 34424 6816
rect 32948 6738 32998 6792
rect 34470 6766 34530 7096
rect 34592 7056 34638 7068
rect 32670 6691 32766 6738
rect 32670 6657 32726 6691
rect 32760 6657 32766 6691
rect 32670 6619 32766 6657
rect 32670 6585 32726 6619
rect 32760 6585 32766 6619
rect 32816 6691 32862 6738
rect 32816 6657 32822 6691
rect 32856 6657 32862 6691
rect 32816 6619 32862 6657
rect 32816 6598 32822 6619
rect 32670 6538 32766 6585
rect 32806 6590 32822 6598
rect 32856 6598 32862 6619
rect 32912 6691 32998 6738
rect 34002 6746 34530 6766
rect 34002 6712 34014 6746
rect 34048 6732 34530 6746
rect 34048 6712 34060 6732
rect 34002 6698 34060 6712
rect 32912 6657 32918 6691
rect 32952 6657 32998 6691
rect 32912 6619 32998 6657
rect 32856 6590 32872 6598
rect 32806 6538 32814 6590
rect 32866 6538 32872 6590
rect 32912 6585 32918 6619
rect 32952 6585 32998 6619
rect 33074 6659 33140 6672
rect 33074 6625 33090 6659
rect 33124 6625 33140 6659
rect 33468 6652 33536 6654
rect 33074 6614 33140 6625
rect 33384 6648 33536 6652
rect 33384 6642 33477 6648
rect 33384 6608 33404 6642
rect 33438 6608 33477 6642
rect 33384 6602 33477 6608
rect 33468 6596 33477 6602
rect 33529 6596 33536 6648
rect 33468 6590 33536 6596
rect 33572 6636 33646 6660
rect 33572 6602 33600 6636
rect 33634 6602 33646 6636
rect 32912 6542 32998 6585
rect 33572 6582 33646 6602
rect 33770 6652 33842 6664
rect 33770 6600 33781 6652
rect 33833 6600 33842 6652
rect 34316 6659 34382 6668
rect 34316 6625 34332 6659
rect 34366 6625 34382 6659
rect 34316 6612 34382 6625
rect 33770 6596 33842 6600
rect 32912 6538 32958 6542
rect 32806 6530 32872 6538
rect 33040 6531 33086 6578
rect 32582 6491 32820 6500
rect 32582 6468 32774 6491
rect 32482 6442 32488 6459
rect 31240 6376 31312 6404
rect 32394 6378 32440 6425
rect 32470 6436 32488 6442
rect 32522 6442 32528 6459
rect 32580 6457 32774 6468
rect 32808 6457 32820 6491
rect 33040 6497 33046 6531
rect 33080 6497 33086 6531
rect 33040 6464 33086 6497
rect 32522 6436 32536 6442
rect 32470 6384 32476 6436
rect 32528 6384 32536 6436
rect 32470 6378 32536 6384
rect 32580 6440 32820 6457
rect 30928 6328 31018 6349
rect 31186 6331 31252 6340
rect 31186 6297 31202 6331
rect 31236 6297 31252 6331
rect 31186 6294 31252 6297
rect 30692 6266 31252 6294
rect 30596 6210 30664 6224
rect 30596 6176 30614 6210
rect 30648 6176 30664 6210
rect 30596 6166 30664 6176
rect 30636 5862 30664 6166
rect 30692 6084 30726 6266
rect 31024 6200 31096 6212
rect 31024 6148 31034 6200
rect 31086 6148 31096 6200
rect 31024 6136 31096 6148
rect 30948 6084 31012 6102
rect 30692 6050 30964 6084
rect 30998 6050 31012 6084
rect 30948 6040 31012 6050
rect 31284 6026 31312 6376
rect 31352 6342 31628 6372
rect 31352 6341 31384 6342
rect 31436 6341 31628 6342
rect 31352 6307 31381 6341
rect 31436 6307 31473 6341
rect 31507 6307 31565 6341
rect 31599 6307 31628 6341
rect 31352 6290 31384 6307
rect 31436 6290 31628 6307
rect 31352 6276 31628 6290
rect 31696 6348 32320 6366
rect 31696 6335 32238 6348
rect 31696 6301 31727 6335
rect 31761 6301 31819 6335
rect 31853 6301 31911 6335
rect 31945 6333 32238 6335
rect 32290 6333 32320 6348
rect 31945 6301 32073 6333
rect 31696 6299 32073 6301
rect 32107 6299 32165 6333
rect 32199 6299 32238 6333
rect 32291 6299 32320 6333
rect 31696 6296 32238 6299
rect 32290 6296 32320 6299
rect 31402 6084 31468 6090
rect 31402 6032 31408 6084
rect 31460 6032 31468 6084
rect 31402 6026 31468 6032
rect 31058 6012 31312 6026
rect 30814 6000 30860 6012
rect 30360 5834 30664 5862
rect 30780 5966 30820 6000
rect 30854 5966 30860 6000
rect 30780 5928 30860 5966
rect 30900 6006 30966 6012
rect 30900 5954 30906 6006
rect 30958 5954 30966 6006
rect 30900 5948 30966 5954
rect 31006 6000 31312 6012
rect 31006 5966 31012 6000
rect 31046 5998 31312 6000
rect 31046 5966 31108 5998
rect 30780 5894 30820 5928
rect 30854 5894 30860 5928
rect 30780 5882 30860 5894
rect 30910 5928 30956 5948
rect 30910 5894 30916 5928
rect 30950 5894 30956 5928
rect 30910 5882 30956 5894
rect 31006 5928 31108 5966
rect 31006 5894 31012 5928
rect 31046 5894 31108 5928
rect 31006 5882 31108 5894
rect 31228 5951 31462 5960
rect 31228 5899 31234 5951
rect 31286 5932 31410 5951
rect 31286 5899 31292 5932
rect 31228 5892 31292 5899
rect 31404 5899 31410 5932
rect 31462 5899 31468 5932
rect 31404 5892 31468 5899
rect 30360 5831 30636 5834
rect 30360 5797 30389 5831
rect 30423 5797 30481 5831
rect 30515 5797 30573 5831
rect 30607 5797 30636 5831
rect 30360 5766 30636 5797
rect 30466 5718 30530 5724
rect 30466 5666 30472 5718
rect 30524 5666 30530 5718
rect 30466 5660 30530 5666
rect 30780 5682 30826 5882
rect 30856 5844 30914 5854
rect 30856 5810 30868 5844
rect 30902 5810 30914 5844
rect 30856 5792 30914 5810
rect 30968 5763 31026 5780
rect 30968 5729 30980 5763
rect 31014 5729 31026 5763
rect 30968 5714 31026 5729
rect 31058 5682 31108 5882
rect 31174 5831 31450 5862
rect 31174 5797 31203 5831
rect 31237 5797 31295 5831
rect 31329 5797 31387 5831
rect 31421 5797 31450 5831
rect 31174 5766 31450 5797
rect 30780 5635 30876 5682
rect 30378 5602 30442 5608
rect 30378 5550 30384 5602
rect 30436 5550 30442 5602
rect 30378 5544 30442 5550
rect 30548 5592 30618 5610
rect 30548 5558 30569 5592
rect 30603 5558 30618 5592
rect 30548 5550 30618 5558
rect 30780 5601 30836 5635
rect 30870 5601 30876 5635
rect 30780 5563 30876 5601
rect 30548 5514 30576 5550
rect 30780 5529 30836 5563
rect 30870 5529 30876 5563
rect 30926 5635 30972 5682
rect 30926 5601 30932 5635
rect 30966 5601 30972 5635
rect 30926 5563 30972 5601
rect 30926 5542 30932 5563
rect 30780 5514 30876 5529
rect 30548 5482 30876 5514
rect 30916 5534 30932 5542
rect 30966 5542 30972 5563
rect 31022 5635 31108 5682
rect 31280 5716 31348 5726
rect 31280 5664 31288 5716
rect 31340 5664 31348 5716
rect 31280 5658 31348 5664
rect 31022 5601 31028 5635
rect 31062 5601 31108 5635
rect 31022 5563 31108 5601
rect 30966 5534 30982 5542
rect 30916 5482 30924 5534
rect 30976 5482 30982 5534
rect 31022 5529 31028 5563
rect 31062 5529 31108 5563
rect 31190 5604 31258 5610
rect 31190 5552 31196 5604
rect 31248 5552 31258 5604
rect 31190 5546 31258 5552
rect 31364 5590 31430 5602
rect 31364 5556 31381 5590
rect 31415 5556 31430 5590
rect 31364 5548 31430 5556
rect 31022 5510 31108 5529
rect 31402 5510 31430 5548
rect 31022 5482 31430 5510
rect 30916 5474 30982 5482
rect 31064 5478 31430 5482
rect 30868 5435 30930 5444
rect 30868 5401 30884 5435
rect 30918 5401 30930 5435
rect 30868 5384 30930 5401
rect 30872 5382 30930 5384
rect 30926 5327 31016 5348
rect 30926 5318 30953 5327
rect 29099 5293 30953 5318
rect 30987 5318 31016 5327
rect 31530 5318 31608 6276
rect 31696 6264 32320 6296
rect 32428 6331 32494 6342
rect 32428 6297 32444 6331
rect 32478 6297 32494 6331
rect 32428 6286 32494 6297
rect 32580 6294 32614 6440
rect 32762 6438 32820 6440
rect 33018 6459 33086 6464
rect 33018 6456 33046 6459
rect 33018 6404 33026 6456
rect 33080 6425 33086 6459
rect 33078 6404 33086 6425
rect 32816 6383 32906 6404
rect 33018 6398 33086 6404
rect 32816 6349 32843 6383
rect 32877 6349 32906 6383
rect 33040 6378 33086 6398
rect 33128 6531 33174 6578
rect 33128 6497 33134 6531
rect 33168 6497 33174 6531
rect 33128 6459 33174 6497
rect 33128 6425 33134 6459
rect 33168 6425 33174 6459
rect 33128 6404 33174 6425
rect 34282 6531 34328 6578
rect 34282 6497 34288 6531
rect 34322 6497 34328 6531
rect 34282 6459 34328 6497
rect 34282 6425 34288 6459
rect 34322 6425 34328 6459
rect 34370 6531 34416 6578
rect 34370 6497 34376 6531
rect 34410 6497 34416 6531
rect 34370 6459 34416 6497
rect 34470 6500 34530 6732
rect 34558 7022 34598 7056
rect 34632 7022 34638 7056
rect 34558 6984 34638 7022
rect 34678 7062 34744 7068
rect 34678 7010 34684 7062
rect 34736 7010 34744 7062
rect 34678 7004 34744 7010
rect 34784 7056 34886 7068
rect 34784 7022 34790 7056
rect 34824 7022 34886 7056
rect 34558 6950 34598 6984
rect 34632 6950 34638 6984
rect 34558 6938 34638 6950
rect 34688 6984 34734 7004
rect 34688 6950 34694 6984
rect 34728 6950 34734 6984
rect 34688 6938 34734 6950
rect 34784 6984 34886 7022
rect 34784 6950 34790 6984
rect 34824 6950 34886 6984
rect 34784 6938 34886 6950
rect 34558 6738 34604 6938
rect 34634 6900 34692 6910
rect 34634 6866 34646 6900
rect 34680 6866 34692 6900
rect 34634 6848 34692 6866
rect 34836 6858 34886 6938
rect 35252 6916 35336 7186
rect 34994 6906 35052 6912
rect 34986 6900 35060 6906
rect 34746 6819 34804 6836
rect 34746 6785 34758 6819
rect 34792 6785 34804 6819
rect 34746 6770 34804 6785
rect 34836 6792 34906 6858
rect 34986 6848 34997 6900
rect 35049 6848 35060 6900
rect 34986 6842 35060 6848
rect 35128 6890 35404 6916
rect 35998 6910 36096 7186
rect 35128 6885 35229 6890
rect 35281 6885 35404 6890
rect 35128 6851 35157 6885
rect 35191 6851 35229 6885
rect 35283 6851 35341 6885
rect 35375 6851 35404 6885
rect 34994 6834 35052 6842
rect 35128 6838 35229 6851
rect 35281 6838 35404 6851
rect 35128 6820 35404 6838
rect 35474 6879 36096 6910
rect 35474 6845 35503 6879
rect 35537 6845 35595 6879
rect 35629 6845 35687 6879
rect 35721 6877 36096 6879
rect 35721 6845 35849 6877
rect 35474 6843 35849 6845
rect 35883 6843 35941 6877
rect 35975 6843 36033 6877
rect 36067 6843 36096 6877
rect 36358 7140 36678 7158
rect 36358 7106 36630 7140
rect 36664 7106 36678 7140
rect 36358 7096 36678 7106
rect 35474 6812 36096 6843
rect 36236 6868 36312 6874
rect 36236 6816 36252 6868
rect 36304 6816 36312 6868
rect 36236 6810 36312 6816
rect 34836 6738 34886 6792
rect 36358 6766 36418 7096
rect 36480 7056 36526 7068
rect 34558 6691 34654 6738
rect 34558 6657 34614 6691
rect 34648 6657 34654 6691
rect 34558 6619 34654 6657
rect 34558 6585 34614 6619
rect 34648 6585 34654 6619
rect 34704 6691 34750 6738
rect 34704 6657 34710 6691
rect 34744 6657 34750 6691
rect 34704 6619 34750 6657
rect 34704 6598 34710 6619
rect 34558 6538 34654 6585
rect 34694 6590 34710 6598
rect 34744 6598 34750 6619
rect 34800 6691 34886 6738
rect 35890 6746 36418 6766
rect 35890 6712 35902 6746
rect 35936 6732 36418 6746
rect 35936 6712 35948 6732
rect 35890 6698 35948 6712
rect 34800 6657 34806 6691
rect 34840 6657 34886 6691
rect 34800 6619 34886 6657
rect 34744 6590 34760 6598
rect 34694 6538 34702 6590
rect 34754 6538 34760 6590
rect 34800 6585 34806 6619
rect 34840 6585 34886 6619
rect 34962 6659 35028 6672
rect 34962 6625 34978 6659
rect 35012 6625 35028 6659
rect 35356 6652 35424 6654
rect 34962 6614 35028 6625
rect 35272 6648 35424 6652
rect 35272 6642 35365 6648
rect 35272 6608 35292 6642
rect 35326 6608 35365 6642
rect 35272 6602 35365 6608
rect 35356 6596 35365 6602
rect 35417 6596 35424 6648
rect 35356 6590 35424 6596
rect 35460 6636 35534 6660
rect 35460 6602 35488 6636
rect 35522 6602 35534 6636
rect 34800 6542 34886 6585
rect 35460 6582 35534 6602
rect 35658 6652 35730 6664
rect 35658 6600 35669 6652
rect 35721 6600 35730 6652
rect 36204 6659 36270 6668
rect 36204 6625 36220 6659
rect 36254 6625 36270 6659
rect 36204 6612 36270 6625
rect 35658 6596 35730 6600
rect 34800 6538 34846 6542
rect 34694 6530 34760 6538
rect 34928 6531 34974 6578
rect 34470 6491 34708 6500
rect 34470 6468 34662 6491
rect 34370 6442 34376 6459
rect 33128 6376 33200 6404
rect 34282 6378 34328 6425
rect 34358 6436 34376 6442
rect 34410 6442 34416 6459
rect 34468 6457 34662 6468
rect 34696 6457 34708 6491
rect 34928 6497 34934 6531
rect 34968 6497 34974 6531
rect 34928 6464 34974 6497
rect 34410 6436 34424 6442
rect 34358 6384 34364 6436
rect 34416 6384 34424 6436
rect 34358 6378 34424 6384
rect 34468 6440 34708 6457
rect 32816 6328 32906 6349
rect 33074 6331 33140 6340
rect 33074 6297 33090 6331
rect 33124 6297 33140 6331
rect 33074 6294 33140 6297
rect 32580 6266 33140 6294
rect 32484 6210 32552 6224
rect 32484 6176 32502 6210
rect 32536 6176 32552 6210
rect 32484 6166 32552 6176
rect 32524 5862 32552 6166
rect 32580 6084 32614 6266
rect 32912 6200 32984 6212
rect 32912 6148 32922 6200
rect 32974 6148 32984 6200
rect 32912 6136 32984 6148
rect 32836 6084 32900 6102
rect 32580 6050 32852 6084
rect 32886 6050 32900 6084
rect 32836 6040 32900 6050
rect 33172 6026 33200 6376
rect 33240 6342 33516 6372
rect 33240 6341 33272 6342
rect 33324 6341 33516 6342
rect 33240 6307 33269 6341
rect 33324 6307 33361 6341
rect 33395 6307 33453 6341
rect 33487 6307 33516 6341
rect 33240 6290 33272 6307
rect 33324 6290 33516 6307
rect 33240 6276 33516 6290
rect 33584 6348 34208 6366
rect 33584 6335 34126 6348
rect 33584 6301 33615 6335
rect 33649 6301 33707 6335
rect 33741 6301 33799 6335
rect 33833 6333 34126 6335
rect 34178 6333 34208 6348
rect 33833 6301 33961 6333
rect 33584 6299 33961 6301
rect 33995 6299 34053 6333
rect 34087 6299 34126 6333
rect 34179 6299 34208 6333
rect 33584 6296 34126 6299
rect 34178 6296 34208 6299
rect 33290 6084 33356 6090
rect 33290 6032 33296 6084
rect 33348 6032 33356 6084
rect 33290 6026 33356 6032
rect 32946 6012 33200 6026
rect 32702 6000 32748 6012
rect 32248 5834 32552 5862
rect 32668 5966 32708 6000
rect 32742 5966 32748 6000
rect 32668 5928 32748 5966
rect 32788 6006 32854 6012
rect 32788 5954 32794 6006
rect 32846 5954 32854 6006
rect 32788 5948 32854 5954
rect 32894 6000 33200 6012
rect 32894 5966 32900 6000
rect 32934 5998 33200 6000
rect 32934 5966 32996 5998
rect 32668 5894 32708 5928
rect 32742 5894 32748 5928
rect 32668 5882 32748 5894
rect 32798 5928 32844 5948
rect 32798 5894 32804 5928
rect 32838 5894 32844 5928
rect 32798 5882 32844 5894
rect 32894 5928 32996 5966
rect 32894 5894 32900 5928
rect 32934 5894 32996 5928
rect 32894 5882 32996 5894
rect 33116 5951 33350 5960
rect 33116 5899 33122 5951
rect 33174 5932 33298 5951
rect 33174 5899 33180 5932
rect 33116 5892 33180 5899
rect 33292 5899 33298 5932
rect 33350 5899 33356 5932
rect 33292 5892 33356 5899
rect 32248 5831 32524 5834
rect 32248 5797 32277 5831
rect 32311 5797 32369 5831
rect 32403 5797 32461 5831
rect 32495 5797 32524 5831
rect 32248 5766 32524 5797
rect 32354 5718 32418 5724
rect 32354 5666 32360 5718
rect 32412 5666 32418 5718
rect 32354 5660 32418 5666
rect 32668 5682 32714 5882
rect 32744 5844 32802 5854
rect 32744 5810 32756 5844
rect 32790 5810 32802 5844
rect 32744 5792 32802 5810
rect 32856 5763 32914 5780
rect 32856 5729 32868 5763
rect 32902 5729 32914 5763
rect 32856 5714 32914 5729
rect 32946 5682 32996 5882
rect 33062 5831 33338 5862
rect 33062 5797 33091 5831
rect 33125 5797 33183 5831
rect 33217 5797 33275 5831
rect 33309 5797 33338 5831
rect 33062 5766 33338 5797
rect 32668 5635 32764 5682
rect 32266 5602 32330 5608
rect 32266 5550 32272 5602
rect 32324 5550 32330 5602
rect 32266 5544 32330 5550
rect 32436 5592 32506 5610
rect 32436 5558 32457 5592
rect 32491 5558 32506 5592
rect 32436 5550 32506 5558
rect 32668 5601 32724 5635
rect 32758 5601 32764 5635
rect 32668 5563 32764 5601
rect 32436 5514 32464 5550
rect 32668 5529 32724 5563
rect 32758 5529 32764 5563
rect 32814 5635 32860 5682
rect 32814 5601 32820 5635
rect 32854 5601 32860 5635
rect 32814 5563 32860 5601
rect 32814 5542 32820 5563
rect 32668 5514 32764 5529
rect 32436 5482 32764 5514
rect 32804 5534 32820 5542
rect 32854 5542 32860 5563
rect 32910 5635 32996 5682
rect 33168 5716 33236 5726
rect 33168 5664 33176 5716
rect 33228 5664 33236 5716
rect 33168 5658 33236 5664
rect 32910 5601 32916 5635
rect 32950 5601 32996 5635
rect 32910 5563 32996 5601
rect 32854 5534 32870 5542
rect 32804 5482 32812 5534
rect 32864 5482 32870 5534
rect 32910 5529 32916 5563
rect 32950 5529 32996 5563
rect 33078 5604 33146 5610
rect 33078 5552 33084 5604
rect 33136 5552 33146 5604
rect 33078 5546 33146 5552
rect 33252 5590 33318 5602
rect 33252 5556 33269 5590
rect 33303 5556 33318 5590
rect 33252 5548 33318 5556
rect 32910 5510 32996 5529
rect 33290 5510 33318 5548
rect 32910 5482 33318 5510
rect 32804 5474 32870 5482
rect 32952 5478 33318 5482
rect 32756 5435 32818 5444
rect 32756 5401 32772 5435
rect 32806 5401 32818 5435
rect 32756 5384 32818 5401
rect 32760 5382 32818 5384
rect 32814 5327 32904 5348
rect 32814 5318 32841 5327
rect 30987 5293 32841 5318
rect 32875 5318 32904 5327
rect 33418 5318 33496 6276
rect 33584 6264 34208 6296
rect 34316 6331 34382 6342
rect 34316 6297 34332 6331
rect 34366 6297 34382 6331
rect 34316 6286 34382 6297
rect 34468 6294 34502 6440
rect 34650 6438 34708 6440
rect 34906 6459 34974 6464
rect 34906 6456 34934 6459
rect 34906 6404 34914 6456
rect 34968 6425 34974 6459
rect 34966 6404 34974 6425
rect 34704 6383 34794 6404
rect 34906 6398 34974 6404
rect 34704 6349 34731 6383
rect 34765 6349 34794 6383
rect 34928 6378 34974 6398
rect 35016 6531 35062 6578
rect 35016 6497 35022 6531
rect 35056 6497 35062 6531
rect 35016 6459 35062 6497
rect 35016 6425 35022 6459
rect 35056 6425 35062 6459
rect 35016 6404 35062 6425
rect 36170 6531 36216 6578
rect 36170 6497 36176 6531
rect 36210 6497 36216 6531
rect 36170 6459 36216 6497
rect 36170 6425 36176 6459
rect 36210 6425 36216 6459
rect 36258 6531 36304 6578
rect 36258 6497 36264 6531
rect 36298 6497 36304 6531
rect 36258 6459 36304 6497
rect 36358 6500 36418 6732
rect 36446 7022 36486 7056
rect 36520 7022 36526 7056
rect 36446 6984 36526 7022
rect 36566 7062 36632 7068
rect 36566 7010 36572 7062
rect 36624 7010 36632 7062
rect 36566 7004 36632 7010
rect 36672 7056 36774 7068
rect 36672 7022 36678 7056
rect 36712 7022 36774 7056
rect 36446 6950 36486 6984
rect 36520 6950 36526 6984
rect 36446 6938 36526 6950
rect 36576 6984 36622 7004
rect 36576 6950 36582 6984
rect 36616 6950 36622 6984
rect 36576 6938 36622 6950
rect 36672 6984 36774 7022
rect 36672 6950 36678 6984
rect 36712 6950 36774 6984
rect 36672 6938 36774 6950
rect 36446 6738 36492 6938
rect 36522 6900 36580 6910
rect 36522 6866 36534 6900
rect 36568 6866 36580 6900
rect 36522 6848 36580 6866
rect 36724 6858 36774 6938
rect 37140 6916 37224 7186
rect 36882 6906 36940 6912
rect 36874 6900 36948 6906
rect 36634 6819 36692 6836
rect 36634 6785 36646 6819
rect 36680 6785 36692 6819
rect 36634 6770 36692 6785
rect 36724 6792 36794 6858
rect 36874 6848 36885 6900
rect 36937 6848 36948 6900
rect 36874 6842 36948 6848
rect 37016 6890 37292 6916
rect 37886 6910 37984 7186
rect 37016 6885 37117 6890
rect 37169 6885 37292 6890
rect 37016 6851 37045 6885
rect 37079 6851 37117 6885
rect 37171 6851 37229 6885
rect 37263 6851 37292 6885
rect 36882 6834 36940 6842
rect 37016 6838 37117 6851
rect 37169 6838 37292 6851
rect 37016 6820 37292 6838
rect 37362 6879 37984 6910
rect 37362 6845 37391 6879
rect 37425 6845 37483 6879
rect 37517 6845 37575 6879
rect 37609 6877 37984 6879
rect 37609 6845 37737 6877
rect 37362 6843 37737 6845
rect 37771 6843 37829 6877
rect 37863 6843 37921 6877
rect 37955 6843 37984 6877
rect 38246 7140 38566 7158
rect 38246 7106 38518 7140
rect 38552 7106 38566 7140
rect 38246 7096 38566 7106
rect 37362 6812 37984 6843
rect 38124 6868 38200 6874
rect 38124 6816 38140 6868
rect 38192 6816 38200 6868
rect 38124 6810 38200 6816
rect 36724 6738 36774 6792
rect 38246 6766 38306 7096
rect 38368 7056 38414 7068
rect 36446 6691 36542 6738
rect 36446 6657 36502 6691
rect 36536 6657 36542 6691
rect 36446 6619 36542 6657
rect 36446 6585 36502 6619
rect 36536 6585 36542 6619
rect 36592 6691 36638 6738
rect 36592 6657 36598 6691
rect 36632 6657 36638 6691
rect 36592 6619 36638 6657
rect 36592 6598 36598 6619
rect 36446 6538 36542 6585
rect 36582 6590 36598 6598
rect 36632 6598 36638 6619
rect 36688 6691 36774 6738
rect 37778 6746 38306 6766
rect 37778 6712 37790 6746
rect 37824 6732 38306 6746
rect 37824 6712 37836 6732
rect 37778 6698 37836 6712
rect 36688 6657 36694 6691
rect 36728 6657 36774 6691
rect 36688 6619 36774 6657
rect 36632 6590 36648 6598
rect 36582 6538 36590 6590
rect 36642 6538 36648 6590
rect 36688 6585 36694 6619
rect 36728 6585 36774 6619
rect 36850 6659 36916 6672
rect 36850 6625 36866 6659
rect 36900 6625 36916 6659
rect 37244 6652 37312 6654
rect 36850 6614 36916 6625
rect 37160 6648 37312 6652
rect 37160 6642 37253 6648
rect 37160 6608 37180 6642
rect 37214 6608 37253 6642
rect 37160 6602 37253 6608
rect 37244 6596 37253 6602
rect 37305 6596 37312 6648
rect 37244 6590 37312 6596
rect 37348 6636 37422 6660
rect 37348 6602 37376 6636
rect 37410 6602 37422 6636
rect 36688 6542 36774 6585
rect 37348 6582 37422 6602
rect 37546 6652 37618 6664
rect 37546 6600 37557 6652
rect 37609 6600 37618 6652
rect 38092 6659 38158 6668
rect 38092 6625 38108 6659
rect 38142 6625 38158 6659
rect 38092 6612 38158 6625
rect 37546 6596 37618 6600
rect 36688 6538 36734 6542
rect 36582 6530 36648 6538
rect 36816 6531 36862 6578
rect 36358 6491 36596 6500
rect 36358 6468 36550 6491
rect 36258 6442 36264 6459
rect 35016 6376 35088 6404
rect 36170 6378 36216 6425
rect 36246 6436 36264 6442
rect 36298 6442 36304 6459
rect 36356 6457 36550 6468
rect 36584 6457 36596 6491
rect 36816 6497 36822 6531
rect 36856 6497 36862 6531
rect 36816 6464 36862 6497
rect 36298 6436 36312 6442
rect 36246 6384 36252 6436
rect 36304 6384 36312 6436
rect 36246 6378 36312 6384
rect 36356 6440 36596 6457
rect 34704 6328 34794 6349
rect 34962 6331 35028 6340
rect 34962 6297 34978 6331
rect 35012 6297 35028 6331
rect 34962 6294 35028 6297
rect 34468 6266 35028 6294
rect 34372 6210 34440 6224
rect 34372 6176 34390 6210
rect 34424 6176 34440 6210
rect 34372 6166 34440 6176
rect 34412 5862 34440 6166
rect 34468 6084 34502 6266
rect 34800 6200 34872 6212
rect 34800 6148 34810 6200
rect 34862 6148 34872 6200
rect 34800 6136 34872 6148
rect 34724 6084 34788 6102
rect 34468 6050 34740 6084
rect 34774 6050 34788 6084
rect 34724 6040 34788 6050
rect 35060 6026 35088 6376
rect 35128 6342 35404 6372
rect 35128 6341 35160 6342
rect 35212 6341 35404 6342
rect 35128 6307 35157 6341
rect 35212 6307 35249 6341
rect 35283 6307 35341 6341
rect 35375 6307 35404 6341
rect 35128 6290 35160 6307
rect 35212 6290 35404 6307
rect 35128 6276 35404 6290
rect 35472 6348 36096 6366
rect 35472 6335 36014 6348
rect 35472 6301 35503 6335
rect 35537 6301 35595 6335
rect 35629 6301 35687 6335
rect 35721 6333 36014 6335
rect 36066 6333 36096 6348
rect 35721 6301 35849 6333
rect 35472 6299 35849 6301
rect 35883 6299 35941 6333
rect 35975 6299 36014 6333
rect 36067 6299 36096 6333
rect 35472 6296 36014 6299
rect 36066 6296 36096 6299
rect 35178 6084 35244 6090
rect 35178 6032 35184 6084
rect 35236 6032 35244 6084
rect 35178 6026 35244 6032
rect 34834 6012 35088 6026
rect 34590 6000 34636 6012
rect 34136 5834 34440 5862
rect 34556 5966 34596 6000
rect 34630 5966 34636 6000
rect 34556 5928 34636 5966
rect 34676 6006 34742 6012
rect 34676 5954 34682 6006
rect 34734 5954 34742 6006
rect 34676 5948 34742 5954
rect 34782 6000 35088 6012
rect 34782 5966 34788 6000
rect 34822 5998 35088 6000
rect 34822 5966 34884 5998
rect 34556 5894 34596 5928
rect 34630 5894 34636 5928
rect 34556 5882 34636 5894
rect 34686 5928 34732 5948
rect 34686 5894 34692 5928
rect 34726 5894 34732 5928
rect 34686 5882 34732 5894
rect 34782 5928 34884 5966
rect 34782 5894 34788 5928
rect 34822 5894 34884 5928
rect 34782 5882 34884 5894
rect 35004 5951 35238 5960
rect 35004 5899 35010 5951
rect 35062 5932 35186 5951
rect 35062 5899 35068 5932
rect 35004 5892 35068 5899
rect 35180 5899 35186 5932
rect 35238 5899 35244 5932
rect 35180 5892 35244 5899
rect 34136 5831 34412 5834
rect 34136 5797 34165 5831
rect 34199 5797 34257 5831
rect 34291 5797 34349 5831
rect 34383 5797 34412 5831
rect 34136 5766 34412 5797
rect 34242 5718 34306 5724
rect 34242 5666 34248 5718
rect 34300 5666 34306 5718
rect 34242 5660 34306 5666
rect 34556 5682 34602 5882
rect 34632 5844 34690 5854
rect 34632 5810 34644 5844
rect 34678 5810 34690 5844
rect 34632 5792 34690 5810
rect 34744 5763 34802 5780
rect 34744 5729 34756 5763
rect 34790 5729 34802 5763
rect 34744 5714 34802 5729
rect 34834 5682 34884 5882
rect 34950 5831 35226 5862
rect 34950 5797 34979 5831
rect 35013 5797 35071 5831
rect 35105 5797 35163 5831
rect 35197 5797 35226 5831
rect 34950 5766 35226 5797
rect 34556 5635 34652 5682
rect 34154 5602 34218 5608
rect 34154 5550 34160 5602
rect 34212 5550 34218 5602
rect 34154 5544 34218 5550
rect 34324 5592 34394 5610
rect 34324 5558 34345 5592
rect 34379 5558 34394 5592
rect 34324 5550 34394 5558
rect 34556 5601 34612 5635
rect 34646 5601 34652 5635
rect 34556 5563 34652 5601
rect 34324 5514 34352 5550
rect 34556 5529 34612 5563
rect 34646 5529 34652 5563
rect 34702 5635 34748 5682
rect 34702 5601 34708 5635
rect 34742 5601 34748 5635
rect 34702 5563 34748 5601
rect 34702 5542 34708 5563
rect 34556 5514 34652 5529
rect 34324 5482 34652 5514
rect 34692 5534 34708 5542
rect 34742 5542 34748 5563
rect 34798 5635 34884 5682
rect 35056 5716 35124 5726
rect 35056 5664 35064 5716
rect 35116 5664 35124 5716
rect 35056 5658 35124 5664
rect 34798 5601 34804 5635
rect 34838 5601 34884 5635
rect 34798 5563 34884 5601
rect 34742 5534 34758 5542
rect 34692 5482 34700 5534
rect 34752 5482 34758 5534
rect 34798 5529 34804 5563
rect 34838 5529 34884 5563
rect 34966 5604 35034 5610
rect 34966 5552 34972 5604
rect 35024 5552 35034 5604
rect 34966 5546 35034 5552
rect 35140 5590 35206 5602
rect 35140 5556 35157 5590
rect 35191 5556 35206 5590
rect 35140 5548 35206 5556
rect 34798 5510 34884 5529
rect 35178 5510 35206 5548
rect 34798 5482 35206 5510
rect 34692 5474 34758 5482
rect 34840 5478 35206 5482
rect 34644 5435 34706 5444
rect 34644 5401 34660 5435
rect 34694 5401 34706 5435
rect 34644 5384 34706 5401
rect 34648 5382 34706 5384
rect 34702 5327 34792 5348
rect 34702 5318 34729 5327
rect 32875 5293 34729 5318
rect 34763 5318 34792 5327
rect 35306 5318 35384 6276
rect 35472 6264 36096 6296
rect 36204 6331 36270 6342
rect 36204 6297 36220 6331
rect 36254 6297 36270 6331
rect 36204 6286 36270 6297
rect 36356 6294 36390 6440
rect 36538 6438 36596 6440
rect 36794 6459 36862 6464
rect 36794 6456 36822 6459
rect 36794 6404 36802 6456
rect 36856 6425 36862 6459
rect 36854 6404 36862 6425
rect 36592 6383 36682 6404
rect 36794 6398 36862 6404
rect 36592 6349 36619 6383
rect 36653 6349 36682 6383
rect 36816 6378 36862 6398
rect 36904 6531 36950 6578
rect 36904 6497 36910 6531
rect 36944 6497 36950 6531
rect 36904 6459 36950 6497
rect 36904 6425 36910 6459
rect 36944 6425 36950 6459
rect 36904 6404 36950 6425
rect 38058 6531 38104 6578
rect 38058 6497 38064 6531
rect 38098 6497 38104 6531
rect 38058 6459 38104 6497
rect 38058 6425 38064 6459
rect 38098 6425 38104 6459
rect 38146 6531 38192 6578
rect 38146 6497 38152 6531
rect 38186 6497 38192 6531
rect 38146 6459 38192 6497
rect 38246 6500 38306 6732
rect 38334 7022 38374 7056
rect 38408 7022 38414 7056
rect 38334 6984 38414 7022
rect 38454 7062 38520 7068
rect 38454 7010 38460 7062
rect 38512 7010 38520 7062
rect 38454 7004 38520 7010
rect 38560 7056 38662 7068
rect 38560 7022 38566 7056
rect 38600 7022 38662 7056
rect 38334 6950 38374 6984
rect 38408 6950 38414 6984
rect 38334 6938 38414 6950
rect 38464 6984 38510 7004
rect 38464 6950 38470 6984
rect 38504 6950 38510 6984
rect 38464 6938 38510 6950
rect 38560 6984 38662 7022
rect 38560 6950 38566 6984
rect 38600 6950 38662 6984
rect 38560 6938 38662 6950
rect 38334 6738 38380 6938
rect 38410 6900 38468 6910
rect 38410 6866 38422 6900
rect 38456 6866 38468 6900
rect 38410 6848 38468 6866
rect 38612 6858 38662 6938
rect 39028 6916 39112 7186
rect 38770 6906 38828 6912
rect 38762 6900 38836 6906
rect 38522 6819 38580 6836
rect 38522 6785 38534 6819
rect 38568 6785 38580 6819
rect 38522 6770 38580 6785
rect 38612 6792 38682 6858
rect 38762 6848 38773 6900
rect 38825 6848 38836 6900
rect 38762 6842 38836 6848
rect 38904 6890 39180 6916
rect 39774 6910 39872 7186
rect 38904 6885 39005 6890
rect 39057 6885 39180 6890
rect 38904 6851 38933 6885
rect 38967 6851 39005 6885
rect 39059 6851 39117 6885
rect 39151 6851 39180 6885
rect 38770 6834 38828 6842
rect 38904 6838 39005 6851
rect 39057 6838 39180 6851
rect 38904 6820 39180 6838
rect 39250 6879 39872 6910
rect 39250 6845 39279 6879
rect 39313 6845 39371 6879
rect 39405 6845 39463 6879
rect 39497 6877 39872 6879
rect 39497 6845 39625 6877
rect 39250 6843 39625 6845
rect 39659 6843 39717 6877
rect 39751 6843 39809 6877
rect 39843 6843 39872 6877
rect 40134 7140 40454 7158
rect 40134 7106 40406 7140
rect 40440 7106 40454 7140
rect 40134 7096 40454 7106
rect 39250 6812 39872 6843
rect 40012 6868 40088 6874
rect 40012 6816 40028 6868
rect 40080 6816 40088 6868
rect 40012 6810 40088 6816
rect 38612 6738 38662 6792
rect 40134 6766 40194 7096
rect 40256 7056 40302 7068
rect 38334 6691 38430 6738
rect 38334 6657 38390 6691
rect 38424 6657 38430 6691
rect 38334 6619 38430 6657
rect 38334 6585 38390 6619
rect 38424 6585 38430 6619
rect 38480 6691 38526 6738
rect 38480 6657 38486 6691
rect 38520 6657 38526 6691
rect 38480 6619 38526 6657
rect 38480 6598 38486 6619
rect 38334 6538 38430 6585
rect 38470 6590 38486 6598
rect 38520 6598 38526 6619
rect 38576 6691 38662 6738
rect 39666 6746 40194 6766
rect 39666 6712 39678 6746
rect 39712 6732 40194 6746
rect 39712 6712 39724 6732
rect 39666 6698 39724 6712
rect 38576 6657 38582 6691
rect 38616 6657 38662 6691
rect 38576 6619 38662 6657
rect 38520 6590 38536 6598
rect 38470 6538 38478 6590
rect 38530 6538 38536 6590
rect 38576 6585 38582 6619
rect 38616 6585 38662 6619
rect 38738 6659 38804 6672
rect 38738 6625 38754 6659
rect 38788 6625 38804 6659
rect 39132 6652 39200 6654
rect 38738 6614 38804 6625
rect 39048 6648 39200 6652
rect 39048 6642 39141 6648
rect 39048 6608 39068 6642
rect 39102 6608 39141 6642
rect 39048 6602 39141 6608
rect 39132 6596 39141 6602
rect 39193 6596 39200 6648
rect 39132 6590 39200 6596
rect 39236 6636 39310 6660
rect 39236 6602 39264 6636
rect 39298 6602 39310 6636
rect 38576 6542 38662 6585
rect 39236 6582 39310 6602
rect 39434 6652 39506 6664
rect 39434 6600 39445 6652
rect 39497 6600 39506 6652
rect 39980 6659 40046 6668
rect 39980 6625 39996 6659
rect 40030 6625 40046 6659
rect 39980 6612 40046 6625
rect 39434 6596 39506 6600
rect 38576 6538 38622 6542
rect 38470 6530 38536 6538
rect 38704 6531 38750 6578
rect 38246 6491 38484 6500
rect 38246 6468 38438 6491
rect 38146 6442 38152 6459
rect 36904 6376 36976 6404
rect 38058 6378 38104 6425
rect 38134 6436 38152 6442
rect 38186 6442 38192 6459
rect 38244 6457 38438 6468
rect 38472 6457 38484 6491
rect 38704 6497 38710 6531
rect 38744 6497 38750 6531
rect 38704 6464 38750 6497
rect 38186 6436 38200 6442
rect 38134 6384 38140 6436
rect 38192 6384 38200 6436
rect 38134 6378 38200 6384
rect 38244 6440 38484 6457
rect 36592 6328 36682 6349
rect 36850 6331 36916 6340
rect 36850 6297 36866 6331
rect 36900 6297 36916 6331
rect 36850 6294 36916 6297
rect 36356 6266 36916 6294
rect 36260 6210 36328 6224
rect 36260 6176 36278 6210
rect 36312 6176 36328 6210
rect 36260 6166 36328 6176
rect 36300 5862 36328 6166
rect 36356 6084 36390 6266
rect 36688 6200 36760 6212
rect 36688 6148 36698 6200
rect 36750 6148 36760 6200
rect 36688 6136 36760 6148
rect 36612 6084 36676 6102
rect 36356 6050 36628 6084
rect 36662 6050 36676 6084
rect 36612 6040 36676 6050
rect 36948 6026 36976 6376
rect 37016 6342 37292 6372
rect 37016 6341 37048 6342
rect 37100 6341 37292 6342
rect 37016 6307 37045 6341
rect 37100 6307 37137 6341
rect 37171 6307 37229 6341
rect 37263 6307 37292 6341
rect 37016 6290 37048 6307
rect 37100 6290 37292 6307
rect 37016 6276 37292 6290
rect 37360 6348 37984 6366
rect 37360 6335 37902 6348
rect 37360 6301 37391 6335
rect 37425 6301 37483 6335
rect 37517 6301 37575 6335
rect 37609 6333 37902 6335
rect 37954 6333 37984 6348
rect 37609 6301 37737 6333
rect 37360 6299 37737 6301
rect 37771 6299 37829 6333
rect 37863 6299 37902 6333
rect 37955 6299 37984 6333
rect 37360 6296 37902 6299
rect 37954 6296 37984 6299
rect 37066 6084 37132 6090
rect 37066 6032 37072 6084
rect 37124 6032 37132 6084
rect 37066 6026 37132 6032
rect 36722 6012 36976 6026
rect 36478 6000 36524 6012
rect 36024 5834 36328 5862
rect 36444 5966 36484 6000
rect 36518 5966 36524 6000
rect 36444 5928 36524 5966
rect 36564 6006 36630 6012
rect 36564 5954 36570 6006
rect 36622 5954 36630 6006
rect 36564 5948 36630 5954
rect 36670 6000 36976 6012
rect 36670 5966 36676 6000
rect 36710 5998 36976 6000
rect 36710 5966 36772 5998
rect 36444 5894 36484 5928
rect 36518 5894 36524 5928
rect 36444 5882 36524 5894
rect 36574 5928 36620 5948
rect 36574 5894 36580 5928
rect 36614 5894 36620 5928
rect 36574 5882 36620 5894
rect 36670 5928 36772 5966
rect 36670 5894 36676 5928
rect 36710 5894 36772 5928
rect 36670 5882 36772 5894
rect 36892 5951 37126 5960
rect 36892 5899 36898 5951
rect 36950 5932 37074 5951
rect 36950 5899 36956 5932
rect 36892 5892 36956 5899
rect 37068 5899 37074 5932
rect 37126 5899 37132 5932
rect 37068 5892 37132 5899
rect 36024 5831 36300 5834
rect 36024 5797 36053 5831
rect 36087 5797 36145 5831
rect 36179 5797 36237 5831
rect 36271 5797 36300 5831
rect 36024 5766 36300 5797
rect 36130 5718 36194 5724
rect 36130 5666 36136 5718
rect 36188 5666 36194 5718
rect 36130 5660 36194 5666
rect 36444 5682 36490 5882
rect 36520 5844 36578 5854
rect 36520 5810 36532 5844
rect 36566 5810 36578 5844
rect 36520 5792 36578 5810
rect 36632 5763 36690 5780
rect 36632 5729 36644 5763
rect 36678 5729 36690 5763
rect 36632 5714 36690 5729
rect 36722 5682 36772 5882
rect 36838 5831 37114 5862
rect 36838 5797 36867 5831
rect 36901 5797 36959 5831
rect 36993 5797 37051 5831
rect 37085 5797 37114 5831
rect 36838 5766 37114 5797
rect 36444 5635 36540 5682
rect 36042 5602 36106 5608
rect 36042 5550 36048 5602
rect 36100 5550 36106 5602
rect 36042 5544 36106 5550
rect 36212 5592 36282 5610
rect 36212 5558 36233 5592
rect 36267 5558 36282 5592
rect 36212 5550 36282 5558
rect 36444 5601 36500 5635
rect 36534 5601 36540 5635
rect 36444 5563 36540 5601
rect 36212 5514 36240 5550
rect 36444 5529 36500 5563
rect 36534 5529 36540 5563
rect 36590 5635 36636 5682
rect 36590 5601 36596 5635
rect 36630 5601 36636 5635
rect 36590 5563 36636 5601
rect 36590 5542 36596 5563
rect 36444 5514 36540 5529
rect 36212 5482 36540 5514
rect 36580 5534 36596 5542
rect 36630 5542 36636 5563
rect 36686 5635 36772 5682
rect 36944 5716 37012 5726
rect 36944 5664 36952 5716
rect 37004 5664 37012 5716
rect 36944 5658 37012 5664
rect 36686 5601 36692 5635
rect 36726 5601 36772 5635
rect 36686 5563 36772 5601
rect 36630 5534 36646 5542
rect 36580 5482 36588 5534
rect 36640 5482 36646 5534
rect 36686 5529 36692 5563
rect 36726 5529 36772 5563
rect 36854 5604 36922 5610
rect 36854 5552 36860 5604
rect 36912 5552 36922 5604
rect 36854 5546 36922 5552
rect 37028 5590 37094 5602
rect 37028 5556 37045 5590
rect 37079 5556 37094 5590
rect 37028 5548 37094 5556
rect 36686 5510 36772 5529
rect 37066 5510 37094 5548
rect 36686 5482 37094 5510
rect 36580 5474 36646 5482
rect 36728 5478 37094 5482
rect 36532 5435 36594 5444
rect 36532 5401 36548 5435
rect 36582 5401 36594 5435
rect 36532 5384 36594 5401
rect 36536 5382 36594 5384
rect 36590 5327 36680 5348
rect 36590 5318 36617 5327
rect 34763 5293 36617 5318
rect 36651 5318 36680 5327
rect 37194 5318 37272 6276
rect 37360 6264 37984 6296
rect 38092 6331 38158 6342
rect 38092 6297 38108 6331
rect 38142 6297 38158 6331
rect 38092 6286 38158 6297
rect 38244 6294 38278 6440
rect 38426 6438 38484 6440
rect 38682 6459 38750 6464
rect 38682 6456 38710 6459
rect 38682 6404 38690 6456
rect 38744 6425 38750 6459
rect 38742 6404 38750 6425
rect 38480 6383 38570 6404
rect 38682 6398 38750 6404
rect 38480 6349 38507 6383
rect 38541 6349 38570 6383
rect 38704 6378 38750 6398
rect 38792 6531 38838 6578
rect 38792 6497 38798 6531
rect 38832 6497 38838 6531
rect 38792 6459 38838 6497
rect 38792 6425 38798 6459
rect 38832 6425 38838 6459
rect 38792 6404 38838 6425
rect 39946 6531 39992 6578
rect 39946 6497 39952 6531
rect 39986 6497 39992 6531
rect 39946 6459 39992 6497
rect 39946 6425 39952 6459
rect 39986 6425 39992 6459
rect 40034 6531 40080 6578
rect 40034 6497 40040 6531
rect 40074 6497 40080 6531
rect 40034 6459 40080 6497
rect 40134 6500 40194 6732
rect 40222 7022 40262 7056
rect 40296 7022 40302 7056
rect 40222 6984 40302 7022
rect 40342 7062 40408 7068
rect 40342 7010 40348 7062
rect 40400 7010 40408 7062
rect 40342 7004 40408 7010
rect 40448 7056 40550 7068
rect 40448 7022 40454 7056
rect 40488 7022 40550 7056
rect 40222 6950 40262 6984
rect 40296 6950 40302 6984
rect 40222 6938 40302 6950
rect 40352 6984 40398 7004
rect 40352 6950 40358 6984
rect 40392 6950 40398 6984
rect 40352 6938 40398 6950
rect 40448 6984 40550 7022
rect 40448 6950 40454 6984
rect 40488 6950 40550 6984
rect 40448 6938 40550 6950
rect 40222 6738 40268 6938
rect 40298 6900 40356 6910
rect 40298 6866 40310 6900
rect 40344 6866 40356 6900
rect 40298 6848 40356 6866
rect 40500 6858 40550 6938
rect 40916 6916 41000 7186
rect 40658 6906 40716 6912
rect 40650 6900 40724 6906
rect 40410 6819 40468 6836
rect 40410 6785 40422 6819
rect 40456 6785 40468 6819
rect 40410 6770 40468 6785
rect 40500 6792 40570 6858
rect 40650 6848 40661 6900
rect 40713 6848 40724 6900
rect 40650 6842 40724 6848
rect 40792 6890 41068 6916
rect 41662 6910 41760 7186
rect 40792 6885 40893 6890
rect 40945 6885 41068 6890
rect 40792 6851 40821 6885
rect 40855 6851 40893 6885
rect 40947 6851 41005 6885
rect 41039 6851 41068 6885
rect 40658 6834 40716 6842
rect 40792 6838 40893 6851
rect 40945 6838 41068 6851
rect 40792 6820 41068 6838
rect 41138 6879 41760 6910
rect 41138 6845 41167 6879
rect 41201 6845 41259 6879
rect 41293 6845 41351 6879
rect 41385 6877 41760 6879
rect 41385 6845 41513 6877
rect 41138 6843 41513 6845
rect 41547 6843 41605 6877
rect 41639 6843 41697 6877
rect 41731 6843 41760 6877
rect 42022 7140 42342 7158
rect 42022 7106 42294 7140
rect 42328 7106 42342 7140
rect 42022 7096 42342 7106
rect 41138 6812 41760 6843
rect 41900 6868 41976 6874
rect 41900 6816 41916 6868
rect 41968 6816 41976 6868
rect 41900 6810 41976 6816
rect 40500 6738 40550 6792
rect 42022 6766 42082 7096
rect 42144 7056 42190 7068
rect 40222 6691 40318 6738
rect 40222 6657 40278 6691
rect 40312 6657 40318 6691
rect 40222 6619 40318 6657
rect 40222 6585 40278 6619
rect 40312 6585 40318 6619
rect 40368 6691 40414 6738
rect 40368 6657 40374 6691
rect 40408 6657 40414 6691
rect 40368 6619 40414 6657
rect 40368 6598 40374 6619
rect 40222 6538 40318 6585
rect 40358 6590 40374 6598
rect 40408 6598 40414 6619
rect 40464 6691 40550 6738
rect 41554 6746 42082 6766
rect 41554 6712 41566 6746
rect 41600 6732 42082 6746
rect 41600 6712 41612 6732
rect 41554 6698 41612 6712
rect 40464 6657 40470 6691
rect 40504 6657 40550 6691
rect 40464 6619 40550 6657
rect 40408 6590 40424 6598
rect 40358 6538 40366 6590
rect 40418 6538 40424 6590
rect 40464 6585 40470 6619
rect 40504 6585 40550 6619
rect 40626 6659 40692 6672
rect 40626 6625 40642 6659
rect 40676 6625 40692 6659
rect 41020 6652 41088 6654
rect 40626 6614 40692 6625
rect 40936 6648 41088 6652
rect 40936 6642 41029 6648
rect 40936 6608 40956 6642
rect 40990 6608 41029 6642
rect 40936 6602 41029 6608
rect 41020 6596 41029 6602
rect 41081 6596 41088 6648
rect 41020 6590 41088 6596
rect 41124 6636 41198 6660
rect 41124 6602 41152 6636
rect 41186 6602 41198 6636
rect 40464 6542 40550 6585
rect 41124 6582 41198 6602
rect 41322 6652 41394 6664
rect 41322 6600 41333 6652
rect 41385 6600 41394 6652
rect 41868 6659 41934 6668
rect 41868 6625 41884 6659
rect 41918 6625 41934 6659
rect 41868 6612 41934 6625
rect 41322 6596 41394 6600
rect 40464 6538 40510 6542
rect 40358 6530 40424 6538
rect 40592 6531 40638 6578
rect 40134 6491 40372 6500
rect 40134 6468 40326 6491
rect 40034 6442 40040 6459
rect 38792 6376 38864 6404
rect 39946 6378 39992 6425
rect 40022 6436 40040 6442
rect 40074 6442 40080 6459
rect 40132 6457 40326 6468
rect 40360 6457 40372 6491
rect 40592 6497 40598 6531
rect 40632 6497 40638 6531
rect 40592 6464 40638 6497
rect 40074 6436 40088 6442
rect 40022 6384 40028 6436
rect 40080 6384 40088 6436
rect 40022 6378 40088 6384
rect 40132 6440 40372 6457
rect 38480 6328 38570 6349
rect 38738 6331 38804 6340
rect 38738 6297 38754 6331
rect 38788 6297 38804 6331
rect 38738 6294 38804 6297
rect 38244 6266 38804 6294
rect 38148 6210 38216 6224
rect 38148 6176 38166 6210
rect 38200 6176 38216 6210
rect 38148 6166 38216 6176
rect 38188 5862 38216 6166
rect 38244 6084 38278 6266
rect 38576 6200 38648 6212
rect 38576 6148 38586 6200
rect 38638 6148 38648 6200
rect 38576 6136 38648 6148
rect 38500 6084 38564 6102
rect 38244 6050 38516 6084
rect 38550 6050 38564 6084
rect 38500 6040 38564 6050
rect 38836 6026 38864 6376
rect 38904 6342 39180 6372
rect 38904 6341 38936 6342
rect 38988 6341 39180 6342
rect 38904 6307 38933 6341
rect 38988 6307 39025 6341
rect 39059 6307 39117 6341
rect 39151 6307 39180 6341
rect 38904 6290 38936 6307
rect 38988 6290 39180 6307
rect 38904 6276 39180 6290
rect 39248 6348 39872 6366
rect 39248 6335 39790 6348
rect 39248 6301 39279 6335
rect 39313 6301 39371 6335
rect 39405 6301 39463 6335
rect 39497 6333 39790 6335
rect 39842 6333 39872 6348
rect 39497 6301 39625 6333
rect 39248 6299 39625 6301
rect 39659 6299 39717 6333
rect 39751 6299 39790 6333
rect 39843 6299 39872 6333
rect 39248 6296 39790 6299
rect 39842 6296 39872 6299
rect 38954 6084 39020 6090
rect 38954 6032 38960 6084
rect 39012 6032 39020 6084
rect 38954 6026 39020 6032
rect 38610 6012 38864 6026
rect 38366 6000 38412 6012
rect 37912 5834 38216 5862
rect 38332 5966 38372 6000
rect 38406 5966 38412 6000
rect 38332 5928 38412 5966
rect 38452 6006 38518 6012
rect 38452 5954 38458 6006
rect 38510 5954 38518 6006
rect 38452 5948 38518 5954
rect 38558 6000 38864 6012
rect 38558 5966 38564 6000
rect 38598 5998 38864 6000
rect 38598 5966 38660 5998
rect 38332 5894 38372 5928
rect 38406 5894 38412 5928
rect 38332 5882 38412 5894
rect 38462 5928 38508 5948
rect 38462 5894 38468 5928
rect 38502 5894 38508 5928
rect 38462 5882 38508 5894
rect 38558 5928 38660 5966
rect 38558 5894 38564 5928
rect 38598 5894 38660 5928
rect 38558 5882 38660 5894
rect 38780 5951 39014 5960
rect 38780 5899 38786 5951
rect 38838 5932 38962 5951
rect 38838 5899 38844 5932
rect 38780 5892 38844 5899
rect 38956 5899 38962 5932
rect 39014 5899 39020 5932
rect 38956 5892 39020 5899
rect 37912 5831 38188 5834
rect 37912 5797 37941 5831
rect 37975 5797 38033 5831
rect 38067 5797 38125 5831
rect 38159 5797 38188 5831
rect 37912 5766 38188 5797
rect 38018 5718 38082 5724
rect 38018 5666 38024 5718
rect 38076 5666 38082 5718
rect 38018 5660 38082 5666
rect 38332 5682 38378 5882
rect 38408 5844 38466 5854
rect 38408 5810 38420 5844
rect 38454 5810 38466 5844
rect 38408 5792 38466 5810
rect 38520 5763 38578 5780
rect 38520 5729 38532 5763
rect 38566 5729 38578 5763
rect 38520 5714 38578 5729
rect 38610 5682 38660 5882
rect 38726 5831 39002 5862
rect 38726 5797 38755 5831
rect 38789 5797 38847 5831
rect 38881 5797 38939 5831
rect 38973 5797 39002 5831
rect 38726 5766 39002 5797
rect 38332 5635 38428 5682
rect 37930 5602 37994 5608
rect 37930 5550 37936 5602
rect 37988 5550 37994 5602
rect 37930 5544 37994 5550
rect 38100 5592 38170 5610
rect 38100 5558 38121 5592
rect 38155 5558 38170 5592
rect 38100 5550 38170 5558
rect 38332 5601 38388 5635
rect 38422 5601 38428 5635
rect 38332 5563 38428 5601
rect 38100 5514 38128 5550
rect 38332 5529 38388 5563
rect 38422 5529 38428 5563
rect 38478 5635 38524 5682
rect 38478 5601 38484 5635
rect 38518 5601 38524 5635
rect 38478 5563 38524 5601
rect 38478 5542 38484 5563
rect 38332 5514 38428 5529
rect 38100 5482 38428 5514
rect 38468 5534 38484 5542
rect 38518 5542 38524 5563
rect 38574 5635 38660 5682
rect 38832 5716 38900 5726
rect 38832 5664 38840 5716
rect 38892 5664 38900 5716
rect 38832 5658 38900 5664
rect 38574 5601 38580 5635
rect 38614 5601 38660 5635
rect 38574 5563 38660 5601
rect 38518 5534 38534 5542
rect 38468 5482 38476 5534
rect 38528 5482 38534 5534
rect 38574 5529 38580 5563
rect 38614 5529 38660 5563
rect 38742 5604 38810 5610
rect 38742 5552 38748 5604
rect 38800 5552 38810 5604
rect 38742 5546 38810 5552
rect 38916 5590 38982 5602
rect 38916 5556 38933 5590
rect 38967 5556 38982 5590
rect 38916 5548 38982 5556
rect 38574 5510 38660 5529
rect 38954 5510 38982 5548
rect 38574 5482 38982 5510
rect 38468 5474 38534 5482
rect 38616 5478 38982 5482
rect 38420 5435 38482 5444
rect 38420 5401 38436 5435
rect 38470 5401 38482 5435
rect 38420 5384 38482 5401
rect 38424 5382 38482 5384
rect 38478 5327 38568 5348
rect 38478 5318 38505 5327
rect 36651 5293 38505 5318
rect 38539 5318 38568 5327
rect 39082 5318 39160 6276
rect 39248 6264 39872 6296
rect 39980 6331 40046 6342
rect 39980 6297 39996 6331
rect 40030 6297 40046 6331
rect 39980 6286 40046 6297
rect 40132 6294 40166 6440
rect 40314 6438 40372 6440
rect 40570 6459 40638 6464
rect 40570 6456 40598 6459
rect 40570 6404 40578 6456
rect 40632 6425 40638 6459
rect 40630 6404 40638 6425
rect 40368 6383 40458 6404
rect 40570 6398 40638 6404
rect 40368 6349 40395 6383
rect 40429 6349 40458 6383
rect 40592 6378 40638 6398
rect 40680 6531 40726 6578
rect 40680 6497 40686 6531
rect 40720 6497 40726 6531
rect 40680 6459 40726 6497
rect 40680 6425 40686 6459
rect 40720 6425 40726 6459
rect 40680 6404 40726 6425
rect 41834 6531 41880 6578
rect 41834 6497 41840 6531
rect 41874 6497 41880 6531
rect 41834 6459 41880 6497
rect 41834 6425 41840 6459
rect 41874 6425 41880 6459
rect 41922 6531 41968 6578
rect 41922 6497 41928 6531
rect 41962 6497 41968 6531
rect 41922 6459 41968 6497
rect 42022 6500 42082 6732
rect 42110 7022 42150 7056
rect 42184 7022 42190 7056
rect 42110 6984 42190 7022
rect 42230 7062 42296 7068
rect 42230 7010 42236 7062
rect 42288 7010 42296 7062
rect 42230 7004 42296 7010
rect 42336 7056 42438 7068
rect 42336 7022 42342 7056
rect 42376 7022 42438 7056
rect 42110 6950 42150 6984
rect 42184 6950 42190 6984
rect 42110 6938 42190 6950
rect 42240 6984 42286 7004
rect 42240 6950 42246 6984
rect 42280 6950 42286 6984
rect 42240 6938 42286 6950
rect 42336 6984 42438 7022
rect 42336 6950 42342 6984
rect 42376 6950 42438 6984
rect 42336 6938 42438 6950
rect 42110 6738 42156 6938
rect 42186 6900 42244 6910
rect 42186 6866 42198 6900
rect 42232 6866 42244 6900
rect 42186 6848 42244 6866
rect 42388 6858 42438 6938
rect 42804 6916 42888 7186
rect 42546 6906 42604 6912
rect 42538 6900 42612 6906
rect 42298 6819 42356 6836
rect 42298 6785 42310 6819
rect 42344 6785 42356 6819
rect 42298 6770 42356 6785
rect 42388 6792 42458 6858
rect 42538 6848 42549 6900
rect 42601 6848 42612 6900
rect 42538 6842 42612 6848
rect 42680 6890 42956 6916
rect 43550 6910 43648 7186
rect 42680 6885 42781 6890
rect 42833 6885 42956 6890
rect 42680 6851 42709 6885
rect 42743 6851 42781 6885
rect 42835 6851 42893 6885
rect 42927 6851 42956 6885
rect 42546 6834 42604 6842
rect 42680 6838 42781 6851
rect 42833 6838 42956 6851
rect 42680 6820 42956 6838
rect 43026 6879 43648 6910
rect 43026 6845 43055 6879
rect 43089 6845 43147 6879
rect 43181 6845 43239 6879
rect 43273 6877 43648 6879
rect 43273 6845 43401 6877
rect 43026 6843 43401 6845
rect 43435 6843 43493 6877
rect 43527 6843 43585 6877
rect 43619 6843 43648 6877
rect 43910 7140 44230 7158
rect 43910 7106 44182 7140
rect 44216 7106 44230 7140
rect 43910 7096 44230 7106
rect 43026 6812 43648 6843
rect 43788 6868 43864 6874
rect 43788 6816 43804 6868
rect 43856 6816 43864 6868
rect 43788 6810 43864 6816
rect 42388 6738 42438 6792
rect 43910 6766 43970 7096
rect 44032 7056 44078 7068
rect 42110 6691 42206 6738
rect 42110 6657 42166 6691
rect 42200 6657 42206 6691
rect 42110 6619 42206 6657
rect 42110 6585 42166 6619
rect 42200 6585 42206 6619
rect 42256 6691 42302 6738
rect 42256 6657 42262 6691
rect 42296 6657 42302 6691
rect 42256 6619 42302 6657
rect 42256 6598 42262 6619
rect 42110 6538 42206 6585
rect 42246 6590 42262 6598
rect 42296 6598 42302 6619
rect 42352 6691 42438 6738
rect 43442 6746 43970 6766
rect 43442 6712 43454 6746
rect 43488 6732 43970 6746
rect 43488 6712 43500 6732
rect 43442 6698 43500 6712
rect 42352 6657 42358 6691
rect 42392 6657 42438 6691
rect 42352 6619 42438 6657
rect 42296 6590 42312 6598
rect 42246 6538 42254 6590
rect 42306 6538 42312 6590
rect 42352 6585 42358 6619
rect 42392 6585 42438 6619
rect 42514 6659 42580 6672
rect 42514 6625 42530 6659
rect 42564 6625 42580 6659
rect 42908 6652 42976 6654
rect 42514 6614 42580 6625
rect 42824 6648 42976 6652
rect 42824 6642 42917 6648
rect 42824 6608 42844 6642
rect 42878 6608 42917 6642
rect 42824 6602 42917 6608
rect 42908 6596 42917 6602
rect 42969 6596 42976 6648
rect 42908 6590 42976 6596
rect 43012 6636 43086 6660
rect 43012 6602 43040 6636
rect 43074 6602 43086 6636
rect 42352 6542 42438 6585
rect 43012 6582 43086 6602
rect 43210 6652 43282 6664
rect 43210 6600 43221 6652
rect 43273 6600 43282 6652
rect 43756 6659 43822 6668
rect 43756 6625 43772 6659
rect 43806 6625 43822 6659
rect 43756 6612 43822 6625
rect 43210 6596 43282 6600
rect 42352 6538 42398 6542
rect 42246 6530 42312 6538
rect 42480 6531 42526 6578
rect 42022 6491 42260 6500
rect 42022 6468 42214 6491
rect 41922 6442 41928 6459
rect 40680 6376 40752 6404
rect 41834 6378 41880 6425
rect 41910 6436 41928 6442
rect 41962 6442 41968 6459
rect 42020 6457 42214 6468
rect 42248 6457 42260 6491
rect 42480 6497 42486 6531
rect 42520 6497 42526 6531
rect 42480 6464 42526 6497
rect 41962 6436 41976 6442
rect 41910 6384 41916 6436
rect 41968 6384 41976 6436
rect 41910 6378 41976 6384
rect 42020 6440 42260 6457
rect 40368 6328 40458 6349
rect 40626 6331 40692 6340
rect 40626 6297 40642 6331
rect 40676 6297 40692 6331
rect 40626 6294 40692 6297
rect 40132 6266 40692 6294
rect 40036 6210 40104 6224
rect 40036 6176 40054 6210
rect 40088 6176 40104 6210
rect 40036 6166 40104 6176
rect 40076 5862 40104 6166
rect 40132 6084 40166 6266
rect 40464 6200 40536 6212
rect 40464 6148 40474 6200
rect 40526 6148 40536 6200
rect 40464 6136 40536 6148
rect 40388 6084 40452 6102
rect 40132 6050 40404 6084
rect 40438 6050 40452 6084
rect 40388 6040 40452 6050
rect 40724 6026 40752 6376
rect 40792 6342 41068 6372
rect 40792 6341 40824 6342
rect 40876 6341 41068 6342
rect 40792 6307 40821 6341
rect 40876 6307 40913 6341
rect 40947 6307 41005 6341
rect 41039 6307 41068 6341
rect 40792 6290 40824 6307
rect 40876 6290 41068 6307
rect 40792 6276 41068 6290
rect 41136 6348 41760 6366
rect 41136 6335 41678 6348
rect 41136 6301 41167 6335
rect 41201 6301 41259 6335
rect 41293 6301 41351 6335
rect 41385 6333 41678 6335
rect 41730 6333 41760 6348
rect 41385 6301 41513 6333
rect 41136 6299 41513 6301
rect 41547 6299 41605 6333
rect 41639 6299 41678 6333
rect 41731 6299 41760 6333
rect 41136 6296 41678 6299
rect 41730 6296 41760 6299
rect 40842 6084 40908 6090
rect 40842 6032 40848 6084
rect 40900 6032 40908 6084
rect 40842 6026 40908 6032
rect 40498 6012 40752 6026
rect 40254 6000 40300 6012
rect 39800 5834 40104 5862
rect 40220 5966 40260 6000
rect 40294 5966 40300 6000
rect 40220 5928 40300 5966
rect 40340 6006 40406 6012
rect 40340 5954 40346 6006
rect 40398 5954 40406 6006
rect 40340 5948 40406 5954
rect 40446 6000 40752 6012
rect 40446 5966 40452 6000
rect 40486 5998 40752 6000
rect 40486 5966 40548 5998
rect 40220 5894 40260 5928
rect 40294 5894 40300 5928
rect 40220 5882 40300 5894
rect 40350 5928 40396 5948
rect 40350 5894 40356 5928
rect 40390 5894 40396 5928
rect 40350 5882 40396 5894
rect 40446 5928 40548 5966
rect 40446 5894 40452 5928
rect 40486 5894 40548 5928
rect 40446 5882 40548 5894
rect 40668 5951 40902 5960
rect 40668 5899 40674 5951
rect 40726 5932 40850 5951
rect 40726 5899 40732 5932
rect 40668 5892 40732 5899
rect 40844 5899 40850 5932
rect 40902 5899 40908 5932
rect 40844 5892 40908 5899
rect 39800 5831 40076 5834
rect 39800 5797 39829 5831
rect 39863 5797 39921 5831
rect 39955 5797 40013 5831
rect 40047 5797 40076 5831
rect 39800 5766 40076 5797
rect 39906 5718 39970 5724
rect 39906 5666 39912 5718
rect 39964 5666 39970 5718
rect 39906 5660 39970 5666
rect 40220 5682 40266 5882
rect 40296 5844 40354 5854
rect 40296 5810 40308 5844
rect 40342 5810 40354 5844
rect 40296 5792 40354 5810
rect 40408 5763 40466 5780
rect 40408 5729 40420 5763
rect 40454 5729 40466 5763
rect 40408 5714 40466 5729
rect 40498 5682 40548 5882
rect 40614 5831 40890 5862
rect 40614 5797 40643 5831
rect 40677 5797 40735 5831
rect 40769 5797 40827 5831
rect 40861 5797 40890 5831
rect 40614 5766 40890 5797
rect 40220 5635 40316 5682
rect 39818 5602 39882 5608
rect 39818 5550 39824 5602
rect 39876 5550 39882 5602
rect 39818 5544 39882 5550
rect 39988 5592 40058 5610
rect 39988 5558 40009 5592
rect 40043 5558 40058 5592
rect 39988 5550 40058 5558
rect 40220 5601 40276 5635
rect 40310 5601 40316 5635
rect 40220 5563 40316 5601
rect 39988 5514 40016 5550
rect 40220 5529 40276 5563
rect 40310 5529 40316 5563
rect 40366 5635 40412 5682
rect 40366 5601 40372 5635
rect 40406 5601 40412 5635
rect 40366 5563 40412 5601
rect 40366 5542 40372 5563
rect 40220 5514 40316 5529
rect 39988 5482 40316 5514
rect 40356 5534 40372 5542
rect 40406 5542 40412 5563
rect 40462 5635 40548 5682
rect 40720 5716 40788 5726
rect 40720 5664 40728 5716
rect 40780 5664 40788 5716
rect 40720 5658 40788 5664
rect 40462 5601 40468 5635
rect 40502 5601 40548 5635
rect 40462 5563 40548 5601
rect 40406 5534 40422 5542
rect 40356 5482 40364 5534
rect 40416 5482 40422 5534
rect 40462 5529 40468 5563
rect 40502 5529 40548 5563
rect 40630 5604 40698 5610
rect 40630 5552 40636 5604
rect 40688 5552 40698 5604
rect 40630 5546 40698 5552
rect 40804 5590 40870 5602
rect 40804 5556 40821 5590
rect 40855 5556 40870 5590
rect 40804 5548 40870 5556
rect 40462 5510 40548 5529
rect 40842 5510 40870 5548
rect 40462 5482 40870 5510
rect 40356 5474 40422 5482
rect 40504 5478 40870 5482
rect 40308 5435 40370 5444
rect 40308 5401 40324 5435
rect 40358 5401 40370 5435
rect 40308 5384 40370 5401
rect 40312 5382 40370 5384
rect 40366 5327 40456 5348
rect 40366 5318 40393 5327
rect 38539 5293 40393 5318
rect 40427 5318 40456 5327
rect 40970 5318 41048 6276
rect 41136 6264 41760 6296
rect 41868 6331 41934 6342
rect 41868 6297 41884 6331
rect 41918 6297 41934 6331
rect 41868 6286 41934 6297
rect 42020 6294 42054 6440
rect 42202 6438 42260 6440
rect 42458 6459 42526 6464
rect 42458 6456 42486 6459
rect 42458 6404 42466 6456
rect 42520 6425 42526 6459
rect 42518 6404 42526 6425
rect 42256 6383 42346 6404
rect 42458 6398 42526 6404
rect 42256 6349 42283 6383
rect 42317 6349 42346 6383
rect 42480 6378 42526 6398
rect 42568 6531 42614 6578
rect 42568 6497 42574 6531
rect 42608 6497 42614 6531
rect 42568 6459 42614 6497
rect 42568 6425 42574 6459
rect 42608 6425 42614 6459
rect 42568 6404 42614 6425
rect 43722 6531 43768 6578
rect 43722 6497 43728 6531
rect 43762 6497 43768 6531
rect 43722 6459 43768 6497
rect 43722 6425 43728 6459
rect 43762 6425 43768 6459
rect 43810 6531 43856 6578
rect 43810 6497 43816 6531
rect 43850 6497 43856 6531
rect 43810 6459 43856 6497
rect 43910 6500 43970 6732
rect 43998 7022 44038 7056
rect 44072 7022 44078 7056
rect 43998 6984 44078 7022
rect 44118 7062 44184 7068
rect 44118 7010 44124 7062
rect 44176 7010 44184 7062
rect 44118 7004 44184 7010
rect 44224 7056 44326 7068
rect 44224 7022 44230 7056
rect 44264 7022 44326 7056
rect 43998 6950 44038 6984
rect 44072 6950 44078 6984
rect 43998 6938 44078 6950
rect 44128 6984 44174 7004
rect 44128 6950 44134 6984
rect 44168 6950 44174 6984
rect 44128 6938 44174 6950
rect 44224 6984 44326 7022
rect 44224 6950 44230 6984
rect 44264 6950 44326 6984
rect 44224 6938 44326 6950
rect 43998 6738 44044 6938
rect 44074 6900 44132 6910
rect 44074 6866 44086 6900
rect 44120 6866 44132 6900
rect 44074 6848 44132 6866
rect 44276 6858 44326 6938
rect 44692 6916 44776 7186
rect 44434 6906 44492 6912
rect 44426 6900 44500 6906
rect 44186 6819 44244 6836
rect 44186 6785 44198 6819
rect 44232 6785 44244 6819
rect 44186 6770 44244 6785
rect 44276 6792 44346 6858
rect 44426 6848 44437 6900
rect 44489 6848 44500 6900
rect 44426 6842 44500 6848
rect 44568 6890 44844 6916
rect 45432 6910 45530 7186
rect 44568 6885 44669 6890
rect 44721 6885 44844 6890
rect 44568 6851 44597 6885
rect 44631 6851 44669 6885
rect 44723 6851 44781 6885
rect 44815 6851 44844 6885
rect 44434 6834 44492 6842
rect 44568 6838 44669 6851
rect 44721 6838 44844 6851
rect 44568 6820 44844 6838
rect 44908 6879 45530 6910
rect 44908 6845 44937 6879
rect 44971 6845 45029 6879
rect 45063 6845 45121 6879
rect 45155 6877 45530 6879
rect 45155 6845 45283 6877
rect 44908 6843 45283 6845
rect 45317 6843 45375 6877
rect 45409 6843 45467 6877
rect 45501 6843 45530 6877
rect 45792 7140 46112 7158
rect 45792 7106 46064 7140
rect 46098 7106 46112 7140
rect 45792 7096 46112 7106
rect 44908 6812 45530 6843
rect 45670 6868 45746 6874
rect 45670 6816 45686 6868
rect 45738 6816 45746 6868
rect 45670 6810 45746 6816
rect 44276 6738 44326 6792
rect 45792 6766 45852 7096
rect 45914 7056 45960 7068
rect 43998 6691 44094 6738
rect 43998 6657 44054 6691
rect 44088 6657 44094 6691
rect 43998 6619 44094 6657
rect 43998 6585 44054 6619
rect 44088 6585 44094 6619
rect 44144 6691 44190 6738
rect 44144 6657 44150 6691
rect 44184 6657 44190 6691
rect 44144 6619 44190 6657
rect 44144 6598 44150 6619
rect 43998 6538 44094 6585
rect 44134 6590 44150 6598
rect 44184 6598 44190 6619
rect 44240 6691 44326 6738
rect 45324 6746 45852 6766
rect 45324 6712 45336 6746
rect 45370 6732 45852 6746
rect 45370 6712 45382 6732
rect 45324 6698 45382 6712
rect 44240 6657 44246 6691
rect 44280 6657 44326 6691
rect 44240 6619 44326 6657
rect 44184 6590 44200 6598
rect 44134 6538 44142 6590
rect 44194 6538 44200 6590
rect 44240 6585 44246 6619
rect 44280 6585 44326 6619
rect 44402 6659 44468 6672
rect 44402 6625 44418 6659
rect 44452 6625 44468 6659
rect 44796 6652 44864 6654
rect 44402 6614 44468 6625
rect 44712 6648 44864 6652
rect 44712 6642 44805 6648
rect 44712 6608 44732 6642
rect 44766 6608 44805 6642
rect 44712 6602 44805 6608
rect 44796 6596 44805 6602
rect 44857 6596 44864 6648
rect 44796 6590 44864 6596
rect 44894 6636 44968 6660
rect 44894 6602 44922 6636
rect 44956 6602 44968 6636
rect 44240 6542 44326 6585
rect 44894 6582 44968 6602
rect 45092 6652 45164 6664
rect 45092 6600 45103 6652
rect 45155 6600 45164 6652
rect 45638 6659 45704 6668
rect 45638 6625 45654 6659
rect 45688 6625 45704 6659
rect 45638 6612 45704 6625
rect 45092 6596 45164 6600
rect 44240 6538 44286 6542
rect 44134 6530 44200 6538
rect 44368 6531 44414 6578
rect 43910 6491 44148 6500
rect 43910 6468 44102 6491
rect 43810 6442 43816 6459
rect 42568 6376 42640 6404
rect 43722 6378 43768 6425
rect 43798 6436 43816 6442
rect 43850 6442 43856 6459
rect 43908 6457 44102 6468
rect 44136 6457 44148 6491
rect 44368 6497 44374 6531
rect 44408 6497 44414 6531
rect 44368 6464 44414 6497
rect 43850 6436 43864 6442
rect 43798 6384 43804 6436
rect 43856 6384 43864 6436
rect 43798 6378 43864 6384
rect 43908 6440 44148 6457
rect 42256 6328 42346 6349
rect 42514 6331 42580 6340
rect 42514 6297 42530 6331
rect 42564 6297 42580 6331
rect 42514 6294 42580 6297
rect 42020 6266 42580 6294
rect 41924 6210 41992 6224
rect 41924 6176 41942 6210
rect 41976 6176 41992 6210
rect 41924 6166 41992 6176
rect 41964 5862 41992 6166
rect 42020 6084 42054 6266
rect 42352 6200 42424 6212
rect 42352 6148 42362 6200
rect 42414 6148 42424 6200
rect 42352 6136 42424 6148
rect 42276 6084 42340 6102
rect 42020 6050 42292 6084
rect 42326 6050 42340 6084
rect 42276 6040 42340 6050
rect 42612 6026 42640 6376
rect 42680 6342 42956 6372
rect 42680 6341 42712 6342
rect 42764 6341 42956 6342
rect 42680 6307 42709 6341
rect 42764 6307 42801 6341
rect 42835 6307 42893 6341
rect 42927 6307 42956 6341
rect 42680 6290 42712 6307
rect 42764 6290 42956 6307
rect 42680 6276 42956 6290
rect 43024 6348 43648 6366
rect 43024 6335 43566 6348
rect 43024 6301 43055 6335
rect 43089 6301 43147 6335
rect 43181 6301 43239 6335
rect 43273 6333 43566 6335
rect 43618 6333 43648 6348
rect 43273 6301 43401 6333
rect 43024 6299 43401 6301
rect 43435 6299 43493 6333
rect 43527 6299 43566 6333
rect 43619 6299 43648 6333
rect 43024 6296 43566 6299
rect 43618 6296 43648 6299
rect 42730 6084 42796 6090
rect 42730 6032 42736 6084
rect 42788 6032 42796 6084
rect 42730 6026 42796 6032
rect 42386 6012 42640 6026
rect 42142 6000 42188 6012
rect 41688 5834 41992 5862
rect 42108 5966 42148 6000
rect 42182 5966 42188 6000
rect 42108 5928 42188 5966
rect 42228 6006 42294 6012
rect 42228 5954 42234 6006
rect 42286 5954 42294 6006
rect 42228 5948 42294 5954
rect 42334 6000 42640 6012
rect 42334 5966 42340 6000
rect 42374 5998 42640 6000
rect 42374 5966 42436 5998
rect 42108 5894 42148 5928
rect 42182 5894 42188 5928
rect 42108 5882 42188 5894
rect 42238 5928 42284 5948
rect 42238 5894 42244 5928
rect 42278 5894 42284 5928
rect 42238 5882 42284 5894
rect 42334 5928 42436 5966
rect 42334 5894 42340 5928
rect 42374 5894 42436 5928
rect 42334 5882 42436 5894
rect 42556 5951 42790 5960
rect 42556 5899 42562 5951
rect 42614 5932 42738 5951
rect 42614 5899 42620 5932
rect 42556 5892 42620 5899
rect 42732 5899 42738 5932
rect 42790 5899 42796 5932
rect 42732 5892 42796 5899
rect 41688 5831 41964 5834
rect 41688 5797 41717 5831
rect 41751 5797 41809 5831
rect 41843 5797 41901 5831
rect 41935 5797 41964 5831
rect 41688 5766 41964 5797
rect 41794 5718 41858 5724
rect 41794 5666 41800 5718
rect 41852 5666 41858 5718
rect 41794 5660 41858 5666
rect 42108 5682 42154 5882
rect 42184 5844 42242 5854
rect 42184 5810 42196 5844
rect 42230 5810 42242 5844
rect 42184 5792 42242 5810
rect 42296 5763 42354 5780
rect 42296 5729 42308 5763
rect 42342 5729 42354 5763
rect 42296 5714 42354 5729
rect 42386 5682 42436 5882
rect 42502 5831 42778 5862
rect 42502 5797 42531 5831
rect 42565 5797 42623 5831
rect 42657 5797 42715 5831
rect 42749 5797 42778 5831
rect 42502 5766 42778 5797
rect 42108 5635 42204 5682
rect 41706 5602 41770 5608
rect 41706 5550 41712 5602
rect 41764 5550 41770 5602
rect 41706 5544 41770 5550
rect 41876 5592 41946 5610
rect 41876 5558 41897 5592
rect 41931 5558 41946 5592
rect 41876 5550 41946 5558
rect 42108 5601 42164 5635
rect 42198 5601 42204 5635
rect 42108 5563 42204 5601
rect 41876 5514 41904 5550
rect 42108 5529 42164 5563
rect 42198 5529 42204 5563
rect 42254 5635 42300 5682
rect 42254 5601 42260 5635
rect 42294 5601 42300 5635
rect 42254 5563 42300 5601
rect 42254 5542 42260 5563
rect 42108 5514 42204 5529
rect 41876 5482 42204 5514
rect 42244 5534 42260 5542
rect 42294 5542 42300 5563
rect 42350 5635 42436 5682
rect 42608 5716 42676 5726
rect 42608 5664 42616 5716
rect 42668 5664 42676 5716
rect 42608 5658 42676 5664
rect 42350 5601 42356 5635
rect 42390 5601 42436 5635
rect 42350 5563 42436 5601
rect 42294 5534 42310 5542
rect 42244 5482 42252 5534
rect 42304 5482 42310 5534
rect 42350 5529 42356 5563
rect 42390 5529 42436 5563
rect 42518 5604 42586 5610
rect 42518 5552 42524 5604
rect 42576 5552 42586 5604
rect 42518 5546 42586 5552
rect 42692 5590 42758 5602
rect 42692 5556 42709 5590
rect 42743 5556 42758 5590
rect 42692 5548 42758 5556
rect 42350 5510 42436 5529
rect 42730 5510 42758 5548
rect 42350 5482 42758 5510
rect 42244 5474 42310 5482
rect 42392 5478 42758 5482
rect 42196 5435 42258 5444
rect 42196 5401 42212 5435
rect 42246 5401 42258 5435
rect 42196 5384 42258 5401
rect 42200 5382 42258 5384
rect 42254 5327 42344 5348
rect 42254 5318 42281 5327
rect 40427 5293 42281 5318
rect 42315 5318 42344 5327
rect 42858 5318 42936 6276
rect 43024 6264 43648 6296
rect 43756 6331 43822 6342
rect 43756 6297 43772 6331
rect 43806 6297 43822 6331
rect 43756 6286 43822 6297
rect 43908 6294 43942 6440
rect 44090 6438 44148 6440
rect 44346 6459 44414 6464
rect 44346 6456 44374 6459
rect 44346 6404 44354 6456
rect 44408 6425 44414 6459
rect 44406 6404 44414 6425
rect 44144 6383 44234 6404
rect 44346 6398 44414 6404
rect 44144 6349 44171 6383
rect 44205 6349 44234 6383
rect 44368 6378 44414 6398
rect 44456 6531 44502 6578
rect 44456 6497 44462 6531
rect 44496 6497 44502 6531
rect 44456 6459 44502 6497
rect 44456 6425 44462 6459
rect 44496 6425 44502 6459
rect 44456 6404 44502 6425
rect 45604 6531 45650 6578
rect 45604 6497 45610 6531
rect 45644 6497 45650 6531
rect 45604 6459 45650 6497
rect 45604 6425 45610 6459
rect 45644 6425 45650 6459
rect 45692 6531 45738 6578
rect 45692 6497 45698 6531
rect 45732 6497 45738 6531
rect 45692 6459 45738 6497
rect 45792 6500 45852 6732
rect 45880 7022 45920 7056
rect 45954 7022 45960 7056
rect 45880 6984 45960 7022
rect 46000 7062 46066 7068
rect 46000 7010 46006 7062
rect 46058 7010 46066 7062
rect 46000 7004 46066 7010
rect 46106 7056 46208 7068
rect 46106 7022 46112 7056
rect 46146 7022 46208 7056
rect 45880 6950 45920 6984
rect 45954 6950 45960 6984
rect 45880 6938 45960 6950
rect 46010 6984 46056 7004
rect 46010 6950 46016 6984
rect 46050 6950 46056 6984
rect 46010 6938 46056 6950
rect 46106 6984 46208 7022
rect 46106 6950 46112 6984
rect 46146 6950 46208 6984
rect 46106 6938 46208 6950
rect 45880 6738 45926 6938
rect 45956 6900 46014 6910
rect 45956 6866 45968 6900
rect 46002 6866 46014 6900
rect 45956 6848 46014 6866
rect 46158 6858 46208 6938
rect 46574 6916 46658 7186
rect 46316 6906 46374 6912
rect 46308 6900 46382 6906
rect 46068 6819 46126 6836
rect 46068 6785 46080 6819
rect 46114 6785 46126 6819
rect 46068 6770 46126 6785
rect 46158 6792 46228 6858
rect 46308 6848 46319 6900
rect 46371 6848 46382 6900
rect 46308 6842 46382 6848
rect 46450 6890 46726 6916
rect 47320 6910 47418 7186
rect 46450 6885 46551 6890
rect 46603 6885 46726 6890
rect 46450 6851 46479 6885
rect 46513 6851 46551 6885
rect 46605 6851 46663 6885
rect 46697 6851 46726 6885
rect 46316 6834 46374 6842
rect 46450 6838 46551 6851
rect 46603 6838 46726 6851
rect 46450 6820 46726 6838
rect 46796 6879 47418 6910
rect 46796 6845 46825 6879
rect 46859 6845 46917 6879
rect 46951 6845 47009 6879
rect 47043 6877 47418 6879
rect 47043 6845 47171 6877
rect 46796 6843 47171 6845
rect 47205 6843 47263 6877
rect 47297 6843 47355 6877
rect 47389 6843 47418 6877
rect 47680 7140 48000 7158
rect 47680 7106 47952 7140
rect 47986 7106 48000 7140
rect 47680 7096 48000 7106
rect 46796 6812 47418 6843
rect 47558 6868 47634 6874
rect 47558 6816 47574 6868
rect 47626 6816 47634 6868
rect 47558 6810 47634 6816
rect 46158 6738 46208 6792
rect 47680 6766 47740 7096
rect 47802 7056 47848 7068
rect 45880 6691 45976 6738
rect 45880 6657 45936 6691
rect 45970 6657 45976 6691
rect 45880 6619 45976 6657
rect 45880 6585 45936 6619
rect 45970 6585 45976 6619
rect 46026 6691 46072 6738
rect 46026 6657 46032 6691
rect 46066 6657 46072 6691
rect 46026 6619 46072 6657
rect 46026 6598 46032 6619
rect 45880 6538 45976 6585
rect 46016 6590 46032 6598
rect 46066 6598 46072 6619
rect 46122 6691 46208 6738
rect 47212 6746 47740 6766
rect 47212 6712 47224 6746
rect 47258 6732 47740 6746
rect 47258 6712 47270 6732
rect 47212 6698 47270 6712
rect 46122 6657 46128 6691
rect 46162 6657 46208 6691
rect 46122 6619 46208 6657
rect 46066 6590 46082 6598
rect 46016 6538 46024 6590
rect 46076 6538 46082 6590
rect 46122 6585 46128 6619
rect 46162 6585 46208 6619
rect 46284 6659 46350 6672
rect 46284 6625 46300 6659
rect 46334 6625 46350 6659
rect 46678 6652 46746 6654
rect 46284 6614 46350 6625
rect 46594 6648 46746 6652
rect 46594 6642 46687 6648
rect 46594 6608 46614 6642
rect 46648 6608 46687 6642
rect 46594 6602 46687 6608
rect 46678 6596 46687 6602
rect 46739 6596 46746 6648
rect 46678 6590 46746 6596
rect 46782 6636 46856 6660
rect 46782 6602 46810 6636
rect 46844 6602 46856 6636
rect 46122 6542 46208 6585
rect 46782 6582 46856 6602
rect 46980 6652 47052 6664
rect 46980 6600 46991 6652
rect 47043 6600 47052 6652
rect 47526 6659 47592 6668
rect 47526 6625 47542 6659
rect 47576 6625 47592 6659
rect 47526 6612 47592 6625
rect 46980 6596 47052 6600
rect 46122 6538 46168 6542
rect 46016 6530 46082 6538
rect 46250 6531 46296 6578
rect 45792 6491 46030 6500
rect 45792 6468 45984 6491
rect 45692 6442 45698 6459
rect 44456 6376 44528 6404
rect 45604 6378 45650 6425
rect 45680 6436 45698 6442
rect 45732 6442 45738 6459
rect 45790 6457 45984 6468
rect 46018 6457 46030 6491
rect 46250 6497 46256 6531
rect 46290 6497 46296 6531
rect 46250 6464 46296 6497
rect 45732 6436 45746 6442
rect 45680 6384 45686 6436
rect 45738 6384 45746 6436
rect 45680 6378 45746 6384
rect 45790 6440 46030 6457
rect 44144 6328 44234 6349
rect 44402 6331 44468 6340
rect 44402 6297 44418 6331
rect 44452 6297 44468 6331
rect 44402 6294 44468 6297
rect 43908 6266 44468 6294
rect 43812 6210 43880 6224
rect 43812 6176 43830 6210
rect 43864 6176 43880 6210
rect 43812 6166 43880 6176
rect 43852 5862 43880 6166
rect 43908 6084 43942 6266
rect 44240 6200 44312 6212
rect 44240 6148 44250 6200
rect 44302 6148 44312 6200
rect 44240 6136 44312 6148
rect 44164 6084 44228 6102
rect 43908 6050 44180 6084
rect 44214 6050 44228 6084
rect 44164 6040 44228 6050
rect 44500 6026 44528 6376
rect 44568 6342 44844 6372
rect 44568 6341 44600 6342
rect 44652 6341 44844 6342
rect 44568 6307 44597 6341
rect 44652 6307 44689 6341
rect 44723 6307 44781 6341
rect 44815 6307 44844 6341
rect 44568 6290 44600 6307
rect 44652 6290 44844 6307
rect 44568 6276 44844 6290
rect 44906 6348 45530 6366
rect 44906 6335 45448 6348
rect 44906 6301 44937 6335
rect 44971 6301 45029 6335
rect 45063 6301 45121 6335
rect 45155 6333 45448 6335
rect 45500 6333 45530 6348
rect 45155 6301 45283 6333
rect 44906 6299 45283 6301
rect 45317 6299 45375 6333
rect 45409 6299 45448 6333
rect 45501 6299 45530 6333
rect 44906 6296 45448 6299
rect 45500 6296 45530 6299
rect 44618 6084 44684 6090
rect 44618 6032 44624 6084
rect 44676 6032 44684 6084
rect 44618 6026 44684 6032
rect 44274 6012 44528 6026
rect 44030 6000 44076 6012
rect 43576 5834 43880 5862
rect 43996 5966 44036 6000
rect 44070 5966 44076 6000
rect 43996 5928 44076 5966
rect 44116 6006 44182 6012
rect 44116 5954 44122 6006
rect 44174 5954 44182 6006
rect 44116 5948 44182 5954
rect 44222 6000 44528 6012
rect 44222 5966 44228 6000
rect 44262 5998 44528 6000
rect 44262 5966 44324 5998
rect 43996 5894 44036 5928
rect 44070 5894 44076 5928
rect 43996 5882 44076 5894
rect 44126 5928 44172 5948
rect 44126 5894 44132 5928
rect 44166 5894 44172 5928
rect 44126 5882 44172 5894
rect 44222 5928 44324 5966
rect 44222 5894 44228 5928
rect 44262 5894 44324 5928
rect 44222 5882 44324 5894
rect 44444 5951 44678 5960
rect 44444 5899 44450 5951
rect 44502 5932 44626 5951
rect 44502 5899 44508 5932
rect 44444 5892 44508 5899
rect 44620 5899 44626 5932
rect 44678 5899 44684 5932
rect 44620 5892 44684 5899
rect 43576 5831 43852 5834
rect 43576 5797 43605 5831
rect 43639 5797 43697 5831
rect 43731 5797 43789 5831
rect 43823 5797 43852 5831
rect 43576 5766 43852 5797
rect 43682 5718 43746 5724
rect 43682 5666 43688 5718
rect 43740 5666 43746 5718
rect 43682 5660 43746 5666
rect 43996 5682 44042 5882
rect 44072 5844 44130 5854
rect 44072 5810 44084 5844
rect 44118 5810 44130 5844
rect 44072 5792 44130 5810
rect 44184 5763 44242 5780
rect 44184 5729 44196 5763
rect 44230 5729 44242 5763
rect 44184 5714 44242 5729
rect 44274 5682 44324 5882
rect 44390 5831 44666 5862
rect 44390 5797 44419 5831
rect 44453 5797 44511 5831
rect 44545 5797 44603 5831
rect 44637 5797 44666 5831
rect 44390 5766 44666 5797
rect 43996 5635 44092 5682
rect 43594 5602 43658 5608
rect 43594 5550 43600 5602
rect 43652 5550 43658 5602
rect 43594 5544 43658 5550
rect 43764 5592 43834 5610
rect 43764 5558 43785 5592
rect 43819 5558 43834 5592
rect 43764 5550 43834 5558
rect 43996 5601 44052 5635
rect 44086 5601 44092 5635
rect 43996 5563 44092 5601
rect 43764 5514 43792 5550
rect 43996 5529 44052 5563
rect 44086 5529 44092 5563
rect 44142 5635 44188 5682
rect 44142 5601 44148 5635
rect 44182 5601 44188 5635
rect 44142 5563 44188 5601
rect 44142 5542 44148 5563
rect 43996 5514 44092 5529
rect 43764 5482 44092 5514
rect 44132 5534 44148 5542
rect 44182 5542 44188 5563
rect 44238 5635 44324 5682
rect 44496 5716 44564 5726
rect 44496 5664 44504 5716
rect 44556 5664 44564 5716
rect 44496 5658 44564 5664
rect 44238 5601 44244 5635
rect 44278 5601 44324 5635
rect 44238 5563 44324 5601
rect 44182 5534 44198 5542
rect 44132 5482 44140 5534
rect 44192 5482 44198 5534
rect 44238 5529 44244 5563
rect 44278 5529 44324 5563
rect 44406 5604 44474 5610
rect 44406 5552 44412 5604
rect 44464 5552 44474 5604
rect 44406 5546 44474 5552
rect 44580 5590 44646 5602
rect 44580 5556 44597 5590
rect 44631 5556 44646 5590
rect 44580 5548 44646 5556
rect 44238 5510 44324 5529
rect 44618 5510 44646 5548
rect 44238 5482 44646 5510
rect 44132 5474 44198 5482
rect 44280 5478 44646 5482
rect 44084 5435 44146 5444
rect 44084 5401 44100 5435
rect 44134 5401 44146 5435
rect 44084 5384 44146 5401
rect 44088 5382 44146 5384
rect 44142 5327 44232 5348
rect 44142 5318 44169 5327
rect 42315 5293 44169 5318
rect 44203 5318 44232 5327
rect 44746 5318 44824 6276
rect 44906 6264 45530 6296
rect 45638 6331 45704 6342
rect 45638 6297 45654 6331
rect 45688 6297 45704 6331
rect 45638 6286 45704 6297
rect 45790 6294 45824 6440
rect 45972 6438 46030 6440
rect 46228 6459 46296 6464
rect 46228 6456 46256 6459
rect 46228 6404 46236 6456
rect 46290 6425 46296 6459
rect 46288 6404 46296 6425
rect 46026 6383 46116 6404
rect 46228 6398 46296 6404
rect 46026 6349 46053 6383
rect 46087 6349 46116 6383
rect 46250 6378 46296 6398
rect 46338 6531 46384 6578
rect 46338 6497 46344 6531
rect 46378 6497 46384 6531
rect 46338 6459 46384 6497
rect 46338 6425 46344 6459
rect 46378 6425 46384 6459
rect 46338 6404 46384 6425
rect 47492 6531 47538 6578
rect 47492 6497 47498 6531
rect 47532 6497 47538 6531
rect 47492 6459 47538 6497
rect 47492 6425 47498 6459
rect 47532 6425 47538 6459
rect 47580 6531 47626 6578
rect 47580 6497 47586 6531
rect 47620 6497 47626 6531
rect 47580 6459 47626 6497
rect 47680 6500 47740 6732
rect 47768 7022 47808 7056
rect 47842 7022 47848 7056
rect 47768 6984 47848 7022
rect 47888 7062 47954 7068
rect 47888 7010 47894 7062
rect 47946 7010 47954 7062
rect 47888 7004 47954 7010
rect 47994 7056 48096 7068
rect 47994 7022 48000 7056
rect 48034 7022 48096 7056
rect 47768 6950 47808 6984
rect 47842 6950 47848 6984
rect 47768 6938 47848 6950
rect 47898 6984 47944 7004
rect 47898 6950 47904 6984
rect 47938 6950 47944 6984
rect 47898 6938 47944 6950
rect 47994 6984 48096 7022
rect 47994 6950 48000 6984
rect 48034 6950 48096 6984
rect 47994 6938 48096 6950
rect 47768 6738 47814 6938
rect 47844 6900 47902 6910
rect 47844 6866 47856 6900
rect 47890 6866 47902 6900
rect 47844 6848 47902 6866
rect 48046 6858 48096 6938
rect 48462 6916 48546 7186
rect 48204 6906 48262 6912
rect 48196 6900 48270 6906
rect 47956 6819 48014 6836
rect 47956 6785 47968 6819
rect 48002 6785 48014 6819
rect 47956 6770 48014 6785
rect 48046 6792 48116 6858
rect 48196 6848 48207 6900
rect 48259 6848 48270 6900
rect 48196 6842 48270 6848
rect 48338 6890 48614 6916
rect 49208 6910 49306 7186
rect 48338 6885 48439 6890
rect 48491 6885 48614 6890
rect 48338 6851 48367 6885
rect 48401 6851 48439 6885
rect 48493 6851 48551 6885
rect 48585 6851 48614 6885
rect 48204 6834 48262 6842
rect 48338 6838 48439 6851
rect 48491 6838 48614 6851
rect 48338 6820 48614 6838
rect 48684 6879 49306 6910
rect 48684 6845 48713 6879
rect 48747 6845 48805 6879
rect 48839 6845 48897 6879
rect 48931 6877 49306 6879
rect 48931 6845 49059 6877
rect 48684 6843 49059 6845
rect 49093 6843 49151 6877
rect 49185 6843 49243 6877
rect 49277 6843 49306 6877
rect 49568 7140 49888 7158
rect 49568 7106 49840 7140
rect 49874 7106 49888 7140
rect 49568 7096 49888 7106
rect 48684 6812 49306 6843
rect 49446 6868 49522 6874
rect 49446 6816 49462 6868
rect 49514 6816 49522 6868
rect 49446 6810 49522 6816
rect 48046 6738 48096 6792
rect 49568 6766 49628 7096
rect 49690 7056 49736 7068
rect 47768 6691 47864 6738
rect 47768 6657 47824 6691
rect 47858 6657 47864 6691
rect 47768 6619 47864 6657
rect 47768 6585 47824 6619
rect 47858 6585 47864 6619
rect 47914 6691 47960 6738
rect 47914 6657 47920 6691
rect 47954 6657 47960 6691
rect 47914 6619 47960 6657
rect 47914 6598 47920 6619
rect 47768 6538 47864 6585
rect 47904 6590 47920 6598
rect 47954 6598 47960 6619
rect 48010 6691 48096 6738
rect 49100 6746 49628 6766
rect 49100 6712 49112 6746
rect 49146 6732 49628 6746
rect 49146 6712 49158 6732
rect 49100 6698 49158 6712
rect 48010 6657 48016 6691
rect 48050 6657 48096 6691
rect 48010 6619 48096 6657
rect 47954 6590 47970 6598
rect 47904 6538 47912 6590
rect 47964 6538 47970 6590
rect 48010 6585 48016 6619
rect 48050 6585 48096 6619
rect 48172 6659 48238 6672
rect 48172 6625 48188 6659
rect 48222 6625 48238 6659
rect 48566 6652 48634 6654
rect 48172 6614 48238 6625
rect 48482 6648 48634 6652
rect 48482 6642 48575 6648
rect 48482 6608 48502 6642
rect 48536 6608 48575 6642
rect 48482 6602 48575 6608
rect 48566 6596 48575 6602
rect 48627 6596 48634 6648
rect 48566 6590 48634 6596
rect 48670 6636 48744 6660
rect 48670 6602 48698 6636
rect 48732 6602 48744 6636
rect 48010 6542 48096 6585
rect 48670 6582 48744 6602
rect 48868 6652 48940 6664
rect 48868 6600 48879 6652
rect 48931 6600 48940 6652
rect 49414 6659 49480 6668
rect 49414 6625 49430 6659
rect 49464 6625 49480 6659
rect 49414 6612 49480 6625
rect 48868 6596 48940 6600
rect 48010 6538 48056 6542
rect 47904 6530 47970 6538
rect 48138 6531 48184 6578
rect 47680 6491 47918 6500
rect 47680 6468 47872 6491
rect 47580 6442 47586 6459
rect 46338 6376 46410 6404
rect 47492 6378 47538 6425
rect 47568 6436 47586 6442
rect 47620 6442 47626 6459
rect 47678 6457 47872 6468
rect 47906 6457 47918 6491
rect 48138 6497 48144 6531
rect 48178 6497 48184 6531
rect 48138 6464 48184 6497
rect 47620 6436 47634 6442
rect 47568 6384 47574 6436
rect 47626 6384 47634 6436
rect 47568 6378 47634 6384
rect 47678 6440 47918 6457
rect 46026 6328 46116 6349
rect 46284 6331 46350 6340
rect 46284 6297 46300 6331
rect 46334 6297 46350 6331
rect 46284 6294 46350 6297
rect 45790 6266 46350 6294
rect 45694 6210 45762 6224
rect 45694 6176 45712 6210
rect 45746 6176 45762 6210
rect 45694 6166 45762 6176
rect 45734 5862 45762 6166
rect 45790 6084 45824 6266
rect 46122 6200 46194 6212
rect 46122 6148 46132 6200
rect 46184 6148 46194 6200
rect 46122 6136 46194 6148
rect 46046 6084 46110 6102
rect 45790 6050 46062 6084
rect 46096 6050 46110 6084
rect 46046 6040 46110 6050
rect 46382 6026 46410 6376
rect 46450 6342 46726 6372
rect 46450 6341 46482 6342
rect 46534 6341 46726 6342
rect 46450 6307 46479 6341
rect 46534 6307 46571 6341
rect 46605 6307 46663 6341
rect 46697 6307 46726 6341
rect 46450 6290 46482 6307
rect 46534 6290 46726 6307
rect 46450 6276 46726 6290
rect 46794 6348 47418 6366
rect 46794 6335 47336 6348
rect 46794 6301 46825 6335
rect 46859 6301 46917 6335
rect 46951 6301 47009 6335
rect 47043 6333 47336 6335
rect 47388 6333 47418 6348
rect 47043 6301 47171 6333
rect 46794 6299 47171 6301
rect 47205 6299 47263 6333
rect 47297 6299 47336 6333
rect 47389 6299 47418 6333
rect 46794 6296 47336 6299
rect 47388 6296 47418 6299
rect 46500 6084 46566 6090
rect 46500 6032 46506 6084
rect 46558 6032 46566 6084
rect 46500 6026 46566 6032
rect 46156 6012 46410 6026
rect 45912 6000 45958 6012
rect 45458 5834 45762 5862
rect 45878 5966 45918 6000
rect 45952 5966 45958 6000
rect 45878 5928 45958 5966
rect 45998 6006 46064 6012
rect 45998 5954 46004 6006
rect 46056 5954 46064 6006
rect 45998 5948 46064 5954
rect 46104 6000 46410 6012
rect 46104 5966 46110 6000
rect 46144 5998 46410 6000
rect 46144 5966 46206 5998
rect 45878 5894 45918 5928
rect 45952 5894 45958 5928
rect 45878 5882 45958 5894
rect 46008 5928 46054 5948
rect 46008 5894 46014 5928
rect 46048 5894 46054 5928
rect 46008 5882 46054 5894
rect 46104 5928 46206 5966
rect 46104 5894 46110 5928
rect 46144 5894 46206 5928
rect 46104 5882 46206 5894
rect 46326 5951 46560 5960
rect 46326 5899 46332 5951
rect 46384 5932 46508 5951
rect 46384 5899 46390 5932
rect 46326 5892 46390 5899
rect 46502 5899 46508 5932
rect 46560 5899 46566 5932
rect 46502 5892 46566 5899
rect 45458 5831 45734 5834
rect 45458 5797 45487 5831
rect 45521 5797 45579 5831
rect 45613 5797 45671 5831
rect 45705 5797 45734 5831
rect 45458 5766 45734 5797
rect 45564 5718 45628 5724
rect 45564 5666 45570 5718
rect 45622 5666 45628 5718
rect 45564 5660 45628 5666
rect 45878 5682 45924 5882
rect 45954 5844 46012 5854
rect 45954 5810 45966 5844
rect 46000 5810 46012 5844
rect 45954 5792 46012 5810
rect 46066 5763 46124 5780
rect 46066 5729 46078 5763
rect 46112 5729 46124 5763
rect 46066 5714 46124 5729
rect 46156 5682 46206 5882
rect 46272 5831 46548 5862
rect 46272 5797 46301 5831
rect 46335 5797 46393 5831
rect 46427 5797 46485 5831
rect 46519 5797 46548 5831
rect 46272 5766 46548 5797
rect 45878 5635 45974 5682
rect 45476 5602 45540 5608
rect 45476 5550 45482 5602
rect 45534 5550 45540 5602
rect 45476 5544 45540 5550
rect 45646 5592 45716 5610
rect 45646 5558 45667 5592
rect 45701 5558 45716 5592
rect 45646 5550 45716 5558
rect 45878 5601 45934 5635
rect 45968 5601 45974 5635
rect 45878 5563 45974 5601
rect 45646 5514 45674 5550
rect 45878 5529 45934 5563
rect 45968 5529 45974 5563
rect 46024 5635 46070 5682
rect 46024 5601 46030 5635
rect 46064 5601 46070 5635
rect 46024 5563 46070 5601
rect 46024 5542 46030 5563
rect 45878 5514 45974 5529
rect 45646 5482 45974 5514
rect 46014 5534 46030 5542
rect 46064 5542 46070 5563
rect 46120 5635 46206 5682
rect 46378 5716 46446 5726
rect 46378 5664 46386 5716
rect 46438 5664 46446 5716
rect 46378 5658 46446 5664
rect 46120 5601 46126 5635
rect 46160 5601 46206 5635
rect 46120 5563 46206 5601
rect 46064 5534 46080 5542
rect 46014 5482 46022 5534
rect 46074 5482 46080 5534
rect 46120 5529 46126 5563
rect 46160 5529 46206 5563
rect 46288 5604 46356 5610
rect 46288 5552 46294 5604
rect 46346 5552 46356 5604
rect 46288 5546 46356 5552
rect 46462 5590 46528 5602
rect 46462 5556 46479 5590
rect 46513 5556 46528 5590
rect 46462 5548 46528 5556
rect 46120 5510 46206 5529
rect 46500 5510 46528 5548
rect 46120 5482 46528 5510
rect 46014 5474 46080 5482
rect 46162 5478 46528 5482
rect 45966 5435 46028 5444
rect 45966 5401 45982 5435
rect 46016 5401 46028 5435
rect 45966 5384 46028 5401
rect 45970 5382 46028 5384
rect 46024 5327 46114 5348
rect 46024 5318 46051 5327
rect 44203 5293 46051 5318
rect 46085 5318 46114 5327
rect 46628 5318 46706 6276
rect 46794 6264 47418 6296
rect 47526 6331 47592 6342
rect 47526 6297 47542 6331
rect 47576 6297 47592 6331
rect 47526 6286 47592 6297
rect 47678 6294 47712 6440
rect 47860 6438 47918 6440
rect 48116 6459 48184 6464
rect 48116 6456 48144 6459
rect 48116 6404 48124 6456
rect 48178 6425 48184 6459
rect 48176 6404 48184 6425
rect 47914 6383 48004 6404
rect 48116 6398 48184 6404
rect 47914 6349 47941 6383
rect 47975 6349 48004 6383
rect 48138 6378 48184 6398
rect 48226 6531 48272 6578
rect 48226 6497 48232 6531
rect 48266 6497 48272 6531
rect 48226 6459 48272 6497
rect 48226 6425 48232 6459
rect 48266 6425 48272 6459
rect 48226 6404 48272 6425
rect 49380 6531 49426 6578
rect 49380 6497 49386 6531
rect 49420 6497 49426 6531
rect 49380 6459 49426 6497
rect 49380 6425 49386 6459
rect 49420 6425 49426 6459
rect 49468 6531 49514 6578
rect 49468 6497 49474 6531
rect 49508 6497 49514 6531
rect 49468 6459 49514 6497
rect 49568 6500 49628 6732
rect 49656 7022 49696 7056
rect 49730 7022 49736 7056
rect 49656 6984 49736 7022
rect 49776 7062 49842 7068
rect 49776 7010 49782 7062
rect 49834 7010 49842 7062
rect 49776 7004 49842 7010
rect 49882 7056 49984 7068
rect 49882 7022 49888 7056
rect 49922 7022 49984 7056
rect 49656 6950 49696 6984
rect 49730 6950 49736 6984
rect 49656 6938 49736 6950
rect 49786 6984 49832 7004
rect 49786 6950 49792 6984
rect 49826 6950 49832 6984
rect 49786 6938 49832 6950
rect 49882 6984 49984 7022
rect 49882 6950 49888 6984
rect 49922 6950 49984 6984
rect 49882 6938 49984 6950
rect 49656 6738 49702 6938
rect 49732 6900 49790 6910
rect 49732 6866 49744 6900
rect 49778 6866 49790 6900
rect 49732 6848 49790 6866
rect 49934 6858 49984 6938
rect 50350 6916 50434 7186
rect 50092 6906 50150 6912
rect 50084 6900 50158 6906
rect 49844 6819 49902 6836
rect 49844 6785 49856 6819
rect 49890 6785 49902 6819
rect 49844 6770 49902 6785
rect 49934 6792 50004 6858
rect 50084 6848 50095 6900
rect 50147 6848 50158 6900
rect 50084 6842 50158 6848
rect 50226 6890 50502 6916
rect 51096 6910 51194 7186
rect 50226 6885 50327 6890
rect 50379 6885 50502 6890
rect 50226 6851 50255 6885
rect 50289 6851 50327 6885
rect 50381 6851 50439 6885
rect 50473 6851 50502 6885
rect 50092 6834 50150 6842
rect 50226 6838 50327 6851
rect 50379 6838 50502 6851
rect 50226 6820 50502 6838
rect 50572 6879 51194 6910
rect 50572 6845 50601 6879
rect 50635 6845 50693 6879
rect 50727 6845 50785 6879
rect 50819 6877 51194 6879
rect 50819 6845 50947 6877
rect 50572 6843 50947 6845
rect 50981 6843 51039 6877
rect 51073 6843 51131 6877
rect 51165 6843 51194 6877
rect 51456 7140 51776 7158
rect 51456 7106 51728 7140
rect 51762 7106 51776 7140
rect 51456 7096 51776 7106
rect 50572 6812 51194 6843
rect 51334 6868 51410 6874
rect 51334 6816 51350 6868
rect 51402 6816 51410 6868
rect 51334 6810 51410 6816
rect 49934 6738 49984 6792
rect 51456 6766 51516 7096
rect 51578 7056 51624 7068
rect 49656 6691 49752 6738
rect 49656 6657 49712 6691
rect 49746 6657 49752 6691
rect 49656 6619 49752 6657
rect 49656 6585 49712 6619
rect 49746 6585 49752 6619
rect 49802 6691 49848 6738
rect 49802 6657 49808 6691
rect 49842 6657 49848 6691
rect 49802 6619 49848 6657
rect 49802 6598 49808 6619
rect 49656 6538 49752 6585
rect 49792 6590 49808 6598
rect 49842 6598 49848 6619
rect 49898 6691 49984 6738
rect 50988 6746 51516 6766
rect 50988 6712 51000 6746
rect 51034 6732 51516 6746
rect 51034 6712 51046 6732
rect 50988 6698 51046 6712
rect 49898 6657 49904 6691
rect 49938 6657 49984 6691
rect 49898 6619 49984 6657
rect 49842 6590 49858 6598
rect 49792 6538 49800 6590
rect 49852 6538 49858 6590
rect 49898 6585 49904 6619
rect 49938 6585 49984 6619
rect 50060 6659 50126 6672
rect 50060 6625 50076 6659
rect 50110 6625 50126 6659
rect 50454 6652 50522 6654
rect 50060 6614 50126 6625
rect 50370 6648 50522 6652
rect 50370 6642 50463 6648
rect 50370 6608 50390 6642
rect 50424 6608 50463 6642
rect 50370 6602 50463 6608
rect 50454 6596 50463 6602
rect 50515 6596 50522 6648
rect 50454 6590 50522 6596
rect 50558 6636 50632 6660
rect 50558 6602 50586 6636
rect 50620 6602 50632 6636
rect 49898 6542 49984 6585
rect 50558 6582 50632 6602
rect 50756 6652 50828 6664
rect 50756 6600 50767 6652
rect 50819 6600 50828 6652
rect 51302 6659 51368 6668
rect 51302 6625 51318 6659
rect 51352 6625 51368 6659
rect 51302 6612 51368 6625
rect 50756 6596 50828 6600
rect 49898 6538 49944 6542
rect 49792 6530 49858 6538
rect 50026 6531 50072 6578
rect 49568 6491 49806 6500
rect 49568 6468 49760 6491
rect 49468 6442 49474 6459
rect 48226 6376 48298 6404
rect 49380 6378 49426 6425
rect 49456 6436 49474 6442
rect 49508 6442 49514 6459
rect 49566 6457 49760 6468
rect 49794 6457 49806 6491
rect 50026 6497 50032 6531
rect 50066 6497 50072 6531
rect 50026 6464 50072 6497
rect 49508 6436 49522 6442
rect 49456 6384 49462 6436
rect 49514 6384 49522 6436
rect 49456 6378 49522 6384
rect 49566 6440 49806 6457
rect 47914 6328 48004 6349
rect 48172 6331 48238 6340
rect 48172 6297 48188 6331
rect 48222 6297 48238 6331
rect 48172 6294 48238 6297
rect 47678 6266 48238 6294
rect 47582 6210 47650 6224
rect 47582 6176 47600 6210
rect 47634 6176 47650 6210
rect 47582 6166 47650 6176
rect 47622 5862 47650 6166
rect 47678 6084 47712 6266
rect 48010 6200 48082 6212
rect 48010 6148 48020 6200
rect 48072 6148 48082 6200
rect 48010 6136 48082 6148
rect 47934 6084 47998 6102
rect 47678 6050 47950 6084
rect 47984 6050 47998 6084
rect 47934 6040 47998 6050
rect 48270 6026 48298 6376
rect 48338 6342 48614 6372
rect 48338 6341 48370 6342
rect 48422 6341 48614 6342
rect 48338 6307 48367 6341
rect 48422 6307 48459 6341
rect 48493 6307 48551 6341
rect 48585 6307 48614 6341
rect 48338 6290 48370 6307
rect 48422 6290 48614 6307
rect 48338 6276 48614 6290
rect 48682 6348 49306 6366
rect 48682 6335 49224 6348
rect 48682 6301 48713 6335
rect 48747 6301 48805 6335
rect 48839 6301 48897 6335
rect 48931 6333 49224 6335
rect 49276 6333 49306 6348
rect 48931 6301 49059 6333
rect 48682 6299 49059 6301
rect 49093 6299 49151 6333
rect 49185 6299 49224 6333
rect 49277 6299 49306 6333
rect 48682 6296 49224 6299
rect 49276 6296 49306 6299
rect 48388 6084 48454 6090
rect 48388 6032 48394 6084
rect 48446 6032 48454 6084
rect 48388 6026 48454 6032
rect 48044 6012 48298 6026
rect 47800 6000 47846 6012
rect 47346 5834 47650 5862
rect 47766 5966 47806 6000
rect 47840 5966 47846 6000
rect 47766 5928 47846 5966
rect 47886 6006 47952 6012
rect 47886 5954 47892 6006
rect 47944 5954 47952 6006
rect 47886 5948 47952 5954
rect 47992 6000 48298 6012
rect 47992 5966 47998 6000
rect 48032 5998 48298 6000
rect 48032 5966 48094 5998
rect 47766 5894 47806 5928
rect 47840 5894 47846 5928
rect 47766 5882 47846 5894
rect 47896 5928 47942 5948
rect 47896 5894 47902 5928
rect 47936 5894 47942 5928
rect 47896 5882 47942 5894
rect 47992 5928 48094 5966
rect 47992 5894 47998 5928
rect 48032 5894 48094 5928
rect 47992 5882 48094 5894
rect 48214 5951 48448 5960
rect 48214 5899 48220 5951
rect 48272 5932 48396 5951
rect 48272 5899 48278 5932
rect 48214 5892 48278 5899
rect 48390 5899 48396 5932
rect 48448 5899 48454 5932
rect 48390 5892 48454 5899
rect 47346 5831 47622 5834
rect 47346 5797 47375 5831
rect 47409 5797 47467 5831
rect 47501 5797 47559 5831
rect 47593 5797 47622 5831
rect 47346 5766 47622 5797
rect 47452 5718 47516 5724
rect 47452 5666 47458 5718
rect 47510 5666 47516 5718
rect 47452 5660 47516 5666
rect 47766 5682 47812 5882
rect 47842 5844 47900 5854
rect 47842 5810 47854 5844
rect 47888 5810 47900 5844
rect 47842 5792 47900 5810
rect 47954 5763 48012 5780
rect 47954 5729 47966 5763
rect 48000 5729 48012 5763
rect 47954 5714 48012 5729
rect 48044 5682 48094 5882
rect 48160 5831 48436 5862
rect 48160 5797 48189 5831
rect 48223 5797 48281 5831
rect 48315 5797 48373 5831
rect 48407 5797 48436 5831
rect 48160 5766 48436 5797
rect 47766 5635 47862 5682
rect 47364 5602 47428 5608
rect 47364 5550 47370 5602
rect 47422 5550 47428 5602
rect 47364 5544 47428 5550
rect 47534 5592 47604 5610
rect 47534 5558 47555 5592
rect 47589 5558 47604 5592
rect 47534 5550 47604 5558
rect 47766 5601 47822 5635
rect 47856 5601 47862 5635
rect 47766 5563 47862 5601
rect 47534 5514 47562 5550
rect 47766 5529 47822 5563
rect 47856 5529 47862 5563
rect 47912 5635 47958 5682
rect 47912 5601 47918 5635
rect 47952 5601 47958 5635
rect 47912 5563 47958 5601
rect 47912 5542 47918 5563
rect 47766 5514 47862 5529
rect 47534 5482 47862 5514
rect 47902 5534 47918 5542
rect 47952 5542 47958 5563
rect 48008 5635 48094 5682
rect 48266 5716 48334 5726
rect 48266 5664 48274 5716
rect 48326 5664 48334 5716
rect 48266 5658 48334 5664
rect 48008 5601 48014 5635
rect 48048 5601 48094 5635
rect 48008 5563 48094 5601
rect 47952 5534 47968 5542
rect 47902 5482 47910 5534
rect 47962 5482 47968 5534
rect 48008 5529 48014 5563
rect 48048 5529 48094 5563
rect 48176 5604 48244 5610
rect 48176 5552 48182 5604
rect 48234 5552 48244 5604
rect 48176 5546 48244 5552
rect 48350 5590 48416 5602
rect 48350 5556 48367 5590
rect 48401 5556 48416 5590
rect 48350 5548 48416 5556
rect 48008 5510 48094 5529
rect 48388 5510 48416 5548
rect 48008 5482 48416 5510
rect 47902 5474 47968 5482
rect 48050 5478 48416 5482
rect 47854 5435 47916 5444
rect 47854 5401 47870 5435
rect 47904 5401 47916 5435
rect 47854 5384 47916 5401
rect 47858 5382 47916 5384
rect 47912 5327 48002 5348
rect 47912 5318 47939 5327
rect 46085 5293 47939 5318
rect 47973 5318 48002 5327
rect 48516 5318 48594 6276
rect 48682 6264 49306 6296
rect 49414 6331 49480 6342
rect 49414 6297 49430 6331
rect 49464 6297 49480 6331
rect 49414 6286 49480 6297
rect 49566 6294 49600 6440
rect 49748 6438 49806 6440
rect 50004 6459 50072 6464
rect 50004 6456 50032 6459
rect 50004 6404 50012 6456
rect 50066 6425 50072 6459
rect 50064 6404 50072 6425
rect 49802 6383 49892 6404
rect 50004 6398 50072 6404
rect 49802 6349 49829 6383
rect 49863 6349 49892 6383
rect 50026 6378 50072 6398
rect 50114 6531 50160 6578
rect 50114 6497 50120 6531
rect 50154 6497 50160 6531
rect 50114 6459 50160 6497
rect 50114 6425 50120 6459
rect 50154 6425 50160 6459
rect 50114 6404 50160 6425
rect 51268 6531 51314 6578
rect 51268 6497 51274 6531
rect 51308 6497 51314 6531
rect 51268 6459 51314 6497
rect 51268 6425 51274 6459
rect 51308 6425 51314 6459
rect 51356 6531 51402 6578
rect 51356 6497 51362 6531
rect 51396 6497 51402 6531
rect 51356 6459 51402 6497
rect 51456 6500 51516 6732
rect 51544 7022 51584 7056
rect 51618 7022 51624 7056
rect 51544 6984 51624 7022
rect 51664 7062 51730 7068
rect 51664 7010 51670 7062
rect 51722 7010 51730 7062
rect 51664 7004 51730 7010
rect 51770 7056 51872 7068
rect 51770 7022 51776 7056
rect 51810 7022 51872 7056
rect 51544 6950 51584 6984
rect 51618 6950 51624 6984
rect 51544 6938 51624 6950
rect 51674 6984 51720 7004
rect 51674 6950 51680 6984
rect 51714 6950 51720 6984
rect 51674 6938 51720 6950
rect 51770 6984 51872 7022
rect 51770 6950 51776 6984
rect 51810 6950 51872 6984
rect 51770 6938 51872 6950
rect 51544 6738 51590 6938
rect 51620 6900 51678 6910
rect 51620 6866 51632 6900
rect 51666 6866 51678 6900
rect 51620 6848 51678 6866
rect 51822 6858 51872 6938
rect 52238 6916 52322 7186
rect 51980 6906 52038 6912
rect 51972 6900 52046 6906
rect 51732 6819 51790 6836
rect 51732 6785 51744 6819
rect 51778 6785 51790 6819
rect 51732 6770 51790 6785
rect 51822 6792 51892 6858
rect 51972 6848 51983 6900
rect 52035 6848 52046 6900
rect 51972 6842 52046 6848
rect 52114 6890 52390 6916
rect 52984 6910 53082 7186
rect 52114 6885 52215 6890
rect 52267 6885 52390 6890
rect 52114 6851 52143 6885
rect 52177 6851 52215 6885
rect 52269 6851 52327 6885
rect 52361 6851 52390 6885
rect 51980 6834 52038 6842
rect 52114 6838 52215 6851
rect 52267 6838 52390 6851
rect 52114 6820 52390 6838
rect 52460 6879 53082 6910
rect 52460 6845 52489 6879
rect 52523 6845 52581 6879
rect 52615 6845 52673 6879
rect 52707 6877 53082 6879
rect 52707 6845 52835 6877
rect 52460 6843 52835 6845
rect 52869 6843 52927 6877
rect 52961 6843 53019 6877
rect 53053 6843 53082 6877
rect 53344 7140 53664 7158
rect 53344 7106 53616 7140
rect 53650 7106 53664 7140
rect 53344 7096 53664 7106
rect 52460 6812 53082 6843
rect 53222 6868 53298 6874
rect 53222 6816 53238 6868
rect 53290 6816 53298 6868
rect 53222 6810 53298 6816
rect 51822 6738 51872 6792
rect 53344 6766 53404 7096
rect 53466 7056 53512 7068
rect 51544 6691 51640 6738
rect 51544 6657 51600 6691
rect 51634 6657 51640 6691
rect 51544 6619 51640 6657
rect 51544 6585 51600 6619
rect 51634 6585 51640 6619
rect 51690 6691 51736 6738
rect 51690 6657 51696 6691
rect 51730 6657 51736 6691
rect 51690 6619 51736 6657
rect 51690 6598 51696 6619
rect 51544 6538 51640 6585
rect 51680 6590 51696 6598
rect 51730 6598 51736 6619
rect 51786 6691 51872 6738
rect 52876 6746 53404 6766
rect 52876 6712 52888 6746
rect 52922 6732 53404 6746
rect 52922 6712 52934 6732
rect 52876 6698 52934 6712
rect 51786 6657 51792 6691
rect 51826 6657 51872 6691
rect 51786 6619 51872 6657
rect 51730 6590 51746 6598
rect 51680 6538 51688 6590
rect 51740 6538 51746 6590
rect 51786 6585 51792 6619
rect 51826 6585 51872 6619
rect 51948 6659 52014 6672
rect 51948 6625 51964 6659
rect 51998 6625 52014 6659
rect 52342 6652 52410 6654
rect 51948 6614 52014 6625
rect 52258 6648 52410 6652
rect 52258 6642 52351 6648
rect 52258 6608 52278 6642
rect 52312 6608 52351 6642
rect 52258 6602 52351 6608
rect 52342 6596 52351 6602
rect 52403 6596 52410 6648
rect 52342 6590 52410 6596
rect 52446 6636 52520 6660
rect 52446 6602 52474 6636
rect 52508 6602 52520 6636
rect 51786 6542 51872 6585
rect 52446 6582 52520 6602
rect 52644 6652 52716 6664
rect 52644 6600 52655 6652
rect 52707 6600 52716 6652
rect 53190 6659 53256 6668
rect 53190 6625 53206 6659
rect 53240 6625 53256 6659
rect 53190 6612 53256 6625
rect 52644 6596 52716 6600
rect 51786 6538 51832 6542
rect 51680 6530 51746 6538
rect 51914 6531 51960 6578
rect 51456 6491 51694 6500
rect 51456 6468 51648 6491
rect 51356 6442 51362 6459
rect 50114 6376 50186 6404
rect 51268 6378 51314 6425
rect 51344 6436 51362 6442
rect 51396 6442 51402 6459
rect 51454 6457 51648 6468
rect 51682 6457 51694 6491
rect 51914 6497 51920 6531
rect 51954 6497 51960 6531
rect 51914 6464 51960 6497
rect 51396 6436 51410 6442
rect 51344 6384 51350 6436
rect 51402 6384 51410 6436
rect 51344 6378 51410 6384
rect 51454 6440 51694 6457
rect 49802 6328 49892 6349
rect 50060 6331 50126 6340
rect 50060 6297 50076 6331
rect 50110 6297 50126 6331
rect 50060 6294 50126 6297
rect 49566 6266 50126 6294
rect 49470 6210 49538 6224
rect 49470 6176 49488 6210
rect 49522 6176 49538 6210
rect 49470 6166 49538 6176
rect 49510 5862 49538 6166
rect 49566 6084 49600 6266
rect 49898 6200 49970 6212
rect 49898 6148 49908 6200
rect 49960 6148 49970 6200
rect 49898 6136 49970 6148
rect 49822 6084 49886 6102
rect 49566 6050 49838 6084
rect 49872 6050 49886 6084
rect 49822 6040 49886 6050
rect 50158 6026 50186 6376
rect 50226 6342 50502 6372
rect 50226 6341 50258 6342
rect 50310 6341 50502 6342
rect 50226 6307 50255 6341
rect 50310 6307 50347 6341
rect 50381 6307 50439 6341
rect 50473 6307 50502 6341
rect 50226 6290 50258 6307
rect 50310 6290 50502 6307
rect 50226 6276 50502 6290
rect 50570 6348 51194 6366
rect 50570 6335 51112 6348
rect 50570 6301 50601 6335
rect 50635 6301 50693 6335
rect 50727 6301 50785 6335
rect 50819 6333 51112 6335
rect 51164 6333 51194 6348
rect 50819 6301 50947 6333
rect 50570 6299 50947 6301
rect 50981 6299 51039 6333
rect 51073 6299 51112 6333
rect 51165 6299 51194 6333
rect 50570 6296 51112 6299
rect 51164 6296 51194 6299
rect 50276 6084 50342 6090
rect 50276 6032 50282 6084
rect 50334 6032 50342 6084
rect 50276 6026 50342 6032
rect 49932 6012 50186 6026
rect 49688 6000 49734 6012
rect 49234 5834 49538 5862
rect 49654 5966 49694 6000
rect 49728 5966 49734 6000
rect 49654 5928 49734 5966
rect 49774 6006 49840 6012
rect 49774 5954 49780 6006
rect 49832 5954 49840 6006
rect 49774 5948 49840 5954
rect 49880 6000 50186 6012
rect 49880 5966 49886 6000
rect 49920 5998 50186 6000
rect 49920 5966 49982 5998
rect 49654 5894 49694 5928
rect 49728 5894 49734 5928
rect 49654 5882 49734 5894
rect 49784 5928 49830 5948
rect 49784 5894 49790 5928
rect 49824 5894 49830 5928
rect 49784 5882 49830 5894
rect 49880 5928 49982 5966
rect 49880 5894 49886 5928
rect 49920 5894 49982 5928
rect 49880 5882 49982 5894
rect 50102 5951 50336 5960
rect 50102 5899 50108 5951
rect 50160 5932 50284 5951
rect 50160 5899 50166 5932
rect 50102 5892 50166 5899
rect 50278 5899 50284 5932
rect 50336 5899 50342 5932
rect 50278 5892 50342 5899
rect 49234 5831 49510 5834
rect 49234 5797 49263 5831
rect 49297 5797 49355 5831
rect 49389 5797 49447 5831
rect 49481 5797 49510 5831
rect 49234 5766 49510 5797
rect 49340 5718 49404 5724
rect 49340 5666 49346 5718
rect 49398 5666 49404 5718
rect 49340 5660 49404 5666
rect 49654 5682 49700 5882
rect 49730 5844 49788 5854
rect 49730 5810 49742 5844
rect 49776 5810 49788 5844
rect 49730 5792 49788 5810
rect 49842 5763 49900 5780
rect 49842 5729 49854 5763
rect 49888 5729 49900 5763
rect 49842 5714 49900 5729
rect 49932 5682 49982 5882
rect 50048 5831 50324 5862
rect 50048 5797 50077 5831
rect 50111 5797 50169 5831
rect 50203 5797 50261 5831
rect 50295 5797 50324 5831
rect 50048 5766 50324 5797
rect 49654 5635 49750 5682
rect 49252 5602 49316 5608
rect 49252 5550 49258 5602
rect 49310 5550 49316 5602
rect 49252 5544 49316 5550
rect 49422 5592 49492 5610
rect 49422 5558 49443 5592
rect 49477 5558 49492 5592
rect 49422 5550 49492 5558
rect 49654 5601 49710 5635
rect 49744 5601 49750 5635
rect 49654 5563 49750 5601
rect 49422 5514 49450 5550
rect 49654 5529 49710 5563
rect 49744 5529 49750 5563
rect 49800 5635 49846 5682
rect 49800 5601 49806 5635
rect 49840 5601 49846 5635
rect 49800 5563 49846 5601
rect 49800 5542 49806 5563
rect 49654 5514 49750 5529
rect 49422 5482 49750 5514
rect 49790 5534 49806 5542
rect 49840 5542 49846 5563
rect 49896 5635 49982 5682
rect 50154 5716 50222 5726
rect 50154 5664 50162 5716
rect 50214 5664 50222 5716
rect 50154 5658 50222 5664
rect 49896 5601 49902 5635
rect 49936 5601 49982 5635
rect 49896 5563 49982 5601
rect 49840 5534 49856 5542
rect 49790 5482 49798 5534
rect 49850 5482 49856 5534
rect 49896 5529 49902 5563
rect 49936 5529 49982 5563
rect 50064 5604 50132 5610
rect 50064 5552 50070 5604
rect 50122 5552 50132 5604
rect 50064 5546 50132 5552
rect 50238 5590 50304 5602
rect 50238 5556 50255 5590
rect 50289 5556 50304 5590
rect 50238 5548 50304 5556
rect 49896 5510 49982 5529
rect 50276 5510 50304 5548
rect 49896 5482 50304 5510
rect 49790 5474 49856 5482
rect 49938 5478 50304 5482
rect 49742 5435 49804 5444
rect 49742 5401 49758 5435
rect 49792 5401 49804 5435
rect 49742 5384 49804 5401
rect 49746 5382 49804 5384
rect 49800 5327 49890 5348
rect 49800 5318 49827 5327
rect 47973 5293 49827 5318
rect 49861 5318 49890 5327
rect 50404 5318 50482 6276
rect 50570 6264 51194 6296
rect 51302 6331 51368 6342
rect 51302 6297 51318 6331
rect 51352 6297 51368 6331
rect 51302 6286 51368 6297
rect 51454 6294 51488 6440
rect 51636 6438 51694 6440
rect 51892 6459 51960 6464
rect 51892 6456 51920 6459
rect 51892 6404 51900 6456
rect 51954 6425 51960 6459
rect 51952 6404 51960 6425
rect 51690 6383 51780 6404
rect 51892 6398 51960 6404
rect 51690 6349 51717 6383
rect 51751 6349 51780 6383
rect 51914 6378 51960 6398
rect 52002 6531 52048 6578
rect 52002 6497 52008 6531
rect 52042 6497 52048 6531
rect 52002 6459 52048 6497
rect 52002 6425 52008 6459
rect 52042 6425 52048 6459
rect 52002 6404 52048 6425
rect 53156 6531 53202 6578
rect 53156 6497 53162 6531
rect 53196 6497 53202 6531
rect 53156 6459 53202 6497
rect 53156 6425 53162 6459
rect 53196 6425 53202 6459
rect 53244 6531 53290 6578
rect 53244 6497 53250 6531
rect 53284 6497 53290 6531
rect 53244 6459 53290 6497
rect 53344 6500 53404 6732
rect 53432 7022 53472 7056
rect 53506 7022 53512 7056
rect 53432 6984 53512 7022
rect 53552 7062 53618 7068
rect 53552 7010 53558 7062
rect 53610 7010 53618 7062
rect 53552 7004 53618 7010
rect 53658 7056 53760 7068
rect 53658 7022 53664 7056
rect 53698 7022 53760 7056
rect 53432 6950 53472 6984
rect 53506 6950 53512 6984
rect 53432 6938 53512 6950
rect 53562 6984 53608 7004
rect 53562 6950 53568 6984
rect 53602 6950 53608 6984
rect 53562 6938 53608 6950
rect 53658 6984 53760 7022
rect 53658 6950 53664 6984
rect 53698 6950 53760 6984
rect 53658 6938 53760 6950
rect 53432 6738 53478 6938
rect 53508 6900 53566 6910
rect 53508 6866 53520 6900
rect 53554 6866 53566 6900
rect 53508 6848 53566 6866
rect 53710 6858 53760 6938
rect 54126 6916 54210 7186
rect 53868 6906 53926 6912
rect 53860 6900 53934 6906
rect 53620 6819 53678 6836
rect 53620 6785 53632 6819
rect 53666 6785 53678 6819
rect 53620 6770 53678 6785
rect 53710 6792 53780 6858
rect 53860 6848 53871 6900
rect 53923 6848 53934 6900
rect 53860 6842 53934 6848
rect 54002 6890 54278 6916
rect 54872 6910 54970 7186
rect 54002 6885 54103 6890
rect 54155 6885 54278 6890
rect 54002 6851 54031 6885
rect 54065 6851 54103 6885
rect 54157 6851 54215 6885
rect 54249 6851 54278 6885
rect 53868 6834 53926 6842
rect 54002 6838 54103 6851
rect 54155 6838 54278 6851
rect 54002 6820 54278 6838
rect 54348 6879 54970 6910
rect 54348 6845 54377 6879
rect 54411 6845 54469 6879
rect 54503 6845 54561 6879
rect 54595 6877 54970 6879
rect 54595 6845 54723 6877
rect 54348 6843 54723 6845
rect 54757 6843 54815 6877
rect 54849 6843 54907 6877
rect 54941 6843 54970 6877
rect 55232 7140 55552 7158
rect 55232 7106 55504 7140
rect 55538 7106 55552 7140
rect 55232 7096 55552 7106
rect 54348 6812 54970 6843
rect 55110 6868 55186 6874
rect 55110 6816 55126 6868
rect 55178 6816 55186 6868
rect 55110 6810 55186 6816
rect 53710 6738 53760 6792
rect 55232 6766 55292 7096
rect 55354 7056 55400 7068
rect 53432 6691 53528 6738
rect 53432 6657 53488 6691
rect 53522 6657 53528 6691
rect 53432 6619 53528 6657
rect 53432 6585 53488 6619
rect 53522 6585 53528 6619
rect 53578 6691 53624 6738
rect 53578 6657 53584 6691
rect 53618 6657 53624 6691
rect 53578 6619 53624 6657
rect 53578 6598 53584 6619
rect 53432 6538 53528 6585
rect 53568 6590 53584 6598
rect 53618 6598 53624 6619
rect 53674 6691 53760 6738
rect 54764 6746 55292 6766
rect 54764 6712 54776 6746
rect 54810 6732 55292 6746
rect 54810 6712 54822 6732
rect 54764 6698 54822 6712
rect 53674 6657 53680 6691
rect 53714 6657 53760 6691
rect 53674 6619 53760 6657
rect 53618 6590 53634 6598
rect 53568 6538 53576 6590
rect 53628 6538 53634 6590
rect 53674 6585 53680 6619
rect 53714 6585 53760 6619
rect 53836 6659 53902 6672
rect 53836 6625 53852 6659
rect 53886 6625 53902 6659
rect 54230 6652 54298 6654
rect 53836 6614 53902 6625
rect 54146 6648 54298 6652
rect 54146 6642 54239 6648
rect 54146 6608 54166 6642
rect 54200 6608 54239 6642
rect 54146 6602 54239 6608
rect 54230 6596 54239 6602
rect 54291 6596 54298 6648
rect 54230 6590 54298 6596
rect 54334 6636 54408 6660
rect 54334 6602 54362 6636
rect 54396 6602 54408 6636
rect 53674 6542 53760 6585
rect 54334 6582 54408 6602
rect 54532 6652 54604 6664
rect 54532 6600 54543 6652
rect 54595 6600 54604 6652
rect 55078 6659 55144 6668
rect 55078 6625 55094 6659
rect 55128 6625 55144 6659
rect 55078 6612 55144 6625
rect 54532 6596 54604 6600
rect 53674 6538 53720 6542
rect 53568 6530 53634 6538
rect 53802 6531 53848 6578
rect 53344 6491 53582 6500
rect 53344 6468 53536 6491
rect 53244 6442 53250 6459
rect 52002 6376 52074 6404
rect 53156 6378 53202 6425
rect 53232 6436 53250 6442
rect 53284 6442 53290 6459
rect 53342 6457 53536 6468
rect 53570 6457 53582 6491
rect 53802 6497 53808 6531
rect 53842 6497 53848 6531
rect 53802 6464 53848 6497
rect 53284 6436 53298 6442
rect 53232 6384 53238 6436
rect 53290 6384 53298 6436
rect 53232 6378 53298 6384
rect 53342 6440 53582 6457
rect 51690 6328 51780 6349
rect 51948 6331 52014 6340
rect 51948 6297 51964 6331
rect 51998 6297 52014 6331
rect 51948 6294 52014 6297
rect 51454 6266 52014 6294
rect 51358 6210 51426 6224
rect 51358 6176 51376 6210
rect 51410 6176 51426 6210
rect 51358 6166 51426 6176
rect 51398 5862 51426 6166
rect 51454 6084 51488 6266
rect 51786 6200 51858 6212
rect 51786 6148 51796 6200
rect 51848 6148 51858 6200
rect 51786 6136 51858 6148
rect 51710 6084 51774 6102
rect 51454 6050 51726 6084
rect 51760 6050 51774 6084
rect 51710 6040 51774 6050
rect 52046 6026 52074 6376
rect 52114 6342 52390 6372
rect 52114 6341 52146 6342
rect 52198 6341 52390 6342
rect 52114 6307 52143 6341
rect 52198 6307 52235 6341
rect 52269 6307 52327 6341
rect 52361 6307 52390 6341
rect 52114 6290 52146 6307
rect 52198 6290 52390 6307
rect 52114 6276 52390 6290
rect 52458 6348 53082 6366
rect 52458 6335 53000 6348
rect 52458 6301 52489 6335
rect 52523 6301 52581 6335
rect 52615 6301 52673 6335
rect 52707 6333 53000 6335
rect 53052 6333 53082 6348
rect 52707 6301 52835 6333
rect 52458 6299 52835 6301
rect 52869 6299 52927 6333
rect 52961 6299 53000 6333
rect 53053 6299 53082 6333
rect 52458 6296 53000 6299
rect 53052 6296 53082 6299
rect 52164 6084 52230 6090
rect 52164 6032 52170 6084
rect 52222 6032 52230 6084
rect 52164 6026 52230 6032
rect 51820 6012 52074 6026
rect 51576 6000 51622 6012
rect 51122 5834 51426 5862
rect 51542 5966 51582 6000
rect 51616 5966 51622 6000
rect 51542 5928 51622 5966
rect 51662 6006 51728 6012
rect 51662 5954 51668 6006
rect 51720 5954 51728 6006
rect 51662 5948 51728 5954
rect 51768 6000 52074 6012
rect 51768 5966 51774 6000
rect 51808 5998 52074 6000
rect 51808 5966 51870 5998
rect 51542 5894 51582 5928
rect 51616 5894 51622 5928
rect 51542 5882 51622 5894
rect 51672 5928 51718 5948
rect 51672 5894 51678 5928
rect 51712 5894 51718 5928
rect 51672 5882 51718 5894
rect 51768 5928 51870 5966
rect 51768 5894 51774 5928
rect 51808 5894 51870 5928
rect 51768 5882 51870 5894
rect 51990 5951 52224 5960
rect 51990 5899 51996 5951
rect 52048 5932 52172 5951
rect 52048 5899 52054 5932
rect 51990 5892 52054 5899
rect 52166 5899 52172 5932
rect 52224 5899 52230 5932
rect 52166 5892 52230 5899
rect 51122 5831 51398 5834
rect 51122 5797 51151 5831
rect 51185 5797 51243 5831
rect 51277 5797 51335 5831
rect 51369 5797 51398 5831
rect 51122 5766 51398 5797
rect 51228 5718 51292 5724
rect 51228 5666 51234 5718
rect 51286 5666 51292 5718
rect 51228 5660 51292 5666
rect 51542 5682 51588 5882
rect 51618 5844 51676 5854
rect 51618 5810 51630 5844
rect 51664 5810 51676 5844
rect 51618 5792 51676 5810
rect 51730 5763 51788 5780
rect 51730 5729 51742 5763
rect 51776 5729 51788 5763
rect 51730 5714 51788 5729
rect 51820 5682 51870 5882
rect 51936 5831 52212 5862
rect 51936 5797 51965 5831
rect 51999 5797 52057 5831
rect 52091 5797 52149 5831
rect 52183 5797 52212 5831
rect 51936 5766 52212 5797
rect 51542 5635 51638 5682
rect 51140 5602 51204 5608
rect 51140 5550 51146 5602
rect 51198 5550 51204 5602
rect 51140 5544 51204 5550
rect 51310 5592 51380 5610
rect 51310 5558 51331 5592
rect 51365 5558 51380 5592
rect 51310 5550 51380 5558
rect 51542 5601 51598 5635
rect 51632 5601 51638 5635
rect 51542 5563 51638 5601
rect 51310 5514 51338 5550
rect 51542 5529 51598 5563
rect 51632 5529 51638 5563
rect 51688 5635 51734 5682
rect 51688 5601 51694 5635
rect 51728 5601 51734 5635
rect 51688 5563 51734 5601
rect 51688 5542 51694 5563
rect 51542 5514 51638 5529
rect 51310 5482 51638 5514
rect 51678 5534 51694 5542
rect 51728 5542 51734 5563
rect 51784 5635 51870 5682
rect 52042 5716 52110 5726
rect 52042 5664 52050 5716
rect 52102 5664 52110 5716
rect 52042 5658 52110 5664
rect 51784 5601 51790 5635
rect 51824 5601 51870 5635
rect 51784 5563 51870 5601
rect 51728 5534 51744 5542
rect 51678 5482 51686 5534
rect 51738 5482 51744 5534
rect 51784 5529 51790 5563
rect 51824 5529 51870 5563
rect 51952 5604 52020 5610
rect 51952 5552 51958 5604
rect 52010 5552 52020 5604
rect 51952 5546 52020 5552
rect 52126 5590 52192 5602
rect 52126 5556 52143 5590
rect 52177 5556 52192 5590
rect 52126 5548 52192 5556
rect 51784 5510 51870 5529
rect 52164 5510 52192 5548
rect 51784 5482 52192 5510
rect 51678 5474 51744 5482
rect 51826 5478 52192 5482
rect 51630 5435 51692 5444
rect 51630 5401 51646 5435
rect 51680 5401 51692 5435
rect 51630 5384 51692 5401
rect 51634 5382 51692 5384
rect 51688 5327 51778 5348
rect 51688 5318 51715 5327
rect 49861 5293 51715 5318
rect 51749 5318 51778 5327
rect 52292 5318 52370 6276
rect 52458 6264 53082 6296
rect 53190 6331 53256 6342
rect 53190 6297 53206 6331
rect 53240 6297 53256 6331
rect 53190 6286 53256 6297
rect 53342 6294 53376 6440
rect 53524 6438 53582 6440
rect 53780 6459 53848 6464
rect 53780 6456 53808 6459
rect 53780 6404 53788 6456
rect 53842 6425 53848 6459
rect 53840 6404 53848 6425
rect 53578 6383 53668 6404
rect 53780 6398 53848 6404
rect 53578 6349 53605 6383
rect 53639 6349 53668 6383
rect 53802 6378 53848 6398
rect 53890 6531 53936 6578
rect 53890 6497 53896 6531
rect 53930 6497 53936 6531
rect 53890 6459 53936 6497
rect 53890 6425 53896 6459
rect 53930 6425 53936 6459
rect 53890 6404 53936 6425
rect 55044 6531 55090 6578
rect 55044 6497 55050 6531
rect 55084 6497 55090 6531
rect 55044 6459 55090 6497
rect 55044 6425 55050 6459
rect 55084 6425 55090 6459
rect 55132 6531 55178 6578
rect 55132 6497 55138 6531
rect 55172 6497 55178 6531
rect 55132 6459 55178 6497
rect 55232 6500 55292 6732
rect 55320 7022 55360 7056
rect 55394 7022 55400 7056
rect 55320 6984 55400 7022
rect 55440 7062 55506 7068
rect 55440 7010 55446 7062
rect 55498 7010 55506 7062
rect 55440 7004 55506 7010
rect 55546 7056 55648 7068
rect 55546 7022 55552 7056
rect 55586 7022 55648 7056
rect 55320 6950 55360 6984
rect 55394 6950 55400 6984
rect 55320 6938 55400 6950
rect 55450 6984 55496 7004
rect 55450 6950 55456 6984
rect 55490 6950 55496 6984
rect 55450 6938 55496 6950
rect 55546 6984 55648 7022
rect 55546 6950 55552 6984
rect 55586 6950 55648 6984
rect 55546 6938 55648 6950
rect 55320 6738 55366 6938
rect 55396 6900 55454 6910
rect 55396 6866 55408 6900
rect 55442 6866 55454 6900
rect 55396 6848 55454 6866
rect 55598 6858 55648 6938
rect 56014 6916 56098 7186
rect 55756 6906 55814 6912
rect 55748 6900 55822 6906
rect 55508 6819 55566 6836
rect 55508 6785 55520 6819
rect 55554 6785 55566 6819
rect 55508 6770 55566 6785
rect 55598 6792 55668 6858
rect 55748 6848 55759 6900
rect 55811 6848 55822 6900
rect 55748 6842 55822 6848
rect 55890 6890 56166 6916
rect 56760 6910 56858 7186
rect 55890 6885 55991 6890
rect 56043 6885 56166 6890
rect 55890 6851 55919 6885
rect 55953 6851 55991 6885
rect 56045 6851 56103 6885
rect 56137 6851 56166 6885
rect 55756 6834 55814 6842
rect 55890 6838 55991 6851
rect 56043 6838 56166 6851
rect 55890 6820 56166 6838
rect 56236 6879 56858 6910
rect 56236 6845 56265 6879
rect 56299 6845 56357 6879
rect 56391 6845 56449 6879
rect 56483 6877 56858 6879
rect 56483 6845 56611 6877
rect 56236 6843 56611 6845
rect 56645 6843 56703 6877
rect 56737 6843 56795 6877
rect 56829 6843 56858 6877
rect 57120 7140 57440 7158
rect 57120 7106 57392 7140
rect 57426 7106 57440 7140
rect 57120 7096 57440 7106
rect 56236 6812 56858 6843
rect 56998 6868 57074 6874
rect 56998 6816 57014 6868
rect 57066 6816 57074 6868
rect 56998 6810 57074 6816
rect 55598 6738 55648 6792
rect 57120 6766 57180 7096
rect 57242 7056 57288 7068
rect 55320 6691 55416 6738
rect 55320 6657 55376 6691
rect 55410 6657 55416 6691
rect 55320 6619 55416 6657
rect 55320 6585 55376 6619
rect 55410 6585 55416 6619
rect 55466 6691 55512 6738
rect 55466 6657 55472 6691
rect 55506 6657 55512 6691
rect 55466 6619 55512 6657
rect 55466 6598 55472 6619
rect 55320 6538 55416 6585
rect 55456 6590 55472 6598
rect 55506 6598 55512 6619
rect 55562 6691 55648 6738
rect 56652 6746 57180 6766
rect 56652 6712 56664 6746
rect 56698 6732 57180 6746
rect 56698 6712 56710 6732
rect 56652 6698 56710 6712
rect 55562 6657 55568 6691
rect 55602 6657 55648 6691
rect 55562 6619 55648 6657
rect 55506 6590 55522 6598
rect 55456 6538 55464 6590
rect 55516 6538 55522 6590
rect 55562 6585 55568 6619
rect 55602 6585 55648 6619
rect 55724 6659 55790 6672
rect 55724 6625 55740 6659
rect 55774 6625 55790 6659
rect 56118 6652 56186 6654
rect 55724 6614 55790 6625
rect 56034 6648 56186 6652
rect 56034 6642 56127 6648
rect 56034 6608 56054 6642
rect 56088 6608 56127 6642
rect 56034 6602 56127 6608
rect 56118 6596 56127 6602
rect 56179 6596 56186 6648
rect 56118 6590 56186 6596
rect 56222 6636 56296 6660
rect 56222 6602 56250 6636
rect 56284 6602 56296 6636
rect 55562 6542 55648 6585
rect 56222 6582 56296 6602
rect 56420 6652 56492 6664
rect 56420 6600 56431 6652
rect 56483 6600 56492 6652
rect 56966 6659 57032 6668
rect 56966 6625 56982 6659
rect 57016 6625 57032 6659
rect 56966 6612 57032 6625
rect 56420 6596 56492 6600
rect 55562 6538 55608 6542
rect 55456 6530 55522 6538
rect 55690 6531 55736 6578
rect 55232 6491 55470 6500
rect 55232 6468 55424 6491
rect 55132 6442 55138 6459
rect 53890 6376 53962 6404
rect 55044 6378 55090 6425
rect 55120 6436 55138 6442
rect 55172 6442 55178 6459
rect 55230 6457 55424 6468
rect 55458 6457 55470 6491
rect 55690 6497 55696 6531
rect 55730 6497 55736 6531
rect 55690 6464 55736 6497
rect 55172 6436 55186 6442
rect 55120 6384 55126 6436
rect 55178 6384 55186 6436
rect 55120 6378 55186 6384
rect 55230 6440 55470 6457
rect 53578 6328 53668 6349
rect 53836 6331 53902 6340
rect 53836 6297 53852 6331
rect 53886 6297 53902 6331
rect 53836 6294 53902 6297
rect 53342 6266 53902 6294
rect 53246 6210 53314 6224
rect 53246 6176 53264 6210
rect 53298 6176 53314 6210
rect 53246 6166 53314 6176
rect 53286 5862 53314 6166
rect 53342 6084 53376 6266
rect 53674 6200 53746 6212
rect 53674 6148 53684 6200
rect 53736 6148 53746 6200
rect 53674 6136 53746 6148
rect 53598 6084 53662 6102
rect 53342 6050 53614 6084
rect 53648 6050 53662 6084
rect 53598 6040 53662 6050
rect 53934 6026 53962 6376
rect 54002 6342 54278 6372
rect 54002 6341 54034 6342
rect 54086 6341 54278 6342
rect 54002 6307 54031 6341
rect 54086 6307 54123 6341
rect 54157 6307 54215 6341
rect 54249 6307 54278 6341
rect 54002 6290 54034 6307
rect 54086 6290 54278 6307
rect 54002 6276 54278 6290
rect 54346 6348 54970 6366
rect 54346 6335 54888 6348
rect 54346 6301 54377 6335
rect 54411 6301 54469 6335
rect 54503 6301 54561 6335
rect 54595 6333 54888 6335
rect 54940 6333 54970 6348
rect 54595 6301 54723 6333
rect 54346 6299 54723 6301
rect 54757 6299 54815 6333
rect 54849 6299 54888 6333
rect 54941 6299 54970 6333
rect 54346 6296 54888 6299
rect 54940 6296 54970 6299
rect 54052 6084 54118 6090
rect 54052 6032 54058 6084
rect 54110 6032 54118 6084
rect 54052 6026 54118 6032
rect 53708 6012 53962 6026
rect 53464 6000 53510 6012
rect 53010 5834 53314 5862
rect 53430 5966 53470 6000
rect 53504 5966 53510 6000
rect 53430 5928 53510 5966
rect 53550 6006 53616 6012
rect 53550 5954 53556 6006
rect 53608 5954 53616 6006
rect 53550 5948 53616 5954
rect 53656 6000 53962 6012
rect 53656 5966 53662 6000
rect 53696 5998 53962 6000
rect 53696 5966 53758 5998
rect 53430 5894 53470 5928
rect 53504 5894 53510 5928
rect 53430 5882 53510 5894
rect 53560 5928 53606 5948
rect 53560 5894 53566 5928
rect 53600 5894 53606 5928
rect 53560 5882 53606 5894
rect 53656 5928 53758 5966
rect 53656 5894 53662 5928
rect 53696 5894 53758 5928
rect 53656 5882 53758 5894
rect 53878 5951 54112 5960
rect 53878 5899 53884 5951
rect 53936 5932 54060 5951
rect 53936 5899 53942 5932
rect 53878 5892 53942 5899
rect 54054 5899 54060 5932
rect 54112 5899 54118 5932
rect 54054 5892 54118 5899
rect 53010 5831 53286 5834
rect 53010 5797 53039 5831
rect 53073 5797 53131 5831
rect 53165 5797 53223 5831
rect 53257 5797 53286 5831
rect 53010 5766 53286 5797
rect 53116 5718 53180 5724
rect 53116 5666 53122 5718
rect 53174 5666 53180 5718
rect 53116 5660 53180 5666
rect 53430 5682 53476 5882
rect 53506 5844 53564 5854
rect 53506 5810 53518 5844
rect 53552 5810 53564 5844
rect 53506 5792 53564 5810
rect 53618 5763 53676 5780
rect 53618 5729 53630 5763
rect 53664 5729 53676 5763
rect 53618 5714 53676 5729
rect 53708 5682 53758 5882
rect 53824 5831 54100 5862
rect 53824 5797 53853 5831
rect 53887 5797 53945 5831
rect 53979 5797 54037 5831
rect 54071 5797 54100 5831
rect 53824 5766 54100 5797
rect 53430 5635 53526 5682
rect 53028 5602 53092 5608
rect 53028 5550 53034 5602
rect 53086 5550 53092 5602
rect 53028 5544 53092 5550
rect 53198 5592 53268 5610
rect 53198 5558 53219 5592
rect 53253 5558 53268 5592
rect 53198 5550 53268 5558
rect 53430 5601 53486 5635
rect 53520 5601 53526 5635
rect 53430 5563 53526 5601
rect 53198 5514 53226 5550
rect 53430 5529 53486 5563
rect 53520 5529 53526 5563
rect 53576 5635 53622 5682
rect 53576 5601 53582 5635
rect 53616 5601 53622 5635
rect 53576 5563 53622 5601
rect 53576 5542 53582 5563
rect 53430 5514 53526 5529
rect 53198 5482 53526 5514
rect 53566 5534 53582 5542
rect 53616 5542 53622 5563
rect 53672 5635 53758 5682
rect 53930 5716 53998 5726
rect 53930 5664 53938 5716
rect 53990 5664 53998 5716
rect 53930 5658 53998 5664
rect 53672 5601 53678 5635
rect 53712 5601 53758 5635
rect 53672 5563 53758 5601
rect 53616 5534 53632 5542
rect 53566 5482 53574 5534
rect 53626 5482 53632 5534
rect 53672 5529 53678 5563
rect 53712 5529 53758 5563
rect 53840 5604 53908 5610
rect 53840 5552 53846 5604
rect 53898 5552 53908 5604
rect 53840 5546 53908 5552
rect 54014 5590 54080 5602
rect 54014 5556 54031 5590
rect 54065 5556 54080 5590
rect 54014 5548 54080 5556
rect 53672 5510 53758 5529
rect 54052 5510 54080 5548
rect 53672 5482 54080 5510
rect 53566 5474 53632 5482
rect 53714 5478 54080 5482
rect 53518 5435 53580 5444
rect 53518 5401 53534 5435
rect 53568 5401 53580 5435
rect 53518 5384 53580 5401
rect 53522 5382 53580 5384
rect 53576 5327 53666 5348
rect 53576 5318 53603 5327
rect 51749 5293 53603 5318
rect 53637 5318 53666 5327
rect 54180 5318 54258 6276
rect 54346 6264 54970 6296
rect 55078 6331 55144 6342
rect 55078 6297 55094 6331
rect 55128 6297 55144 6331
rect 55078 6286 55144 6297
rect 55230 6294 55264 6440
rect 55412 6438 55470 6440
rect 55668 6459 55736 6464
rect 55668 6456 55696 6459
rect 55668 6404 55676 6456
rect 55730 6425 55736 6459
rect 55728 6404 55736 6425
rect 55466 6383 55556 6404
rect 55668 6398 55736 6404
rect 55466 6349 55493 6383
rect 55527 6349 55556 6383
rect 55690 6378 55736 6398
rect 55778 6531 55824 6578
rect 55778 6497 55784 6531
rect 55818 6497 55824 6531
rect 55778 6459 55824 6497
rect 55778 6425 55784 6459
rect 55818 6425 55824 6459
rect 55778 6404 55824 6425
rect 56932 6531 56978 6578
rect 56932 6497 56938 6531
rect 56972 6497 56978 6531
rect 56932 6459 56978 6497
rect 56932 6425 56938 6459
rect 56972 6425 56978 6459
rect 57020 6531 57066 6578
rect 57020 6497 57026 6531
rect 57060 6497 57066 6531
rect 57020 6459 57066 6497
rect 57120 6500 57180 6732
rect 57208 7022 57248 7056
rect 57282 7022 57288 7056
rect 57208 6984 57288 7022
rect 57328 7062 57394 7068
rect 57328 7010 57334 7062
rect 57386 7010 57394 7062
rect 57328 7004 57394 7010
rect 57434 7056 57536 7068
rect 57434 7022 57440 7056
rect 57474 7022 57536 7056
rect 57208 6950 57248 6984
rect 57282 6950 57288 6984
rect 57208 6938 57288 6950
rect 57338 6984 57384 7004
rect 57338 6950 57344 6984
rect 57378 6950 57384 6984
rect 57338 6938 57384 6950
rect 57434 6984 57536 7022
rect 57434 6950 57440 6984
rect 57474 6950 57536 6984
rect 57434 6938 57536 6950
rect 57208 6738 57254 6938
rect 57284 6900 57342 6910
rect 57284 6866 57296 6900
rect 57330 6866 57342 6900
rect 57284 6848 57342 6866
rect 57486 6858 57536 6938
rect 57902 6916 57986 7186
rect 57644 6906 57702 6912
rect 57636 6900 57710 6906
rect 57396 6819 57454 6836
rect 57396 6785 57408 6819
rect 57442 6785 57454 6819
rect 57396 6770 57454 6785
rect 57486 6792 57556 6858
rect 57636 6848 57647 6900
rect 57699 6848 57710 6900
rect 57636 6842 57710 6848
rect 57778 6890 58054 6916
rect 58648 6910 58746 7186
rect 57778 6885 57879 6890
rect 57931 6885 58054 6890
rect 57778 6851 57807 6885
rect 57841 6851 57879 6885
rect 57933 6851 57991 6885
rect 58025 6851 58054 6885
rect 57644 6834 57702 6842
rect 57778 6838 57879 6851
rect 57931 6838 58054 6851
rect 57778 6820 58054 6838
rect 58124 6879 58746 6910
rect 58124 6845 58153 6879
rect 58187 6845 58245 6879
rect 58279 6845 58337 6879
rect 58371 6877 58746 6879
rect 58371 6845 58499 6877
rect 58124 6843 58499 6845
rect 58533 6843 58591 6877
rect 58625 6843 58683 6877
rect 58717 6843 58746 6877
rect 59008 7140 59328 7158
rect 59008 7106 59280 7140
rect 59314 7106 59328 7140
rect 59008 7096 59328 7106
rect 58124 6812 58746 6843
rect 58886 6868 58962 6874
rect 58886 6816 58902 6868
rect 58954 6816 58962 6868
rect 58886 6810 58962 6816
rect 57486 6738 57536 6792
rect 59008 6766 59068 7096
rect 59130 7056 59176 7068
rect 57208 6691 57304 6738
rect 57208 6657 57264 6691
rect 57298 6657 57304 6691
rect 57208 6619 57304 6657
rect 57208 6585 57264 6619
rect 57298 6585 57304 6619
rect 57354 6691 57400 6738
rect 57354 6657 57360 6691
rect 57394 6657 57400 6691
rect 57354 6619 57400 6657
rect 57354 6598 57360 6619
rect 57208 6538 57304 6585
rect 57344 6590 57360 6598
rect 57394 6598 57400 6619
rect 57450 6691 57536 6738
rect 58540 6746 59068 6766
rect 58540 6712 58552 6746
rect 58586 6732 59068 6746
rect 58586 6712 58598 6732
rect 58540 6698 58598 6712
rect 57450 6657 57456 6691
rect 57490 6657 57536 6691
rect 57450 6619 57536 6657
rect 57394 6590 57410 6598
rect 57344 6538 57352 6590
rect 57404 6538 57410 6590
rect 57450 6585 57456 6619
rect 57490 6585 57536 6619
rect 57612 6659 57678 6672
rect 57612 6625 57628 6659
rect 57662 6625 57678 6659
rect 58006 6652 58074 6654
rect 57612 6614 57678 6625
rect 57922 6648 58074 6652
rect 57922 6642 58015 6648
rect 57922 6608 57942 6642
rect 57976 6608 58015 6642
rect 57922 6602 58015 6608
rect 58006 6596 58015 6602
rect 58067 6596 58074 6648
rect 58006 6590 58074 6596
rect 58110 6636 58184 6660
rect 58110 6602 58138 6636
rect 58172 6602 58184 6636
rect 57450 6542 57536 6585
rect 58110 6582 58184 6602
rect 58308 6652 58380 6664
rect 58308 6600 58319 6652
rect 58371 6600 58380 6652
rect 58854 6659 58920 6668
rect 58854 6625 58870 6659
rect 58904 6625 58920 6659
rect 58854 6612 58920 6625
rect 58308 6596 58380 6600
rect 57450 6538 57496 6542
rect 57344 6530 57410 6538
rect 57578 6531 57624 6578
rect 57120 6491 57358 6500
rect 57120 6468 57312 6491
rect 57020 6442 57026 6459
rect 55778 6376 55850 6404
rect 56932 6378 56978 6425
rect 57008 6436 57026 6442
rect 57060 6442 57066 6459
rect 57118 6457 57312 6468
rect 57346 6457 57358 6491
rect 57578 6497 57584 6531
rect 57618 6497 57624 6531
rect 57578 6464 57624 6497
rect 57060 6436 57074 6442
rect 57008 6384 57014 6436
rect 57066 6384 57074 6436
rect 57008 6378 57074 6384
rect 57118 6440 57358 6457
rect 55466 6328 55556 6349
rect 55724 6331 55790 6340
rect 55724 6297 55740 6331
rect 55774 6297 55790 6331
rect 55724 6294 55790 6297
rect 55230 6266 55790 6294
rect 55134 6210 55202 6224
rect 55134 6176 55152 6210
rect 55186 6176 55202 6210
rect 55134 6166 55202 6176
rect 55174 5862 55202 6166
rect 55230 6084 55264 6266
rect 55562 6200 55634 6212
rect 55562 6148 55572 6200
rect 55624 6148 55634 6200
rect 55562 6136 55634 6148
rect 55486 6084 55550 6102
rect 55230 6050 55502 6084
rect 55536 6050 55550 6084
rect 55486 6040 55550 6050
rect 55822 6026 55850 6376
rect 55890 6342 56166 6372
rect 55890 6341 55922 6342
rect 55974 6341 56166 6342
rect 55890 6307 55919 6341
rect 55974 6307 56011 6341
rect 56045 6307 56103 6341
rect 56137 6307 56166 6341
rect 55890 6290 55922 6307
rect 55974 6290 56166 6307
rect 55890 6276 56166 6290
rect 56234 6348 56858 6366
rect 56234 6335 56776 6348
rect 56234 6301 56265 6335
rect 56299 6301 56357 6335
rect 56391 6301 56449 6335
rect 56483 6333 56776 6335
rect 56828 6333 56858 6348
rect 56483 6301 56611 6333
rect 56234 6299 56611 6301
rect 56645 6299 56703 6333
rect 56737 6299 56776 6333
rect 56829 6299 56858 6333
rect 56234 6296 56776 6299
rect 56828 6296 56858 6299
rect 55940 6084 56006 6090
rect 55940 6032 55946 6084
rect 55998 6032 56006 6084
rect 55940 6026 56006 6032
rect 55596 6012 55850 6026
rect 55352 6000 55398 6012
rect 54898 5834 55202 5862
rect 55318 5966 55358 6000
rect 55392 5966 55398 6000
rect 55318 5928 55398 5966
rect 55438 6006 55504 6012
rect 55438 5954 55444 6006
rect 55496 5954 55504 6006
rect 55438 5948 55504 5954
rect 55544 6000 55850 6012
rect 55544 5966 55550 6000
rect 55584 5998 55850 6000
rect 55584 5966 55646 5998
rect 55318 5894 55358 5928
rect 55392 5894 55398 5928
rect 55318 5882 55398 5894
rect 55448 5928 55494 5948
rect 55448 5894 55454 5928
rect 55488 5894 55494 5928
rect 55448 5882 55494 5894
rect 55544 5928 55646 5966
rect 55544 5894 55550 5928
rect 55584 5894 55646 5928
rect 55544 5882 55646 5894
rect 55766 5951 56000 5960
rect 55766 5899 55772 5951
rect 55824 5932 55948 5951
rect 55824 5899 55830 5932
rect 55766 5892 55830 5899
rect 55942 5899 55948 5932
rect 56000 5899 56006 5932
rect 55942 5892 56006 5899
rect 54898 5831 55174 5834
rect 54898 5797 54927 5831
rect 54961 5797 55019 5831
rect 55053 5797 55111 5831
rect 55145 5797 55174 5831
rect 54898 5766 55174 5797
rect 55004 5718 55068 5724
rect 55004 5666 55010 5718
rect 55062 5666 55068 5718
rect 55004 5660 55068 5666
rect 55318 5682 55364 5882
rect 55394 5844 55452 5854
rect 55394 5810 55406 5844
rect 55440 5810 55452 5844
rect 55394 5792 55452 5810
rect 55506 5763 55564 5780
rect 55506 5729 55518 5763
rect 55552 5729 55564 5763
rect 55506 5714 55564 5729
rect 55596 5682 55646 5882
rect 55712 5831 55988 5862
rect 55712 5797 55741 5831
rect 55775 5797 55833 5831
rect 55867 5797 55925 5831
rect 55959 5797 55988 5831
rect 55712 5766 55988 5797
rect 55318 5635 55414 5682
rect 54916 5602 54980 5608
rect 54916 5550 54922 5602
rect 54974 5550 54980 5602
rect 54916 5544 54980 5550
rect 55086 5592 55156 5610
rect 55086 5558 55107 5592
rect 55141 5558 55156 5592
rect 55086 5550 55156 5558
rect 55318 5601 55374 5635
rect 55408 5601 55414 5635
rect 55318 5563 55414 5601
rect 55086 5514 55114 5550
rect 55318 5529 55374 5563
rect 55408 5529 55414 5563
rect 55464 5635 55510 5682
rect 55464 5601 55470 5635
rect 55504 5601 55510 5635
rect 55464 5563 55510 5601
rect 55464 5542 55470 5563
rect 55318 5514 55414 5529
rect 55086 5482 55414 5514
rect 55454 5534 55470 5542
rect 55504 5542 55510 5563
rect 55560 5635 55646 5682
rect 55818 5716 55886 5726
rect 55818 5664 55826 5716
rect 55878 5664 55886 5716
rect 55818 5658 55886 5664
rect 55560 5601 55566 5635
rect 55600 5601 55646 5635
rect 55560 5563 55646 5601
rect 55504 5534 55520 5542
rect 55454 5482 55462 5534
rect 55514 5482 55520 5534
rect 55560 5529 55566 5563
rect 55600 5529 55646 5563
rect 55728 5604 55796 5610
rect 55728 5552 55734 5604
rect 55786 5552 55796 5604
rect 55728 5546 55796 5552
rect 55902 5590 55968 5602
rect 55902 5556 55919 5590
rect 55953 5556 55968 5590
rect 55902 5548 55968 5556
rect 55560 5510 55646 5529
rect 55940 5510 55968 5548
rect 55560 5482 55968 5510
rect 55454 5474 55520 5482
rect 55602 5478 55968 5482
rect 55406 5435 55468 5444
rect 55406 5401 55422 5435
rect 55456 5401 55468 5435
rect 55406 5384 55468 5401
rect 55410 5382 55468 5384
rect 55464 5327 55554 5348
rect 55464 5318 55491 5327
rect 53637 5293 55491 5318
rect 55525 5318 55554 5327
rect 56068 5318 56146 6276
rect 56234 6264 56858 6296
rect 56966 6331 57032 6342
rect 56966 6297 56982 6331
rect 57016 6297 57032 6331
rect 56966 6286 57032 6297
rect 57118 6294 57152 6440
rect 57300 6438 57358 6440
rect 57556 6459 57624 6464
rect 57556 6456 57584 6459
rect 57556 6404 57564 6456
rect 57618 6425 57624 6459
rect 57616 6404 57624 6425
rect 57354 6383 57444 6404
rect 57556 6398 57624 6404
rect 57354 6349 57381 6383
rect 57415 6349 57444 6383
rect 57578 6378 57624 6398
rect 57666 6531 57712 6578
rect 57666 6497 57672 6531
rect 57706 6497 57712 6531
rect 57666 6459 57712 6497
rect 57666 6425 57672 6459
rect 57706 6425 57712 6459
rect 57666 6404 57712 6425
rect 58820 6531 58866 6578
rect 58820 6497 58826 6531
rect 58860 6497 58866 6531
rect 58820 6459 58866 6497
rect 58820 6425 58826 6459
rect 58860 6425 58866 6459
rect 58908 6531 58954 6578
rect 58908 6497 58914 6531
rect 58948 6497 58954 6531
rect 58908 6459 58954 6497
rect 59008 6500 59068 6732
rect 59096 7022 59136 7056
rect 59170 7022 59176 7056
rect 59096 6984 59176 7022
rect 59216 7062 59282 7068
rect 59216 7010 59222 7062
rect 59274 7010 59282 7062
rect 59216 7004 59282 7010
rect 59322 7056 59424 7068
rect 59322 7022 59328 7056
rect 59362 7022 59424 7056
rect 59096 6950 59136 6984
rect 59170 6950 59176 6984
rect 59096 6938 59176 6950
rect 59226 6984 59272 7004
rect 59226 6950 59232 6984
rect 59266 6950 59272 6984
rect 59226 6938 59272 6950
rect 59322 6984 59424 7022
rect 59322 6950 59328 6984
rect 59362 6950 59424 6984
rect 59322 6938 59424 6950
rect 59096 6738 59142 6938
rect 59172 6900 59230 6910
rect 59172 6866 59184 6900
rect 59218 6866 59230 6900
rect 59172 6848 59230 6866
rect 59374 6858 59424 6938
rect 59790 6916 59874 7186
rect 59532 6906 59590 6912
rect 59524 6900 59598 6906
rect 59284 6819 59342 6836
rect 59284 6785 59296 6819
rect 59330 6785 59342 6819
rect 59284 6770 59342 6785
rect 59374 6792 59444 6858
rect 59524 6848 59535 6900
rect 59587 6848 59598 6900
rect 59524 6842 59598 6848
rect 59666 6890 59942 6916
rect 59666 6885 59767 6890
rect 59819 6885 59942 6890
rect 59666 6851 59695 6885
rect 59729 6851 59767 6885
rect 59821 6851 59879 6885
rect 59913 6851 59942 6885
rect 59532 6834 59590 6842
rect 59666 6838 59767 6851
rect 59819 6838 59942 6851
rect 59666 6820 59942 6838
rect 59374 6738 59424 6792
rect 59096 6691 59192 6738
rect 59096 6657 59152 6691
rect 59186 6657 59192 6691
rect 59096 6619 59192 6657
rect 59096 6585 59152 6619
rect 59186 6585 59192 6619
rect 59242 6691 59288 6738
rect 59242 6657 59248 6691
rect 59282 6657 59288 6691
rect 59242 6619 59288 6657
rect 59242 6598 59248 6619
rect 59096 6538 59192 6585
rect 59232 6590 59248 6598
rect 59282 6598 59288 6619
rect 59338 6691 59424 6738
rect 59338 6657 59344 6691
rect 59378 6657 59424 6691
rect 59338 6619 59424 6657
rect 59282 6590 59298 6598
rect 59232 6538 59240 6590
rect 59292 6538 59298 6590
rect 59338 6585 59344 6619
rect 59378 6585 59424 6619
rect 59500 6659 59566 6672
rect 59500 6625 59516 6659
rect 59550 6625 59566 6659
rect 59894 6652 59962 6654
rect 59500 6614 59566 6625
rect 59810 6648 59962 6652
rect 59810 6642 59903 6648
rect 59810 6608 59830 6642
rect 59864 6608 59903 6642
rect 59810 6602 59903 6608
rect 59894 6596 59903 6602
rect 59955 6596 59962 6648
rect 59894 6590 59962 6596
rect 59338 6542 59424 6585
rect 59338 6538 59384 6542
rect 59232 6530 59298 6538
rect 59466 6531 59512 6578
rect 59008 6491 59246 6500
rect 59008 6468 59200 6491
rect 58908 6442 58914 6459
rect 57666 6376 57738 6404
rect 58820 6378 58866 6425
rect 58896 6436 58914 6442
rect 58948 6442 58954 6459
rect 59006 6457 59200 6468
rect 59234 6457 59246 6491
rect 59466 6497 59472 6531
rect 59506 6497 59512 6531
rect 59466 6464 59512 6497
rect 58948 6436 58962 6442
rect 58896 6384 58902 6436
rect 58954 6384 58962 6436
rect 58896 6378 58962 6384
rect 59006 6440 59246 6457
rect 57354 6328 57444 6349
rect 57612 6331 57678 6340
rect 57612 6297 57628 6331
rect 57662 6297 57678 6331
rect 57612 6294 57678 6297
rect 57118 6266 57678 6294
rect 57022 6210 57090 6224
rect 57022 6176 57040 6210
rect 57074 6176 57090 6210
rect 57022 6166 57090 6176
rect 57062 5862 57090 6166
rect 57118 6084 57152 6266
rect 57450 6200 57522 6212
rect 57450 6148 57460 6200
rect 57512 6148 57522 6200
rect 57450 6136 57522 6148
rect 57374 6084 57438 6102
rect 57118 6050 57390 6084
rect 57424 6050 57438 6084
rect 57374 6040 57438 6050
rect 57710 6026 57738 6376
rect 57778 6342 58054 6372
rect 57778 6341 57810 6342
rect 57862 6341 58054 6342
rect 57778 6307 57807 6341
rect 57862 6307 57899 6341
rect 57933 6307 57991 6341
rect 58025 6307 58054 6341
rect 57778 6290 57810 6307
rect 57862 6290 58054 6307
rect 57778 6276 58054 6290
rect 58122 6348 58746 6366
rect 58122 6335 58664 6348
rect 58122 6301 58153 6335
rect 58187 6301 58245 6335
rect 58279 6301 58337 6335
rect 58371 6333 58664 6335
rect 58716 6333 58746 6348
rect 58371 6301 58499 6333
rect 58122 6299 58499 6301
rect 58533 6299 58591 6333
rect 58625 6299 58664 6333
rect 58717 6299 58746 6333
rect 58122 6296 58664 6299
rect 58716 6296 58746 6299
rect 57828 6084 57894 6090
rect 57828 6032 57834 6084
rect 57886 6032 57894 6084
rect 57828 6026 57894 6032
rect 57484 6012 57738 6026
rect 57240 6000 57286 6012
rect 56786 5834 57090 5862
rect 57206 5966 57246 6000
rect 57280 5966 57286 6000
rect 57206 5928 57286 5966
rect 57326 6006 57392 6012
rect 57326 5954 57332 6006
rect 57384 5954 57392 6006
rect 57326 5948 57392 5954
rect 57432 6000 57738 6012
rect 57432 5966 57438 6000
rect 57472 5998 57738 6000
rect 57472 5966 57534 5998
rect 57206 5894 57246 5928
rect 57280 5894 57286 5928
rect 57206 5882 57286 5894
rect 57336 5928 57382 5948
rect 57336 5894 57342 5928
rect 57376 5894 57382 5928
rect 57336 5882 57382 5894
rect 57432 5928 57534 5966
rect 57432 5894 57438 5928
rect 57472 5894 57534 5928
rect 57432 5882 57534 5894
rect 57654 5951 57888 5960
rect 57654 5899 57660 5951
rect 57712 5932 57836 5951
rect 57712 5899 57718 5932
rect 57654 5892 57718 5899
rect 57830 5899 57836 5932
rect 57888 5899 57894 5932
rect 57830 5892 57894 5899
rect 56786 5831 57062 5834
rect 56786 5797 56815 5831
rect 56849 5797 56907 5831
rect 56941 5797 56999 5831
rect 57033 5797 57062 5831
rect 56786 5766 57062 5797
rect 56892 5718 56956 5724
rect 56892 5666 56898 5718
rect 56950 5666 56956 5718
rect 56892 5660 56956 5666
rect 57206 5682 57252 5882
rect 57282 5844 57340 5854
rect 57282 5810 57294 5844
rect 57328 5810 57340 5844
rect 57282 5792 57340 5810
rect 57394 5763 57452 5780
rect 57394 5729 57406 5763
rect 57440 5729 57452 5763
rect 57394 5714 57452 5729
rect 57484 5682 57534 5882
rect 57600 5831 57876 5862
rect 57600 5797 57629 5831
rect 57663 5797 57721 5831
rect 57755 5797 57813 5831
rect 57847 5797 57876 5831
rect 57600 5766 57876 5797
rect 57206 5635 57302 5682
rect 56804 5602 56868 5608
rect 56804 5550 56810 5602
rect 56862 5550 56868 5602
rect 56804 5544 56868 5550
rect 56974 5592 57044 5610
rect 56974 5558 56995 5592
rect 57029 5558 57044 5592
rect 56974 5550 57044 5558
rect 57206 5601 57262 5635
rect 57296 5601 57302 5635
rect 57206 5563 57302 5601
rect 56974 5514 57002 5550
rect 57206 5529 57262 5563
rect 57296 5529 57302 5563
rect 57352 5635 57398 5682
rect 57352 5601 57358 5635
rect 57392 5601 57398 5635
rect 57352 5563 57398 5601
rect 57352 5542 57358 5563
rect 57206 5514 57302 5529
rect 56974 5482 57302 5514
rect 57342 5534 57358 5542
rect 57392 5542 57398 5563
rect 57448 5635 57534 5682
rect 57706 5716 57774 5726
rect 57706 5664 57714 5716
rect 57766 5664 57774 5716
rect 57706 5658 57774 5664
rect 57448 5601 57454 5635
rect 57488 5601 57534 5635
rect 57448 5563 57534 5601
rect 57392 5534 57408 5542
rect 57342 5482 57350 5534
rect 57402 5482 57408 5534
rect 57448 5529 57454 5563
rect 57488 5529 57534 5563
rect 57616 5604 57684 5610
rect 57616 5552 57622 5604
rect 57674 5552 57684 5604
rect 57616 5546 57684 5552
rect 57790 5590 57856 5602
rect 57790 5556 57807 5590
rect 57841 5556 57856 5590
rect 57790 5548 57856 5556
rect 57448 5510 57534 5529
rect 57828 5510 57856 5548
rect 57448 5482 57856 5510
rect 57342 5474 57408 5482
rect 57490 5478 57856 5482
rect 57294 5435 57356 5444
rect 57294 5401 57310 5435
rect 57344 5401 57356 5435
rect 57294 5384 57356 5401
rect 57298 5382 57356 5384
rect 57352 5327 57442 5348
rect 57352 5318 57379 5327
rect 55525 5293 57379 5318
rect 57413 5318 57442 5327
rect 57956 5318 58034 6276
rect 58122 6264 58746 6296
rect 58854 6331 58920 6342
rect 58854 6297 58870 6331
rect 58904 6297 58920 6331
rect 58854 6286 58920 6297
rect 59006 6294 59040 6440
rect 59188 6438 59246 6440
rect 59444 6459 59512 6464
rect 59444 6456 59472 6459
rect 59444 6404 59452 6456
rect 59506 6425 59512 6459
rect 59504 6404 59512 6425
rect 59242 6383 59332 6404
rect 59444 6398 59512 6404
rect 59242 6349 59269 6383
rect 59303 6349 59332 6383
rect 59466 6378 59512 6398
rect 59554 6531 59600 6578
rect 59554 6497 59560 6531
rect 59594 6497 59600 6531
rect 59554 6459 59600 6497
rect 59554 6425 59560 6459
rect 59594 6425 59600 6459
rect 59554 6404 59600 6425
rect 59554 6376 59626 6404
rect 59242 6328 59332 6349
rect 59500 6331 59566 6340
rect 59500 6297 59516 6331
rect 59550 6297 59566 6331
rect 59500 6294 59566 6297
rect 59006 6266 59566 6294
rect 58910 6210 58978 6224
rect 58910 6176 58928 6210
rect 58962 6176 58978 6210
rect 58910 6166 58978 6176
rect 58950 5862 58978 6166
rect 59006 6084 59040 6266
rect 59338 6200 59410 6212
rect 59338 6148 59348 6200
rect 59400 6148 59410 6200
rect 59338 6136 59410 6148
rect 59262 6084 59326 6102
rect 59006 6050 59278 6084
rect 59312 6050 59326 6084
rect 59262 6040 59326 6050
rect 59598 6026 59626 6376
rect 59666 6342 59942 6372
rect 59666 6341 59698 6342
rect 59750 6341 59942 6342
rect 59666 6307 59695 6341
rect 59750 6307 59787 6341
rect 59821 6307 59879 6341
rect 59913 6307 59942 6341
rect 59666 6290 59698 6307
rect 59750 6290 59942 6307
rect 59666 6276 59942 6290
rect 59716 6084 59782 6090
rect 59716 6032 59722 6084
rect 59774 6032 59782 6084
rect 59716 6026 59782 6032
rect 59372 6012 59626 6026
rect 59128 6000 59174 6012
rect 58674 5834 58978 5862
rect 59094 5966 59134 6000
rect 59168 5966 59174 6000
rect 59094 5928 59174 5966
rect 59214 6006 59280 6012
rect 59214 5954 59220 6006
rect 59272 5954 59280 6006
rect 59214 5948 59280 5954
rect 59320 6000 59626 6012
rect 59320 5966 59326 6000
rect 59360 5998 59626 6000
rect 59360 5966 59422 5998
rect 59094 5894 59134 5928
rect 59168 5894 59174 5928
rect 59094 5882 59174 5894
rect 59224 5928 59270 5948
rect 59224 5894 59230 5928
rect 59264 5894 59270 5928
rect 59224 5882 59270 5894
rect 59320 5928 59422 5966
rect 59320 5894 59326 5928
rect 59360 5894 59422 5928
rect 59320 5882 59422 5894
rect 59542 5951 59776 5960
rect 59542 5899 59548 5951
rect 59600 5932 59724 5951
rect 59600 5899 59606 5932
rect 59542 5892 59606 5899
rect 59718 5899 59724 5932
rect 59776 5899 59782 5932
rect 59718 5892 59782 5899
rect 58674 5831 58950 5834
rect 58674 5797 58703 5831
rect 58737 5797 58795 5831
rect 58829 5797 58887 5831
rect 58921 5797 58950 5831
rect 58674 5766 58950 5797
rect 58780 5718 58844 5724
rect 58780 5666 58786 5718
rect 58838 5666 58844 5718
rect 58780 5660 58844 5666
rect 59094 5682 59140 5882
rect 59170 5844 59228 5854
rect 59170 5810 59182 5844
rect 59216 5810 59228 5844
rect 59170 5792 59228 5810
rect 59282 5763 59340 5780
rect 59282 5729 59294 5763
rect 59328 5729 59340 5763
rect 59282 5714 59340 5729
rect 59372 5682 59422 5882
rect 59488 5831 59764 5862
rect 59488 5797 59517 5831
rect 59551 5797 59609 5831
rect 59643 5797 59701 5831
rect 59735 5797 59764 5831
rect 59488 5766 59764 5797
rect 59094 5635 59190 5682
rect 58692 5602 58756 5608
rect 58692 5550 58698 5602
rect 58750 5550 58756 5602
rect 58692 5544 58756 5550
rect 58862 5592 58932 5610
rect 58862 5558 58883 5592
rect 58917 5558 58932 5592
rect 58862 5550 58932 5558
rect 59094 5601 59150 5635
rect 59184 5601 59190 5635
rect 59094 5563 59190 5601
rect 58862 5514 58890 5550
rect 59094 5529 59150 5563
rect 59184 5529 59190 5563
rect 59240 5635 59286 5682
rect 59240 5601 59246 5635
rect 59280 5601 59286 5635
rect 59240 5563 59286 5601
rect 59240 5542 59246 5563
rect 59094 5514 59190 5529
rect 58862 5482 59190 5514
rect 59230 5534 59246 5542
rect 59280 5542 59286 5563
rect 59336 5635 59422 5682
rect 59594 5716 59662 5726
rect 59594 5664 59602 5716
rect 59654 5664 59662 5716
rect 59594 5658 59662 5664
rect 59336 5601 59342 5635
rect 59376 5601 59422 5635
rect 59336 5563 59422 5601
rect 59280 5534 59296 5542
rect 59230 5482 59238 5534
rect 59290 5482 59296 5534
rect 59336 5529 59342 5563
rect 59376 5529 59422 5563
rect 59504 5604 59572 5610
rect 59504 5552 59510 5604
rect 59562 5552 59572 5604
rect 59504 5546 59572 5552
rect 59678 5590 59744 5602
rect 59678 5556 59695 5590
rect 59729 5556 59744 5590
rect 59678 5548 59744 5556
rect 59336 5510 59422 5529
rect 59716 5510 59744 5548
rect 59336 5482 59744 5510
rect 59230 5474 59296 5482
rect 59378 5478 59744 5482
rect 59182 5435 59244 5444
rect 59182 5401 59198 5435
rect 59232 5401 59244 5435
rect 59182 5384 59244 5401
rect 59186 5382 59244 5384
rect 59240 5327 59330 5348
rect 59240 5318 59267 5327
rect 57413 5293 59267 5318
rect 59301 5318 59330 5327
rect 59844 5318 59922 6276
rect 59301 5293 59982 5318
rect -430 5287 59982 5293
rect -430 5253 187 5287
rect 221 5253 279 5287
rect 313 5253 371 5287
rect 405 5253 1001 5287
rect 1035 5253 1093 5287
rect 1127 5253 1185 5287
rect 1219 5253 2075 5287
rect 2109 5253 2167 5287
rect 2201 5253 2259 5287
rect 2293 5253 2889 5287
rect 2923 5253 2981 5287
rect 3015 5253 3073 5287
rect 3107 5253 3963 5287
rect 3997 5253 4055 5287
rect 4089 5253 4147 5287
rect 4181 5253 4777 5287
rect 4811 5253 4869 5287
rect 4903 5253 4961 5287
rect 4995 5253 5851 5287
rect 5885 5253 5943 5287
rect 5977 5253 6035 5287
rect 6069 5253 6665 5287
rect 6699 5253 6757 5287
rect 6791 5253 6849 5287
rect 6883 5253 7739 5287
rect 7773 5253 7831 5287
rect 7865 5253 7923 5287
rect 7957 5253 8553 5287
rect 8587 5253 8645 5287
rect 8679 5253 8737 5287
rect 8771 5253 9627 5287
rect 9661 5253 9719 5287
rect 9753 5253 9811 5287
rect 9845 5253 10441 5287
rect 10475 5253 10533 5287
rect 10567 5253 10625 5287
rect 10659 5253 11515 5287
rect 11549 5253 11607 5287
rect 11641 5253 11699 5287
rect 11733 5253 12329 5287
rect 12363 5253 12421 5287
rect 12455 5253 12513 5287
rect 12547 5253 13403 5287
rect 13437 5253 13495 5287
rect 13529 5253 13587 5287
rect 13621 5253 14217 5287
rect 14251 5253 14309 5287
rect 14343 5253 14401 5287
rect 14435 5253 15285 5287
rect 15319 5253 15377 5287
rect 15411 5253 15469 5287
rect 15503 5253 16099 5287
rect 16133 5253 16191 5287
rect 16225 5253 16283 5287
rect 16317 5253 17173 5287
rect 17207 5253 17265 5287
rect 17299 5253 17357 5287
rect 17391 5253 17987 5287
rect 18021 5253 18079 5287
rect 18113 5253 18171 5287
rect 18205 5253 19061 5287
rect 19095 5253 19153 5287
rect 19187 5253 19245 5287
rect 19279 5253 19875 5287
rect 19909 5253 19967 5287
rect 20001 5253 20059 5287
rect 20093 5253 20949 5287
rect 20983 5253 21041 5287
rect 21075 5253 21133 5287
rect 21167 5253 21763 5287
rect 21797 5253 21855 5287
rect 21889 5253 21947 5287
rect 21981 5253 22837 5287
rect 22871 5253 22929 5287
rect 22963 5253 23021 5287
rect 23055 5253 23651 5287
rect 23685 5253 23743 5287
rect 23777 5253 23835 5287
rect 23869 5253 24725 5287
rect 24759 5253 24817 5287
rect 24851 5253 24909 5287
rect 24943 5253 25539 5287
rect 25573 5253 25631 5287
rect 25665 5253 25723 5287
rect 25757 5253 26613 5287
rect 26647 5253 26705 5287
rect 26739 5253 26797 5287
rect 26831 5253 27427 5287
rect 27461 5253 27519 5287
rect 27553 5253 27611 5287
rect 27645 5253 28501 5287
rect 28535 5253 28593 5287
rect 28627 5253 28685 5287
rect 28719 5253 29315 5287
rect 29349 5253 29407 5287
rect 29441 5253 29499 5287
rect 29533 5253 30389 5287
rect 30423 5253 30481 5287
rect 30515 5253 30573 5287
rect 30607 5253 31203 5287
rect 31237 5253 31295 5287
rect 31329 5253 31387 5287
rect 31421 5253 32277 5287
rect 32311 5253 32369 5287
rect 32403 5253 32461 5287
rect 32495 5253 33091 5287
rect 33125 5253 33183 5287
rect 33217 5253 33275 5287
rect 33309 5253 34165 5287
rect 34199 5253 34257 5287
rect 34291 5253 34349 5287
rect 34383 5253 34979 5287
rect 35013 5253 35071 5287
rect 35105 5253 35163 5287
rect 35197 5253 36053 5287
rect 36087 5253 36145 5287
rect 36179 5253 36237 5287
rect 36271 5253 36867 5287
rect 36901 5253 36959 5287
rect 36993 5253 37051 5287
rect 37085 5253 37941 5287
rect 37975 5253 38033 5287
rect 38067 5253 38125 5287
rect 38159 5253 38755 5287
rect 38789 5253 38847 5287
rect 38881 5253 38939 5287
rect 38973 5253 39829 5287
rect 39863 5253 39921 5287
rect 39955 5253 40013 5287
rect 40047 5253 40643 5287
rect 40677 5253 40735 5287
rect 40769 5253 40827 5287
rect 40861 5253 41717 5287
rect 41751 5253 41809 5287
rect 41843 5253 41901 5287
rect 41935 5253 42531 5287
rect 42565 5253 42623 5287
rect 42657 5253 42715 5287
rect 42749 5253 43605 5287
rect 43639 5253 43697 5287
rect 43731 5253 43789 5287
rect 43823 5253 44419 5287
rect 44453 5253 44511 5287
rect 44545 5253 44603 5287
rect 44637 5253 45487 5287
rect 45521 5253 45579 5287
rect 45613 5253 45671 5287
rect 45705 5253 46301 5287
rect 46335 5253 46393 5287
rect 46427 5253 46485 5287
rect 46519 5253 47375 5287
rect 47409 5253 47467 5287
rect 47501 5253 47559 5287
rect 47593 5253 48189 5287
rect 48223 5253 48281 5287
rect 48315 5253 48373 5287
rect 48407 5253 49263 5287
rect 49297 5253 49355 5287
rect 49389 5253 49447 5287
rect 49481 5253 50077 5287
rect 50111 5253 50169 5287
rect 50203 5253 50261 5287
rect 50295 5253 51151 5287
rect 51185 5253 51243 5287
rect 51277 5253 51335 5287
rect 51369 5253 51965 5287
rect 51999 5253 52057 5287
rect 52091 5253 52149 5287
rect 52183 5253 53039 5287
rect 53073 5253 53131 5287
rect 53165 5253 53223 5287
rect 53257 5253 53853 5287
rect 53887 5253 53945 5287
rect 53979 5253 54037 5287
rect 54071 5253 54927 5287
rect 54961 5253 55019 5287
rect 55053 5253 55111 5287
rect 55145 5253 55741 5287
rect 55775 5253 55833 5287
rect 55867 5253 55925 5287
rect 55959 5253 56815 5287
rect 56849 5253 56907 5287
rect 56941 5253 56999 5287
rect 57033 5253 57629 5287
rect 57663 5253 57721 5287
rect 57755 5253 57813 5287
rect 57847 5253 58703 5287
rect 58737 5253 58795 5287
rect 58829 5253 58887 5287
rect 58921 5253 59517 5287
rect 59551 5253 59609 5287
rect 59643 5253 59701 5287
rect 59735 5253 59982 5287
rect -430 5252 59982 5253
rect -430 5136 -377 5252
rect -69 5136 1511 5252
rect 1819 5136 3399 5252
rect 3707 5136 5287 5252
rect 5595 5209 7175 5252
rect 5595 5175 5693 5209
rect 5727 5175 5785 5209
rect 5819 5175 5877 5209
rect 5911 5175 5969 5209
rect 6003 5175 6061 5209
rect 6095 5175 6153 5209
rect 6187 5175 6245 5209
rect 6279 5175 6337 5209
rect 6371 5175 6429 5209
rect 6463 5175 6521 5209
rect 6555 5175 6613 5209
rect 6647 5175 6705 5209
rect 6739 5175 6797 5209
rect 6831 5175 6889 5209
rect 6923 5175 6981 5209
rect 7015 5175 7073 5209
rect 7107 5175 7175 5209
rect 5595 5136 7175 5175
rect 7483 5207 9063 5252
rect 7483 5173 7575 5207
rect 7609 5173 7667 5207
rect 7701 5173 7759 5207
rect 7793 5173 7851 5207
rect 7885 5173 7943 5207
rect 7977 5173 8035 5207
rect 8069 5173 8127 5207
rect 8161 5173 8219 5207
rect 8253 5173 8311 5207
rect 8345 5173 8403 5207
rect 8437 5173 8495 5207
rect 8529 5173 8587 5207
rect 8621 5173 8679 5207
rect 8713 5173 8771 5207
rect 8805 5173 8863 5207
rect 8897 5173 8955 5207
rect 8989 5173 9063 5207
rect 7483 5136 9063 5173
rect 9371 5136 10951 5252
rect 11259 5136 12839 5252
rect 13147 5136 14721 5252
rect 15029 5136 16609 5252
rect 16917 5136 18497 5252
rect 18805 5136 20385 5252
rect 20693 5209 22273 5252
rect 20693 5175 20791 5209
rect 20825 5175 20883 5209
rect 20917 5175 20975 5209
rect 21009 5175 21067 5209
rect 21101 5175 21159 5209
rect 21193 5175 21251 5209
rect 21285 5175 21343 5209
rect 21377 5175 21435 5209
rect 21469 5175 21527 5209
rect 21561 5175 21619 5209
rect 21653 5175 21711 5209
rect 21745 5175 21803 5209
rect 21837 5175 21895 5209
rect 21929 5175 21987 5209
rect 22021 5175 22079 5209
rect 22113 5175 22171 5209
rect 22205 5175 22273 5209
rect 20693 5136 22273 5175
rect 22581 5207 24161 5252
rect 22581 5173 22673 5207
rect 22707 5173 22765 5207
rect 22799 5173 22857 5207
rect 22891 5173 22949 5207
rect 22983 5173 23041 5207
rect 23075 5173 23133 5207
rect 23167 5173 23225 5207
rect 23259 5173 23317 5207
rect 23351 5173 23409 5207
rect 23443 5173 23501 5207
rect 23535 5173 23593 5207
rect 23627 5173 23685 5207
rect 23719 5173 23777 5207
rect 23811 5173 23869 5207
rect 23903 5173 23961 5207
rect 23995 5173 24053 5207
rect 24087 5173 24161 5207
rect 22581 5136 24161 5173
rect 24469 5136 26049 5252
rect 26357 5136 27937 5252
rect 28245 5136 29825 5252
rect 30133 5136 31713 5252
rect 32021 5136 33601 5252
rect 33909 5136 35489 5252
rect 35797 5209 37377 5252
rect 35797 5175 35895 5209
rect 35929 5175 35987 5209
rect 36021 5175 36079 5209
rect 36113 5175 36171 5209
rect 36205 5175 36263 5209
rect 36297 5175 36355 5209
rect 36389 5175 36447 5209
rect 36481 5175 36539 5209
rect 36573 5175 36631 5209
rect 36665 5175 36723 5209
rect 36757 5175 36815 5209
rect 36849 5175 36907 5209
rect 36941 5175 36999 5209
rect 37033 5175 37091 5209
rect 37125 5175 37183 5209
rect 37217 5175 37275 5209
rect 37309 5175 37377 5209
rect 35797 5136 37377 5175
rect 37685 5207 39265 5252
rect 37685 5173 37777 5207
rect 37811 5173 37869 5207
rect 37903 5173 37961 5207
rect 37995 5173 38053 5207
rect 38087 5173 38145 5207
rect 38179 5173 38237 5207
rect 38271 5173 38329 5207
rect 38363 5173 38421 5207
rect 38455 5173 38513 5207
rect 38547 5173 38605 5207
rect 38639 5173 38697 5207
rect 38731 5173 38789 5207
rect 38823 5173 38881 5207
rect 38915 5173 38973 5207
rect 39007 5173 39065 5207
rect 39099 5173 39157 5207
rect 39191 5173 39265 5207
rect 37685 5136 39265 5173
rect 39573 5136 41153 5252
rect 41461 5136 43041 5252
rect 43349 5136 44923 5252
rect 45231 5136 46811 5252
rect 47119 5136 48699 5252
rect 49007 5136 50587 5252
rect 50895 5209 52475 5252
rect 50895 5175 50993 5209
rect 51027 5175 51085 5209
rect 51119 5175 51177 5209
rect 51211 5175 51269 5209
rect 51303 5175 51361 5209
rect 51395 5175 51453 5209
rect 51487 5175 51545 5209
rect 51579 5175 51637 5209
rect 51671 5175 51729 5209
rect 51763 5175 51821 5209
rect 51855 5175 51913 5209
rect 51947 5175 52005 5209
rect 52039 5175 52097 5209
rect 52131 5175 52189 5209
rect 52223 5175 52281 5209
rect 52315 5175 52373 5209
rect 52407 5175 52475 5209
rect 50895 5136 52475 5175
rect 52783 5207 54363 5252
rect 52783 5173 52875 5207
rect 52909 5173 52967 5207
rect 53001 5173 53059 5207
rect 53093 5173 53151 5207
rect 53185 5173 53243 5207
rect 53277 5173 53335 5207
rect 53369 5173 53427 5207
rect 53461 5173 53519 5207
rect 53553 5173 53611 5207
rect 53645 5173 53703 5207
rect 53737 5173 53795 5207
rect 53829 5173 53887 5207
rect 53921 5173 53979 5207
rect 54013 5173 54071 5207
rect 54105 5173 54163 5207
rect 54197 5173 54255 5207
rect 54289 5173 54363 5207
rect 52783 5136 54363 5173
rect 54671 5136 56251 5252
rect 56559 5136 58139 5252
rect 58447 5136 59982 5252
rect -430 5064 59982 5136
rect 5765 5019 7021 5034
rect 5765 5005 5864 5019
rect 5765 4971 5799 5005
rect 5833 4971 5864 5005
rect 5765 4967 5864 4971
rect 5916 5009 5979 5019
rect 5916 4975 5962 5009
rect 5916 4967 5979 4975
rect 6031 4967 6106 5019
rect 6158 5007 6223 5019
rect 6166 4973 6223 5007
rect 6158 4967 6223 4973
rect 6275 5007 6337 5019
rect 6275 4973 6297 5007
rect 6331 4973 6337 5007
rect 6275 4967 6337 4973
rect 6389 5018 7021 5019
rect 6389 4967 6456 5018
rect 5765 4966 6456 4967
rect 6508 4966 6554 5018
rect 6606 4996 6650 5018
rect 6606 4966 6637 4996
rect 6702 4966 6758 5018
rect 6810 5001 6857 5018
rect 6833 4967 6857 5001
rect 6810 4966 6857 4967
rect 6909 4966 6951 5018
rect 7003 5002 7021 5018
rect 7006 4968 7021 5002
rect 7003 4966 7021 4968
rect 5765 4959 6466 4966
rect 6500 4962 6637 4966
rect 6671 4962 7021 4966
rect 6500 4959 7021 4962
rect 5765 4950 7021 4959
rect 7640 5017 8907 5032
rect 7640 4965 7665 5017
rect 7717 4965 7761 5017
rect 7813 5016 8907 5017
rect 7813 5003 7850 5016
rect 7813 4969 7845 5003
rect 7813 4965 7850 4969
rect 7640 4964 7850 4965
rect 7902 4964 7950 5016
rect 8002 5012 8047 5016
rect 8002 4978 8015 5012
rect 8099 5010 8184 5016
rect 8002 4964 8047 4978
rect 8099 4976 8183 5010
rect 8099 4964 8184 4976
rect 8236 4964 8338 5016
rect 8390 5014 8907 5016
rect 8390 4964 8464 5014
rect 8516 5002 8566 5014
rect 8549 4968 8566 5002
rect 7640 4963 8350 4964
rect 8384 4963 8464 4964
rect 7640 4962 8464 4963
rect 8516 4962 8566 4968
rect 8618 4962 8673 5014
rect 8725 5012 8907 5014
rect 8725 4962 8785 5012
rect 7640 4960 8785 4962
rect 8837 5001 8907 5012
rect 8837 4967 8851 5001
rect 8885 4967 8907 5001
rect 8837 4960 8907 4967
rect 7640 4948 8907 4960
rect 6168 4900 8859 4906
rect 6168 4866 6318 4900
rect 6352 4866 6426 4900
rect 6460 4866 6534 4900
rect 6568 4866 6642 4900
rect 6676 4866 6750 4900
rect 6784 4866 6858 4900
rect 6892 4866 6966 4900
rect 7000 4866 7074 4900
rect 7108 4866 7930 4900
rect 7964 4866 8081 4900
rect 8115 4866 8178 4900
rect 8212 4866 8275 4900
rect 8309 4866 8372 4900
rect 8406 4866 8469 4900
rect 8503 4866 8566 4900
rect 8600 4866 8663 4900
rect 8697 4866 8760 4900
rect 8794 4866 8859 4900
rect 6168 4860 8859 4866
rect 7230 4813 7428 4860
rect 7230 4761 7264 4813
rect 7316 4812 7428 4813
rect 7316 4761 7345 4812
rect 7230 4760 7345 4761
rect 7397 4760 7428 4812
rect 7230 4746 7428 4760
rect 14423 4747 14678 5064
rect 20882 5021 22108 5034
rect 20882 5020 21676 5021
rect 20882 4968 20891 5020
rect 20943 4968 20988 5020
rect 21040 4998 21085 5020
rect 21040 4968 21060 4998
rect 21137 4968 21191 5020
rect 21243 5000 21296 5020
rect 21264 4968 21296 5000
rect 21348 5006 21413 5020
rect 21465 5019 21676 5020
rect 21348 4972 21400 5006
rect 21348 4968 21413 4972
rect 21465 4968 21547 5019
rect 21599 5018 21676 5019
rect 20882 4962 20901 4968
rect 20935 4964 21060 4968
rect 21094 4966 21230 4968
rect 21264 4967 21547 4968
rect 21264 4966 21554 4967
rect 21606 4969 21676 5018
rect 21728 5003 21792 5021
rect 21728 4969 21733 5003
rect 21767 4969 21792 5003
rect 21844 4969 21898 5021
rect 21950 4969 22005 5021
rect 22057 4997 22108 5021
rect 22057 4969 22060 4997
rect 21606 4966 21900 4969
rect 21094 4964 21564 4966
rect 20935 4962 21564 4964
rect 20882 4959 21564 4962
rect 21598 4963 21900 4966
rect 21934 4963 22060 4969
rect 22094 4963 22108 4997
rect 21598 4959 22108 4963
rect 20882 4950 22108 4959
rect 22761 5018 23998 5032
rect 22761 5017 23565 5018
rect 22761 4994 22780 5017
rect 22761 4960 22774 4994
rect 22832 4965 22877 5017
rect 22929 4996 22974 5017
rect 22929 4965 22944 4996
rect 23026 4965 23080 5017
rect 23132 5002 23185 5017
rect 23144 4968 23185 5002
rect 23132 4965 23185 4968
rect 23237 5001 23302 5017
rect 23354 5016 23565 5017
rect 23237 4967 23279 5001
rect 23237 4965 23302 4967
rect 23354 4965 23436 5016
rect 22808 4962 22944 4965
rect 22978 4964 23436 4965
rect 23488 4966 23565 5016
rect 23617 4999 23681 5018
rect 23617 4966 23619 4999
rect 23488 4965 23619 4966
rect 23653 4966 23681 4999
rect 23733 4997 23787 5018
rect 23733 4966 23783 4997
rect 23839 4966 23894 5018
rect 23946 4995 23998 5018
rect 23946 4966 23949 4995
rect 23653 4965 23783 4966
rect 23488 4964 23783 4965
rect 22978 4963 23448 4964
rect 23482 4963 23783 4964
rect 23817 4963 23949 4966
rect 22978 4962 23949 4963
rect 22808 4961 23949 4962
rect 23983 4961 23998 4995
rect 22808 4960 23998 4961
rect 22761 4948 23998 4960
rect 21206 4900 24010 4906
rect 21206 4866 21458 4900
rect 21492 4866 21577 4900
rect 21611 4866 21696 4900
rect 21730 4866 21815 4900
rect 21849 4866 21934 4900
rect 21968 4866 22053 4900
rect 22087 4866 22172 4900
rect 22206 4866 23028 4900
rect 23062 4866 23132 4900
rect 23166 4866 23248 4900
rect 23282 4866 23361 4900
rect 23395 4866 23474 4900
rect 23508 4866 23587 4900
rect 23621 4866 23700 4900
rect 23734 4866 23813 4900
rect 23847 4866 23926 4900
rect 23960 4866 24010 4900
rect 21206 4860 24010 4866
rect 22334 4810 22540 4860
rect 22334 4758 22380 4810
rect 22432 4758 22475 4810
rect 22527 4758 22540 4810
rect 22334 4748 22540 4758
rect 30359 4770 30693 5064
rect 35967 5019 37223 5034
rect 35967 5005 36066 5019
rect 35967 4971 36001 5005
rect 36035 4971 36066 5005
rect 35967 4967 36066 4971
rect 36118 5009 36181 5019
rect 36118 4975 36164 5009
rect 36118 4967 36181 4975
rect 36233 4967 36308 5019
rect 36360 5007 36425 5019
rect 36368 4973 36425 5007
rect 36360 4967 36425 4973
rect 36477 5007 36539 5019
rect 36477 4973 36499 5007
rect 36533 4973 36539 5007
rect 36477 4967 36539 4973
rect 36591 5018 37223 5019
rect 36591 4967 36658 5018
rect 35967 4966 36658 4967
rect 36710 4966 36756 5018
rect 36808 4996 36852 5018
rect 36808 4966 36839 4996
rect 36904 4966 36960 5018
rect 37012 5001 37059 5018
rect 37035 4967 37059 5001
rect 37012 4966 37059 4967
rect 37111 4966 37153 5018
rect 37205 5002 37223 5018
rect 37208 4968 37223 5002
rect 37205 4966 37223 4968
rect 35967 4959 36668 4966
rect 36702 4962 36839 4966
rect 36873 4962 37223 4966
rect 36702 4959 37223 4962
rect 35967 4950 37223 4959
rect 37842 5017 39109 5032
rect 37842 4965 37867 5017
rect 37919 4965 37963 5017
rect 38015 5016 39109 5017
rect 38015 5003 38052 5016
rect 38015 4969 38047 5003
rect 38015 4965 38052 4969
rect 37842 4964 38052 4965
rect 38104 4964 38152 5016
rect 38204 5012 38249 5016
rect 38204 4978 38217 5012
rect 38301 5010 38386 5016
rect 38204 4964 38249 4978
rect 38301 4976 38385 5010
rect 38301 4964 38386 4976
rect 38438 4964 38540 5016
rect 38592 5014 39109 5016
rect 38592 4964 38666 5014
rect 38718 5002 38768 5014
rect 38751 4968 38768 5002
rect 37842 4963 38552 4964
rect 38586 4963 38666 4964
rect 37842 4962 38666 4963
rect 38718 4962 38768 4968
rect 38820 4962 38875 5014
rect 38927 5012 39109 5014
rect 38927 4962 38987 5012
rect 37842 4960 38987 4962
rect 39039 5001 39109 5012
rect 39039 4967 39053 5001
rect 39087 4967 39109 5001
rect 39039 4960 39109 4967
rect 37842 4948 39109 4960
rect 36370 4900 39061 4906
rect 36370 4866 36520 4900
rect 36554 4866 36628 4900
rect 36662 4866 36736 4900
rect 36770 4866 36844 4900
rect 36878 4866 36952 4900
rect 36986 4866 37060 4900
rect 37094 4866 37168 4900
rect 37202 4866 37276 4900
rect 37310 4866 38132 4900
rect 38166 4866 38283 4900
rect 38317 4866 38380 4900
rect 38414 4866 38477 4900
rect 38511 4866 38574 4900
rect 38608 4866 38671 4900
rect 38705 4866 38768 4900
rect 38802 4866 38865 4900
rect 38899 4866 38962 4900
rect 38996 4866 39061 4900
rect 36370 4860 39061 4866
rect 5664 4690 7136 4696
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14678 4747
rect 30359 4718 30402 4770
rect 30454 4718 30515 4770
rect 30567 4718 30616 4770
rect 30668 4718 30693 4770
rect 37432 4812 37630 4860
rect 37432 4760 37457 4812
rect 37509 4760 37559 4812
rect 37611 4760 37630 4812
rect 37432 4746 37630 4760
rect 44563 4747 44790 5064
rect 51084 5021 52310 5034
rect 51084 5020 51878 5021
rect 51084 4968 51093 5020
rect 51145 4968 51190 5020
rect 51242 4998 51287 5020
rect 51242 4968 51262 4998
rect 51339 4968 51393 5020
rect 51445 5000 51498 5020
rect 51466 4968 51498 5000
rect 51550 5006 51615 5020
rect 51667 5019 51878 5020
rect 51550 4972 51602 5006
rect 51550 4968 51615 4972
rect 51667 4968 51749 5019
rect 51801 5018 51878 5019
rect 51084 4962 51103 4968
rect 51137 4964 51262 4968
rect 51296 4966 51432 4968
rect 51466 4967 51749 4968
rect 51466 4966 51756 4967
rect 51808 4969 51878 5018
rect 51930 5003 51994 5021
rect 51930 4969 51935 5003
rect 51969 4969 51994 5003
rect 52046 4969 52100 5021
rect 52152 4969 52207 5021
rect 52259 4997 52310 5021
rect 52259 4969 52262 4997
rect 51808 4966 52102 4969
rect 51296 4964 51766 4966
rect 51137 4962 51766 4964
rect 51084 4959 51766 4962
rect 51800 4963 52102 4966
rect 52136 4963 52262 4969
rect 52296 4963 52310 4997
rect 51800 4959 52310 4963
rect 51084 4950 52310 4959
rect 52963 5018 54200 5032
rect 52963 5017 53767 5018
rect 52963 4994 52982 5017
rect 52963 4960 52976 4994
rect 53034 4965 53079 5017
rect 53131 4996 53176 5017
rect 53131 4965 53146 4996
rect 53228 4965 53282 5017
rect 53334 5002 53387 5017
rect 53346 4968 53387 5002
rect 53334 4965 53387 4968
rect 53439 5001 53504 5017
rect 53556 5016 53767 5017
rect 53439 4967 53481 5001
rect 53439 4965 53504 4967
rect 53556 4965 53638 5016
rect 53010 4962 53146 4965
rect 53180 4964 53638 4965
rect 53690 4966 53767 5016
rect 53819 4999 53883 5018
rect 53819 4966 53821 4999
rect 53690 4965 53821 4966
rect 53855 4966 53883 4999
rect 53935 4997 53989 5018
rect 53935 4966 53985 4997
rect 54041 4966 54096 5018
rect 54148 4995 54200 5018
rect 54148 4966 54151 4995
rect 53855 4965 53985 4966
rect 53690 4964 53985 4965
rect 53180 4963 53650 4964
rect 53684 4963 53985 4964
rect 54019 4963 54151 4966
rect 53180 4962 54151 4963
rect 53010 4961 54151 4962
rect 54185 4961 54200 4995
rect 53010 4960 54200 4961
rect 52963 4948 54200 4960
rect 51408 4900 54212 4906
rect 51408 4866 51660 4900
rect 51694 4866 51779 4900
rect 51813 4866 51898 4900
rect 51932 4866 52017 4900
rect 52051 4866 52136 4900
rect 52170 4866 52255 4900
rect 52289 4866 52374 4900
rect 52408 4866 53230 4900
rect 53264 4866 53334 4900
rect 53368 4866 53450 4900
rect 53484 4866 53563 4900
rect 53597 4866 53676 4900
rect 53710 4866 53789 4900
rect 53823 4866 53902 4900
rect 53936 4866 54015 4900
rect 54049 4866 54128 4900
rect 54162 4866 54212 4900
rect 51408 4860 54212 4866
rect 52536 4812 52742 4860
rect 7546 4690 9018 4694
rect 5664 4670 9018 4690
rect 5664 4669 6581 4670
rect 5664 4667 6379 4669
rect 5664 4665 6272 4667
rect 6324 4665 6379 4667
rect 6431 4665 6481 4669
rect 6533 4665 6581 4669
rect 6633 4665 9018 4670
rect 14423 4665 14678 4695
rect 20762 4673 22234 4696
rect 22644 4673 24116 4694
rect 30359 4674 30693 4718
rect 35866 4681 37338 4696
rect 44563 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 52529 4785 52742 4812
rect 52529 4733 52575 4785
rect 52627 4733 52670 4785
rect 52722 4748 52742 4785
rect 52722 4733 52735 4748
rect 52529 4723 52735 4733
rect 37748 4681 39220 4694
rect 35866 4674 39220 4681
rect 20762 4665 21302 4673
rect 21354 4665 21405 4673
rect 21457 4665 21488 4673
rect 21540 4665 21589 4673
rect 21641 4665 21676 4673
rect 21728 4665 24116 4673
rect 5664 4631 5693 4665
rect 5727 4631 5785 4665
rect 5819 4631 5877 4665
rect 5911 4631 5969 4665
rect 6003 4631 6061 4665
rect 6095 4631 6153 4665
rect 6187 4631 6245 4665
rect 6324 4631 6337 4665
rect 6371 4631 6379 4665
rect 6463 4631 6481 4665
rect 6555 4631 6581 4665
rect 6647 4631 6705 4665
rect 6739 4631 6797 4665
rect 6831 4631 6889 4665
rect 6923 4631 6981 4665
rect 7015 4631 7073 4665
rect 7107 4663 9018 4665
rect 7107 4631 7575 4663
rect 5664 4615 6272 4631
rect 6324 4617 6379 4631
rect 6431 4617 6481 4631
rect 6533 4618 6581 4631
rect 6633 4629 7575 4631
rect 7609 4629 7667 4663
rect 7701 4629 7759 4663
rect 7793 4629 7851 4663
rect 7885 4629 7943 4663
rect 7977 4629 8035 4663
rect 8069 4629 8127 4663
rect 8161 4629 8219 4663
rect 8253 4629 8311 4663
rect 8345 4629 8403 4663
rect 8437 4629 8495 4663
rect 8529 4629 8587 4663
rect 8621 4629 8679 4663
rect 8713 4629 8771 4663
rect 8805 4629 8863 4663
rect 8897 4629 8955 4663
rect 8989 4629 9018 4663
rect 6633 4618 9018 4629
rect 6533 4617 9018 4618
rect 6324 4615 9018 4617
rect 5664 4606 9018 4615
rect 5664 4600 7136 4606
rect 7546 4598 9018 4606
rect 20762 4631 20791 4665
rect 20825 4631 20883 4665
rect 20917 4631 20975 4665
rect 21009 4631 21067 4665
rect 21101 4631 21159 4665
rect 21193 4631 21251 4665
rect 21285 4631 21302 4665
rect 21377 4631 21405 4665
rect 21469 4631 21488 4665
rect 21561 4631 21589 4665
rect 21653 4631 21676 4665
rect 21745 4631 21803 4665
rect 21837 4631 21895 4665
rect 21929 4631 21987 4665
rect 22021 4631 22079 4665
rect 22113 4631 22171 4665
rect 22205 4663 24116 4665
rect 22205 4631 22673 4663
rect 20762 4621 21302 4631
rect 21354 4621 21405 4631
rect 21457 4621 21488 4631
rect 21540 4621 21589 4631
rect 21641 4621 21676 4631
rect 21728 4629 22673 4631
rect 22707 4629 22765 4663
rect 22799 4629 22857 4663
rect 22891 4629 22949 4663
rect 22983 4629 23041 4663
rect 23075 4629 23133 4663
rect 23167 4629 23225 4663
rect 23259 4629 23317 4663
rect 23351 4629 23409 4663
rect 23443 4629 23501 4663
rect 23535 4629 23593 4663
rect 23627 4629 23685 4663
rect 23719 4629 23777 4663
rect 23811 4629 23869 4663
rect 23903 4629 23961 4663
rect 23995 4629 24053 4663
rect 24087 4629 24116 4663
rect 21728 4621 24116 4629
rect 20762 4615 24116 4621
rect 20762 4600 22234 4615
rect 22644 4598 24116 4615
rect 35866 4669 36607 4674
rect 35866 4665 36434 4669
rect 35866 4631 35895 4665
rect 35929 4631 35987 4665
rect 36021 4631 36079 4665
rect 36113 4631 36171 4665
rect 36205 4631 36263 4665
rect 36297 4631 36355 4665
rect 36389 4631 36434 4665
rect 35866 4617 36434 4631
rect 36486 4617 36522 4669
rect 36574 4622 36607 4669
rect 36659 4665 39220 4674
rect 36665 4631 36723 4665
rect 36757 4631 36815 4665
rect 36849 4631 36907 4665
rect 36941 4631 36999 4665
rect 37033 4631 37091 4665
rect 37125 4631 37183 4665
rect 37217 4631 37275 4665
rect 37309 4663 39220 4665
rect 37309 4631 37777 4663
rect 36659 4629 37777 4631
rect 37811 4629 37869 4663
rect 37903 4629 37961 4663
rect 37995 4629 38053 4663
rect 38087 4629 38145 4663
rect 38179 4629 38237 4663
rect 38271 4629 38329 4663
rect 38363 4629 38421 4663
rect 38455 4629 38513 4663
rect 38547 4629 38605 4663
rect 38639 4629 38697 4663
rect 38731 4629 38789 4663
rect 38823 4629 38881 4663
rect 38915 4629 38973 4663
rect 39007 4629 39065 4663
rect 39099 4629 39157 4663
rect 39191 4629 39220 4663
rect 44563 4661 44790 4695
rect 50964 4687 52436 4696
rect 52846 4687 54318 4694
rect 50964 4666 54318 4687
rect 50964 4665 53350 4666
rect 36659 4623 39220 4629
rect 36659 4622 37338 4623
rect 36574 4617 37338 4622
rect 35866 4600 37338 4617
rect 37748 4598 39220 4623
rect 50964 4631 50993 4665
rect 51027 4631 51085 4665
rect 51119 4631 51177 4665
rect 51211 4631 51269 4665
rect 51303 4631 51361 4665
rect 51395 4631 51453 4665
rect 51487 4631 51545 4665
rect 51579 4631 51637 4665
rect 51671 4631 51729 4665
rect 51763 4631 51821 4665
rect 51855 4631 51913 4665
rect 51947 4631 52005 4665
rect 52039 4631 52097 4665
rect 52131 4631 52189 4665
rect 52223 4631 52281 4665
rect 52315 4631 52373 4665
rect 52407 4663 53350 4665
rect 53402 4663 53444 4666
rect 53496 4663 53521 4666
rect 53573 4665 53675 4666
rect 52407 4631 52875 4663
rect 50964 4629 52875 4631
rect 52909 4629 52967 4663
rect 53001 4629 53059 4663
rect 53093 4629 53151 4663
rect 53185 4629 53243 4663
rect 53277 4629 53335 4663
rect 53402 4629 53427 4663
rect 53496 4629 53519 4663
rect 50964 4600 52436 4629
rect 52846 4614 53350 4629
rect 53402 4614 53444 4629
rect 53496 4614 53521 4629
rect 53573 4614 53601 4665
rect 52846 4613 53601 4614
rect 53653 4614 53675 4665
rect 53727 4663 54318 4666
rect 53737 4629 53795 4663
rect 53829 4629 53887 4663
rect 53921 4629 53979 4663
rect 54013 4629 54071 4663
rect 54105 4629 54163 4663
rect 54197 4629 54255 4663
rect 54289 4629 54318 4663
rect 53727 4614 54318 4629
rect 53653 4613 54318 4614
rect 52846 4598 54318 4613
rect 30027 4150 32062 4163
rect 30027 4147 30517 4150
rect 30027 4132 30414 4147
rect 30027 4098 30056 4132
rect 30090 4098 30148 4132
rect 30182 4098 30240 4132
rect 30274 4098 30332 4132
rect 30366 4098 30414 4132
rect 30466 4098 30517 4147
rect 30569 4132 30618 4150
rect 30569 4098 30584 4132
rect 30670 4132 32062 4150
rect 30670 4098 30676 4132
rect 30710 4098 30768 4132
rect 30802 4098 30860 4132
rect 30894 4098 30952 4132
rect 30986 4098 31044 4132
rect 31078 4098 31136 4132
rect 31170 4098 31228 4132
rect 31262 4098 31320 4132
rect 31354 4098 31412 4132
rect 31446 4098 31504 4132
rect 31538 4098 31596 4132
rect 31630 4098 31688 4132
rect 31722 4098 31780 4132
rect 31814 4098 31872 4132
rect 31906 4098 31964 4132
rect 31998 4098 32062 4132
rect 30027 4095 30414 4098
rect 30466 4095 32062 4098
rect 30027 4067 32062 4095
rect 43381 3932 44853 3947
rect 45311 3932 46783 3947
rect 43381 3923 46783 3932
rect 43381 3922 44690 3923
rect 43381 3916 44600 3922
rect 30408 3862 30487 3890
rect 30408 3828 30423 3862
rect 30457 3834 30487 3862
rect 43381 3882 43410 3916
rect 43444 3882 43502 3916
rect 43536 3882 43594 3916
rect 43628 3882 43686 3916
rect 43720 3882 43778 3916
rect 43812 3882 43870 3916
rect 43904 3882 43962 3916
rect 43996 3882 44054 3916
rect 44088 3882 44146 3916
rect 44180 3882 44238 3916
rect 44272 3882 44330 3916
rect 44364 3882 44422 3916
rect 44456 3882 44514 3916
rect 44548 3882 44600 3916
rect 43381 3870 44600 3882
rect 44652 3871 44690 3922
rect 44742 3916 46783 3923
rect 44742 3882 44790 3916
rect 44824 3882 45340 3916
rect 45374 3882 45432 3916
rect 45466 3882 45524 3916
rect 45558 3882 45616 3916
rect 45650 3882 45708 3916
rect 45742 3882 45800 3916
rect 45834 3882 45892 3916
rect 45926 3882 45984 3916
rect 46018 3882 46076 3916
rect 46110 3882 46168 3916
rect 46202 3882 46260 3916
rect 46294 3882 46352 3916
rect 46386 3882 46444 3916
rect 46478 3882 46536 3916
rect 46570 3882 46628 3916
rect 46662 3882 46720 3916
rect 46754 3882 46783 3916
rect 44742 3874 46783 3882
rect 44742 3871 44853 3874
rect 44652 3870 44853 3871
rect 43381 3851 44853 3870
rect 45311 3851 46783 3874
rect 30457 3828 31406 3834
rect 30408 3826 31406 3828
rect 30408 3792 30606 3826
rect 30640 3792 30694 3826
rect 30728 3792 30782 3826
rect 30816 3792 30870 3826
rect 30904 3792 30958 3826
rect 30992 3792 31046 3826
rect 31080 3792 31134 3826
rect 31168 3792 31222 3826
rect 31256 3792 31310 3826
rect 31344 3792 31406 3826
rect 13239 3770 14711 3787
rect 13239 3756 14467 3770
rect 14519 3756 14590 3770
rect 13239 3722 13268 3756
rect 13302 3722 13360 3756
rect 13394 3722 13452 3756
rect 13486 3722 13544 3756
rect 13578 3722 13636 3756
rect 13670 3722 13728 3756
rect 13762 3722 13820 3756
rect 13854 3722 13912 3756
rect 13946 3722 14004 3756
rect 14038 3722 14096 3756
rect 14130 3722 14188 3756
rect 14222 3722 14280 3756
rect 14314 3722 14372 3756
rect 14406 3722 14464 3756
rect 14519 3722 14556 3756
rect 13239 3718 14467 3722
rect 14519 3718 14590 3722
rect 14642 3768 14711 3770
rect 15169 3768 16641 3787
rect 14642 3756 16641 3768
rect 14642 3722 14648 3756
rect 14682 3722 15198 3756
rect 15232 3722 15290 3756
rect 15324 3722 15382 3756
rect 15416 3722 15474 3756
rect 15508 3722 15566 3756
rect 15600 3722 15658 3756
rect 15692 3722 15750 3756
rect 15784 3722 15842 3756
rect 15876 3722 15934 3756
rect 15968 3722 16026 3756
rect 16060 3722 16118 3756
rect 16152 3722 16210 3756
rect 16244 3722 16302 3756
rect 16336 3722 16394 3756
rect 16428 3722 16486 3756
rect 16520 3722 16578 3756
rect 16612 3722 16641 3756
rect 30408 3786 31406 3792
rect 30408 3782 30490 3786
rect 30408 3748 30423 3782
rect 30457 3748 30490 3782
rect 30408 3730 30490 3748
rect 30979 3741 31924 3754
rect 14642 3718 16641 3722
rect 13239 3710 16641 3718
rect 13239 3691 14711 3710
rect 15169 3691 16641 3710
rect 30979 3724 31195 3741
rect 30979 3690 31029 3724
rect 31063 3690 31195 3724
rect 30979 3686 31195 3690
rect 31247 3689 31355 3741
rect 31407 3689 31488 3741
rect 31540 3724 31601 3741
rect 31564 3690 31601 3724
rect 31540 3689 31601 3690
rect 31653 3726 31924 3741
rect 31653 3725 31864 3726
rect 31653 3691 31700 3725
rect 31734 3692 31864 3725
rect 31898 3692 31924 3726
rect 31734 3691 31924 3692
rect 31653 3689 31924 3691
rect 31229 3686 31924 3689
rect 30979 3671 31924 3686
rect 37381 3723 52816 3733
rect 37381 3721 44018 3723
rect 37381 3714 43682 3721
rect 37381 3713 37563 3714
rect 37381 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3669 43514 3714
rect 43548 3676 43682 3714
rect 43716 3711 44018 3721
rect 43716 3676 43850 3711
rect 43548 3669 43850 3676
rect 37615 3666 43850 3669
rect 43884 3678 44018 3711
rect 44052 3721 44350 3723
rect 44052 3678 44184 3721
rect 43884 3676 44184 3678
rect 44218 3678 44350 3721
rect 44384 3678 44518 3723
rect 44552 3721 45780 3723
rect 44552 3678 44692 3721
rect 44218 3676 44692 3678
rect 44726 3719 45780 3721
rect 44726 3715 45610 3719
rect 44726 3676 45448 3715
rect 43884 3670 45448 3676
rect 45482 3674 45610 3715
rect 45644 3678 45780 3719
rect 45814 3719 52816 3723
rect 45814 3678 45944 3719
rect 45644 3674 45944 3678
rect 45978 3674 46114 3719
rect 46148 3715 46450 3719
rect 46148 3674 46282 3715
rect 45482 3670 46282 3674
rect 46316 3674 46450 3715
rect 46484 3715 52816 3719
rect 46484 3674 46624 3715
rect 46316 3670 46624 3674
rect 46658 3714 52816 3715
rect 46658 3709 52664 3714
rect 46658 3670 52573 3709
rect 43884 3666 52573 3670
rect 37615 3662 52573 3666
rect 37512 3661 52573 3662
rect 37381 3657 52573 3661
rect 52625 3662 52664 3709
rect 52716 3662 52816 3714
rect 52625 3657 52816 3662
rect 37381 3652 52816 3657
rect 30027 3600 32062 3619
rect 30027 3597 30577 3600
rect 30027 3595 30466 3597
rect 30027 3588 30370 3595
rect 7224 3563 22590 3573
rect 7224 3561 13876 3563
rect 7224 3558 13540 3561
rect 7224 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3554 13540 3558
rect 7413 3509 13372 3554
rect 13406 3516 13540 3554
rect 13574 3551 13876 3561
rect 13574 3516 13708 3551
rect 13406 3509 13708 3516
rect 7413 3506 13708 3509
rect 13742 3518 13876 3551
rect 13910 3561 14208 3563
rect 13910 3518 14042 3561
rect 13742 3516 14042 3518
rect 14076 3518 14208 3561
rect 14242 3518 14376 3563
rect 14410 3561 15638 3563
rect 14410 3518 14550 3561
rect 14076 3516 14550 3518
rect 14584 3559 15638 3561
rect 14584 3555 15468 3559
rect 14584 3516 15306 3555
rect 13742 3510 15306 3516
rect 15340 3514 15468 3555
rect 15502 3518 15638 3559
rect 15672 3559 22590 3563
rect 15672 3518 15802 3559
rect 15502 3514 15802 3518
rect 15836 3514 15972 3559
rect 16006 3555 16308 3559
rect 16006 3514 16140 3555
rect 15340 3510 16140 3514
rect 16174 3514 16308 3555
rect 16342 3556 22590 3559
rect 16342 3555 22475 3556
rect 16342 3514 16482 3555
rect 16174 3510 16482 3514
rect 16516 3549 22475 3555
rect 16516 3510 22376 3549
rect 13742 3506 22376 3510
rect 7224 3497 22376 3506
rect 22428 3504 22475 3549
rect 22527 3504 22590 3556
rect 30027 3554 30056 3588
rect 30090 3554 30148 3588
rect 30182 3554 30240 3588
rect 30274 3554 30332 3588
rect 30366 3554 30370 3588
rect 30027 3543 30370 3554
rect 30422 3588 30466 3595
rect 30422 3554 30424 3588
rect 30458 3554 30466 3588
rect 30422 3545 30466 3554
rect 30518 3548 30577 3597
rect 30629 3597 32062 3600
rect 30629 3548 30669 3597
rect 30721 3588 32062 3597
rect 30721 3554 30768 3588
rect 30802 3554 30860 3588
rect 30894 3554 30952 3588
rect 30986 3554 31044 3588
rect 31078 3554 31136 3588
rect 31170 3554 31228 3588
rect 31262 3554 31320 3588
rect 31354 3554 31412 3588
rect 31446 3554 31504 3588
rect 31538 3554 31596 3588
rect 31630 3554 31688 3588
rect 31722 3554 31780 3588
rect 31814 3554 31872 3588
rect 31906 3554 31964 3588
rect 31998 3554 32062 3588
rect 43682 3612 46285 3618
rect 43682 3578 43714 3612
rect 43748 3578 43814 3612
rect 43848 3578 43914 3612
rect 43948 3578 44014 3612
rect 44048 3578 44114 3612
rect 44148 3578 44214 3612
rect 44248 3578 44314 3612
rect 44348 3578 44414 3612
rect 44448 3578 45374 3612
rect 45408 3578 45474 3612
rect 45508 3578 45574 3612
rect 45608 3578 45674 3612
rect 45708 3578 45774 3612
rect 45808 3578 45874 3612
rect 45908 3578 45974 3612
rect 46008 3578 46074 3612
rect 46108 3578 46285 3612
rect 43682 3573 46285 3578
rect 43682 3570 45128 3573
rect 30518 3545 30669 3548
rect 30721 3545 32062 3554
rect 30422 3543 32062 3545
rect 30027 3523 32062 3543
rect 44978 3569 45128 3570
rect 22428 3497 22590 3504
rect 7224 3492 22590 3497
rect 44978 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3570 46285 3573
rect 45180 3521 45206 3570
rect 45075 3517 45206 3521
rect 44978 3478 45206 3517
rect 13540 3452 16143 3458
rect 13540 3418 13572 3452
rect 13606 3418 13672 3452
rect 13706 3418 13772 3452
rect 13806 3418 13872 3452
rect 13906 3418 13972 3452
rect 14006 3418 14072 3452
rect 14106 3418 14172 3452
rect 14206 3418 14272 3452
rect 14306 3418 15232 3452
rect 15266 3418 15332 3452
rect 15366 3418 15432 3452
rect 15466 3418 15532 3452
rect 15566 3418 15632 3452
rect 15666 3418 15732 3452
rect 15766 3418 15832 3452
rect 15866 3418 15932 3452
rect 15966 3418 16143 3452
rect 13540 3413 16143 3418
rect 13540 3410 14986 3413
rect 14836 3409 14986 3410
rect 14836 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3410 16143 3413
rect 15038 3361 15064 3410
rect 14933 3357 15064 3361
rect 14836 3318 15064 3357
rect 43381 3384 44853 3403
rect 45311 3384 46783 3403
rect 43381 3383 46783 3384
rect 43381 3382 46127 3383
rect 43381 3372 46035 3382
rect 46087 3372 46127 3382
rect 46179 3382 46783 3383
rect 46179 3372 46217 3382
rect 46269 3381 46783 3382
rect 46269 3372 46305 3381
rect 46357 3372 46783 3381
rect 43381 3338 43410 3372
rect 43444 3338 43502 3372
rect 43536 3338 43594 3372
rect 43628 3338 43686 3372
rect 43720 3338 43778 3372
rect 43812 3338 43870 3372
rect 43904 3338 43962 3372
rect 43996 3338 44054 3372
rect 44088 3338 44146 3372
rect 44180 3338 44238 3372
rect 44272 3338 44330 3372
rect 44364 3338 44422 3372
rect 44456 3338 44514 3372
rect 44548 3338 44606 3372
rect 44640 3338 44698 3372
rect 44732 3338 44790 3372
rect 44824 3338 45340 3372
rect 45374 3338 45432 3372
rect 45466 3338 45524 3372
rect 45558 3338 45616 3372
rect 45650 3338 45708 3372
rect 45742 3338 45800 3372
rect 45834 3338 45892 3372
rect 45926 3338 45984 3372
rect 46018 3338 46035 3372
rect 46110 3338 46127 3372
rect 46202 3338 46217 3372
rect 46294 3338 46305 3372
rect 46386 3338 46444 3372
rect 46478 3338 46536 3372
rect 46570 3338 46628 3372
rect 46662 3338 46720 3372
rect 46754 3338 46783 3372
rect 43381 3330 46035 3338
rect 46087 3331 46127 3338
rect 46179 3331 46217 3338
rect 46087 3330 46217 3331
rect 46269 3330 46305 3338
rect 43381 3329 46305 3330
rect 46357 3329 46783 3338
rect 43381 3326 46783 3329
rect 43381 3307 44853 3326
rect 45311 3307 46783 3326
rect 13202 3243 13253 3244
rect 13202 3230 14711 3243
rect 15169 3230 16641 3243
rect 13202 3222 16641 3230
rect 13202 3221 13857 3222
rect 13202 3212 13680 3221
rect 13732 3212 13764 3221
rect 13202 3178 13268 3212
rect 13302 3178 13360 3212
rect 13394 3178 13452 3212
rect 13486 3178 13544 3212
rect 13578 3178 13636 3212
rect 13670 3178 13680 3212
rect 13762 3178 13764 3212
rect 13202 3169 13680 3178
rect 13732 3169 13764 3178
rect 13816 3212 13857 3221
rect 13816 3178 13820 3212
rect 13854 3178 13857 3212
rect 13816 3170 13857 3178
rect 13909 3212 16641 3222
rect 13909 3178 13912 3212
rect 13946 3178 14004 3212
rect 14038 3178 14096 3212
rect 14130 3178 14188 3212
rect 14222 3178 14280 3212
rect 14314 3178 14372 3212
rect 14406 3178 14464 3212
rect 14498 3178 14556 3212
rect 14590 3178 14648 3212
rect 14682 3178 15198 3212
rect 15232 3178 15290 3212
rect 15324 3178 15382 3212
rect 15416 3178 15474 3212
rect 15508 3178 15566 3212
rect 15600 3178 15658 3212
rect 15692 3178 15750 3212
rect 15784 3178 15842 3212
rect 15876 3178 15934 3212
rect 15968 3178 16026 3212
rect 16060 3178 16118 3212
rect 16152 3178 16210 3212
rect 16244 3178 16302 3212
rect 16336 3178 16394 3212
rect 16428 3178 16486 3212
rect 16520 3178 16578 3212
rect 16612 3178 16641 3212
rect 13909 3172 16641 3178
rect 13909 3170 14711 3172
rect 13816 3169 14711 3170
rect 13202 3147 14711 3169
rect 15169 3147 16641 3172
rect 19721 3175 45232 3219
rect 19721 3173 45120 3175
rect 19721 3121 31184 3173
rect 31236 3121 31328 3173
rect 31380 3121 31472 3173
rect 31524 3172 45120 3173
rect 31524 3121 45031 3172
rect 19721 3120 45031 3121
rect 45083 3123 45120 3172
rect 45172 3123 45232 3175
rect 45083 3120 45232 3123
rect 19721 3096 45232 3120
rect 19721 3089 45031 3096
rect 19721 3037 31183 3089
rect 31235 3037 31327 3089
rect 31379 3037 31471 3089
rect 31523 3044 45031 3089
rect 45083 3044 45124 3096
rect 45176 3044 45232 3096
rect 31523 3037 45232 3044
rect 14848 3013 45232 3037
rect 14848 2992 19927 3013
rect 14848 2940 14885 2992
rect 14937 2987 19927 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 19927 2987
rect 14848 2914 19927 2935
rect 14848 2912 14979 2914
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 19927 2914
rect 14937 2860 19927 2862
rect 5664 2820 7136 2842
rect 7546 2820 9018 2840
rect 14848 2831 19927 2860
rect 20762 2832 22234 2842
rect 22644 2832 24116 2840
rect 5664 2817 9018 2820
rect 5664 2811 6266 2817
rect 6318 2811 6364 2817
rect 6416 2811 6459 2817
rect 6511 2811 6564 2817
rect 6616 2811 9018 2817
rect 5664 2777 5693 2811
rect 5727 2777 5785 2811
rect 5819 2777 5877 2811
rect 5911 2777 5969 2811
rect 6003 2777 6061 2811
rect 6095 2777 6153 2811
rect 6187 2777 6245 2811
rect 6318 2777 6337 2811
rect 6416 2777 6429 2811
rect 6511 2777 6521 2811
rect 6555 2777 6564 2811
rect 6647 2777 6705 2811
rect 6739 2777 6797 2811
rect 6831 2777 6889 2811
rect 6923 2777 6981 2811
rect 7015 2777 7073 2811
rect 7107 2809 9018 2811
rect 7107 2777 7575 2809
rect 5664 2765 6266 2777
rect 6318 2765 6364 2777
rect 6416 2765 6459 2777
rect 6511 2765 6564 2777
rect 6616 2775 7575 2777
rect 7609 2775 7667 2809
rect 7701 2775 7759 2809
rect 7793 2775 7851 2809
rect 7885 2775 7943 2809
rect 7977 2775 8035 2809
rect 8069 2775 8127 2809
rect 8161 2775 8219 2809
rect 8253 2775 8311 2809
rect 8345 2775 8403 2809
rect 8437 2775 8495 2809
rect 8529 2775 8587 2809
rect 8621 2775 8679 2809
rect 8713 2775 8771 2809
rect 8805 2775 8863 2809
rect 8897 2775 8955 2809
rect 8989 2775 9018 2809
rect 6616 2765 9018 2775
rect 5664 2762 9018 2765
rect 5664 2746 7136 2762
rect 7546 2744 9018 2762
rect 20762 2822 24116 2832
rect 20762 2811 21316 2822
rect 21368 2811 21416 2822
rect 21468 2811 21515 2822
rect 20762 2777 20791 2811
rect 20825 2777 20883 2811
rect 20917 2777 20975 2811
rect 21009 2777 21067 2811
rect 21101 2777 21159 2811
rect 21193 2777 21251 2811
rect 21285 2777 21316 2811
rect 21377 2777 21416 2811
rect 21469 2777 21515 2811
rect 20762 2770 21316 2777
rect 21368 2770 21416 2777
rect 21468 2770 21515 2777
rect 21567 2770 21618 2822
rect 21670 2811 24116 2822
rect 21670 2777 21711 2811
rect 21745 2777 21803 2811
rect 21837 2777 21895 2811
rect 21929 2777 21987 2811
rect 22021 2777 22079 2811
rect 22113 2777 22171 2811
rect 22205 2809 24116 2811
rect 22205 2777 22673 2809
rect 21670 2775 22673 2777
rect 22707 2775 22765 2809
rect 22799 2775 22857 2809
rect 22891 2775 22949 2809
rect 22983 2775 23041 2809
rect 23075 2775 23133 2809
rect 23167 2775 23225 2809
rect 23259 2775 23317 2809
rect 23351 2775 23409 2809
rect 23443 2775 23501 2809
rect 23535 2775 23593 2809
rect 23627 2775 23685 2809
rect 23719 2775 23777 2809
rect 23811 2775 23869 2809
rect 23903 2775 23961 2809
rect 23995 2775 24053 2809
rect 24087 2775 24116 2809
rect 21670 2774 24116 2775
rect 21670 2770 22234 2774
rect 20762 2746 22234 2770
rect 22644 2744 24116 2774
rect 35866 2832 37338 2842
rect 37748 2832 39220 2840
rect 35866 2816 39220 2832
rect 35866 2811 36424 2816
rect 36476 2811 36512 2816
rect 36564 2812 39220 2816
rect 36564 2811 36610 2812
rect 36662 2811 39220 2812
rect 35866 2777 35895 2811
rect 35929 2777 35987 2811
rect 36021 2777 36079 2811
rect 36113 2777 36171 2811
rect 36205 2777 36263 2811
rect 36297 2777 36355 2811
rect 36389 2777 36424 2811
rect 36481 2777 36512 2811
rect 36573 2777 36610 2811
rect 36665 2777 36723 2811
rect 36757 2777 36815 2811
rect 36849 2777 36907 2811
rect 36941 2777 36999 2811
rect 37033 2777 37091 2811
rect 37125 2777 37183 2811
rect 37217 2777 37275 2811
rect 37309 2809 39220 2811
rect 37309 2777 37777 2809
rect 35866 2764 36424 2777
rect 36476 2764 36512 2777
rect 36564 2764 36610 2777
rect 35866 2760 36610 2764
rect 36662 2775 37777 2777
rect 37811 2775 37869 2809
rect 37903 2775 37961 2809
rect 37995 2775 38053 2809
rect 38087 2775 38145 2809
rect 38179 2775 38237 2809
rect 38271 2775 38329 2809
rect 38363 2775 38421 2809
rect 38455 2775 38513 2809
rect 38547 2775 38605 2809
rect 38639 2775 38697 2809
rect 38731 2775 38789 2809
rect 38823 2775 38881 2809
rect 38915 2775 38973 2809
rect 39007 2775 39065 2809
rect 39099 2775 39157 2809
rect 39191 2775 39220 2809
rect 36662 2774 39220 2775
rect 36662 2760 37338 2774
rect 35866 2746 37338 2760
rect 37748 2744 39220 2774
rect 50964 2823 52436 2842
rect 52846 2823 54318 2840
rect 50964 2813 54318 2823
rect 50964 2811 53346 2813
rect 50964 2777 50993 2811
rect 51027 2777 51085 2811
rect 51119 2777 51177 2811
rect 51211 2777 51269 2811
rect 51303 2777 51361 2811
rect 51395 2777 51453 2811
rect 51487 2777 51545 2811
rect 51579 2777 51637 2811
rect 51671 2777 51729 2811
rect 51763 2777 51821 2811
rect 51855 2777 51913 2811
rect 51947 2777 52005 2811
rect 52039 2777 52097 2811
rect 52131 2777 52189 2811
rect 52223 2777 52281 2811
rect 52315 2777 52373 2811
rect 52407 2809 53346 2811
rect 53398 2809 53434 2813
rect 52407 2777 52875 2809
rect 50964 2775 52875 2777
rect 52909 2775 52967 2809
rect 53001 2775 53059 2809
rect 53093 2775 53151 2809
rect 53185 2775 53243 2809
rect 53277 2775 53335 2809
rect 53398 2775 53427 2809
rect 50964 2765 53346 2775
rect 50964 2746 52436 2765
rect 52846 2761 53346 2765
rect 53398 2761 53434 2775
rect 53486 2761 53517 2813
rect 53569 2761 53604 2813
rect 53656 2809 54318 2813
rect 53656 2775 53703 2809
rect 53737 2775 53795 2809
rect 53829 2775 53887 2809
rect 53921 2775 53979 2809
rect 54013 2775 54071 2809
rect 54105 2775 54163 2809
rect 54197 2775 54255 2809
rect 54289 2775 54318 2809
rect 53656 2761 54318 2775
rect 52846 2744 54318 2761
rect 7240 2675 7446 2692
rect 7240 2623 7265 2675
rect 7317 2673 7446 2675
rect 7317 2623 7345 2673
rect 7240 2621 7345 2623
rect 7397 2621 7446 2673
rect 7240 2580 7446 2621
rect 22352 2690 22550 2694
rect 22352 2638 22381 2690
rect 22433 2638 22464 2690
rect 22516 2638 22550 2690
rect 22352 2580 22550 2638
rect 37442 2680 37648 2692
rect 37442 2628 37459 2680
rect 37511 2628 37550 2680
rect 37602 2628 37648 2680
rect 52554 2669 52752 2694
rect 37442 2580 37648 2628
rect 52547 2665 52752 2669
rect 52547 2613 52576 2665
rect 52628 2613 52659 2665
rect 52711 2613 52752 2665
rect 52547 2580 52752 2613
rect 5770 2574 8574 2580
rect 5770 2540 5820 2574
rect 5854 2540 5933 2574
rect 5967 2540 6046 2574
rect 6080 2540 6159 2574
rect 6193 2540 6272 2574
rect 6306 2540 6385 2574
rect 6419 2540 6498 2574
rect 6532 2540 6614 2574
rect 6648 2540 6718 2574
rect 6752 2540 7574 2574
rect 7608 2540 7693 2574
rect 7727 2540 7812 2574
rect 7846 2540 7931 2574
rect 7965 2540 8050 2574
rect 8084 2540 8169 2574
rect 8203 2540 8288 2574
rect 8322 2540 8574 2574
rect 5770 2534 8574 2540
rect 20921 2574 23612 2580
rect 20921 2540 20986 2574
rect 21020 2540 21083 2574
rect 21117 2540 21180 2574
rect 21214 2540 21277 2574
rect 21311 2540 21374 2574
rect 21408 2540 21471 2574
rect 21505 2540 21568 2574
rect 21602 2540 21665 2574
rect 21699 2540 21816 2574
rect 21850 2540 22672 2574
rect 22706 2540 22780 2574
rect 22814 2540 22888 2574
rect 22922 2540 22996 2574
rect 23030 2540 23104 2574
rect 23138 2540 23212 2574
rect 23246 2540 23320 2574
rect 23354 2540 23428 2574
rect 23462 2540 23612 2574
rect 20921 2534 23612 2540
rect 35972 2574 38776 2580
rect 35972 2540 36022 2574
rect 36056 2540 36135 2574
rect 36169 2540 36248 2574
rect 36282 2540 36361 2574
rect 36395 2540 36474 2574
rect 36508 2540 36587 2574
rect 36621 2540 36700 2574
rect 36734 2540 36816 2574
rect 36850 2540 36920 2574
rect 36954 2540 37776 2574
rect 37810 2540 37895 2574
rect 37929 2540 38014 2574
rect 38048 2540 38133 2574
rect 38167 2540 38252 2574
rect 38286 2540 38371 2574
rect 38405 2540 38490 2574
rect 38524 2540 38776 2574
rect 35972 2534 38776 2540
rect 51123 2574 53814 2580
rect 51123 2540 51188 2574
rect 51222 2540 51285 2574
rect 51319 2540 51382 2574
rect 51416 2540 51479 2574
rect 51513 2540 51576 2574
rect 51610 2540 51673 2574
rect 51707 2540 51770 2574
rect 51804 2540 51867 2574
rect 51901 2540 52018 2574
rect 52052 2540 52874 2574
rect 52908 2540 52982 2574
rect 53016 2540 53090 2574
rect 53124 2540 53198 2574
rect 53232 2540 53306 2574
rect 53340 2540 53414 2574
rect 53448 2540 53522 2574
rect 53556 2540 53630 2574
rect 53664 2540 53814 2574
rect 51123 2534 53814 2540
rect 5782 2480 7019 2492
rect 5782 2479 6972 2480
rect 5782 2445 5797 2479
rect 5831 2478 6972 2479
rect 5831 2477 6802 2478
rect 5831 2474 5963 2477
rect 5997 2476 6298 2477
rect 6332 2476 6802 2477
rect 5997 2475 6292 2476
rect 5997 2474 6127 2475
rect 5831 2445 5834 2474
rect 5782 2422 5834 2445
rect 5886 2422 5941 2474
rect 5997 2443 6047 2474
rect 5993 2422 6047 2443
rect 6099 2441 6127 2474
rect 6161 2474 6292 2475
rect 6161 2441 6163 2474
rect 6099 2422 6163 2441
rect 6215 2424 6292 2474
rect 6344 2475 6802 2476
rect 6836 2475 6972 2478
rect 6344 2424 6426 2475
rect 6478 2473 6543 2475
rect 6501 2439 6543 2473
rect 6215 2423 6426 2424
rect 6478 2423 6543 2439
rect 6595 2472 6648 2475
rect 6595 2438 6636 2472
rect 6595 2423 6648 2438
rect 6700 2423 6754 2475
rect 6836 2444 6851 2475
rect 6806 2423 6851 2444
rect 6903 2423 6948 2475
rect 7006 2446 7019 2480
rect 7000 2423 7019 2446
rect 6215 2422 7019 2423
rect 5782 2408 7019 2422
rect 7672 2481 8898 2490
rect 7672 2477 8182 2481
rect 7672 2443 7686 2477
rect 7720 2471 7846 2477
rect 7880 2474 8182 2477
rect 8216 2478 8898 2481
rect 8216 2476 8845 2478
rect 8216 2474 8686 2476
rect 7880 2471 8174 2474
rect 7720 2443 7723 2471
rect 7672 2419 7723 2443
rect 7775 2419 7830 2471
rect 7882 2419 7936 2471
rect 7988 2437 8013 2471
rect 8047 2437 8052 2471
rect 7988 2419 8052 2437
rect 8104 2422 8174 2471
rect 8226 2473 8516 2474
rect 8233 2472 8516 2473
rect 8550 2472 8686 2474
rect 8720 2472 8845 2476
rect 8879 2472 8898 2478
rect 8104 2421 8181 2422
rect 8233 2421 8315 2472
rect 8367 2468 8432 2472
rect 8380 2434 8432 2468
rect 8104 2420 8315 2421
rect 8367 2420 8432 2434
rect 8484 2440 8516 2472
rect 8484 2420 8537 2440
rect 8589 2420 8643 2472
rect 8720 2442 8740 2472
rect 8695 2420 8740 2442
rect 8792 2420 8837 2472
rect 8889 2420 8898 2472
rect 8104 2419 8898 2420
rect 7672 2406 8898 2419
rect 20873 2480 22140 2492
rect 20873 2473 20943 2480
rect 20873 2439 20895 2473
rect 20929 2439 20943 2473
rect 20873 2428 20943 2439
rect 20995 2478 22140 2480
rect 20995 2428 21055 2478
rect 20873 2426 21055 2428
rect 21107 2426 21162 2478
rect 21214 2472 21264 2478
rect 21316 2477 22140 2478
rect 21316 2476 21396 2477
rect 21430 2476 22140 2477
rect 21214 2438 21231 2472
rect 21214 2426 21264 2438
rect 21316 2426 21390 2476
rect 20873 2424 21390 2426
rect 21442 2424 21544 2476
rect 21596 2464 21681 2476
rect 21597 2430 21681 2464
rect 21733 2462 21778 2476
rect 21596 2424 21681 2430
rect 21765 2428 21778 2462
rect 21733 2424 21778 2428
rect 21830 2424 21878 2476
rect 21930 2475 22140 2476
rect 21930 2471 21967 2475
rect 21935 2437 21967 2471
rect 21930 2424 21967 2437
rect 20873 2423 21967 2424
rect 22019 2423 22063 2475
rect 22115 2423 22140 2475
rect 20873 2408 22140 2423
rect 22759 2481 24015 2490
rect 22759 2478 23280 2481
rect 22759 2474 23109 2478
rect 23143 2474 23280 2478
rect 23314 2474 24015 2481
rect 22759 2472 22777 2474
rect 22759 2438 22774 2472
rect 22759 2422 22777 2438
rect 22829 2422 22871 2474
rect 22923 2473 22970 2474
rect 22923 2439 22947 2473
rect 22923 2422 22970 2439
rect 23022 2422 23078 2474
rect 23143 2444 23174 2474
rect 23130 2422 23174 2444
rect 23226 2422 23272 2474
rect 23324 2473 24015 2474
rect 23324 2422 23391 2473
rect 22759 2421 23391 2422
rect 23443 2467 23505 2473
rect 23443 2433 23449 2467
rect 23483 2433 23505 2467
rect 23443 2421 23505 2433
rect 23557 2467 23622 2473
rect 23557 2433 23614 2467
rect 23557 2421 23622 2433
rect 23674 2421 23749 2473
rect 23801 2465 23864 2473
rect 23818 2431 23864 2465
rect 23801 2421 23864 2431
rect 23916 2469 24015 2473
rect 23916 2435 23947 2469
rect 23981 2435 24015 2469
rect 23916 2421 24015 2435
rect 22759 2406 24015 2421
rect 35984 2480 37221 2492
rect 35984 2479 37174 2480
rect 35984 2445 35999 2479
rect 36033 2478 37174 2479
rect 36033 2477 37004 2478
rect 36033 2474 36165 2477
rect 36199 2476 36500 2477
rect 36534 2476 37004 2477
rect 36199 2475 36494 2476
rect 36199 2474 36329 2475
rect 36033 2445 36036 2474
rect 35984 2422 36036 2445
rect 36088 2422 36143 2474
rect 36199 2443 36249 2474
rect 36195 2422 36249 2443
rect 36301 2441 36329 2474
rect 36363 2474 36494 2475
rect 36363 2441 36365 2474
rect 36301 2422 36365 2441
rect 36417 2424 36494 2474
rect 36546 2475 37004 2476
rect 37038 2475 37174 2478
rect 36546 2424 36628 2475
rect 36680 2473 36745 2475
rect 36703 2439 36745 2473
rect 36417 2423 36628 2424
rect 36680 2423 36745 2439
rect 36797 2472 36850 2475
rect 36797 2438 36838 2472
rect 36797 2423 36850 2438
rect 36902 2423 36956 2475
rect 37038 2444 37053 2475
rect 37008 2423 37053 2444
rect 37105 2423 37150 2475
rect 37208 2446 37221 2480
rect 37202 2423 37221 2446
rect 36417 2422 37221 2423
rect 35984 2408 37221 2422
rect 37874 2481 39100 2490
rect 37874 2477 38384 2481
rect 37874 2443 37888 2477
rect 37922 2471 38048 2477
rect 38082 2474 38384 2477
rect 38418 2478 39100 2481
rect 38418 2476 39047 2478
rect 38418 2474 38888 2476
rect 38082 2471 38376 2474
rect 37922 2443 37925 2471
rect 37874 2419 37925 2443
rect 37977 2419 38032 2471
rect 38084 2419 38138 2471
rect 38190 2437 38215 2471
rect 38249 2437 38254 2471
rect 38190 2419 38254 2437
rect 38306 2422 38376 2471
rect 38428 2473 38718 2474
rect 38435 2472 38718 2473
rect 38752 2472 38888 2474
rect 38922 2472 39047 2476
rect 39081 2472 39100 2478
rect 38306 2421 38383 2422
rect 38435 2421 38517 2472
rect 38569 2468 38634 2472
rect 38582 2434 38634 2468
rect 38306 2420 38517 2421
rect 38569 2420 38634 2434
rect 38686 2440 38718 2472
rect 38686 2420 38739 2440
rect 38791 2420 38845 2472
rect 38922 2442 38942 2472
rect 38897 2420 38942 2442
rect 38994 2420 39039 2472
rect 39091 2420 39100 2472
rect 38306 2419 39100 2420
rect 37874 2406 39100 2419
rect 51075 2480 52342 2492
rect 51075 2473 51145 2480
rect 51075 2439 51097 2473
rect 51131 2439 51145 2473
rect 51075 2428 51145 2439
rect 51197 2478 52342 2480
rect 51197 2428 51257 2478
rect 51075 2426 51257 2428
rect 51309 2426 51364 2478
rect 51416 2472 51466 2478
rect 51518 2477 52342 2478
rect 51518 2476 51598 2477
rect 51632 2476 52342 2477
rect 51416 2438 51433 2472
rect 51416 2426 51466 2438
rect 51518 2426 51592 2476
rect 51075 2424 51592 2426
rect 51644 2424 51746 2476
rect 51798 2464 51883 2476
rect 51799 2430 51883 2464
rect 51935 2462 51980 2476
rect 51798 2424 51883 2430
rect 51967 2428 51980 2462
rect 51935 2424 51980 2428
rect 52032 2424 52080 2476
rect 52132 2475 52342 2476
rect 52132 2471 52169 2475
rect 52137 2437 52169 2471
rect 52132 2424 52169 2437
rect 51075 2423 52169 2424
rect 52221 2423 52265 2475
rect 52317 2423 52342 2475
rect 51075 2408 52342 2423
rect 52961 2481 54217 2490
rect 52961 2478 53482 2481
rect 52961 2474 53311 2478
rect 53345 2474 53482 2478
rect 53516 2474 54217 2481
rect 52961 2472 52979 2474
rect 52961 2438 52976 2472
rect 52961 2422 52979 2438
rect 53031 2422 53073 2474
rect 53125 2473 53172 2474
rect 53125 2439 53149 2473
rect 53125 2422 53172 2439
rect 53224 2422 53280 2474
rect 53345 2444 53376 2474
rect 53332 2422 53376 2444
rect 53428 2422 53474 2474
rect 53526 2473 54217 2474
rect 53526 2422 53593 2473
rect 52961 2421 53593 2422
rect 53645 2467 53707 2473
rect 53645 2433 53651 2467
rect 53685 2433 53707 2467
rect 53645 2421 53707 2433
rect 53759 2467 53824 2473
rect 53759 2433 53816 2467
rect 53759 2421 53824 2433
rect 53876 2421 53951 2473
rect 54003 2465 54066 2473
rect 54020 2431 54066 2465
rect 54003 2421 54066 2431
rect 54118 2469 54217 2473
rect 54118 2435 54149 2469
rect 54183 2435 54217 2469
rect 54118 2421 54217 2435
rect 52961 2406 54217 2421
rect 0 2304 60412 2376
rect 0 2188 1535 2304
rect 1843 2188 3423 2304
rect 3731 2188 5311 2304
rect 5619 2267 7199 2304
rect 5619 2233 5693 2267
rect 5727 2233 5785 2267
rect 5819 2233 5877 2267
rect 5911 2233 5969 2267
rect 6003 2233 6061 2267
rect 6095 2233 6153 2267
rect 6187 2233 6245 2267
rect 6279 2233 6337 2267
rect 6371 2233 6429 2267
rect 6463 2233 6521 2267
rect 6555 2233 6613 2267
rect 6647 2233 6705 2267
rect 6739 2233 6797 2267
rect 6831 2233 6889 2267
rect 6923 2233 6981 2267
rect 7015 2233 7073 2267
rect 7107 2233 7199 2267
rect 5619 2188 7199 2233
rect 7507 2265 9087 2304
rect 7507 2231 7575 2265
rect 7609 2231 7667 2265
rect 7701 2231 7759 2265
rect 7793 2231 7851 2265
rect 7885 2231 7943 2265
rect 7977 2231 8035 2265
rect 8069 2231 8127 2265
rect 8161 2231 8219 2265
rect 8253 2231 8311 2265
rect 8345 2231 8403 2265
rect 8437 2231 8495 2265
rect 8529 2231 8587 2265
rect 8621 2231 8679 2265
rect 8713 2231 8771 2265
rect 8805 2231 8863 2265
rect 8897 2231 8955 2265
rect 8989 2231 9087 2265
rect 7507 2188 9087 2231
rect 9395 2188 10975 2304
rect 11283 2188 12863 2304
rect 13171 2188 14751 2304
rect 15059 2188 16633 2304
rect 16941 2188 18521 2304
rect 18829 2188 20409 2304
rect 20717 2267 22297 2304
rect 20717 2233 20791 2267
rect 20825 2233 20883 2267
rect 20917 2233 20975 2267
rect 21009 2233 21067 2267
rect 21101 2233 21159 2267
rect 21193 2233 21251 2267
rect 21285 2233 21343 2267
rect 21377 2233 21435 2267
rect 21469 2233 21527 2267
rect 21561 2233 21619 2267
rect 21653 2233 21711 2267
rect 21745 2233 21803 2267
rect 21837 2233 21895 2267
rect 21929 2233 21987 2267
rect 22021 2233 22079 2267
rect 22113 2233 22171 2267
rect 22205 2233 22297 2267
rect 20717 2188 22297 2233
rect 22605 2265 24185 2304
rect 22605 2231 22673 2265
rect 22707 2231 22765 2265
rect 22799 2231 22857 2265
rect 22891 2231 22949 2265
rect 22983 2231 23041 2265
rect 23075 2231 23133 2265
rect 23167 2231 23225 2265
rect 23259 2231 23317 2265
rect 23351 2231 23409 2265
rect 23443 2231 23501 2265
rect 23535 2231 23593 2265
rect 23627 2231 23685 2265
rect 23719 2231 23777 2265
rect 23811 2231 23869 2265
rect 23903 2231 23961 2265
rect 23995 2231 24053 2265
rect 24087 2231 24185 2265
rect 22605 2188 24185 2231
rect 24493 2188 26073 2304
rect 26381 2188 27961 2304
rect 28269 2188 29849 2304
rect 30157 2188 31737 2304
rect 32045 2188 33625 2304
rect 33933 2188 35513 2304
rect 35821 2267 37401 2304
rect 35821 2233 35895 2267
rect 35929 2233 35987 2267
rect 36021 2233 36079 2267
rect 36113 2233 36171 2267
rect 36205 2233 36263 2267
rect 36297 2233 36355 2267
rect 36389 2233 36447 2267
rect 36481 2233 36539 2267
rect 36573 2233 36631 2267
rect 36665 2233 36723 2267
rect 36757 2233 36815 2267
rect 36849 2233 36907 2267
rect 36941 2233 36999 2267
rect 37033 2233 37091 2267
rect 37125 2233 37183 2267
rect 37217 2233 37275 2267
rect 37309 2233 37401 2267
rect 35821 2188 37401 2233
rect 37709 2265 39289 2304
rect 37709 2231 37777 2265
rect 37811 2231 37869 2265
rect 37903 2231 37961 2265
rect 37995 2231 38053 2265
rect 38087 2231 38145 2265
rect 38179 2231 38237 2265
rect 38271 2231 38329 2265
rect 38363 2231 38421 2265
rect 38455 2231 38513 2265
rect 38547 2231 38605 2265
rect 38639 2231 38697 2265
rect 38731 2231 38789 2265
rect 38823 2231 38881 2265
rect 38915 2231 38973 2265
rect 39007 2231 39065 2265
rect 39099 2231 39157 2265
rect 39191 2231 39289 2265
rect 37709 2188 39289 2231
rect 39597 2188 41177 2304
rect 41485 2188 43065 2304
rect 43373 2188 44953 2304
rect 45261 2188 46835 2304
rect 47143 2188 48723 2304
rect 49031 2188 50611 2304
rect 50919 2267 52499 2304
rect 50919 2233 50993 2267
rect 51027 2233 51085 2267
rect 51119 2233 51177 2267
rect 51211 2233 51269 2267
rect 51303 2233 51361 2267
rect 51395 2233 51453 2267
rect 51487 2233 51545 2267
rect 51579 2233 51637 2267
rect 51671 2233 51729 2267
rect 51763 2233 51821 2267
rect 51855 2233 51913 2267
rect 51947 2233 52005 2267
rect 52039 2233 52097 2267
rect 52131 2233 52189 2267
rect 52223 2233 52281 2267
rect 52315 2233 52373 2267
rect 52407 2233 52499 2267
rect 50919 2188 52499 2233
rect 52807 2265 54387 2304
rect 52807 2231 52875 2265
rect 52909 2231 52967 2265
rect 53001 2231 53059 2265
rect 53093 2231 53151 2265
rect 53185 2231 53243 2265
rect 53277 2231 53335 2265
rect 53369 2231 53427 2265
rect 53461 2231 53519 2265
rect 53553 2231 53611 2265
rect 53645 2231 53703 2265
rect 53737 2231 53795 2265
rect 53829 2231 53887 2265
rect 53921 2231 53979 2265
rect 54013 2231 54071 2265
rect 54105 2231 54163 2265
rect 54197 2231 54255 2265
rect 54289 2231 54387 2265
rect 52807 2188 54387 2231
rect 54695 2188 56275 2304
rect 56583 2188 58163 2304
rect 58471 2188 60051 2304
rect 60359 2188 60412 2304
rect 0 2187 60412 2188
rect 0 2153 247 2187
rect 281 2153 339 2187
rect 373 2153 431 2187
rect 465 2153 1061 2187
rect 1095 2153 1153 2187
rect 1187 2153 1245 2187
rect 1279 2153 2135 2187
rect 2169 2153 2227 2187
rect 2261 2153 2319 2187
rect 2353 2153 2949 2187
rect 2983 2153 3041 2187
rect 3075 2153 3133 2187
rect 3167 2153 4023 2187
rect 4057 2153 4115 2187
rect 4149 2153 4207 2187
rect 4241 2153 4837 2187
rect 4871 2153 4929 2187
rect 4963 2153 5021 2187
rect 5055 2153 5911 2187
rect 5945 2153 6003 2187
rect 6037 2153 6095 2187
rect 6129 2153 6725 2187
rect 6759 2153 6817 2187
rect 6851 2153 6909 2187
rect 6943 2153 7799 2187
rect 7833 2153 7891 2187
rect 7925 2153 7983 2187
rect 8017 2153 8613 2187
rect 8647 2153 8705 2187
rect 8739 2153 8797 2187
rect 8831 2153 9687 2187
rect 9721 2153 9779 2187
rect 9813 2153 9871 2187
rect 9905 2153 10501 2187
rect 10535 2153 10593 2187
rect 10627 2153 10685 2187
rect 10719 2153 11575 2187
rect 11609 2153 11667 2187
rect 11701 2153 11759 2187
rect 11793 2153 12389 2187
rect 12423 2153 12481 2187
rect 12515 2153 12573 2187
rect 12607 2153 13463 2187
rect 13497 2153 13555 2187
rect 13589 2153 13647 2187
rect 13681 2153 14277 2187
rect 14311 2153 14369 2187
rect 14403 2153 14461 2187
rect 14495 2153 15345 2187
rect 15379 2153 15437 2187
rect 15471 2153 15529 2187
rect 15563 2153 16159 2187
rect 16193 2153 16251 2187
rect 16285 2153 16343 2187
rect 16377 2153 17233 2187
rect 17267 2153 17325 2187
rect 17359 2153 17417 2187
rect 17451 2153 18047 2187
rect 18081 2153 18139 2187
rect 18173 2153 18231 2187
rect 18265 2153 19121 2187
rect 19155 2153 19213 2187
rect 19247 2153 19305 2187
rect 19339 2153 19935 2187
rect 19969 2153 20027 2187
rect 20061 2153 20119 2187
rect 20153 2153 21009 2187
rect 21043 2153 21101 2187
rect 21135 2153 21193 2187
rect 21227 2153 21823 2187
rect 21857 2153 21915 2187
rect 21949 2153 22007 2187
rect 22041 2153 22897 2187
rect 22931 2153 22989 2187
rect 23023 2153 23081 2187
rect 23115 2153 23711 2187
rect 23745 2153 23803 2187
rect 23837 2153 23895 2187
rect 23929 2153 24785 2187
rect 24819 2153 24877 2187
rect 24911 2153 24969 2187
rect 25003 2153 25599 2187
rect 25633 2153 25691 2187
rect 25725 2153 25783 2187
rect 25817 2153 26673 2187
rect 26707 2153 26765 2187
rect 26799 2153 26857 2187
rect 26891 2153 27487 2187
rect 27521 2153 27579 2187
rect 27613 2153 27671 2187
rect 27705 2153 28561 2187
rect 28595 2153 28653 2187
rect 28687 2153 28745 2187
rect 28779 2153 29375 2187
rect 29409 2153 29467 2187
rect 29501 2153 29559 2187
rect 29593 2153 30449 2187
rect 30483 2153 30541 2187
rect 30575 2153 30633 2187
rect 30667 2153 31263 2187
rect 31297 2153 31355 2187
rect 31389 2153 31447 2187
rect 31481 2153 32337 2187
rect 32371 2153 32429 2187
rect 32463 2153 32521 2187
rect 32555 2153 33151 2187
rect 33185 2153 33243 2187
rect 33277 2153 33335 2187
rect 33369 2153 34225 2187
rect 34259 2153 34317 2187
rect 34351 2153 34409 2187
rect 34443 2153 35039 2187
rect 35073 2153 35131 2187
rect 35165 2153 35223 2187
rect 35257 2153 36113 2187
rect 36147 2153 36205 2187
rect 36239 2153 36297 2187
rect 36331 2153 36927 2187
rect 36961 2153 37019 2187
rect 37053 2153 37111 2187
rect 37145 2153 38001 2187
rect 38035 2153 38093 2187
rect 38127 2153 38185 2187
rect 38219 2153 38815 2187
rect 38849 2153 38907 2187
rect 38941 2153 38999 2187
rect 39033 2153 39889 2187
rect 39923 2153 39981 2187
rect 40015 2153 40073 2187
rect 40107 2153 40703 2187
rect 40737 2153 40795 2187
rect 40829 2153 40887 2187
rect 40921 2153 41777 2187
rect 41811 2153 41869 2187
rect 41903 2153 41961 2187
rect 41995 2153 42591 2187
rect 42625 2153 42683 2187
rect 42717 2153 42775 2187
rect 42809 2153 43665 2187
rect 43699 2153 43757 2187
rect 43791 2153 43849 2187
rect 43883 2153 44479 2187
rect 44513 2153 44571 2187
rect 44605 2153 44663 2187
rect 44697 2153 45547 2187
rect 45581 2153 45639 2187
rect 45673 2153 45731 2187
rect 45765 2153 46361 2187
rect 46395 2153 46453 2187
rect 46487 2153 46545 2187
rect 46579 2153 47435 2187
rect 47469 2153 47527 2187
rect 47561 2153 47619 2187
rect 47653 2153 48249 2187
rect 48283 2153 48341 2187
rect 48375 2153 48433 2187
rect 48467 2153 49323 2187
rect 49357 2153 49415 2187
rect 49449 2153 49507 2187
rect 49541 2153 50137 2187
rect 50171 2153 50229 2187
rect 50263 2153 50321 2187
rect 50355 2153 51211 2187
rect 51245 2153 51303 2187
rect 51337 2153 51395 2187
rect 51429 2153 52025 2187
rect 52059 2153 52117 2187
rect 52151 2153 52209 2187
rect 52243 2153 53099 2187
rect 53133 2153 53191 2187
rect 53225 2153 53283 2187
rect 53317 2153 53913 2187
rect 53947 2153 54005 2187
rect 54039 2153 54097 2187
rect 54131 2153 54987 2187
rect 55021 2153 55079 2187
rect 55113 2153 55171 2187
rect 55205 2153 55801 2187
rect 55835 2153 55893 2187
rect 55927 2153 55985 2187
rect 56019 2153 56875 2187
rect 56909 2153 56967 2187
rect 57001 2153 57059 2187
rect 57093 2153 57689 2187
rect 57723 2153 57781 2187
rect 57815 2153 57873 2187
rect 57907 2153 58763 2187
rect 58797 2153 58855 2187
rect 58889 2153 58947 2187
rect 58981 2153 59577 2187
rect 59611 2153 59669 2187
rect 59703 2153 59761 2187
rect 59795 2153 60412 2187
rect 0 2147 60412 2153
rect 0 2122 681 2147
rect 60 1164 138 2122
rect 652 2113 681 2122
rect 715 2122 2569 2147
rect 715 2113 742 2122
rect 652 2092 742 2113
rect 738 2056 796 2058
rect 738 2039 800 2056
rect 738 2005 750 2039
rect 784 2005 800 2039
rect 738 1996 800 2005
rect 238 1958 604 1962
rect 686 1958 752 1966
rect 238 1930 646 1958
rect 238 1892 266 1930
rect 560 1911 646 1930
rect 238 1884 304 1892
rect 238 1850 253 1884
rect 287 1850 304 1884
rect 238 1838 304 1850
rect 410 1888 478 1894
rect 410 1836 420 1888
rect 472 1836 478 1888
rect 410 1830 478 1836
rect 560 1877 606 1911
rect 640 1877 646 1911
rect 686 1906 692 1958
rect 744 1906 752 1958
rect 686 1898 702 1906
rect 560 1839 646 1877
rect 560 1805 606 1839
rect 640 1805 646 1839
rect 320 1776 388 1782
rect 320 1724 328 1776
rect 380 1724 388 1776
rect 320 1714 388 1724
rect 560 1758 646 1805
rect 696 1877 702 1898
rect 736 1898 752 1906
rect 792 1926 1120 1958
rect 792 1911 888 1926
rect 736 1877 742 1898
rect 696 1839 742 1877
rect 696 1805 702 1839
rect 736 1805 742 1839
rect 696 1758 742 1805
rect 792 1877 798 1911
rect 832 1877 888 1911
rect 1092 1890 1120 1926
rect 792 1839 888 1877
rect 792 1805 798 1839
rect 832 1805 888 1839
rect 1050 1882 1120 1890
rect 1050 1848 1065 1882
rect 1099 1848 1120 1882
rect 1050 1830 1120 1848
rect 1226 1890 1290 1896
rect 1226 1838 1232 1890
rect 1284 1838 1290 1890
rect 1226 1832 1290 1838
rect 792 1758 888 1805
rect 218 1643 494 1674
rect 218 1609 247 1643
rect 281 1609 339 1643
rect 373 1609 431 1643
rect 465 1609 494 1643
rect 218 1578 494 1609
rect 560 1558 610 1758
rect 642 1711 700 1726
rect 642 1677 654 1711
rect 688 1677 700 1711
rect 642 1660 700 1677
rect 754 1630 812 1648
rect 754 1596 766 1630
rect 800 1596 812 1630
rect 754 1586 812 1596
rect 842 1558 888 1758
rect 1138 1774 1202 1780
rect 1138 1722 1144 1774
rect 1196 1722 1202 1774
rect 1138 1716 1202 1722
rect 1032 1643 1308 1674
rect 1032 1609 1061 1643
rect 1095 1609 1153 1643
rect 1187 1609 1245 1643
rect 1279 1609 1308 1643
rect 1032 1606 1308 1609
rect 200 1541 264 1548
rect 200 1508 206 1541
rect 258 1508 264 1541
rect 376 1541 440 1548
rect 376 1508 382 1541
rect 258 1489 382 1508
rect 434 1489 440 1541
rect 206 1480 440 1489
rect 560 1546 662 1558
rect 560 1512 622 1546
rect 656 1512 662 1546
rect 560 1474 662 1512
rect 712 1546 758 1558
rect 712 1512 718 1546
rect 752 1512 758 1546
rect 712 1492 758 1512
rect 808 1546 888 1558
rect 808 1512 814 1546
rect 848 1512 888 1546
rect 560 1442 622 1474
rect 356 1440 622 1442
rect 656 1440 662 1474
rect 356 1428 662 1440
rect 702 1486 768 1492
rect 702 1434 710 1486
rect 762 1434 768 1486
rect 702 1428 768 1434
rect 808 1474 888 1512
rect 808 1440 814 1474
rect 848 1440 888 1474
rect 1004 1578 1308 1606
rect 808 1428 854 1440
rect 356 1414 610 1428
rect 200 1408 266 1414
rect 200 1356 208 1408
rect 260 1356 266 1408
rect 200 1350 266 1356
rect 40 1150 316 1164
rect 40 1133 232 1150
rect 284 1133 316 1150
rect 40 1099 69 1133
rect 103 1099 161 1133
rect 195 1099 232 1133
rect 287 1099 316 1133
rect 40 1098 232 1099
rect 284 1098 316 1099
rect 40 1068 316 1098
rect 356 1064 384 1414
rect 656 1390 720 1400
rect 656 1356 670 1390
rect 704 1356 976 1390
rect 656 1338 720 1356
rect 572 1292 644 1304
rect 572 1240 582 1292
rect 634 1240 644 1292
rect 572 1228 644 1240
rect 942 1174 976 1356
rect 1004 1274 1032 1578
rect 1004 1264 1072 1274
rect 1004 1230 1020 1264
rect 1054 1230 1072 1264
rect 1004 1216 1072 1230
rect 416 1146 976 1174
rect 416 1143 482 1146
rect 416 1109 432 1143
rect 466 1109 482 1143
rect 416 1100 482 1109
rect 650 1091 740 1112
rect 356 1036 428 1064
rect 382 1015 428 1036
rect 382 981 388 1015
rect 422 981 428 1015
rect 382 943 428 981
rect 382 909 388 943
rect 422 909 428 943
rect 382 862 428 909
rect 470 1042 516 1062
rect 650 1057 679 1091
rect 713 1057 740 1091
rect 470 1036 538 1042
rect 650 1036 740 1057
rect 470 1015 478 1036
rect 470 981 476 1015
rect 530 984 538 1036
rect 510 981 538 984
rect 470 976 538 981
rect 736 1000 794 1002
rect 942 1000 976 1146
rect 1062 1143 1128 1154
rect 1062 1109 1078 1143
rect 1112 1109 1128 1143
rect 1062 1098 1128 1109
rect 1236 1144 1860 1176
rect 1948 1164 2026 2122
rect 2540 2113 2569 2122
rect 2603 2122 4457 2147
rect 2603 2113 2630 2122
rect 2540 2092 2630 2113
rect 2626 2056 2684 2058
rect 2626 2039 2688 2056
rect 2626 2005 2638 2039
rect 2672 2005 2688 2039
rect 2626 1996 2688 2005
rect 2126 1958 2492 1962
rect 2574 1958 2640 1966
rect 2126 1930 2534 1958
rect 2126 1892 2154 1930
rect 2448 1911 2534 1930
rect 2126 1884 2192 1892
rect 2126 1850 2141 1884
rect 2175 1850 2192 1884
rect 2126 1838 2192 1850
rect 2298 1888 2366 1894
rect 2298 1836 2308 1888
rect 2360 1836 2366 1888
rect 2298 1830 2366 1836
rect 2448 1877 2494 1911
rect 2528 1877 2534 1911
rect 2574 1906 2580 1958
rect 2632 1906 2640 1958
rect 2574 1898 2590 1906
rect 2448 1839 2534 1877
rect 2448 1805 2494 1839
rect 2528 1805 2534 1839
rect 2208 1776 2276 1782
rect 2208 1724 2216 1776
rect 2268 1724 2276 1776
rect 2208 1714 2276 1724
rect 2448 1758 2534 1805
rect 2584 1877 2590 1898
rect 2624 1898 2640 1906
rect 2680 1926 3008 1958
rect 2680 1911 2776 1926
rect 2624 1877 2630 1898
rect 2584 1839 2630 1877
rect 2584 1805 2590 1839
rect 2624 1805 2630 1839
rect 2584 1758 2630 1805
rect 2680 1877 2686 1911
rect 2720 1877 2776 1911
rect 2980 1890 3008 1926
rect 2680 1839 2776 1877
rect 2680 1805 2686 1839
rect 2720 1805 2776 1839
rect 2938 1882 3008 1890
rect 2938 1848 2953 1882
rect 2987 1848 3008 1882
rect 2938 1830 3008 1848
rect 3114 1890 3178 1896
rect 3114 1838 3120 1890
rect 3172 1838 3178 1890
rect 3114 1832 3178 1838
rect 2680 1758 2776 1805
rect 2106 1643 2382 1674
rect 2106 1609 2135 1643
rect 2169 1609 2227 1643
rect 2261 1609 2319 1643
rect 2353 1609 2382 1643
rect 2106 1578 2382 1609
rect 2448 1558 2498 1758
rect 2530 1711 2588 1726
rect 2530 1677 2542 1711
rect 2576 1677 2588 1711
rect 2530 1660 2588 1677
rect 2642 1630 2700 1648
rect 2642 1596 2654 1630
rect 2688 1596 2700 1630
rect 2642 1586 2700 1596
rect 2730 1558 2776 1758
rect 3026 1774 3090 1780
rect 3026 1722 3032 1774
rect 3084 1722 3090 1774
rect 3026 1716 3090 1722
rect 2920 1643 3196 1674
rect 2920 1609 2949 1643
rect 2983 1609 3041 1643
rect 3075 1609 3133 1643
rect 3167 1609 3196 1643
rect 2920 1606 3196 1609
rect 2088 1541 2152 1548
rect 2088 1508 2094 1541
rect 2146 1508 2152 1541
rect 2264 1541 2328 1548
rect 2264 1508 2270 1541
rect 2146 1489 2270 1508
rect 2322 1489 2328 1541
rect 2094 1480 2328 1489
rect 2448 1546 2550 1558
rect 2448 1512 2510 1546
rect 2544 1512 2550 1546
rect 2448 1474 2550 1512
rect 2600 1546 2646 1558
rect 2600 1512 2606 1546
rect 2640 1512 2646 1546
rect 2600 1492 2646 1512
rect 2696 1546 2776 1558
rect 2696 1512 2702 1546
rect 2736 1512 2776 1546
rect 2448 1442 2510 1474
rect 2244 1440 2510 1442
rect 2544 1440 2550 1474
rect 2244 1428 2550 1440
rect 2590 1486 2656 1492
rect 2590 1434 2598 1486
rect 2650 1434 2656 1486
rect 2590 1428 2656 1434
rect 2696 1474 2776 1512
rect 2696 1440 2702 1474
rect 2736 1440 2776 1474
rect 2892 1578 3196 1606
rect 2696 1428 2742 1440
rect 2244 1414 2498 1428
rect 2088 1408 2154 1414
rect 2088 1356 2096 1408
rect 2148 1356 2154 1408
rect 2088 1350 2154 1356
rect 1236 1141 1266 1144
rect 1318 1141 1860 1144
rect 1236 1107 1265 1141
rect 1318 1107 1357 1141
rect 1391 1107 1449 1141
rect 1483 1139 1860 1141
rect 1483 1107 1611 1139
rect 1236 1092 1266 1107
rect 1318 1105 1611 1107
rect 1645 1105 1703 1139
rect 1737 1105 1795 1139
rect 1829 1105 1860 1139
rect 1318 1092 1860 1105
rect 1236 1074 1860 1092
rect 1928 1150 2204 1164
rect 1928 1133 2120 1150
rect 2172 1133 2204 1150
rect 1928 1099 1957 1133
rect 1991 1099 2049 1133
rect 2083 1099 2120 1133
rect 2175 1099 2204 1133
rect 1928 1098 2120 1099
rect 2172 1098 2204 1099
rect 1928 1068 2204 1098
rect 2244 1064 2272 1414
rect 2544 1390 2608 1400
rect 2544 1356 2558 1390
rect 2592 1356 2864 1390
rect 2544 1338 2608 1356
rect 2460 1292 2532 1304
rect 2460 1240 2470 1292
rect 2522 1240 2532 1292
rect 2460 1228 2532 1240
rect 2830 1174 2864 1356
rect 2892 1274 2920 1578
rect 2892 1264 2960 1274
rect 2892 1230 2908 1264
rect 2942 1230 2960 1264
rect 2892 1216 2960 1230
rect 2304 1146 2864 1174
rect 2304 1143 2370 1146
rect 2304 1109 2320 1143
rect 2354 1109 2370 1143
rect 2304 1100 2370 1109
rect 2538 1091 2628 1112
rect 736 983 976 1000
rect 1020 1056 1086 1062
rect 1020 1004 1028 1056
rect 1080 1004 1086 1056
rect 1020 998 1034 1004
rect 470 943 516 976
rect 470 909 476 943
rect 510 909 516 943
rect 736 949 748 983
rect 782 972 976 983
rect 1028 981 1034 998
rect 1068 998 1086 1004
rect 1116 1015 1162 1062
rect 2244 1036 2316 1064
rect 1068 981 1074 998
rect 782 949 974 972
rect 736 940 974 949
rect 470 862 516 909
rect 684 902 750 910
rect 598 898 644 902
rect 558 855 644 898
rect 20 844 88 850
rect 20 792 27 844
rect 79 838 88 844
rect 79 832 172 838
rect 79 798 118 832
rect 152 798 172 832
rect 79 792 172 798
rect 20 788 172 792
rect 416 815 482 826
rect 20 786 88 788
rect 416 781 432 815
rect 466 781 482 815
rect 416 768 482 781
rect 558 821 604 855
rect 638 821 644 855
rect 684 850 690 902
rect 742 850 750 902
rect 684 842 700 850
rect 558 783 644 821
rect 558 749 604 783
rect 638 749 644 783
rect 558 702 644 749
rect 694 821 700 842
rect 734 842 750 850
rect 790 855 886 902
rect 734 821 740 842
rect 694 783 740 821
rect 694 749 700 783
rect 734 749 740 783
rect 694 702 740 749
rect 790 821 796 855
rect 830 821 886 855
rect 790 783 886 821
rect 790 749 796 783
rect 830 749 886 783
rect 790 702 886 749
rect 558 648 608 702
rect 40 602 316 620
rect 40 589 163 602
rect 215 589 316 602
rect 392 598 450 606
rect 40 555 69 589
rect 103 555 161 589
rect 215 555 253 589
rect 287 555 316 589
rect 40 550 163 555
rect 215 550 316 555
rect 40 524 316 550
rect 384 592 458 598
rect 384 540 395 592
rect 447 540 458 592
rect 538 582 608 648
rect 640 655 698 670
rect 640 621 652 655
rect 686 621 698 655
rect 640 604 698 621
rect 384 534 458 540
rect 392 528 450 534
rect 108 254 192 524
rect 558 502 608 582
rect 752 574 810 592
rect 752 540 764 574
rect 798 540 810 574
rect 752 530 810 540
rect 840 502 886 702
rect 558 490 660 502
rect 558 456 620 490
rect 654 456 660 490
rect 558 418 660 456
rect 710 490 756 502
rect 710 456 716 490
rect 750 456 756 490
rect 710 436 756 456
rect 806 490 886 502
rect 806 456 812 490
rect 846 456 886 490
rect 558 384 620 418
rect 654 384 660 418
rect 558 372 660 384
rect 700 430 766 436
rect 700 378 708 430
rect 760 378 766 430
rect 700 372 766 378
rect 806 418 886 456
rect 806 384 812 418
rect 846 384 886 418
rect 914 708 974 940
rect 1028 943 1074 981
rect 1028 909 1034 943
rect 1068 909 1074 943
rect 1028 862 1074 909
rect 1116 981 1122 1015
rect 1156 981 1162 1015
rect 1116 943 1162 981
rect 1116 909 1122 943
rect 1156 909 1162 943
rect 1116 862 1162 909
rect 2270 1015 2316 1036
rect 2270 981 2276 1015
rect 2310 981 2316 1015
rect 2270 943 2316 981
rect 2270 909 2276 943
rect 2310 909 2316 943
rect 2270 862 2316 909
rect 2358 1042 2404 1062
rect 2538 1057 2567 1091
rect 2601 1057 2628 1091
rect 2358 1036 2426 1042
rect 2538 1036 2628 1057
rect 2358 1015 2366 1036
rect 2358 981 2364 1015
rect 2418 984 2426 1036
rect 2398 981 2426 984
rect 2358 976 2426 981
rect 2624 1000 2682 1002
rect 2830 1000 2864 1146
rect 2950 1143 3016 1154
rect 2950 1109 2966 1143
rect 3000 1109 3016 1143
rect 2950 1098 3016 1109
rect 3124 1144 3748 1176
rect 3836 1164 3914 2122
rect 4428 2113 4457 2122
rect 4491 2122 6345 2147
rect 4491 2113 4518 2122
rect 4428 2092 4518 2113
rect 4514 2056 4572 2058
rect 4514 2039 4576 2056
rect 4514 2005 4526 2039
rect 4560 2005 4576 2039
rect 4514 1996 4576 2005
rect 4014 1958 4380 1962
rect 4462 1958 4528 1966
rect 4014 1930 4422 1958
rect 4014 1892 4042 1930
rect 4336 1911 4422 1930
rect 4014 1884 4080 1892
rect 4014 1850 4029 1884
rect 4063 1850 4080 1884
rect 4014 1838 4080 1850
rect 4186 1888 4254 1894
rect 4186 1836 4196 1888
rect 4248 1836 4254 1888
rect 4186 1830 4254 1836
rect 4336 1877 4382 1911
rect 4416 1877 4422 1911
rect 4462 1906 4468 1958
rect 4520 1906 4528 1958
rect 4462 1898 4478 1906
rect 4336 1839 4422 1877
rect 4336 1805 4382 1839
rect 4416 1805 4422 1839
rect 4096 1776 4164 1782
rect 4096 1724 4104 1776
rect 4156 1724 4164 1776
rect 4096 1714 4164 1724
rect 4336 1758 4422 1805
rect 4472 1877 4478 1898
rect 4512 1898 4528 1906
rect 4568 1926 4896 1958
rect 4568 1911 4664 1926
rect 4512 1877 4518 1898
rect 4472 1839 4518 1877
rect 4472 1805 4478 1839
rect 4512 1805 4518 1839
rect 4472 1758 4518 1805
rect 4568 1877 4574 1911
rect 4608 1877 4664 1911
rect 4868 1890 4896 1926
rect 4568 1839 4664 1877
rect 4568 1805 4574 1839
rect 4608 1805 4664 1839
rect 4826 1882 4896 1890
rect 4826 1848 4841 1882
rect 4875 1848 4896 1882
rect 4826 1830 4896 1848
rect 5002 1890 5066 1896
rect 5002 1838 5008 1890
rect 5060 1838 5066 1890
rect 5002 1832 5066 1838
rect 4568 1758 4664 1805
rect 3994 1643 4270 1674
rect 3994 1609 4023 1643
rect 4057 1609 4115 1643
rect 4149 1609 4207 1643
rect 4241 1609 4270 1643
rect 3994 1578 4270 1609
rect 4336 1558 4386 1758
rect 4418 1711 4476 1726
rect 4418 1677 4430 1711
rect 4464 1677 4476 1711
rect 4418 1660 4476 1677
rect 4530 1630 4588 1648
rect 4530 1596 4542 1630
rect 4576 1596 4588 1630
rect 4530 1586 4588 1596
rect 4618 1558 4664 1758
rect 4914 1774 4978 1780
rect 4914 1722 4920 1774
rect 4972 1722 4978 1774
rect 4914 1716 4978 1722
rect 4808 1643 5084 1674
rect 4808 1609 4837 1643
rect 4871 1609 4929 1643
rect 4963 1609 5021 1643
rect 5055 1609 5084 1643
rect 4808 1606 5084 1609
rect 3976 1541 4040 1548
rect 3976 1508 3982 1541
rect 4034 1508 4040 1541
rect 4152 1541 4216 1548
rect 4152 1508 4158 1541
rect 4034 1489 4158 1508
rect 4210 1489 4216 1541
rect 3982 1480 4216 1489
rect 4336 1546 4438 1558
rect 4336 1512 4398 1546
rect 4432 1512 4438 1546
rect 4336 1474 4438 1512
rect 4488 1546 4534 1558
rect 4488 1512 4494 1546
rect 4528 1512 4534 1546
rect 4488 1492 4534 1512
rect 4584 1546 4664 1558
rect 4584 1512 4590 1546
rect 4624 1512 4664 1546
rect 4336 1442 4398 1474
rect 4132 1440 4398 1442
rect 4432 1440 4438 1474
rect 4132 1428 4438 1440
rect 4478 1486 4544 1492
rect 4478 1434 4486 1486
rect 4538 1434 4544 1486
rect 4478 1428 4544 1434
rect 4584 1474 4664 1512
rect 4584 1440 4590 1474
rect 4624 1440 4664 1474
rect 4780 1578 5084 1606
rect 4584 1428 4630 1440
rect 4132 1414 4386 1428
rect 3976 1408 4042 1414
rect 3976 1356 3984 1408
rect 4036 1356 4042 1408
rect 3976 1350 4042 1356
rect 3124 1141 3154 1144
rect 3206 1141 3748 1144
rect 3124 1107 3153 1141
rect 3206 1107 3245 1141
rect 3279 1107 3337 1141
rect 3371 1139 3748 1141
rect 3371 1107 3499 1139
rect 3124 1092 3154 1107
rect 3206 1105 3499 1107
rect 3533 1105 3591 1139
rect 3625 1105 3683 1139
rect 3717 1105 3748 1139
rect 3206 1092 3748 1105
rect 3124 1074 3748 1092
rect 3816 1150 4092 1164
rect 3816 1133 4008 1150
rect 4060 1133 4092 1150
rect 3816 1099 3845 1133
rect 3879 1099 3937 1133
rect 3971 1099 4008 1133
rect 4063 1099 4092 1133
rect 3816 1098 4008 1099
rect 4060 1098 4092 1099
rect 3816 1068 4092 1098
rect 4132 1064 4160 1414
rect 4432 1390 4496 1400
rect 4432 1356 4446 1390
rect 4480 1356 4752 1390
rect 4432 1338 4496 1356
rect 4348 1292 4420 1304
rect 4348 1240 4358 1292
rect 4410 1240 4420 1292
rect 4348 1228 4420 1240
rect 4718 1174 4752 1356
rect 4780 1274 4808 1578
rect 4780 1264 4848 1274
rect 4780 1230 4796 1264
rect 4830 1230 4848 1264
rect 4780 1216 4848 1230
rect 4192 1146 4752 1174
rect 4192 1143 4258 1146
rect 4192 1109 4208 1143
rect 4242 1109 4258 1143
rect 4192 1100 4258 1109
rect 4426 1091 4516 1112
rect 2624 983 2864 1000
rect 2908 1056 2974 1062
rect 2908 1004 2916 1056
rect 2968 1004 2974 1056
rect 2908 998 2922 1004
rect 2358 943 2404 976
rect 2358 909 2364 943
rect 2398 909 2404 943
rect 2624 949 2636 983
rect 2670 972 2864 983
rect 2916 981 2922 998
rect 2956 998 2974 1004
rect 3004 1015 3050 1062
rect 4132 1036 4204 1064
rect 2956 981 2962 998
rect 2670 949 2862 972
rect 2624 940 2862 949
rect 2358 862 2404 909
rect 2572 902 2638 910
rect 2486 898 2532 902
rect 1602 840 1674 844
rect 1062 815 1128 828
rect 1062 781 1078 815
rect 1112 781 1128 815
rect 1062 772 1128 781
rect 1602 788 1611 840
rect 1663 788 1674 840
rect 1602 776 1674 788
rect 1798 838 1872 858
rect 2446 855 2532 898
rect 1798 804 1810 838
rect 1844 804 1872 838
rect 1798 780 1872 804
rect 1908 844 1976 850
rect 1908 792 1915 844
rect 1967 838 1976 844
rect 1967 832 2060 838
rect 1967 798 2006 832
rect 2040 798 2060 832
rect 1967 792 2060 798
rect 1908 788 2060 792
rect 2304 815 2370 826
rect 1908 786 1976 788
rect 2304 781 2320 815
rect 2354 781 2370 815
rect 2304 768 2370 781
rect 2446 821 2492 855
rect 2526 821 2532 855
rect 2572 850 2578 902
rect 2630 850 2638 902
rect 2572 842 2588 850
rect 2446 783 2532 821
rect 2446 749 2492 783
rect 2526 749 2532 783
rect 1384 728 1442 742
rect 1384 708 1396 728
rect 914 694 1396 708
rect 1430 694 1442 728
rect 914 674 1442 694
rect 2446 702 2532 749
rect 2582 821 2588 842
rect 2622 842 2638 850
rect 2678 855 2774 902
rect 2622 821 2628 842
rect 2582 783 2628 821
rect 2582 749 2588 783
rect 2622 749 2628 783
rect 2582 702 2628 749
rect 2678 821 2684 855
rect 2718 821 2774 855
rect 2678 783 2774 821
rect 2678 749 2684 783
rect 2718 749 2774 783
rect 2678 702 2774 749
rect 806 372 852 384
rect 914 344 974 674
rect 2446 648 2496 702
rect 1020 624 1096 630
rect 1020 572 1028 624
rect 1080 572 1096 624
rect 1020 566 1096 572
rect 1236 597 1858 628
rect 654 334 974 344
rect 654 300 668 334
rect 702 300 974 334
rect 654 282 974 300
rect 1236 563 1265 597
rect 1299 563 1357 597
rect 1391 563 1449 597
rect 1483 595 1858 597
rect 1483 563 1611 595
rect 1236 561 1611 563
rect 1645 561 1703 595
rect 1737 561 1795 595
rect 1829 561 1858 595
rect 1236 530 1858 561
rect 1928 602 2204 620
rect 1928 589 2051 602
rect 2103 589 2204 602
rect 2280 598 2338 606
rect 1928 555 1957 589
rect 1991 555 2049 589
rect 2103 555 2141 589
rect 2175 555 2204 589
rect 1928 550 2051 555
rect 2103 550 2204 555
rect 1236 254 1334 530
rect 1928 524 2204 550
rect 2272 592 2346 598
rect 2272 540 2283 592
rect 2335 540 2346 592
rect 2426 582 2496 648
rect 2528 655 2586 670
rect 2528 621 2540 655
rect 2574 621 2586 655
rect 2528 604 2586 621
rect 2272 534 2346 540
rect 2280 528 2338 534
rect 1996 254 2080 524
rect 2446 502 2496 582
rect 2640 574 2698 592
rect 2640 540 2652 574
rect 2686 540 2698 574
rect 2640 530 2698 540
rect 2728 502 2774 702
rect 2446 490 2548 502
rect 2446 456 2508 490
rect 2542 456 2548 490
rect 2446 418 2548 456
rect 2598 490 2644 502
rect 2598 456 2604 490
rect 2638 456 2644 490
rect 2598 436 2644 456
rect 2694 490 2774 502
rect 2694 456 2700 490
rect 2734 456 2774 490
rect 2446 384 2508 418
rect 2542 384 2548 418
rect 2446 372 2548 384
rect 2588 430 2654 436
rect 2588 378 2596 430
rect 2648 378 2654 430
rect 2588 372 2654 378
rect 2694 418 2774 456
rect 2694 384 2700 418
rect 2734 384 2774 418
rect 2802 708 2862 940
rect 2916 943 2962 981
rect 2916 909 2922 943
rect 2956 909 2962 943
rect 2916 862 2962 909
rect 3004 981 3010 1015
rect 3044 981 3050 1015
rect 3004 943 3050 981
rect 3004 909 3010 943
rect 3044 909 3050 943
rect 3004 862 3050 909
rect 4158 1015 4204 1036
rect 4158 981 4164 1015
rect 4198 981 4204 1015
rect 4158 943 4204 981
rect 4158 909 4164 943
rect 4198 909 4204 943
rect 4158 862 4204 909
rect 4246 1042 4292 1062
rect 4426 1057 4455 1091
rect 4489 1057 4516 1091
rect 4246 1036 4314 1042
rect 4426 1036 4516 1057
rect 4246 1015 4254 1036
rect 4246 981 4252 1015
rect 4306 984 4314 1036
rect 4286 981 4314 984
rect 4246 976 4314 981
rect 4512 1000 4570 1002
rect 4718 1000 4752 1146
rect 4838 1143 4904 1154
rect 4838 1109 4854 1143
rect 4888 1109 4904 1143
rect 4838 1098 4904 1109
rect 5012 1144 5636 1176
rect 5724 1164 5802 2122
rect 6316 2113 6345 2122
rect 6379 2122 8233 2147
rect 6379 2113 6406 2122
rect 6316 2092 6406 2113
rect 6402 2056 6460 2058
rect 6402 2039 6464 2056
rect 6402 2005 6414 2039
rect 6448 2005 6464 2039
rect 6402 1996 6464 2005
rect 5902 1958 6268 1962
rect 6350 1958 6416 1966
rect 5902 1930 6310 1958
rect 5902 1892 5930 1930
rect 6224 1911 6310 1930
rect 5902 1884 5968 1892
rect 5902 1850 5917 1884
rect 5951 1850 5968 1884
rect 5902 1838 5968 1850
rect 6074 1888 6142 1894
rect 6074 1836 6084 1888
rect 6136 1836 6142 1888
rect 6074 1830 6142 1836
rect 6224 1877 6270 1911
rect 6304 1877 6310 1911
rect 6350 1906 6356 1958
rect 6408 1906 6416 1958
rect 6350 1898 6366 1906
rect 6224 1839 6310 1877
rect 6224 1805 6270 1839
rect 6304 1805 6310 1839
rect 5984 1776 6052 1782
rect 5984 1724 5992 1776
rect 6044 1724 6052 1776
rect 5984 1714 6052 1724
rect 6224 1758 6310 1805
rect 6360 1877 6366 1898
rect 6400 1898 6416 1906
rect 6456 1926 6784 1958
rect 6456 1911 6552 1926
rect 6400 1877 6406 1898
rect 6360 1839 6406 1877
rect 6360 1805 6366 1839
rect 6400 1805 6406 1839
rect 6360 1758 6406 1805
rect 6456 1877 6462 1911
rect 6496 1877 6552 1911
rect 6756 1890 6784 1926
rect 6456 1839 6552 1877
rect 6456 1805 6462 1839
rect 6496 1805 6552 1839
rect 6714 1882 6784 1890
rect 6714 1848 6729 1882
rect 6763 1848 6784 1882
rect 6714 1830 6784 1848
rect 6890 1890 6954 1896
rect 6890 1838 6896 1890
rect 6948 1838 6954 1890
rect 6890 1832 6954 1838
rect 6456 1758 6552 1805
rect 5882 1643 6158 1674
rect 5882 1609 5911 1643
rect 5945 1609 6003 1643
rect 6037 1609 6095 1643
rect 6129 1609 6158 1643
rect 5882 1578 6158 1609
rect 6224 1558 6274 1758
rect 6306 1711 6364 1726
rect 6306 1677 6318 1711
rect 6352 1677 6364 1711
rect 6306 1660 6364 1677
rect 6418 1630 6476 1648
rect 6418 1596 6430 1630
rect 6464 1596 6476 1630
rect 6418 1586 6476 1596
rect 6506 1558 6552 1758
rect 6802 1774 6866 1780
rect 6802 1722 6808 1774
rect 6860 1722 6866 1774
rect 6802 1716 6866 1722
rect 6696 1643 6972 1674
rect 6696 1609 6725 1643
rect 6759 1609 6817 1643
rect 6851 1609 6909 1643
rect 6943 1609 6972 1643
rect 6696 1606 6972 1609
rect 5864 1541 5928 1548
rect 5864 1508 5870 1541
rect 5922 1508 5928 1541
rect 6040 1541 6104 1548
rect 6040 1508 6046 1541
rect 5922 1489 6046 1508
rect 6098 1489 6104 1541
rect 5870 1480 6104 1489
rect 6224 1546 6326 1558
rect 6224 1512 6286 1546
rect 6320 1512 6326 1546
rect 6224 1474 6326 1512
rect 6376 1546 6422 1558
rect 6376 1512 6382 1546
rect 6416 1512 6422 1546
rect 6376 1492 6422 1512
rect 6472 1546 6552 1558
rect 6472 1512 6478 1546
rect 6512 1512 6552 1546
rect 6224 1442 6286 1474
rect 6020 1440 6286 1442
rect 6320 1440 6326 1474
rect 6020 1428 6326 1440
rect 6366 1486 6432 1492
rect 6366 1434 6374 1486
rect 6426 1434 6432 1486
rect 6366 1428 6432 1434
rect 6472 1474 6552 1512
rect 6472 1440 6478 1474
rect 6512 1440 6552 1474
rect 6668 1578 6972 1606
rect 6472 1428 6518 1440
rect 6020 1414 6274 1428
rect 5864 1408 5930 1414
rect 5864 1356 5872 1408
rect 5924 1356 5930 1408
rect 5864 1350 5930 1356
rect 5012 1141 5042 1144
rect 5094 1141 5636 1144
rect 5012 1107 5041 1141
rect 5094 1107 5133 1141
rect 5167 1107 5225 1141
rect 5259 1139 5636 1141
rect 5259 1107 5387 1139
rect 5012 1092 5042 1107
rect 5094 1105 5387 1107
rect 5421 1105 5479 1139
rect 5513 1105 5571 1139
rect 5605 1105 5636 1139
rect 5094 1092 5636 1105
rect 5012 1074 5636 1092
rect 5704 1150 5980 1164
rect 5704 1133 5896 1150
rect 5948 1133 5980 1150
rect 5704 1099 5733 1133
rect 5767 1099 5825 1133
rect 5859 1099 5896 1133
rect 5951 1099 5980 1133
rect 5704 1098 5896 1099
rect 5948 1098 5980 1099
rect 5704 1068 5980 1098
rect 6020 1064 6048 1414
rect 6320 1390 6384 1400
rect 6320 1356 6334 1390
rect 6368 1356 6640 1390
rect 6320 1338 6384 1356
rect 6236 1292 6308 1304
rect 6236 1240 6246 1292
rect 6298 1240 6308 1292
rect 6236 1228 6308 1240
rect 6606 1174 6640 1356
rect 6668 1274 6696 1578
rect 6668 1264 6736 1274
rect 6668 1230 6684 1264
rect 6718 1230 6736 1264
rect 6668 1216 6736 1230
rect 6080 1146 6640 1174
rect 6080 1143 6146 1146
rect 6080 1109 6096 1143
rect 6130 1109 6146 1143
rect 6080 1100 6146 1109
rect 6314 1091 6404 1112
rect 4512 983 4752 1000
rect 4796 1056 4862 1062
rect 4796 1004 4804 1056
rect 4856 1004 4862 1056
rect 4796 998 4810 1004
rect 4246 943 4292 976
rect 4246 909 4252 943
rect 4286 909 4292 943
rect 4512 949 4524 983
rect 4558 972 4752 983
rect 4804 981 4810 998
rect 4844 998 4862 1004
rect 4892 1015 4938 1062
rect 6020 1036 6092 1064
rect 4844 981 4850 998
rect 4558 949 4750 972
rect 4512 940 4750 949
rect 4246 862 4292 909
rect 4460 902 4526 910
rect 4374 898 4420 902
rect 3490 840 3562 844
rect 2950 815 3016 828
rect 2950 781 2966 815
rect 3000 781 3016 815
rect 2950 772 3016 781
rect 3490 788 3499 840
rect 3551 788 3562 840
rect 3490 776 3562 788
rect 3686 838 3760 858
rect 4334 855 4420 898
rect 3686 804 3698 838
rect 3732 804 3760 838
rect 3686 780 3760 804
rect 3796 844 3864 850
rect 3796 792 3803 844
rect 3855 838 3864 844
rect 3855 832 3948 838
rect 3855 798 3894 832
rect 3928 798 3948 832
rect 3855 792 3948 798
rect 3796 788 3948 792
rect 4192 815 4258 826
rect 3796 786 3864 788
rect 4192 781 4208 815
rect 4242 781 4258 815
rect 4192 768 4258 781
rect 4334 821 4380 855
rect 4414 821 4420 855
rect 4460 850 4466 902
rect 4518 850 4526 902
rect 4460 842 4476 850
rect 4334 783 4420 821
rect 4334 749 4380 783
rect 4414 749 4420 783
rect 3272 728 3330 742
rect 3272 708 3284 728
rect 2802 694 3284 708
rect 3318 694 3330 728
rect 2802 674 3330 694
rect 4334 702 4420 749
rect 4470 821 4476 842
rect 4510 842 4526 850
rect 4566 855 4662 902
rect 4510 821 4516 842
rect 4470 783 4516 821
rect 4470 749 4476 783
rect 4510 749 4516 783
rect 4470 702 4516 749
rect 4566 821 4572 855
rect 4606 821 4662 855
rect 4566 783 4662 821
rect 4566 749 4572 783
rect 4606 749 4662 783
rect 4566 702 4662 749
rect 2694 372 2740 384
rect 2802 344 2862 674
rect 4334 648 4384 702
rect 2908 624 2984 630
rect 2908 572 2916 624
rect 2968 572 2984 624
rect 2908 566 2984 572
rect 3124 597 3746 628
rect 2542 334 2862 344
rect 2542 300 2556 334
rect 2590 300 2862 334
rect 2542 282 2862 300
rect 3124 563 3153 597
rect 3187 563 3245 597
rect 3279 563 3337 597
rect 3371 595 3746 597
rect 3371 563 3499 595
rect 3124 561 3499 563
rect 3533 561 3591 595
rect 3625 561 3683 595
rect 3717 561 3746 595
rect 3124 530 3746 561
rect 3816 602 4092 620
rect 3816 589 3939 602
rect 3991 589 4092 602
rect 4168 598 4226 606
rect 3816 555 3845 589
rect 3879 555 3937 589
rect 3991 555 4029 589
rect 4063 555 4092 589
rect 3816 550 3939 555
rect 3991 550 4092 555
rect 3124 254 3222 530
rect 3816 524 4092 550
rect 4160 592 4234 598
rect 4160 540 4171 592
rect 4223 540 4234 592
rect 4314 582 4384 648
rect 4416 655 4474 670
rect 4416 621 4428 655
rect 4462 621 4474 655
rect 4416 604 4474 621
rect 4160 534 4234 540
rect 4168 528 4226 534
rect 3884 254 3968 524
rect 4334 502 4384 582
rect 4528 574 4586 592
rect 4528 540 4540 574
rect 4574 540 4586 574
rect 4528 530 4586 540
rect 4616 502 4662 702
rect 4334 490 4436 502
rect 4334 456 4396 490
rect 4430 456 4436 490
rect 4334 418 4436 456
rect 4486 490 4532 502
rect 4486 456 4492 490
rect 4526 456 4532 490
rect 4486 436 4532 456
rect 4582 490 4662 502
rect 4582 456 4588 490
rect 4622 456 4662 490
rect 4334 384 4396 418
rect 4430 384 4436 418
rect 4334 372 4436 384
rect 4476 430 4542 436
rect 4476 378 4484 430
rect 4536 378 4542 430
rect 4476 372 4542 378
rect 4582 418 4662 456
rect 4582 384 4588 418
rect 4622 384 4662 418
rect 4690 708 4750 940
rect 4804 943 4850 981
rect 4804 909 4810 943
rect 4844 909 4850 943
rect 4804 862 4850 909
rect 4892 981 4898 1015
rect 4932 981 4938 1015
rect 4892 943 4938 981
rect 4892 909 4898 943
rect 4932 909 4938 943
rect 4892 862 4938 909
rect 6046 1015 6092 1036
rect 6046 981 6052 1015
rect 6086 981 6092 1015
rect 6046 943 6092 981
rect 6046 909 6052 943
rect 6086 909 6092 943
rect 6046 862 6092 909
rect 6134 1042 6180 1062
rect 6314 1057 6343 1091
rect 6377 1057 6404 1091
rect 6134 1036 6202 1042
rect 6314 1036 6404 1057
rect 6134 1015 6142 1036
rect 6134 981 6140 1015
rect 6194 984 6202 1036
rect 6174 981 6202 984
rect 6134 976 6202 981
rect 6400 1000 6458 1002
rect 6606 1000 6640 1146
rect 6726 1143 6792 1154
rect 6726 1109 6742 1143
rect 6776 1109 6792 1143
rect 6726 1098 6792 1109
rect 6900 1144 7524 1176
rect 7612 1164 7690 2122
rect 8204 2113 8233 2122
rect 8267 2122 10121 2147
rect 8267 2113 8294 2122
rect 8204 2092 8294 2113
rect 8290 2056 8348 2058
rect 8290 2039 8352 2056
rect 8290 2005 8302 2039
rect 8336 2005 8352 2039
rect 8290 1996 8352 2005
rect 7790 1958 8156 1962
rect 8238 1958 8304 1966
rect 7790 1930 8198 1958
rect 7790 1892 7818 1930
rect 8112 1911 8198 1930
rect 7790 1884 7856 1892
rect 7790 1850 7805 1884
rect 7839 1850 7856 1884
rect 7790 1838 7856 1850
rect 7962 1888 8030 1894
rect 7962 1836 7972 1888
rect 8024 1836 8030 1888
rect 7962 1830 8030 1836
rect 8112 1877 8158 1911
rect 8192 1877 8198 1911
rect 8238 1906 8244 1958
rect 8296 1906 8304 1958
rect 8238 1898 8254 1906
rect 8112 1839 8198 1877
rect 8112 1805 8158 1839
rect 8192 1805 8198 1839
rect 7872 1776 7940 1782
rect 7872 1724 7880 1776
rect 7932 1724 7940 1776
rect 7872 1714 7940 1724
rect 8112 1758 8198 1805
rect 8248 1877 8254 1898
rect 8288 1898 8304 1906
rect 8344 1926 8672 1958
rect 8344 1911 8440 1926
rect 8288 1877 8294 1898
rect 8248 1839 8294 1877
rect 8248 1805 8254 1839
rect 8288 1805 8294 1839
rect 8248 1758 8294 1805
rect 8344 1877 8350 1911
rect 8384 1877 8440 1911
rect 8644 1890 8672 1926
rect 8344 1839 8440 1877
rect 8344 1805 8350 1839
rect 8384 1805 8440 1839
rect 8602 1882 8672 1890
rect 8602 1848 8617 1882
rect 8651 1848 8672 1882
rect 8602 1830 8672 1848
rect 8778 1890 8842 1896
rect 8778 1838 8784 1890
rect 8836 1838 8842 1890
rect 8778 1832 8842 1838
rect 8344 1758 8440 1805
rect 7770 1643 8046 1674
rect 7770 1609 7799 1643
rect 7833 1609 7891 1643
rect 7925 1609 7983 1643
rect 8017 1609 8046 1643
rect 7770 1578 8046 1609
rect 8112 1558 8162 1758
rect 8194 1711 8252 1726
rect 8194 1677 8206 1711
rect 8240 1677 8252 1711
rect 8194 1660 8252 1677
rect 8306 1630 8364 1648
rect 8306 1596 8318 1630
rect 8352 1596 8364 1630
rect 8306 1586 8364 1596
rect 8394 1558 8440 1758
rect 8690 1774 8754 1780
rect 8690 1722 8696 1774
rect 8748 1722 8754 1774
rect 8690 1716 8754 1722
rect 8584 1643 8860 1674
rect 8584 1609 8613 1643
rect 8647 1609 8705 1643
rect 8739 1609 8797 1643
rect 8831 1609 8860 1643
rect 8584 1606 8860 1609
rect 7752 1541 7816 1548
rect 7752 1508 7758 1541
rect 7810 1508 7816 1541
rect 7928 1541 7992 1548
rect 7928 1508 7934 1541
rect 7810 1489 7934 1508
rect 7986 1489 7992 1541
rect 7758 1480 7992 1489
rect 8112 1546 8214 1558
rect 8112 1512 8174 1546
rect 8208 1512 8214 1546
rect 8112 1474 8214 1512
rect 8264 1546 8310 1558
rect 8264 1512 8270 1546
rect 8304 1512 8310 1546
rect 8264 1492 8310 1512
rect 8360 1546 8440 1558
rect 8360 1512 8366 1546
rect 8400 1512 8440 1546
rect 8112 1442 8174 1474
rect 7908 1440 8174 1442
rect 8208 1440 8214 1474
rect 7908 1428 8214 1440
rect 8254 1486 8320 1492
rect 8254 1434 8262 1486
rect 8314 1434 8320 1486
rect 8254 1428 8320 1434
rect 8360 1474 8440 1512
rect 8360 1440 8366 1474
rect 8400 1440 8440 1474
rect 8556 1578 8860 1606
rect 8360 1428 8406 1440
rect 7908 1414 8162 1428
rect 7752 1408 7818 1414
rect 7752 1356 7760 1408
rect 7812 1356 7818 1408
rect 7752 1350 7818 1356
rect 6900 1141 6930 1144
rect 6982 1141 7524 1144
rect 6900 1107 6929 1141
rect 6982 1107 7021 1141
rect 7055 1107 7113 1141
rect 7147 1139 7524 1141
rect 7147 1107 7275 1139
rect 6900 1092 6930 1107
rect 6982 1105 7275 1107
rect 7309 1105 7367 1139
rect 7401 1105 7459 1139
rect 7493 1105 7524 1139
rect 6982 1092 7524 1105
rect 6900 1074 7524 1092
rect 7592 1150 7868 1164
rect 7592 1133 7784 1150
rect 7836 1133 7868 1150
rect 7592 1099 7621 1133
rect 7655 1099 7713 1133
rect 7747 1099 7784 1133
rect 7839 1099 7868 1133
rect 7592 1098 7784 1099
rect 7836 1098 7868 1099
rect 7592 1068 7868 1098
rect 7908 1064 7936 1414
rect 8208 1390 8272 1400
rect 8208 1356 8222 1390
rect 8256 1356 8528 1390
rect 8208 1338 8272 1356
rect 8124 1292 8196 1304
rect 8124 1240 8134 1292
rect 8186 1240 8196 1292
rect 8124 1228 8196 1240
rect 8494 1174 8528 1356
rect 8556 1274 8584 1578
rect 8556 1264 8624 1274
rect 8556 1230 8572 1264
rect 8606 1230 8624 1264
rect 8556 1216 8624 1230
rect 7968 1146 8528 1174
rect 7968 1143 8034 1146
rect 7968 1109 7984 1143
rect 8018 1109 8034 1143
rect 7968 1100 8034 1109
rect 8202 1091 8292 1112
rect 6400 983 6640 1000
rect 6684 1056 6750 1062
rect 6684 1004 6692 1056
rect 6744 1004 6750 1056
rect 6684 998 6698 1004
rect 6134 943 6180 976
rect 6134 909 6140 943
rect 6174 909 6180 943
rect 6400 949 6412 983
rect 6446 972 6640 983
rect 6692 981 6698 998
rect 6732 998 6750 1004
rect 6780 1015 6826 1062
rect 7908 1036 7980 1064
rect 6732 981 6738 998
rect 6446 949 6638 972
rect 6400 940 6638 949
rect 6134 862 6180 909
rect 6348 902 6414 910
rect 6262 898 6308 902
rect 5378 840 5450 844
rect 4838 815 4904 828
rect 4838 781 4854 815
rect 4888 781 4904 815
rect 4838 772 4904 781
rect 5378 788 5387 840
rect 5439 788 5450 840
rect 5378 776 5450 788
rect 5574 838 5648 858
rect 6222 855 6308 898
rect 5574 804 5586 838
rect 5620 804 5648 838
rect 5574 780 5648 804
rect 5684 844 5752 850
rect 5684 792 5691 844
rect 5743 838 5752 844
rect 5743 832 5836 838
rect 5743 798 5782 832
rect 5816 798 5836 832
rect 5743 792 5836 798
rect 5684 788 5836 792
rect 6080 815 6146 826
rect 5684 786 5752 788
rect 6080 781 6096 815
rect 6130 781 6146 815
rect 6080 768 6146 781
rect 6222 821 6268 855
rect 6302 821 6308 855
rect 6348 850 6354 902
rect 6406 850 6414 902
rect 6348 842 6364 850
rect 6222 783 6308 821
rect 6222 749 6268 783
rect 6302 749 6308 783
rect 5160 728 5218 742
rect 5160 708 5172 728
rect 4690 694 5172 708
rect 5206 694 5218 728
rect 4690 674 5218 694
rect 6222 702 6308 749
rect 6358 821 6364 842
rect 6398 842 6414 850
rect 6454 855 6550 902
rect 6398 821 6404 842
rect 6358 783 6404 821
rect 6358 749 6364 783
rect 6398 749 6404 783
rect 6358 702 6404 749
rect 6454 821 6460 855
rect 6494 821 6550 855
rect 6454 783 6550 821
rect 6454 749 6460 783
rect 6494 749 6550 783
rect 6454 702 6550 749
rect 4582 372 4628 384
rect 4690 344 4750 674
rect 6222 648 6272 702
rect 4796 624 4872 630
rect 4796 572 4804 624
rect 4856 572 4872 624
rect 4796 566 4872 572
rect 5012 597 5634 628
rect 4430 334 4750 344
rect 4430 300 4444 334
rect 4478 300 4750 334
rect 4430 282 4750 300
rect 5012 563 5041 597
rect 5075 563 5133 597
rect 5167 563 5225 597
rect 5259 595 5634 597
rect 5259 563 5387 595
rect 5012 561 5387 563
rect 5421 561 5479 595
rect 5513 561 5571 595
rect 5605 561 5634 595
rect 5012 530 5634 561
rect 5704 602 5980 620
rect 5704 589 5827 602
rect 5879 589 5980 602
rect 6056 598 6114 606
rect 5704 555 5733 589
rect 5767 555 5825 589
rect 5879 555 5917 589
rect 5951 555 5980 589
rect 5704 550 5827 555
rect 5879 550 5980 555
rect 5012 254 5110 530
rect 5704 524 5980 550
rect 6048 592 6122 598
rect 6048 540 6059 592
rect 6111 540 6122 592
rect 6202 582 6272 648
rect 6304 655 6362 670
rect 6304 621 6316 655
rect 6350 621 6362 655
rect 6304 604 6362 621
rect 6048 534 6122 540
rect 6056 528 6114 534
rect 5772 254 5856 524
rect 6222 502 6272 582
rect 6416 574 6474 592
rect 6416 540 6428 574
rect 6462 540 6474 574
rect 6416 530 6474 540
rect 6504 502 6550 702
rect 6222 490 6324 502
rect 6222 456 6284 490
rect 6318 456 6324 490
rect 6222 418 6324 456
rect 6374 490 6420 502
rect 6374 456 6380 490
rect 6414 456 6420 490
rect 6374 436 6420 456
rect 6470 490 6550 502
rect 6470 456 6476 490
rect 6510 456 6550 490
rect 6222 384 6284 418
rect 6318 384 6324 418
rect 6222 372 6324 384
rect 6364 430 6430 436
rect 6364 378 6372 430
rect 6424 378 6430 430
rect 6364 372 6430 378
rect 6470 418 6550 456
rect 6470 384 6476 418
rect 6510 384 6550 418
rect 6578 708 6638 940
rect 6692 943 6738 981
rect 6692 909 6698 943
rect 6732 909 6738 943
rect 6692 862 6738 909
rect 6780 981 6786 1015
rect 6820 981 6826 1015
rect 6780 943 6826 981
rect 6780 909 6786 943
rect 6820 909 6826 943
rect 6780 862 6826 909
rect 7934 1015 7980 1036
rect 7934 981 7940 1015
rect 7974 981 7980 1015
rect 7934 943 7980 981
rect 7934 909 7940 943
rect 7974 909 7980 943
rect 7934 862 7980 909
rect 8022 1042 8068 1062
rect 8202 1057 8231 1091
rect 8265 1057 8292 1091
rect 8022 1036 8090 1042
rect 8202 1036 8292 1057
rect 8022 1015 8030 1036
rect 8022 981 8028 1015
rect 8082 984 8090 1036
rect 8062 981 8090 984
rect 8022 976 8090 981
rect 8288 1000 8346 1002
rect 8494 1000 8528 1146
rect 8614 1143 8680 1154
rect 8614 1109 8630 1143
rect 8664 1109 8680 1143
rect 8614 1098 8680 1109
rect 8788 1144 9412 1176
rect 9500 1164 9578 2122
rect 10092 2113 10121 2122
rect 10155 2122 12009 2147
rect 10155 2113 10182 2122
rect 10092 2092 10182 2113
rect 10178 2056 10236 2058
rect 10178 2039 10240 2056
rect 10178 2005 10190 2039
rect 10224 2005 10240 2039
rect 10178 1996 10240 2005
rect 9678 1958 10044 1962
rect 10126 1958 10192 1966
rect 9678 1930 10086 1958
rect 9678 1892 9706 1930
rect 10000 1911 10086 1930
rect 9678 1884 9744 1892
rect 9678 1850 9693 1884
rect 9727 1850 9744 1884
rect 9678 1838 9744 1850
rect 9850 1888 9918 1894
rect 9850 1836 9860 1888
rect 9912 1836 9918 1888
rect 9850 1830 9918 1836
rect 10000 1877 10046 1911
rect 10080 1877 10086 1911
rect 10126 1906 10132 1958
rect 10184 1906 10192 1958
rect 10126 1898 10142 1906
rect 10000 1839 10086 1877
rect 10000 1805 10046 1839
rect 10080 1805 10086 1839
rect 9760 1776 9828 1782
rect 9760 1724 9768 1776
rect 9820 1724 9828 1776
rect 9760 1714 9828 1724
rect 10000 1758 10086 1805
rect 10136 1877 10142 1898
rect 10176 1898 10192 1906
rect 10232 1926 10560 1958
rect 10232 1911 10328 1926
rect 10176 1877 10182 1898
rect 10136 1839 10182 1877
rect 10136 1805 10142 1839
rect 10176 1805 10182 1839
rect 10136 1758 10182 1805
rect 10232 1877 10238 1911
rect 10272 1877 10328 1911
rect 10532 1890 10560 1926
rect 10232 1839 10328 1877
rect 10232 1805 10238 1839
rect 10272 1805 10328 1839
rect 10490 1882 10560 1890
rect 10490 1848 10505 1882
rect 10539 1848 10560 1882
rect 10490 1830 10560 1848
rect 10666 1890 10730 1896
rect 10666 1838 10672 1890
rect 10724 1838 10730 1890
rect 10666 1832 10730 1838
rect 10232 1758 10328 1805
rect 9658 1643 9934 1674
rect 9658 1609 9687 1643
rect 9721 1609 9779 1643
rect 9813 1609 9871 1643
rect 9905 1609 9934 1643
rect 9658 1578 9934 1609
rect 10000 1558 10050 1758
rect 10082 1711 10140 1726
rect 10082 1677 10094 1711
rect 10128 1677 10140 1711
rect 10082 1660 10140 1677
rect 10194 1630 10252 1648
rect 10194 1596 10206 1630
rect 10240 1596 10252 1630
rect 10194 1586 10252 1596
rect 10282 1558 10328 1758
rect 10578 1774 10642 1780
rect 10578 1722 10584 1774
rect 10636 1722 10642 1774
rect 10578 1716 10642 1722
rect 10472 1643 10748 1674
rect 10472 1609 10501 1643
rect 10535 1609 10593 1643
rect 10627 1609 10685 1643
rect 10719 1609 10748 1643
rect 10472 1606 10748 1609
rect 9640 1541 9704 1548
rect 9640 1508 9646 1541
rect 9698 1508 9704 1541
rect 9816 1541 9880 1548
rect 9816 1508 9822 1541
rect 9698 1489 9822 1508
rect 9874 1489 9880 1541
rect 9646 1480 9880 1489
rect 10000 1546 10102 1558
rect 10000 1512 10062 1546
rect 10096 1512 10102 1546
rect 10000 1474 10102 1512
rect 10152 1546 10198 1558
rect 10152 1512 10158 1546
rect 10192 1512 10198 1546
rect 10152 1492 10198 1512
rect 10248 1546 10328 1558
rect 10248 1512 10254 1546
rect 10288 1512 10328 1546
rect 10000 1442 10062 1474
rect 9796 1440 10062 1442
rect 10096 1440 10102 1474
rect 9796 1428 10102 1440
rect 10142 1486 10208 1492
rect 10142 1434 10150 1486
rect 10202 1434 10208 1486
rect 10142 1428 10208 1434
rect 10248 1474 10328 1512
rect 10248 1440 10254 1474
rect 10288 1440 10328 1474
rect 10444 1578 10748 1606
rect 10248 1428 10294 1440
rect 9796 1414 10050 1428
rect 9640 1408 9706 1414
rect 9640 1356 9648 1408
rect 9700 1356 9706 1408
rect 9640 1350 9706 1356
rect 8788 1141 8818 1144
rect 8870 1141 9412 1144
rect 8788 1107 8817 1141
rect 8870 1107 8909 1141
rect 8943 1107 9001 1141
rect 9035 1139 9412 1141
rect 9035 1107 9163 1139
rect 8788 1092 8818 1107
rect 8870 1105 9163 1107
rect 9197 1105 9255 1139
rect 9289 1105 9347 1139
rect 9381 1105 9412 1139
rect 8870 1092 9412 1105
rect 8788 1074 9412 1092
rect 9480 1150 9756 1164
rect 9480 1133 9672 1150
rect 9724 1133 9756 1150
rect 9480 1099 9509 1133
rect 9543 1099 9601 1133
rect 9635 1099 9672 1133
rect 9727 1099 9756 1133
rect 9480 1098 9672 1099
rect 9724 1098 9756 1099
rect 9480 1068 9756 1098
rect 9796 1064 9824 1414
rect 10096 1390 10160 1400
rect 10096 1356 10110 1390
rect 10144 1356 10416 1390
rect 10096 1338 10160 1356
rect 10012 1292 10084 1304
rect 10012 1240 10022 1292
rect 10074 1240 10084 1292
rect 10012 1228 10084 1240
rect 10382 1174 10416 1356
rect 10444 1274 10472 1578
rect 10444 1264 10512 1274
rect 10444 1230 10460 1264
rect 10494 1230 10512 1264
rect 10444 1216 10512 1230
rect 9856 1146 10416 1174
rect 9856 1143 9922 1146
rect 9856 1109 9872 1143
rect 9906 1109 9922 1143
rect 9856 1100 9922 1109
rect 10090 1091 10180 1112
rect 8288 983 8528 1000
rect 8572 1056 8638 1062
rect 8572 1004 8580 1056
rect 8632 1004 8638 1056
rect 8572 998 8586 1004
rect 8022 943 8068 976
rect 8022 909 8028 943
rect 8062 909 8068 943
rect 8288 949 8300 983
rect 8334 972 8528 983
rect 8580 981 8586 998
rect 8620 998 8638 1004
rect 8668 1015 8714 1062
rect 9796 1036 9868 1064
rect 8620 981 8626 998
rect 8334 949 8526 972
rect 8288 940 8526 949
rect 8022 862 8068 909
rect 8236 902 8302 910
rect 8150 898 8196 902
rect 7266 840 7338 844
rect 6726 815 6792 828
rect 6726 781 6742 815
rect 6776 781 6792 815
rect 6726 772 6792 781
rect 7266 788 7275 840
rect 7327 788 7338 840
rect 7266 776 7338 788
rect 7462 838 7536 858
rect 8110 855 8196 898
rect 7462 804 7474 838
rect 7508 804 7536 838
rect 7462 780 7536 804
rect 7572 844 7640 850
rect 7572 792 7579 844
rect 7631 838 7640 844
rect 7631 832 7724 838
rect 7631 798 7670 832
rect 7704 798 7724 832
rect 7631 792 7724 798
rect 7572 788 7724 792
rect 7968 815 8034 826
rect 7572 786 7640 788
rect 7968 781 7984 815
rect 8018 781 8034 815
rect 7968 768 8034 781
rect 8110 821 8156 855
rect 8190 821 8196 855
rect 8236 850 8242 902
rect 8294 850 8302 902
rect 8236 842 8252 850
rect 8110 783 8196 821
rect 8110 749 8156 783
rect 8190 749 8196 783
rect 7048 728 7106 742
rect 7048 708 7060 728
rect 6578 694 7060 708
rect 7094 694 7106 728
rect 6578 674 7106 694
rect 8110 702 8196 749
rect 8246 821 8252 842
rect 8286 842 8302 850
rect 8342 855 8438 902
rect 8286 821 8292 842
rect 8246 783 8292 821
rect 8246 749 8252 783
rect 8286 749 8292 783
rect 8246 702 8292 749
rect 8342 821 8348 855
rect 8382 821 8438 855
rect 8342 783 8438 821
rect 8342 749 8348 783
rect 8382 749 8438 783
rect 8342 702 8438 749
rect 6470 372 6516 384
rect 6578 344 6638 674
rect 8110 648 8160 702
rect 6684 624 6760 630
rect 6684 572 6692 624
rect 6744 572 6760 624
rect 6684 566 6760 572
rect 6900 597 7522 628
rect 6318 334 6638 344
rect 6318 300 6332 334
rect 6366 300 6638 334
rect 6318 282 6638 300
rect 6900 563 6929 597
rect 6963 563 7021 597
rect 7055 563 7113 597
rect 7147 595 7522 597
rect 7147 563 7275 595
rect 6900 561 7275 563
rect 7309 561 7367 595
rect 7401 561 7459 595
rect 7493 561 7522 595
rect 6900 530 7522 561
rect 7592 602 7868 620
rect 7592 589 7715 602
rect 7767 589 7868 602
rect 7944 598 8002 606
rect 7592 555 7621 589
rect 7655 555 7713 589
rect 7767 555 7805 589
rect 7839 555 7868 589
rect 7592 550 7715 555
rect 7767 550 7868 555
rect 6900 254 6998 530
rect 7592 524 7868 550
rect 7936 592 8010 598
rect 7936 540 7947 592
rect 7999 540 8010 592
rect 8090 582 8160 648
rect 8192 655 8250 670
rect 8192 621 8204 655
rect 8238 621 8250 655
rect 8192 604 8250 621
rect 7936 534 8010 540
rect 7944 528 8002 534
rect 7660 254 7744 524
rect 8110 502 8160 582
rect 8304 574 8362 592
rect 8304 540 8316 574
rect 8350 540 8362 574
rect 8304 530 8362 540
rect 8392 502 8438 702
rect 8110 490 8212 502
rect 8110 456 8172 490
rect 8206 456 8212 490
rect 8110 418 8212 456
rect 8262 490 8308 502
rect 8262 456 8268 490
rect 8302 456 8308 490
rect 8262 436 8308 456
rect 8358 490 8438 502
rect 8358 456 8364 490
rect 8398 456 8438 490
rect 8110 384 8172 418
rect 8206 384 8212 418
rect 8110 372 8212 384
rect 8252 430 8318 436
rect 8252 378 8260 430
rect 8312 378 8318 430
rect 8252 372 8318 378
rect 8358 418 8438 456
rect 8358 384 8364 418
rect 8398 384 8438 418
rect 8466 708 8526 940
rect 8580 943 8626 981
rect 8580 909 8586 943
rect 8620 909 8626 943
rect 8580 862 8626 909
rect 8668 981 8674 1015
rect 8708 981 8714 1015
rect 8668 943 8714 981
rect 8668 909 8674 943
rect 8708 909 8714 943
rect 8668 862 8714 909
rect 9822 1015 9868 1036
rect 9822 981 9828 1015
rect 9862 981 9868 1015
rect 9822 943 9868 981
rect 9822 909 9828 943
rect 9862 909 9868 943
rect 9822 862 9868 909
rect 9910 1042 9956 1062
rect 10090 1057 10119 1091
rect 10153 1057 10180 1091
rect 9910 1036 9978 1042
rect 10090 1036 10180 1057
rect 9910 1015 9918 1036
rect 9910 981 9916 1015
rect 9970 984 9978 1036
rect 9950 981 9978 984
rect 9910 976 9978 981
rect 10176 1000 10234 1002
rect 10382 1000 10416 1146
rect 10502 1143 10568 1154
rect 10502 1109 10518 1143
rect 10552 1109 10568 1143
rect 10502 1098 10568 1109
rect 10676 1144 11300 1176
rect 11388 1164 11466 2122
rect 11980 2113 12009 2122
rect 12043 2122 13897 2147
rect 12043 2113 12070 2122
rect 11980 2092 12070 2113
rect 12066 2056 12124 2058
rect 12066 2039 12128 2056
rect 12066 2005 12078 2039
rect 12112 2005 12128 2039
rect 12066 1996 12128 2005
rect 11566 1958 11932 1962
rect 12014 1958 12080 1966
rect 11566 1930 11974 1958
rect 11566 1892 11594 1930
rect 11888 1911 11974 1930
rect 11566 1884 11632 1892
rect 11566 1850 11581 1884
rect 11615 1850 11632 1884
rect 11566 1838 11632 1850
rect 11738 1888 11806 1894
rect 11738 1836 11748 1888
rect 11800 1836 11806 1888
rect 11738 1830 11806 1836
rect 11888 1877 11934 1911
rect 11968 1877 11974 1911
rect 12014 1906 12020 1958
rect 12072 1906 12080 1958
rect 12014 1898 12030 1906
rect 11888 1839 11974 1877
rect 11888 1805 11934 1839
rect 11968 1805 11974 1839
rect 11648 1776 11716 1782
rect 11648 1724 11656 1776
rect 11708 1724 11716 1776
rect 11648 1714 11716 1724
rect 11888 1758 11974 1805
rect 12024 1877 12030 1898
rect 12064 1898 12080 1906
rect 12120 1926 12448 1958
rect 12120 1911 12216 1926
rect 12064 1877 12070 1898
rect 12024 1839 12070 1877
rect 12024 1805 12030 1839
rect 12064 1805 12070 1839
rect 12024 1758 12070 1805
rect 12120 1877 12126 1911
rect 12160 1877 12216 1911
rect 12420 1890 12448 1926
rect 12120 1839 12216 1877
rect 12120 1805 12126 1839
rect 12160 1805 12216 1839
rect 12378 1882 12448 1890
rect 12378 1848 12393 1882
rect 12427 1848 12448 1882
rect 12378 1830 12448 1848
rect 12554 1890 12618 1896
rect 12554 1838 12560 1890
rect 12612 1838 12618 1890
rect 12554 1832 12618 1838
rect 12120 1758 12216 1805
rect 11546 1643 11822 1674
rect 11546 1609 11575 1643
rect 11609 1609 11667 1643
rect 11701 1609 11759 1643
rect 11793 1609 11822 1643
rect 11546 1578 11822 1609
rect 11888 1558 11938 1758
rect 11970 1711 12028 1726
rect 11970 1677 11982 1711
rect 12016 1677 12028 1711
rect 11970 1660 12028 1677
rect 12082 1630 12140 1648
rect 12082 1596 12094 1630
rect 12128 1596 12140 1630
rect 12082 1586 12140 1596
rect 12170 1558 12216 1758
rect 12466 1774 12530 1780
rect 12466 1722 12472 1774
rect 12524 1722 12530 1774
rect 12466 1716 12530 1722
rect 12360 1643 12636 1674
rect 12360 1609 12389 1643
rect 12423 1609 12481 1643
rect 12515 1609 12573 1643
rect 12607 1609 12636 1643
rect 12360 1606 12636 1609
rect 11528 1541 11592 1548
rect 11528 1508 11534 1541
rect 11586 1508 11592 1541
rect 11704 1541 11768 1548
rect 11704 1508 11710 1541
rect 11586 1489 11710 1508
rect 11762 1489 11768 1541
rect 11534 1480 11768 1489
rect 11888 1546 11990 1558
rect 11888 1512 11950 1546
rect 11984 1512 11990 1546
rect 11888 1474 11990 1512
rect 12040 1546 12086 1558
rect 12040 1512 12046 1546
rect 12080 1512 12086 1546
rect 12040 1492 12086 1512
rect 12136 1546 12216 1558
rect 12136 1512 12142 1546
rect 12176 1512 12216 1546
rect 11888 1442 11950 1474
rect 11684 1440 11950 1442
rect 11984 1440 11990 1474
rect 11684 1428 11990 1440
rect 12030 1486 12096 1492
rect 12030 1434 12038 1486
rect 12090 1434 12096 1486
rect 12030 1428 12096 1434
rect 12136 1474 12216 1512
rect 12136 1440 12142 1474
rect 12176 1440 12216 1474
rect 12332 1578 12636 1606
rect 12136 1428 12182 1440
rect 11684 1414 11938 1428
rect 11528 1408 11594 1414
rect 11528 1356 11536 1408
rect 11588 1356 11594 1408
rect 11528 1350 11594 1356
rect 10676 1141 10706 1144
rect 10758 1141 11300 1144
rect 10676 1107 10705 1141
rect 10758 1107 10797 1141
rect 10831 1107 10889 1141
rect 10923 1139 11300 1141
rect 10923 1107 11051 1139
rect 10676 1092 10706 1107
rect 10758 1105 11051 1107
rect 11085 1105 11143 1139
rect 11177 1105 11235 1139
rect 11269 1105 11300 1139
rect 10758 1092 11300 1105
rect 10676 1074 11300 1092
rect 11368 1150 11644 1164
rect 11368 1133 11560 1150
rect 11612 1133 11644 1150
rect 11368 1099 11397 1133
rect 11431 1099 11489 1133
rect 11523 1099 11560 1133
rect 11615 1099 11644 1133
rect 11368 1098 11560 1099
rect 11612 1098 11644 1099
rect 11368 1068 11644 1098
rect 11684 1064 11712 1414
rect 11984 1390 12048 1400
rect 11984 1356 11998 1390
rect 12032 1356 12304 1390
rect 11984 1338 12048 1356
rect 11900 1292 11972 1304
rect 11900 1240 11910 1292
rect 11962 1240 11972 1292
rect 11900 1228 11972 1240
rect 12270 1174 12304 1356
rect 12332 1274 12360 1578
rect 12332 1264 12400 1274
rect 12332 1230 12348 1264
rect 12382 1230 12400 1264
rect 12332 1216 12400 1230
rect 11744 1146 12304 1174
rect 11744 1143 11810 1146
rect 11744 1109 11760 1143
rect 11794 1109 11810 1143
rect 11744 1100 11810 1109
rect 11978 1091 12068 1112
rect 10176 983 10416 1000
rect 10460 1056 10526 1062
rect 10460 1004 10468 1056
rect 10520 1004 10526 1056
rect 10460 998 10474 1004
rect 9910 943 9956 976
rect 9910 909 9916 943
rect 9950 909 9956 943
rect 10176 949 10188 983
rect 10222 972 10416 983
rect 10468 981 10474 998
rect 10508 998 10526 1004
rect 10556 1015 10602 1062
rect 11684 1036 11756 1064
rect 10508 981 10514 998
rect 10222 949 10414 972
rect 10176 940 10414 949
rect 9910 862 9956 909
rect 10124 902 10190 910
rect 10038 898 10084 902
rect 9154 840 9226 844
rect 8614 815 8680 828
rect 8614 781 8630 815
rect 8664 781 8680 815
rect 8614 772 8680 781
rect 9154 788 9163 840
rect 9215 788 9226 840
rect 9154 776 9226 788
rect 9350 838 9424 858
rect 9998 855 10084 898
rect 9350 804 9362 838
rect 9396 804 9424 838
rect 9350 780 9424 804
rect 9460 844 9528 850
rect 9460 792 9467 844
rect 9519 838 9528 844
rect 9519 832 9612 838
rect 9519 798 9558 832
rect 9592 798 9612 832
rect 9519 792 9612 798
rect 9460 788 9612 792
rect 9856 815 9922 826
rect 9460 786 9528 788
rect 9856 781 9872 815
rect 9906 781 9922 815
rect 9856 768 9922 781
rect 9998 821 10044 855
rect 10078 821 10084 855
rect 10124 850 10130 902
rect 10182 850 10190 902
rect 10124 842 10140 850
rect 9998 783 10084 821
rect 9998 749 10044 783
rect 10078 749 10084 783
rect 8936 728 8994 742
rect 8936 708 8948 728
rect 8466 694 8948 708
rect 8982 694 8994 728
rect 8466 674 8994 694
rect 9998 702 10084 749
rect 10134 821 10140 842
rect 10174 842 10190 850
rect 10230 855 10326 902
rect 10174 821 10180 842
rect 10134 783 10180 821
rect 10134 749 10140 783
rect 10174 749 10180 783
rect 10134 702 10180 749
rect 10230 821 10236 855
rect 10270 821 10326 855
rect 10230 783 10326 821
rect 10230 749 10236 783
rect 10270 749 10326 783
rect 10230 702 10326 749
rect 8358 372 8404 384
rect 8466 344 8526 674
rect 9998 648 10048 702
rect 8572 624 8648 630
rect 8572 572 8580 624
rect 8632 572 8648 624
rect 8572 566 8648 572
rect 8788 597 9410 628
rect 8206 334 8526 344
rect 8206 300 8220 334
rect 8254 300 8526 334
rect 8206 282 8526 300
rect 8788 563 8817 597
rect 8851 563 8909 597
rect 8943 563 9001 597
rect 9035 595 9410 597
rect 9035 563 9163 595
rect 8788 561 9163 563
rect 9197 561 9255 595
rect 9289 561 9347 595
rect 9381 561 9410 595
rect 8788 530 9410 561
rect 9480 602 9756 620
rect 9480 589 9603 602
rect 9655 589 9756 602
rect 9832 598 9890 606
rect 9480 555 9509 589
rect 9543 555 9601 589
rect 9655 555 9693 589
rect 9727 555 9756 589
rect 9480 550 9603 555
rect 9655 550 9756 555
rect 8788 254 8886 530
rect 9480 524 9756 550
rect 9824 592 9898 598
rect 9824 540 9835 592
rect 9887 540 9898 592
rect 9978 582 10048 648
rect 10080 655 10138 670
rect 10080 621 10092 655
rect 10126 621 10138 655
rect 10080 604 10138 621
rect 9824 534 9898 540
rect 9832 528 9890 534
rect 9548 254 9632 524
rect 9998 502 10048 582
rect 10192 574 10250 592
rect 10192 540 10204 574
rect 10238 540 10250 574
rect 10192 530 10250 540
rect 10280 502 10326 702
rect 9998 490 10100 502
rect 9998 456 10060 490
rect 10094 456 10100 490
rect 9998 418 10100 456
rect 10150 490 10196 502
rect 10150 456 10156 490
rect 10190 456 10196 490
rect 10150 436 10196 456
rect 10246 490 10326 502
rect 10246 456 10252 490
rect 10286 456 10326 490
rect 9998 384 10060 418
rect 10094 384 10100 418
rect 9998 372 10100 384
rect 10140 430 10206 436
rect 10140 378 10148 430
rect 10200 378 10206 430
rect 10140 372 10206 378
rect 10246 418 10326 456
rect 10246 384 10252 418
rect 10286 384 10326 418
rect 10354 708 10414 940
rect 10468 943 10514 981
rect 10468 909 10474 943
rect 10508 909 10514 943
rect 10468 862 10514 909
rect 10556 981 10562 1015
rect 10596 981 10602 1015
rect 10556 943 10602 981
rect 10556 909 10562 943
rect 10596 909 10602 943
rect 10556 862 10602 909
rect 11710 1015 11756 1036
rect 11710 981 11716 1015
rect 11750 981 11756 1015
rect 11710 943 11756 981
rect 11710 909 11716 943
rect 11750 909 11756 943
rect 11710 862 11756 909
rect 11798 1042 11844 1062
rect 11978 1057 12007 1091
rect 12041 1057 12068 1091
rect 11798 1036 11866 1042
rect 11978 1036 12068 1057
rect 11798 1015 11806 1036
rect 11798 981 11804 1015
rect 11858 984 11866 1036
rect 11838 981 11866 984
rect 11798 976 11866 981
rect 12064 1000 12122 1002
rect 12270 1000 12304 1146
rect 12390 1143 12456 1154
rect 12390 1109 12406 1143
rect 12440 1109 12456 1143
rect 12390 1098 12456 1109
rect 12564 1144 13188 1176
rect 13276 1164 13354 2122
rect 13868 2113 13897 2122
rect 13931 2122 15779 2147
rect 13931 2113 13958 2122
rect 13868 2092 13958 2113
rect 13954 2056 14012 2058
rect 13954 2039 14016 2056
rect 13954 2005 13966 2039
rect 14000 2005 14016 2039
rect 13954 1996 14016 2005
rect 13454 1958 13820 1962
rect 13902 1958 13968 1966
rect 13454 1930 13862 1958
rect 13454 1892 13482 1930
rect 13776 1911 13862 1930
rect 13454 1884 13520 1892
rect 13454 1850 13469 1884
rect 13503 1850 13520 1884
rect 13454 1838 13520 1850
rect 13626 1888 13694 1894
rect 13626 1836 13636 1888
rect 13688 1836 13694 1888
rect 13626 1830 13694 1836
rect 13776 1877 13822 1911
rect 13856 1877 13862 1911
rect 13902 1906 13908 1958
rect 13960 1906 13968 1958
rect 13902 1898 13918 1906
rect 13776 1839 13862 1877
rect 13776 1805 13822 1839
rect 13856 1805 13862 1839
rect 13536 1776 13604 1782
rect 13536 1724 13544 1776
rect 13596 1724 13604 1776
rect 13536 1714 13604 1724
rect 13776 1758 13862 1805
rect 13912 1877 13918 1898
rect 13952 1898 13968 1906
rect 14008 1926 14336 1958
rect 14008 1911 14104 1926
rect 13952 1877 13958 1898
rect 13912 1839 13958 1877
rect 13912 1805 13918 1839
rect 13952 1805 13958 1839
rect 13912 1758 13958 1805
rect 14008 1877 14014 1911
rect 14048 1877 14104 1911
rect 14308 1890 14336 1926
rect 14008 1839 14104 1877
rect 14008 1805 14014 1839
rect 14048 1805 14104 1839
rect 14266 1882 14336 1890
rect 14266 1848 14281 1882
rect 14315 1848 14336 1882
rect 14266 1830 14336 1848
rect 14442 1890 14506 1896
rect 14442 1838 14448 1890
rect 14500 1838 14506 1890
rect 14442 1832 14506 1838
rect 14008 1758 14104 1805
rect 13434 1643 13710 1674
rect 13434 1609 13463 1643
rect 13497 1609 13555 1643
rect 13589 1609 13647 1643
rect 13681 1609 13710 1643
rect 13434 1578 13710 1609
rect 13776 1558 13826 1758
rect 13858 1711 13916 1726
rect 13858 1677 13870 1711
rect 13904 1677 13916 1711
rect 13858 1660 13916 1677
rect 13970 1630 14028 1648
rect 13970 1596 13982 1630
rect 14016 1596 14028 1630
rect 13970 1586 14028 1596
rect 14058 1558 14104 1758
rect 14354 1774 14418 1780
rect 14354 1722 14360 1774
rect 14412 1722 14418 1774
rect 14354 1716 14418 1722
rect 14248 1643 14524 1674
rect 14248 1609 14277 1643
rect 14311 1609 14369 1643
rect 14403 1609 14461 1643
rect 14495 1609 14524 1643
rect 14248 1606 14524 1609
rect 13416 1541 13480 1548
rect 13416 1508 13422 1541
rect 13474 1508 13480 1541
rect 13592 1541 13656 1548
rect 13592 1508 13598 1541
rect 13474 1489 13598 1508
rect 13650 1489 13656 1541
rect 13422 1480 13656 1489
rect 13776 1546 13878 1558
rect 13776 1512 13838 1546
rect 13872 1512 13878 1546
rect 13776 1474 13878 1512
rect 13928 1546 13974 1558
rect 13928 1512 13934 1546
rect 13968 1512 13974 1546
rect 13928 1492 13974 1512
rect 14024 1546 14104 1558
rect 14024 1512 14030 1546
rect 14064 1512 14104 1546
rect 13776 1442 13838 1474
rect 13572 1440 13838 1442
rect 13872 1440 13878 1474
rect 13572 1428 13878 1440
rect 13918 1486 13984 1492
rect 13918 1434 13926 1486
rect 13978 1434 13984 1486
rect 13918 1428 13984 1434
rect 14024 1474 14104 1512
rect 14024 1440 14030 1474
rect 14064 1440 14104 1474
rect 14220 1578 14524 1606
rect 14024 1428 14070 1440
rect 13572 1414 13826 1428
rect 13416 1408 13482 1414
rect 13416 1356 13424 1408
rect 13476 1356 13482 1408
rect 13416 1350 13482 1356
rect 12564 1141 12594 1144
rect 12646 1141 13188 1144
rect 12564 1107 12593 1141
rect 12646 1107 12685 1141
rect 12719 1107 12777 1141
rect 12811 1139 13188 1141
rect 12811 1107 12939 1139
rect 12564 1092 12594 1107
rect 12646 1105 12939 1107
rect 12973 1105 13031 1139
rect 13065 1105 13123 1139
rect 13157 1105 13188 1139
rect 12646 1092 13188 1105
rect 12564 1074 13188 1092
rect 13256 1150 13532 1164
rect 13256 1133 13448 1150
rect 13500 1133 13532 1150
rect 13256 1099 13285 1133
rect 13319 1099 13377 1133
rect 13411 1099 13448 1133
rect 13503 1099 13532 1133
rect 13256 1098 13448 1099
rect 13500 1098 13532 1099
rect 13256 1068 13532 1098
rect 13572 1064 13600 1414
rect 13872 1390 13936 1400
rect 13872 1356 13886 1390
rect 13920 1356 14192 1390
rect 13872 1338 13936 1356
rect 13788 1292 13860 1304
rect 13788 1240 13798 1292
rect 13850 1240 13860 1292
rect 13788 1228 13860 1240
rect 14158 1174 14192 1356
rect 14220 1274 14248 1578
rect 14220 1264 14288 1274
rect 14220 1230 14236 1264
rect 14270 1230 14288 1264
rect 14220 1216 14288 1230
rect 13632 1146 14192 1174
rect 13632 1143 13698 1146
rect 13632 1109 13648 1143
rect 13682 1109 13698 1143
rect 13632 1100 13698 1109
rect 13866 1091 13956 1112
rect 12064 983 12304 1000
rect 12348 1056 12414 1062
rect 12348 1004 12356 1056
rect 12408 1004 12414 1056
rect 12348 998 12362 1004
rect 11798 943 11844 976
rect 11798 909 11804 943
rect 11838 909 11844 943
rect 12064 949 12076 983
rect 12110 972 12304 983
rect 12356 981 12362 998
rect 12396 998 12414 1004
rect 12444 1015 12490 1062
rect 13572 1036 13644 1064
rect 12396 981 12402 998
rect 12110 949 12302 972
rect 12064 940 12302 949
rect 11798 862 11844 909
rect 12012 902 12078 910
rect 11926 898 11972 902
rect 11042 840 11114 844
rect 10502 815 10568 828
rect 10502 781 10518 815
rect 10552 781 10568 815
rect 10502 772 10568 781
rect 11042 788 11051 840
rect 11103 788 11114 840
rect 11042 776 11114 788
rect 11238 838 11312 858
rect 11886 855 11972 898
rect 11238 804 11250 838
rect 11284 804 11312 838
rect 11238 780 11312 804
rect 11348 844 11416 850
rect 11348 792 11355 844
rect 11407 838 11416 844
rect 11407 832 11500 838
rect 11407 798 11446 832
rect 11480 798 11500 832
rect 11407 792 11500 798
rect 11348 788 11500 792
rect 11744 815 11810 826
rect 11348 786 11416 788
rect 11744 781 11760 815
rect 11794 781 11810 815
rect 11744 768 11810 781
rect 11886 821 11932 855
rect 11966 821 11972 855
rect 12012 850 12018 902
rect 12070 850 12078 902
rect 12012 842 12028 850
rect 11886 783 11972 821
rect 11886 749 11932 783
rect 11966 749 11972 783
rect 10824 728 10882 742
rect 10824 708 10836 728
rect 10354 694 10836 708
rect 10870 694 10882 728
rect 10354 674 10882 694
rect 11886 702 11972 749
rect 12022 821 12028 842
rect 12062 842 12078 850
rect 12118 855 12214 902
rect 12062 821 12068 842
rect 12022 783 12068 821
rect 12022 749 12028 783
rect 12062 749 12068 783
rect 12022 702 12068 749
rect 12118 821 12124 855
rect 12158 821 12214 855
rect 12118 783 12214 821
rect 12118 749 12124 783
rect 12158 749 12214 783
rect 12118 702 12214 749
rect 10246 372 10292 384
rect 10354 344 10414 674
rect 11886 648 11936 702
rect 10460 624 10536 630
rect 10460 572 10468 624
rect 10520 572 10536 624
rect 10460 566 10536 572
rect 10676 597 11298 628
rect 10094 334 10414 344
rect 10094 300 10108 334
rect 10142 300 10414 334
rect 10094 282 10414 300
rect 10676 563 10705 597
rect 10739 563 10797 597
rect 10831 563 10889 597
rect 10923 595 11298 597
rect 10923 563 11051 595
rect 10676 561 11051 563
rect 11085 561 11143 595
rect 11177 561 11235 595
rect 11269 561 11298 595
rect 10676 530 11298 561
rect 11368 602 11644 620
rect 11368 589 11491 602
rect 11543 589 11644 602
rect 11720 598 11778 606
rect 11368 555 11397 589
rect 11431 555 11489 589
rect 11543 555 11581 589
rect 11615 555 11644 589
rect 11368 550 11491 555
rect 11543 550 11644 555
rect 10676 254 10774 530
rect 11368 524 11644 550
rect 11712 592 11786 598
rect 11712 540 11723 592
rect 11775 540 11786 592
rect 11866 582 11936 648
rect 11968 655 12026 670
rect 11968 621 11980 655
rect 12014 621 12026 655
rect 11968 604 12026 621
rect 11712 534 11786 540
rect 11720 528 11778 534
rect 11436 254 11520 524
rect 11886 502 11936 582
rect 12080 574 12138 592
rect 12080 540 12092 574
rect 12126 540 12138 574
rect 12080 530 12138 540
rect 12168 502 12214 702
rect 11886 490 11988 502
rect 11886 456 11948 490
rect 11982 456 11988 490
rect 11886 418 11988 456
rect 12038 490 12084 502
rect 12038 456 12044 490
rect 12078 456 12084 490
rect 12038 436 12084 456
rect 12134 490 12214 502
rect 12134 456 12140 490
rect 12174 456 12214 490
rect 11886 384 11948 418
rect 11982 384 11988 418
rect 11886 372 11988 384
rect 12028 430 12094 436
rect 12028 378 12036 430
rect 12088 378 12094 430
rect 12028 372 12094 378
rect 12134 418 12214 456
rect 12134 384 12140 418
rect 12174 384 12214 418
rect 12242 708 12302 940
rect 12356 943 12402 981
rect 12356 909 12362 943
rect 12396 909 12402 943
rect 12356 862 12402 909
rect 12444 981 12450 1015
rect 12484 981 12490 1015
rect 12444 943 12490 981
rect 12444 909 12450 943
rect 12484 909 12490 943
rect 12444 862 12490 909
rect 13598 1015 13644 1036
rect 13598 981 13604 1015
rect 13638 981 13644 1015
rect 13598 943 13644 981
rect 13598 909 13604 943
rect 13638 909 13644 943
rect 13598 862 13644 909
rect 13686 1042 13732 1062
rect 13866 1057 13895 1091
rect 13929 1057 13956 1091
rect 13686 1036 13754 1042
rect 13866 1036 13956 1057
rect 13686 1015 13694 1036
rect 13686 981 13692 1015
rect 13746 984 13754 1036
rect 13726 981 13754 984
rect 13686 976 13754 981
rect 13952 1000 14010 1002
rect 14158 1000 14192 1146
rect 14278 1143 14344 1154
rect 14278 1109 14294 1143
rect 14328 1109 14344 1143
rect 14278 1098 14344 1109
rect 14452 1144 15076 1176
rect 15158 1164 15236 2122
rect 15750 2113 15779 2122
rect 15813 2122 17667 2147
rect 15813 2113 15840 2122
rect 15750 2092 15840 2113
rect 15836 2056 15894 2058
rect 15836 2039 15898 2056
rect 15836 2005 15848 2039
rect 15882 2005 15898 2039
rect 15836 1996 15898 2005
rect 15336 1958 15702 1962
rect 15784 1958 15850 1966
rect 15336 1930 15744 1958
rect 15336 1892 15364 1930
rect 15658 1911 15744 1930
rect 15336 1884 15402 1892
rect 15336 1850 15351 1884
rect 15385 1850 15402 1884
rect 15336 1838 15402 1850
rect 15508 1888 15576 1894
rect 15508 1836 15518 1888
rect 15570 1836 15576 1888
rect 15508 1830 15576 1836
rect 15658 1877 15704 1911
rect 15738 1877 15744 1911
rect 15784 1906 15790 1958
rect 15842 1906 15850 1958
rect 15784 1898 15800 1906
rect 15658 1839 15744 1877
rect 15658 1805 15704 1839
rect 15738 1805 15744 1839
rect 15418 1776 15486 1782
rect 15418 1724 15426 1776
rect 15478 1724 15486 1776
rect 15418 1714 15486 1724
rect 15658 1758 15744 1805
rect 15794 1877 15800 1898
rect 15834 1898 15850 1906
rect 15890 1926 16218 1958
rect 15890 1911 15986 1926
rect 15834 1877 15840 1898
rect 15794 1839 15840 1877
rect 15794 1805 15800 1839
rect 15834 1805 15840 1839
rect 15794 1758 15840 1805
rect 15890 1877 15896 1911
rect 15930 1877 15986 1911
rect 16190 1890 16218 1926
rect 15890 1839 15986 1877
rect 15890 1805 15896 1839
rect 15930 1805 15986 1839
rect 16148 1882 16218 1890
rect 16148 1848 16163 1882
rect 16197 1848 16218 1882
rect 16148 1830 16218 1848
rect 16324 1890 16388 1896
rect 16324 1838 16330 1890
rect 16382 1838 16388 1890
rect 16324 1832 16388 1838
rect 15890 1758 15986 1805
rect 15316 1643 15592 1674
rect 15316 1609 15345 1643
rect 15379 1609 15437 1643
rect 15471 1609 15529 1643
rect 15563 1609 15592 1643
rect 15316 1578 15592 1609
rect 15658 1558 15708 1758
rect 15740 1711 15798 1726
rect 15740 1677 15752 1711
rect 15786 1677 15798 1711
rect 15740 1660 15798 1677
rect 15852 1630 15910 1648
rect 15852 1596 15864 1630
rect 15898 1596 15910 1630
rect 15852 1586 15910 1596
rect 15940 1558 15986 1758
rect 16236 1774 16300 1780
rect 16236 1722 16242 1774
rect 16294 1722 16300 1774
rect 16236 1716 16300 1722
rect 16130 1643 16406 1674
rect 16130 1609 16159 1643
rect 16193 1609 16251 1643
rect 16285 1609 16343 1643
rect 16377 1609 16406 1643
rect 16130 1606 16406 1609
rect 15298 1541 15362 1548
rect 15298 1508 15304 1541
rect 15356 1508 15362 1541
rect 15474 1541 15538 1548
rect 15474 1508 15480 1541
rect 15356 1489 15480 1508
rect 15532 1489 15538 1541
rect 15304 1480 15538 1489
rect 15658 1546 15760 1558
rect 15658 1512 15720 1546
rect 15754 1512 15760 1546
rect 15658 1474 15760 1512
rect 15810 1546 15856 1558
rect 15810 1512 15816 1546
rect 15850 1512 15856 1546
rect 15810 1492 15856 1512
rect 15906 1546 15986 1558
rect 15906 1512 15912 1546
rect 15946 1512 15986 1546
rect 15658 1442 15720 1474
rect 15454 1440 15720 1442
rect 15754 1440 15760 1474
rect 15454 1428 15760 1440
rect 15800 1486 15866 1492
rect 15800 1434 15808 1486
rect 15860 1434 15866 1486
rect 15800 1428 15866 1434
rect 15906 1474 15986 1512
rect 15906 1440 15912 1474
rect 15946 1440 15986 1474
rect 16102 1578 16406 1606
rect 15906 1428 15952 1440
rect 15454 1414 15708 1428
rect 15298 1408 15364 1414
rect 15298 1356 15306 1408
rect 15358 1356 15364 1408
rect 15298 1350 15364 1356
rect 14452 1141 14482 1144
rect 14534 1141 15076 1144
rect 14452 1107 14481 1141
rect 14534 1107 14573 1141
rect 14607 1107 14665 1141
rect 14699 1139 15076 1141
rect 14699 1107 14827 1139
rect 14452 1092 14482 1107
rect 14534 1105 14827 1107
rect 14861 1105 14919 1139
rect 14953 1105 15011 1139
rect 15045 1105 15076 1139
rect 14534 1092 15076 1105
rect 14452 1074 15076 1092
rect 15138 1150 15414 1164
rect 15138 1133 15330 1150
rect 15382 1133 15414 1150
rect 15138 1099 15167 1133
rect 15201 1099 15259 1133
rect 15293 1099 15330 1133
rect 15385 1099 15414 1133
rect 15138 1098 15330 1099
rect 15382 1098 15414 1099
rect 15138 1068 15414 1098
rect 15454 1064 15482 1414
rect 15754 1390 15818 1400
rect 15754 1356 15768 1390
rect 15802 1356 16074 1390
rect 15754 1338 15818 1356
rect 15670 1292 15742 1304
rect 15670 1240 15680 1292
rect 15732 1240 15742 1292
rect 15670 1228 15742 1240
rect 16040 1174 16074 1356
rect 16102 1274 16130 1578
rect 16102 1264 16170 1274
rect 16102 1230 16118 1264
rect 16152 1230 16170 1264
rect 16102 1216 16170 1230
rect 15514 1146 16074 1174
rect 15514 1143 15580 1146
rect 15514 1109 15530 1143
rect 15564 1109 15580 1143
rect 15514 1100 15580 1109
rect 15748 1091 15838 1112
rect 13952 983 14192 1000
rect 14236 1056 14302 1062
rect 14236 1004 14244 1056
rect 14296 1004 14302 1056
rect 14236 998 14250 1004
rect 13686 943 13732 976
rect 13686 909 13692 943
rect 13726 909 13732 943
rect 13952 949 13964 983
rect 13998 972 14192 983
rect 14244 981 14250 998
rect 14284 998 14302 1004
rect 14332 1015 14378 1062
rect 15454 1036 15526 1064
rect 14284 981 14290 998
rect 13998 949 14190 972
rect 13952 940 14190 949
rect 13686 862 13732 909
rect 13900 902 13966 910
rect 13814 898 13860 902
rect 12930 840 13002 844
rect 12390 815 12456 828
rect 12390 781 12406 815
rect 12440 781 12456 815
rect 12390 772 12456 781
rect 12930 788 12939 840
rect 12991 788 13002 840
rect 12930 776 13002 788
rect 13126 838 13200 858
rect 13774 855 13860 898
rect 13126 804 13138 838
rect 13172 804 13200 838
rect 13126 780 13200 804
rect 13236 844 13304 850
rect 13236 792 13243 844
rect 13295 838 13304 844
rect 13295 832 13388 838
rect 13295 798 13334 832
rect 13368 798 13388 832
rect 13295 792 13388 798
rect 13236 788 13388 792
rect 13632 815 13698 826
rect 13236 786 13304 788
rect 13632 781 13648 815
rect 13682 781 13698 815
rect 13632 768 13698 781
rect 13774 821 13820 855
rect 13854 821 13860 855
rect 13900 850 13906 902
rect 13958 850 13966 902
rect 13900 842 13916 850
rect 13774 783 13860 821
rect 13774 749 13820 783
rect 13854 749 13860 783
rect 12712 728 12770 742
rect 12712 708 12724 728
rect 12242 694 12724 708
rect 12758 694 12770 728
rect 12242 674 12770 694
rect 13774 702 13860 749
rect 13910 821 13916 842
rect 13950 842 13966 850
rect 14006 855 14102 902
rect 13950 821 13956 842
rect 13910 783 13956 821
rect 13910 749 13916 783
rect 13950 749 13956 783
rect 13910 702 13956 749
rect 14006 821 14012 855
rect 14046 821 14102 855
rect 14006 783 14102 821
rect 14006 749 14012 783
rect 14046 749 14102 783
rect 14006 702 14102 749
rect 12134 372 12180 384
rect 12242 344 12302 674
rect 13774 648 13824 702
rect 12348 624 12424 630
rect 12348 572 12356 624
rect 12408 572 12424 624
rect 12348 566 12424 572
rect 12564 597 13186 628
rect 11982 334 12302 344
rect 11982 300 11996 334
rect 12030 300 12302 334
rect 11982 282 12302 300
rect 12564 563 12593 597
rect 12627 563 12685 597
rect 12719 563 12777 597
rect 12811 595 13186 597
rect 12811 563 12939 595
rect 12564 561 12939 563
rect 12973 561 13031 595
rect 13065 561 13123 595
rect 13157 561 13186 595
rect 12564 530 13186 561
rect 13256 602 13532 620
rect 13256 589 13379 602
rect 13431 589 13532 602
rect 13608 598 13666 606
rect 13256 555 13285 589
rect 13319 555 13377 589
rect 13431 555 13469 589
rect 13503 555 13532 589
rect 13256 550 13379 555
rect 13431 550 13532 555
rect 12564 254 12662 530
rect 13256 524 13532 550
rect 13600 592 13674 598
rect 13600 540 13611 592
rect 13663 540 13674 592
rect 13754 582 13824 648
rect 13856 655 13914 670
rect 13856 621 13868 655
rect 13902 621 13914 655
rect 13856 604 13914 621
rect 13600 534 13674 540
rect 13608 528 13666 534
rect 13324 254 13408 524
rect 13774 502 13824 582
rect 13968 574 14026 592
rect 13968 540 13980 574
rect 14014 540 14026 574
rect 13968 530 14026 540
rect 14056 502 14102 702
rect 13774 490 13876 502
rect 13774 456 13836 490
rect 13870 456 13876 490
rect 13774 418 13876 456
rect 13926 490 13972 502
rect 13926 456 13932 490
rect 13966 456 13972 490
rect 13926 436 13972 456
rect 14022 490 14102 502
rect 14022 456 14028 490
rect 14062 456 14102 490
rect 13774 384 13836 418
rect 13870 384 13876 418
rect 13774 372 13876 384
rect 13916 430 13982 436
rect 13916 378 13924 430
rect 13976 378 13982 430
rect 13916 372 13982 378
rect 14022 418 14102 456
rect 14022 384 14028 418
rect 14062 384 14102 418
rect 14130 708 14190 940
rect 14244 943 14290 981
rect 14244 909 14250 943
rect 14284 909 14290 943
rect 14244 862 14290 909
rect 14332 981 14338 1015
rect 14372 981 14378 1015
rect 14332 943 14378 981
rect 14332 909 14338 943
rect 14372 909 14378 943
rect 14332 862 14378 909
rect 15480 1015 15526 1036
rect 15480 981 15486 1015
rect 15520 981 15526 1015
rect 15480 943 15526 981
rect 15480 909 15486 943
rect 15520 909 15526 943
rect 15480 862 15526 909
rect 15568 1042 15614 1062
rect 15748 1057 15777 1091
rect 15811 1057 15838 1091
rect 15568 1036 15636 1042
rect 15748 1036 15838 1057
rect 15568 1015 15576 1036
rect 15568 981 15574 1015
rect 15628 984 15636 1036
rect 15608 981 15636 984
rect 15568 976 15636 981
rect 15834 1000 15892 1002
rect 16040 1000 16074 1146
rect 16160 1143 16226 1154
rect 16160 1109 16176 1143
rect 16210 1109 16226 1143
rect 16160 1098 16226 1109
rect 16334 1144 16958 1176
rect 17046 1164 17124 2122
rect 17638 2113 17667 2122
rect 17701 2122 19555 2147
rect 17701 2113 17728 2122
rect 17638 2092 17728 2113
rect 17724 2056 17782 2058
rect 17724 2039 17786 2056
rect 17724 2005 17736 2039
rect 17770 2005 17786 2039
rect 17724 1996 17786 2005
rect 17224 1958 17590 1962
rect 17672 1958 17738 1966
rect 17224 1930 17632 1958
rect 17224 1892 17252 1930
rect 17546 1911 17632 1930
rect 17224 1884 17290 1892
rect 17224 1850 17239 1884
rect 17273 1850 17290 1884
rect 17224 1838 17290 1850
rect 17396 1888 17464 1894
rect 17396 1836 17406 1888
rect 17458 1836 17464 1888
rect 17396 1830 17464 1836
rect 17546 1877 17592 1911
rect 17626 1877 17632 1911
rect 17672 1906 17678 1958
rect 17730 1906 17738 1958
rect 17672 1898 17688 1906
rect 17546 1839 17632 1877
rect 17546 1805 17592 1839
rect 17626 1805 17632 1839
rect 17306 1776 17374 1782
rect 17306 1724 17314 1776
rect 17366 1724 17374 1776
rect 17306 1714 17374 1724
rect 17546 1758 17632 1805
rect 17682 1877 17688 1898
rect 17722 1898 17738 1906
rect 17778 1926 18106 1958
rect 17778 1911 17874 1926
rect 17722 1877 17728 1898
rect 17682 1839 17728 1877
rect 17682 1805 17688 1839
rect 17722 1805 17728 1839
rect 17682 1758 17728 1805
rect 17778 1877 17784 1911
rect 17818 1877 17874 1911
rect 18078 1890 18106 1926
rect 17778 1839 17874 1877
rect 17778 1805 17784 1839
rect 17818 1805 17874 1839
rect 18036 1882 18106 1890
rect 18036 1848 18051 1882
rect 18085 1848 18106 1882
rect 18036 1830 18106 1848
rect 18212 1890 18276 1896
rect 18212 1838 18218 1890
rect 18270 1838 18276 1890
rect 18212 1832 18276 1838
rect 17778 1758 17874 1805
rect 17204 1643 17480 1674
rect 17204 1609 17233 1643
rect 17267 1609 17325 1643
rect 17359 1609 17417 1643
rect 17451 1609 17480 1643
rect 17204 1578 17480 1609
rect 17546 1558 17596 1758
rect 17628 1711 17686 1726
rect 17628 1677 17640 1711
rect 17674 1677 17686 1711
rect 17628 1660 17686 1677
rect 17740 1630 17798 1648
rect 17740 1596 17752 1630
rect 17786 1596 17798 1630
rect 17740 1586 17798 1596
rect 17828 1558 17874 1758
rect 18124 1774 18188 1780
rect 18124 1722 18130 1774
rect 18182 1722 18188 1774
rect 18124 1716 18188 1722
rect 18018 1643 18294 1674
rect 18018 1609 18047 1643
rect 18081 1609 18139 1643
rect 18173 1609 18231 1643
rect 18265 1609 18294 1643
rect 18018 1606 18294 1609
rect 17186 1541 17250 1548
rect 17186 1508 17192 1541
rect 17244 1508 17250 1541
rect 17362 1541 17426 1548
rect 17362 1508 17368 1541
rect 17244 1489 17368 1508
rect 17420 1489 17426 1541
rect 17192 1480 17426 1489
rect 17546 1546 17648 1558
rect 17546 1512 17608 1546
rect 17642 1512 17648 1546
rect 17546 1474 17648 1512
rect 17698 1546 17744 1558
rect 17698 1512 17704 1546
rect 17738 1512 17744 1546
rect 17698 1492 17744 1512
rect 17794 1546 17874 1558
rect 17794 1512 17800 1546
rect 17834 1512 17874 1546
rect 17546 1442 17608 1474
rect 17342 1440 17608 1442
rect 17642 1440 17648 1474
rect 17342 1428 17648 1440
rect 17688 1486 17754 1492
rect 17688 1434 17696 1486
rect 17748 1434 17754 1486
rect 17688 1428 17754 1434
rect 17794 1474 17874 1512
rect 17794 1440 17800 1474
rect 17834 1440 17874 1474
rect 17990 1578 18294 1606
rect 17794 1428 17840 1440
rect 17342 1414 17596 1428
rect 17186 1408 17252 1414
rect 17186 1356 17194 1408
rect 17246 1356 17252 1408
rect 17186 1350 17252 1356
rect 16334 1141 16364 1144
rect 16416 1141 16958 1144
rect 16334 1107 16363 1141
rect 16416 1107 16455 1141
rect 16489 1107 16547 1141
rect 16581 1139 16958 1141
rect 16581 1107 16709 1139
rect 16334 1092 16364 1107
rect 16416 1105 16709 1107
rect 16743 1105 16801 1139
rect 16835 1105 16893 1139
rect 16927 1105 16958 1139
rect 16416 1092 16958 1105
rect 16334 1074 16958 1092
rect 17026 1150 17302 1164
rect 17026 1133 17218 1150
rect 17270 1133 17302 1150
rect 17026 1099 17055 1133
rect 17089 1099 17147 1133
rect 17181 1099 17218 1133
rect 17273 1099 17302 1133
rect 17026 1098 17218 1099
rect 17270 1098 17302 1099
rect 17026 1068 17302 1098
rect 17342 1064 17370 1414
rect 17642 1390 17706 1400
rect 17642 1356 17656 1390
rect 17690 1356 17962 1390
rect 17642 1338 17706 1356
rect 17558 1292 17630 1304
rect 17558 1240 17568 1292
rect 17620 1240 17630 1292
rect 17558 1228 17630 1240
rect 17928 1174 17962 1356
rect 17990 1274 18018 1578
rect 17990 1264 18058 1274
rect 17990 1230 18006 1264
rect 18040 1230 18058 1264
rect 17990 1216 18058 1230
rect 17402 1146 17962 1174
rect 17402 1143 17468 1146
rect 17402 1109 17418 1143
rect 17452 1109 17468 1143
rect 17402 1100 17468 1109
rect 17636 1091 17726 1112
rect 15834 983 16074 1000
rect 16118 1056 16184 1062
rect 16118 1004 16126 1056
rect 16178 1004 16184 1056
rect 16118 998 16132 1004
rect 15568 943 15614 976
rect 15568 909 15574 943
rect 15608 909 15614 943
rect 15834 949 15846 983
rect 15880 972 16074 983
rect 16126 981 16132 998
rect 16166 998 16184 1004
rect 16214 1015 16260 1062
rect 17342 1036 17414 1064
rect 16166 981 16172 998
rect 15880 949 16072 972
rect 15834 940 16072 949
rect 15568 862 15614 909
rect 15782 902 15848 910
rect 15696 898 15742 902
rect 14818 840 14890 844
rect 14278 815 14344 828
rect 14278 781 14294 815
rect 14328 781 14344 815
rect 14278 772 14344 781
rect 14818 788 14827 840
rect 14879 788 14890 840
rect 14818 776 14890 788
rect 15014 838 15088 858
rect 15656 855 15742 898
rect 15014 804 15026 838
rect 15060 804 15088 838
rect 15014 780 15088 804
rect 15118 844 15186 850
rect 15118 792 15125 844
rect 15177 838 15186 844
rect 15177 832 15270 838
rect 15177 798 15216 832
rect 15250 798 15270 832
rect 15177 792 15270 798
rect 15118 788 15270 792
rect 15514 815 15580 826
rect 15118 786 15186 788
rect 15514 781 15530 815
rect 15564 781 15580 815
rect 15514 768 15580 781
rect 15656 821 15702 855
rect 15736 821 15742 855
rect 15782 850 15788 902
rect 15840 850 15848 902
rect 15782 842 15798 850
rect 15656 783 15742 821
rect 15656 749 15702 783
rect 15736 749 15742 783
rect 14600 728 14658 742
rect 14600 708 14612 728
rect 14130 694 14612 708
rect 14646 694 14658 728
rect 14130 674 14658 694
rect 15656 702 15742 749
rect 15792 821 15798 842
rect 15832 842 15848 850
rect 15888 855 15984 902
rect 15832 821 15838 842
rect 15792 783 15838 821
rect 15792 749 15798 783
rect 15832 749 15838 783
rect 15792 702 15838 749
rect 15888 821 15894 855
rect 15928 821 15984 855
rect 15888 783 15984 821
rect 15888 749 15894 783
rect 15928 749 15984 783
rect 15888 702 15984 749
rect 14022 372 14068 384
rect 14130 344 14190 674
rect 15656 648 15706 702
rect 14236 624 14312 630
rect 14236 572 14244 624
rect 14296 572 14312 624
rect 14236 566 14312 572
rect 14452 597 15074 628
rect 13870 334 14190 344
rect 13870 300 13884 334
rect 13918 300 14190 334
rect 13870 282 14190 300
rect 14452 563 14481 597
rect 14515 563 14573 597
rect 14607 563 14665 597
rect 14699 595 15074 597
rect 14699 563 14827 595
rect 14452 561 14827 563
rect 14861 561 14919 595
rect 14953 561 15011 595
rect 15045 561 15074 595
rect 14452 530 15074 561
rect 15138 602 15414 620
rect 15138 589 15261 602
rect 15313 589 15414 602
rect 15490 598 15548 606
rect 15138 555 15167 589
rect 15201 555 15259 589
rect 15313 555 15351 589
rect 15385 555 15414 589
rect 15138 550 15261 555
rect 15313 550 15414 555
rect 14452 254 14550 530
rect 15138 524 15414 550
rect 15482 592 15556 598
rect 15482 540 15493 592
rect 15545 540 15556 592
rect 15636 582 15706 648
rect 15738 655 15796 670
rect 15738 621 15750 655
rect 15784 621 15796 655
rect 15738 604 15796 621
rect 15482 534 15556 540
rect 15490 528 15548 534
rect 15206 254 15290 524
rect 15656 502 15706 582
rect 15850 574 15908 592
rect 15850 540 15862 574
rect 15896 540 15908 574
rect 15850 530 15908 540
rect 15938 502 15984 702
rect 15656 490 15758 502
rect 15656 456 15718 490
rect 15752 456 15758 490
rect 15656 418 15758 456
rect 15808 490 15854 502
rect 15808 456 15814 490
rect 15848 456 15854 490
rect 15808 436 15854 456
rect 15904 490 15984 502
rect 15904 456 15910 490
rect 15944 456 15984 490
rect 15656 384 15718 418
rect 15752 384 15758 418
rect 15656 372 15758 384
rect 15798 430 15864 436
rect 15798 378 15806 430
rect 15858 378 15864 430
rect 15798 372 15864 378
rect 15904 418 15984 456
rect 15904 384 15910 418
rect 15944 384 15984 418
rect 16012 708 16072 940
rect 16126 943 16172 981
rect 16126 909 16132 943
rect 16166 909 16172 943
rect 16126 862 16172 909
rect 16214 981 16220 1015
rect 16254 981 16260 1015
rect 16214 943 16260 981
rect 16214 909 16220 943
rect 16254 909 16260 943
rect 16214 862 16260 909
rect 17368 1015 17414 1036
rect 17368 981 17374 1015
rect 17408 981 17414 1015
rect 17368 943 17414 981
rect 17368 909 17374 943
rect 17408 909 17414 943
rect 17368 862 17414 909
rect 17456 1042 17502 1062
rect 17636 1057 17665 1091
rect 17699 1057 17726 1091
rect 17456 1036 17524 1042
rect 17636 1036 17726 1057
rect 17456 1015 17464 1036
rect 17456 981 17462 1015
rect 17516 984 17524 1036
rect 17496 981 17524 984
rect 17456 976 17524 981
rect 17722 1000 17780 1002
rect 17928 1000 17962 1146
rect 18048 1143 18114 1154
rect 18048 1109 18064 1143
rect 18098 1109 18114 1143
rect 18048 1098 18114 1109
rect 18222 1144 18846 1176
rect 18934 1164 19012 2122
rect 19526 2113 19555 2122
rect 19589 2122 21443 2147
rect 19589 2113 19616 2122
rect 19526 2092 19616 2113
rect 19612 2056 19670 2058
rect 19612 2039 19674 2056
rect 19612 2005 19624 2039
rect 19658 2005 19674 2039
rect 19612 1996 19674 2005
rect 19112 1958 19478 1962
rect 19560 1958 19626 1966
rect 19112 1930 19520 1958
rect 19112 1892 19140 1930
rect 19434 1911 19520 1930
rect 19112 1884 19178 1892
rect 19112 1850 19127 1884
rect 19161 1850 19178 1884
rect 19112 1838 19178 1850
rect 19284 1888 19352 1894
rect 19284 1836 19294 1888
rect 19346 1836 19352 1888
rect 19284 1830 19352 1836
rect 19434 1877 19480 1911
rect 19514 1877 19520 1911
rect 19560 1906 19566 1958
rect 19618 1906 19626 1958
rect 19560 1898 19576 1906
rect 19434 1839 19520 1877
rect 19434 1805 19480 1839
rect 19514 1805 19520 1839
rect 19194 1776 19262 1782
rect 19194 1724 19202 1776
rect 19254 1724 19262 1776
rect 19194 1714 19262 1724
rect 19434 1758 19520 1805
rect 19570 1877 19576 1898
rect 19610 1898 19626 1906
rect 19666 1926 19994 1958
rect 19666 1911 19762 1926
rect 19610 1877 19616 1898
rect 19570 1839 19616 1877
rect 19570 1805 19576 1839
rect 19610 1805 19616 1839
rect 19570 1758 19616 1805
rect 19666 1877 19672 1911
rect 19706 1877 19762 1911
rect 19966 1890 19994 1926
rect 19666 1839 19762 1877
rect 19666 1805 19672 1839
rect 19706 1805 19762 1839
rect 19924 1882 19994 1890
rect 19924 1848 19939 1882
rect 19973 1848 19994 1882
rect 19924 1830 19994 1848
rect 20100 1890 20164 1896
rect 20100 1838 20106 1890
rect 20158 1838 20164 1890
rect 20100 1832 20164 1838
rect 19666 1758 19762 1805
rect 19092 1643 19368 1674
rect 19092 1609 19121 1643
rect 19155 1609 19213 1643
rect 19247 1609 19305 1643
rect 19339 1609 19368 1643
rect 19092 1578 19368 1609
rect 19434 1558 19484 1758
rect 19516 1711 19574 1726
rect 19516 1677 19528 1711
rect 19562 1677 19574 1711
rect 19516 1660 19574 1677
rect 19628 1630 19686 1648
rect 19628 1596 19640 1630
rect 19674 1596 19686 1630
rect 19628 1586 19686 1596
rect 19716 1558 19762 1758
rect 20012 1774 20076 1780
rect 20012 1722 20018 1774
rect 20070 1722 20076 1774
rect 20012 1716 20076 1722
rect 19906 1643 20182 1674
rect 19906 1609 19935 1643
rect 19969 1609 20027 1643
rect 20061 1609 20119 1643
rect 20153 1609 20182 1643
rect 19906 1606 20182 1609
rect 19074 1541 19138 1548
rect 19074 1508 19080 1541
rect 19132 1508 19138 1541
rect 19250 1541 19314 1548
rect 19250 1508 19256 1541
rect 19132 1489 19256 1508
rect 19308 1489 19314 1541
rect 19080 1480 19314 1489
rect 19434 1546 19536 1558
rect 19434 1512 19496 1546
rect 19530 1512 19536 1546
rect 19434 1474 19536 1512
rect 19586 1546 19632 1558
rect 19586 1512 19592 1546
rect 19626 1512 19632 1546
rect 19586 1492 19632 1512
rect 19682 1546 19762 1558
rect 19682 1512 19688 1546
rect 19722 1512 19762 1546
rect 19434 1442 19496 1474
rect 19230 1440 19496 1442
rect 19530 1440 19536 1474
rect 19230 1428 19536 1440
rect 19576 1486 19642 1492
rect 19576 1434 19584 1486
rect 19636 1434 19642 1486
rect 19576 1428 19642 1434
rect 19682 1474 19762 1512
rect 19682 1440 19688 1474
rect 19722 1440 19762 1474
rect 19878 1578 20182 1606
rect 19682 1428 19728 1440
rect 19230 1414 19484 1428
rect 19074 1408 19140 1414
rect 19074 1356 19082 1408
rect 19134 1356 19140 1408
rect 19074 1350 19140 1356
rect 18222 1141 18252 1144
rect 18304 1141 18846 1144
rect 18222 1107 18251 1141
rect 18304 1107 18343 1141
rect 18377 1107 18435 1141
rect 18469 1139 18846 1141
rect 18469 1107 18597 1139
rect 18222 1092 18252 1107
rect 18304 1105 18597 1107
rect 18631 1105 18689 1139
rect 18723 1105 18781 1139
rect 18815 1105 18846 1139
rect 18304 1092 18846 1105
rect 18222 1074 18846 1092
rect 18914 1150 19190 1164
rect 18914 1133 19106 1150
rect 19158 1133 19190 1150
rect 18914 1099 18943 1133
rect 18977 1099 19035 1133
rect 19069 1099 19106 1133
rect 19161 1099 19190 1133
rect 18914 1098 19106 1099
rect 19158 1098 19190 1099
rect 18914 1068 19190 1098
rect 19230 1064 19258 1414
rect 19530 1390 19594 1400
rect 19530 1356 19544 1390
rect 19578 1356 19850 1390
rect 19530 1338 19594 1356
rect 19446 1292 19518 1304
rect 19446 1240 19456 1292
rect 19508 1240 19518 1292
rect 19446 1228 19518 1240
rect 19816 1174 19850 1356
rect 19878 1274 19906 1578
rect 19878 1264 19946 1274
rect 19878 1230 19894 1264
rect 19928 1230 19946 1264
rect 19878 1216 19946 1230
rect 19290 1146 19850 1174
rect 19290 1143 19356 1146
rect 19290 1109 19306 1143
rect 19340 1109 19356 1143
rect 19290 1100 19356 1109
rect 19524 1091 19614 1112
rect 17722 983 17962 1000
rect 18006 1056 18072 1062
rect 18006 1004 18014 1056
rect 18066 1004 18072 1056
rect 18006 998 18020 1004
rect 17456 943 17502 976
rect 17456 909 17462 943
rect 17496 909 17502 943
rect 17722 949 17734 983
rect 17768 972 17962 983
rect 18014 981 18020 998
rect 18054 998 18072 1004
rect 18102 1015 18148 1062
rect 19230 1036 19302 1064
rect 18054 981 18060 998
rect 17768 949 17960 972
rect 17722 940 17960 949
rect 17456 862 17502 909
rect 17670 902 17736 910
rect 17584 898 17630 902
rect 16700 840 16772 844
rect 16160 815 16226 828
rect 16160 781 16176 815
rect 16210 781 16226 815
rect 16160 772 16226 781
rect 16700 788 16709 840
rect 16761 788 16772 840
rect 16700 776 16772 788
rect 16896 838 16970 858
rect 17544 855 17630 898
rect 16896 804 16908 838
rect 16942 804 16970 838
rect 16896 780 16970 804
rect 17006 844 17074 850
rect 17006 792 17013 844
rect 17065 838 17074 844
rect 17065 832 17158 838
rect 17065 798 17104 832
rect 17138 798 17158 832
rect 17065 792 17158 798
rect 17006 788 17158 792
rect 17402 815 17468 826
rect 17006 786 17074 788
rect 17402 781 17418 815
rect 17452 781 17468 815
rect 17402 768 17468 781
rect 17544 821 17590 855
rect 17624 821 17630 855
rect 17670 850 17676 902
rect 17728 850 17736 902
rect 17670 842 17686 850
rect 17544 783 17630 821
rect 17544 749 17590 783
rect 17624 749 17630 783
rect 16482 728 16540 742
rect 16482 708 16494 728
rect 16012 694 16494 708
rect 16528 694 16540 728
rect 16012 674 16540 694
rect 17544 702 17630 749
rect 17680 821 17686 842
rect 17720 842 17736 850
rect 17776 855 17872 902
rect 17720 821 17726 842
rect 17680 783 17726 821
rect 17680 749 17686 783
rect 17720 749 17726 783
rect 17680 702 17726 749
rect 17776 821 17782 855
rect 17816 821 17872 855
rect 17776 783 17872 821
rect 17776 749 17782 783
rect 17816 749 17872 783
rect 17776 702 17872 749
rect 15904 372 15950 384
rect 16012 344 16072 674
rect 17544 648 17594 702
rect 16118 624 16194 630
rect 16118 572 16126 624
rect 16178 572 16194 624
rect 16118 566 16194 572
rect 16334 597 16956 628
rect 15752 334 16072 344
rect 15752 300 15766 334
rect 15800 300 16072 334
rect 15752 282 16072 300
rect 16334 563 16363 597
rect 16397 563 16455 597
rect 16489 563 16547 597
rect 16581 595 16956 597
rect 16581 563 16709 595
rect 16334 561 16709 563
rect 16743 561 16801 595
rect 16835 561 16893 595
rect 16927 561 16956 595
rect 16334 530 16956 561
rect 17026 602 17302 620
rect 17026 589 17149 602
rect 17201 589 17302 602
rect 17378 598 17436 606
rect 17026 555 17055 589
rect 17089 555 17147 589
rect 17201 555 17239 589
rect 17273 555 17302 589
rect 17026 550 17149 555
rect 17201 550 17302 555
rect 16334 254 16432 530
rect 17026 524 17302 550
rect 17370 592 17444 598
rect 17370 540 17381 592
rect 17433 540 17444 592
rect 17524 582 17594 648
rect 17626 655 17684 670
rect 17626 621 17638 655
rect 17672 621 17684 655
rect 17626 604 17684 621
rect 17370 534 17444 540
rect 17378 528 17436 534
rect 17094 254 17178 524
rect 17544 502 17594 582
rect 17738 574 17796 592
rect 17738 540 17750 574
rect 17784 540 17796 574
rect 17738 530 17796 540
rect 17826 502 17872 702
rect 17544 490 17646 502
rect 17544 456 17606 490
rect 17640 456 17646 490
rect 17544 418 17646 456
rect 17696 490 17742 502
rect 17696 456 17702 490
rect 17736 456 17742 490
rect 17696 436 17742 456
rect 17792 490 17872 502
rect 17792 456 17798 490
rect 17832 456 17872 490
rect 17544 384 17606 418
rect 17640 384 17646 418
rect 17544 372 17646 384
rect 17686 430 17752 436
rect 17686 378 17694 430
rect 17746 378 17752 430
rect 17686 372 17752 378
rect 17792 418 17872 456
rect 17792 384 17798 418
rect 17832 384 17872 418
rect 17900 708 17960 940
rect 18014 943 18060 981
rect 18014 909 18020 943
rect 18054 909 18060 943
rect 18014 862 18060 909
rect 18102 981 18108 1015
rect 18142 981 18148 1015
rect 18102 943 18148 981
rect 18102 909 18108 943
rect 18142 909 18148 943
rect 18102 862 18148 909
rect 19256 1015 19302 1036
rect 19256 981 19262 1015
rect 19296 981 19302 1015
rect 19256 943 19302 981
rect 19256 909 19262 943
rect 19296 909 19302 943
rect 19256 862 19302 909
rect 19344 1042 19390 1062
rect 19524 1057 19553 1091
rect 19587 1057 19614 1091
rect 19344 1036 19412 1042
rect 19524 1036 19614 1057
rect 19344 1015 19352 1036
rect 19344 981 19350 1015
rect 19404 984 19412 1036
rect 19384 981 19412 984
rect 19344 976 19412 981
rect 19610 1000 19668 1002
rect 19816 1000 19850 1146
rect 19936 1143 20002 1154
rect 19936 1109 19952 1143
rect 19986 1109 20002 1143
rect 19936 1098 20002 1109
rect 20110 1144 20734 1176
rect 20822 1164 20900 2122
rect 21414 2113 21443 2122
rect 21477 2122 23331 2147
rect 21477 2113 21504 2122
rect 21414 2092 21504 2113
rect 21500 2056 21558 2058
rect 21500 2039 21562 2056
rect 21500 2005 21512 2039
rect 21546 2005 21562 2039
rect 21500 1996 21562 2005
rect 21000 1958 21366 1962
rect 21448 1958 21514 1966
rect 21000 1930 21408 1958
rect 21000 1892 21028 1930
rect 21322 1911 21408 1930
rect 21000 1884 21066 1892
rect 21000 1850 21015 1884
rect 21049 1850 21066 1884
rect 21000 1838 21066 1850
rect 21172 1888 21240 1894
rect 21172 1836 21182 1888
rect 21234 1836 21240 1888
rect 21172 1830 21240 1836
rect 21322 1877 21368 1911
rect 21402 1877 21408 1911
rect 21448 1906 21454 1958
rect 21506 1906 21514 1958
rect 21448 1898 21464 1906
rect 21322 1839 21408 1877
rect 21322 1805 21368 1839
rect 21402 1805 21408 1839
rect 21082 1776 21150 1782
rect 21082 1724 21090 1776
rect 21142 1724 21150 1776
rect 21082 1714 21150 1724
rect 21322 1758 21408 1805
rect 21458 1877 21464 1898
rect 21498 1898 21514 1906
rect 21554 1926 21882 1958
rect 21554 1911 21650 1926
rect 21498 1877 21504 1898
rect 21458 1839 21504 1877
rect 21458 1805 21464 1839
rect 21498 1805 21504 1839
rect 21458 1758 21504 1805
rect 21554 1877 21560 1911
rect 21594 1877 21650 1911
rect 21854 1890 21882 1926
rect 21554 1839 21650 1877
rect 21554 1805 21560 1839
rect 21594 1805 21650 1839
rect 21812 1882 21882 1890
rect 21812 1848 21827 1882
rect 21861 1848 21882 1882
rect 21812 1830 21882 1848
rect 21988 1890 22052 1896
rect 21988 1838 21994 1890
rect 22046 1838 22052 1890
rect 21988 1832 22052 1838
rect 21554 1758 21650 1805
rect 20980 1643 21256 1674
rect 20980 1609 21009 1643
rect 21043 1609 21101 1643
rect 21135 1609 21193 1643
rect 21227 1609 21256 1643
rect 20980 1578 21256 1609
rect 21322 1558 21372 1758
rect 21404 1711 21462 1726
rect 21404 1677 21416 1711
rect 21450 1677 21462 1711
rect 21404 1660 21462 1677
rect 21516 1630 21574 1648
rect 21516 1596 21528 1630
rect 21562 1596 21574 1630
rect 21516 1586 21574 1596
rect 21604 1558 21650 1758
rect 21900 1774 21964 1780
rect 21900 1722 21906 1774
rect 21958 1722 21964 1774
rect 21900 1716 21964 1722
rect 21794 1643 22070 1674
rect 21794 1609 21823 1643
rect 21857 1609 21915 1643
rect 21949 1609 22007 1643
rect 22041 1609 22070 1643
rect 21794 1606 22070 1609
rect 20962 1541 21026 1548
rect 20962 1508 20968 1541
rect 21020 1508 21026 1541
rect 21138 1541 21202 1548
rect 21138 1508 21144 1541
rect 21020 1489 21144 1508
rect 21196 1489 21202 1541
rect 20968 1480 21202 1489
rect 21322 1546 21424 1558
rect 21322 1512 21384 1546
rect 21418 1512 21424 1546
rect 21322 1474 21424 1512
rect 21474 1546 21520 1558
rect 21474 1512 21480 1546
rect 21514 1512 21520 1546
rect 21474 1492 21520 1512
rect 21570 1546 21650 1558
rect 21570 1512 21576 1546
rect 21610 1512 21650 1546
rect 21322 1442 21384 1474
rect 21118 1440 21384 1442
rect 21418 1440 21424 1474
rect 21118 1428 21424 1440
rect 21464 1486 21530 1492
rect 21464 1434 21472 1486
rect 21524 1434 21530 1486
rect 21464 1428 21530 1434
rect 21570 1474 21650 1512
rect 21570 1440 21576 1474
rect 21610 1440 21650 1474
rect 21766 1578 22070 1606
rect 21570 1428 21616 1440
rect 21118 1414 21372 1428
rect 20962 1408 21028 1414
rect 20962 1356 20970 1408
rect 21022 1356 21028 1408
rect 20962 1350 21028 1356
rect 20110 1141 20140 1144
rect 20192 1141 20734 1144
rect 20110 1107 20139 1141
rect 20192 1107 20231 1141
rect 20265 1107 20323 1141
rect 20357 1139 20734 1141
rect 20357 1107 20485 1139
rect 20110 1092 20140 1107
rect 20192 1105 20485 1107
rect 20519 1105 20577 1139
rect 20611 1105 20669 1139
rect 20703 1105 20734 1139
rect 20192 1092 20734 1105
rect 20110 1074 20734 1092
rect 20802 1150 21078 1164
rect 20802 1133 20994 1150
rect 21046 1133 21078 1150
rect 20802 1099 20831 1133
rect 20865 1099 20923 1133
rect 20957 1099 20994 1133
rect 21049 1099 21078 1133
rect 20802 1098 20994 1099
rect 21046 1098 21078 1099
rect 20802 1068 21078 1098
rect 21118 1064 21146 1414
rect 21418 1390 21482 1400
rect 21418 1356 21432 1390
rect 21466 1356 21738 1390
rect 21418 1338 21482 1356
rect 21334 1292 21406 1304
rect 21334 1240 21344 1292
rect 21396 1240 21406 1292
rect 21334 1228 21406 1240
rect 21704 1174 21738 1356
rect 21766 1274 21794 1578
rect 21766 1264 21834 1274
rect 21766 1230 21782 1264
rect 21816 1230 21834 1264
rect 21766 1216 21834 1230
rect 21178 1146 21738 1174
rect 21178 1143 21244 1146
rect 21178 1109 21194 1143
rect 21228 1109 21244 1143
rect 21178 1100 21244 1109
rect 21412 1091 21502 1112
rect 19610 983 19850 1000
rect 19894 1056 19960 1062
rect 19894 1004 19902 1056
rect 19954 1004 19960 1056
rect 19894 998 19908 1004
rect 19344 943 19390 976
rect 19344 909 19350 943
rect 19384 909 19390 943
rect 19610 949 19622 983
rect 19656 972 19850 983
rect 19902 981 19908 998
rect 19942 998 19960 1004
rect 19990 1015 20036 1062
rect 21118 1036 21190 1064
rect 19942 981 19948 998
rect 19656 949 19848 972
rect 19610 940 19848 949
rect 19344 862 19390 909
rect 19558 902 19624 910
rect 19472 898 19518 902
rect 18588 840 18660 844
rect 18048 815 18114 828
rect 18048 781 18064 815
rect 18098 781 18114 815
rect 18048 772 18114 781
rect 18588 788 18597 840
rect 18649 788 18660 840
rect 18588 776 18660 788
rect 18784 838 18858 858
rect 19432 855 19518 898
rect 18784 804 18796 838
rect 18830 804 18858 838
rect 18784 780 18858 804
rect 18894 844 18962 850
rect 18894 792 18901 844
rect 18953 838 18962 844
rect 18953 832 19046 838
rect 18953 798 18992 832
rect 19026 798 19046 832
rect 18953 792 19046 798
rect 18894 788 19046 792
rect 19290 815 19356 826
rect 18894 786 18962 788
rect 19290 781 19306 815
rect 19340 781 19356 815
rect 19290 768 19356 781
rect 19432 821 19478 855
rect 19512 821 19518 855
rect 19558 850 19564 902
rect 19616 850 19624 902
rect 19558 842 19574 850
rect 19432 783 19518 821
rect 19432 749 19478 783
rect 19512 749 19518 783
rect 18370 728 18428 742
rect 18370 708 18382 728
rect 17900 694 18382 708
rect 18416 694 18428 728
rect 17900 674 18428 694
rect 19432 702 19518 749
rect 19568 821 19574 842
rect 19608 842 19624 850
rect 19664 855 19760 902
rect 19608 821 19614 842
rect 19568 783 19614 821
rect 19568 749 19574 783
rect 19608 749 19614 783
rect 19568 702 19614 749
rect 19664 821 19670 855
rect 19704 821 19760 855
rect 19664 783 19760 821
rect 19664 749 19670 783
rect 19704 749 19760 783
rect 19664 702 19760 749
rect 17792 372 17838 384
rect 17900 344 17960 674
rect 19432 648 19482 702
rect 18006 624 18082 630
rect 18006 572 18014 624
rect 18066 572 18082 624
rect 18006 566 18082 572
rect 18222 597 18844 628
rect 17640 334 17960 344
rect 17640 300 17654 334
rect 17688 300 17960 334
rect 17640 282 17960 300
rect 18222 563 18251 597
rect 18285 563 18343 597
rect 18377 563 18435 597
rect 18469 595 18844 597
rect 18469 563 18597 595
rect 18222 561 18597 563
rect 18631 561 18689 595
rect 18723 561 18781 595
rect 18815 561 18844 595
rect 18222 530 18844 561
rect 18914 602 19190 620
rect 18914 589 19037 602
rect 19089 589 19190 602
rect 19266 598 19324 606
rect 18914 555 18943 589
rect 18977 555 19035 589
rect 19089 555 19127 589
rect 19161 555 19190 589
rect 18914 550 19037 555
rect 19089 550 19190 555
rect 18222 254 18320 530
rect 18914 524 19190 550
rect 19258 592 19332 598
rect 19258 540 19269 592
rect 19321 540 19332 592
rect 19412 582 19482 648
rect 19514 655 19572 670
rect 19514 621 19526 655
rect 19560 621 19572 655
rect 19514 604 19572 621
rect 19258 534 19332 540
rect 19266 528 19324 534
rect 18982 254 19066 524
rect 19432 502 19482 582
rect 19626 574 19684 592
rect 19626 540 19638 574
rect 19672 540 19684 574
rect 19626 530 19684 540
rect 19714 502 19760 702
rect 19432 490 19534 502
rect 19432 456 19494 490
rect 19528 456 19534 490
rect 19432 418 19534 456
rect 19584 490 19630 502
rect 19584 456 19590 490
rect 19624 456 19630 490
rect 19584 436 19630 456
rect 19680 490 19760 502
rect 19680 456 19686 490
rect 19720 456 19760 490
rect 19432 384 19494 418
rect 19528 384 19534 418
rect 19432 372 19534 384
rect 19574 430 19640 436
rect 19574 378 19582 430
rect 19634 378 19640 430
rect 19574 372 19640 378
rect 19680 418 19760 456
rect 19680 384 19686 418
rect 19720 384 19760 418
rect 19788 708 19848 940
rect 19902 943 19948 981
rect 19902 909 19908 943
rect 19942 909 19948 943
rect 19902 862 19948 909
rect 19990 981 19996 1015
rect 20030 981 20036 1015
rect 19990 943 20036 981
rect 19990 909 19996 943
rect 20030 909 20036 943
rect 19990 862 20036 909
rect 21144 1015 21190 1036
rect 21144 981 21150 1015
rect 21184 981 21190 1015
rect 21144 943 21190 981
rect 21144 909 21150 943
rect 21184 909 21190 943
rect 21144 862 21190 909
rect 21232 1042 21278 1062
rect 21412 1057 21441 1091
rect 21475 1057 21502 1091
rect 21232 1036 21300 1042
rect 21412 1036 21502 1057
rect 21232 1015 21240 1036
rect 21232 981 21238 1015
rect 21292 984 21300 1036
rect 21272 981 21300 984
rect 21232 976 21300 981
rect 21498 1000 21556 1002
rect 21704 1000 21738 1146
rect 21824 1143 21890 1154
rect 21824 1109 21840 1143
rect 21874 1109 21890 1143
rect 21824 1098 21890 1109
rect 21998 1144 22622 1176
rect 22710 1164 22788 2122
rect 23302 2113 23331 2122
rect 23365 2122 25219 2147
rect 23365 2113 23392 2122
rect 23302 2092 23392 2113
rect 23388 2056 23446 2058
rect 23388 2039 23450 2056
rect 23388 2005 23400 2039
rect 23434 2005 23450 2039
rect 23388 1996 23450 2005
rect 22888 1958 23254 1962
rect 23336 1958 23402 1966
rect 22888 1930 23296 1958
rect 22888 1892 22916 1930
rect 23210 1911 23296 1930
rect 22888 1884 22954 1892
rect 22888 1850 22903 1884
rect 22937 1850 22954 1884
rect 22888 1838 22954 1850
rect 23060 1888 23128 1894
rect 23060 1836 23070 1888
rect 23122 1836 23128 1888
rect 23060 1830 23128 1836
rect 23210 1877 23256 1911
rect 23290 1877 23296 1911
rect 23336 1906 23342 1958
rect 23394 1906 23402 1958
rect 23336 1898 23352 1906
rect 23210 1839 23296 1877
rect 23210 1805 23256 1839
rect 23290 1805 23296 1839
rect 22970 1776 23038 1782
rect 22970 1724 22978 1776
rect 23030 1724 23038 1776
rect 22970 1714 23038 1724
rect 23210 1758 23296 1805
rect 23346 1877 23352 1898
rect 23386 1898 23402 1906
rect 23442 1926 23770 1958
rect 23442 1911 23538 1926
rect 23386 1877 23392 1898
rect 23346 1839 23392 1877
rect 23346 1805 23352 1839
rect 23386 1805 23392 1839
rect 23346 1758 23392 1805
rect 23442 1877 23448 1911
rect 23482 1877 23538 1911
rect 23742 1890 23770 1926
rect 23442 1839 23538 1877
rect 23442 1805 23448 1839
rect 23482 1805 23538 1839
rect 23700 1882 23770 1890
rect 23700 1848 23715 1882
rect 23749 1848 23770 1882
rect 23700 1830 23770 1848
rect 23876 1890 23940 1896
rect 23876 1838 23882 1890
rect 23934 1838 23940 1890
rect 23876 1832 23940 1838
rect 23442 1758 23538 1805
rect 22868 1643 23144 1674
rect 22868 1609 22897 1643
rect 22931 1609 22989 1643
rect 23023 1609 23081 1643
rect 23115 1609 23144 1643
rect 22868 1578 23144 1609
rect 23210 1558 23260 1758
rect 23292 1711 23350 1726
rect 23292 1677 23304 1711
rect 23338 1677 23350 1711
rect 23292 1660 23350 1677
rect 23404 1630 23462 1648
rect 23404 1596 23416 1630
rect 23450 1596 23462 1630
rect 23404 1586 23462 1596
rect 23492 1558 23538 1758
rect 23788 1774 23852 1780
rect 23788 1722 23794 1774
rect 23846 1722 23852 1774
rect 23788 1716 23852 1722
rect 23682 1643 23958 1674
rect 23682 1609 23711 1643
rect 23745 1609 23803 1643
rect 23837 1609 23895 1643
rect 23929 1609 23958 1643
rect 23682 1606 23958 1609
rect 22850 1541 22914 1548
rect 22850 1508 22856 1541
rect 22908 1508 22914 1541
rect 23026 1541 23090 1548
rect 23026 1508 23032 1541
rect 22908 1489 23032 1508
rect 23084 1489 23090 1541
rect 22856 1480 23090 1489
rect 23210 1546 23312 1558
rect 23210 1512 23272 1546
rect 23306 1512 23312 1546
rect 23210 1474 23312 1512
rect 23362 1546 23408 1558
rect 23362 1512 23368 1546
rect 23402 1512 23408 1546
rect 23362 1492 23408 1512
rect 23458 1546 23538 1558
rect 23458 1512 23464 1546
rect 23498 1512 23538 1546
rect 23210 1442 23272 1474
rect 23006 1440 23272 1442
rect 23306 1440 23312 1474
rect 23006 1428 23312 1440
rect 23352 1486 23418 1492
rect 23352 1434 23360 1486
rect 23412 1434 23418 1486
rect 23352 1428 23418 1434
rect 23458 1474 23538 1512
rect 23458 1440 23464 1474
rect 23498 1440 23538 1474
rect 23654 1578 23958 1606
rect 23458 1428 23504 1440
rect 23006 1414 23260 1428
rect 22850 1408 22916 1414
rect 22850 1356 22858 1408
rect 22910 1356 22916 1408
rect 22850 1350 22916 1356
rect 21998 1141 22028 1144
rect 22080 1141 22622 1144
rect 21998 1107 22027 1141
rect 22080 1107 22119 1141
rect 22153 1107 22211 1141
rect 22245 1139 22622 1141
rect 22245 1107 22373 1139
rect 21998 1092 22028 1107
rect 22080 1105 22373 1107
rect 22407 1105 22465 1139
rect 22499 1105 22557 1139
rect 22591 1105 22622 1139
rect 22080 1092 22622 1105
rect 21998 1074 22622 1092
rect 22690 1150 22966 1164
rect 22690 1133 22882 1150
rect 22934 1133 22966 1150
rect 22690 1099 22719 1133
rect 22753 1099 22811 1133
rect 22845 1099 22882 1133
rect 22937 1099 22966 1133
rect 22690 1098 22882 1099
rect 22934 1098 22966 1099
rect 22690 1068 22966 1098
rect 23006 1064 23034 1414
rect 23306 1390 23370 1400
rect 23306 1356 23320 1390
rect 23354 1356 23626 1390
rect 23306 1338 23370 1356
rect 23222 1292 23294 1304
rect 23222 1240 23232 1292
rect 23284 1240 23294 1292
rect 23222 1228 23294 1240
rect 23592 1174 23626 1356
rect 23654 1274 23682 1578
rect 23654 1264 23722 1274
rect 23654 1230 23670 1264
rect 23704 1230 23722 1264
rect 23654 1216 23722 1230
rect 23066 1146 23626 1174
rect 23066 1143 23132 1146
rect 23066 1109 23082 1143
rect 23116 1109 23132 1143
rect 23066 1100 23132 1109
rect 23300 1091 23390 1112
rect 21498 983 21738 1000
rect 21782 1056 21848 1062
rect 21782 1004 21790 1056
rect 21842 1004 21848 1056
rect 21782 998 21796 1004
rect 21232 943 21278 976
rect 21232 909 21238 943
rect 21272 909 21278 943
rect 21498 949 21510 983
rect 21544 972 21738 983
rect 21790 981 21796 998
rect 21830 998 21848 1004
rect 21878 1015 21924 1062
rect 23006 1036 23078 1064
rect 21830 981 21836 998
rect 21544 949 21736 972
rect 21498 940 21736 949
rect 21232 862 21278 909
rect 21446 902 21512 910
rect 21360 898 21406 902
rect 20476 840 20548 844
rect 19936 815 20002 828
rect 19936 781 19952 815
rect 19986 781 20002 815
rect 19936 772 20002 781
rect 20476 788 20485 840
rect 20537 788 20548 840
rect 20476 776 20548 788
rect 20672 838 20746 858
rect 21320 855 21406 898
rect 20672 804 20684 838
rect 20718 804 20746 838
rect 20672 780 20746 804
rect 20782 844 20850 850
rect 20782 792 20789 844
rect 20841 838 20850 844
rect 20841 832 20934 838
rect 20841 798 20880 832
rect 20914 798 20934 832
rect 20841 792 20934 798
rect 20782 788 20934 792
rect 21178 815 21244 826
rect 20782 786 20850 788
rect 21178 781 21194 815
rect 21228 781 21244 815
rect 21178 768 21244 781
rect 21320 821 21366 855
rect 21400 821 21406 855
rect 21446 850 21452 902
rect 21504 850 21512 902
rect 21446 842 21462 850
rect 21320 783 21406 821
rect 21320 749 21366 783
rect 21400 749 21406 783
rect 20258 728 20316 742
rect 20258 708 20270 728
rect 19788 694 20270 708
rect 20304 694 20316 728
rect 19788 674 20316 694
rect 21320 702 21406 749
rect 21456 821 21462 842
rect 21496 842 21512 850
rect 21552 855 21648 902
rect 21496 821 21502 842
rect 21456 783 21502 821
rect 21456 749 21462 783
rect 21496 749 21502 783
rect 21456 702 21502 749
rect 21552 821 21558 855
rect 21592 821 21648 855
rect 21552 783 21648 821
rect 21552 749 21558 783
rect 21592 749 21648 783
rect 21552 702 21648 749
rect 19680 372 19726 384
rect 19788 344 19848 674
rect 21320 648 21370 702
rect 19894 624 19970 630
rect 19894 572 19902 624
rect 19954 572 19970 624
rect 19894 566 19970 572
rect 20110 597 20732 628
rect 19528 334 19848 344
rect 19528 300 19542 334
rect 19576 300 19848 334
rect 19528 282 19848 300
rect 20110 563 20139 597
rect 20173 563 20231 597
rect 20265 563 20323 597
rect 20357 595 20732 597
rect 20357 563 20485 595
rect 20110 561 20485 563
rect 20519 561 20577 595
rect 20611 561 20669 595
rect 20703 561 20732 595
rect 20110 530 20732 561
rect 20802 602 21078 620
rect 20802 589 20925 602
rect 20977 589 21078 602
rect 21154 598 21212 606
rect 20802 555 20831 589
rect 20865 555 20923 589
rect 20977 555 21015 589
rect 21049 555 21078 589
rect 20802 550 20925 555
rect 20977 550 21078 555
rect 20110 254 20208 530
rect 20802 524 21078 550
rect 21146 592 21220 598
rect 21146 540 21157 592
rect 21209 540 21220 592
rect 21300 582 21370 648
rect 21402 655 21460 670
rect 21402 621 21414 655
rect 21448 621 21460 655
rect 21402 604 21460 621
rect 21146 534 21220 540
rect 21154 528 21212 534
rect 20870 254 20954 524
rect 21320 502 21370 582
rect 21514 574 21572 592
rect 21514 540 21526 574
rect 21560 540 21572 574
rect 21514 530 21572 540
rect 21602 502 21648 702
rect 21320 490 21422 502
rect 21320 456 21382 490
rect 21416 456 21422 490
rect 21320 418 21422 456
rect 21472 490 21518 502
rect 21472 456 21478 490
rect 21512 456 21518 490
rect 21472 436 21518 456
rect 21568 490 21648 502
rect 21568 456 21574 490
rect 21608 456 21648 490
rect 21320 384 21382 418
rect 21416 384 21422 418
rect 21320 372 21422 384
rect 21462 430 21528 436
rect 21462 378 21470 430
rect 21522 378 21528 430
rect 21462 372 21528 378
rect 21568 418 21648 456
rect 21568 384 21574 418
rect 21608 384 21648 418
rect 21676 708 21736 940
rect 21790 943 21836 981
rect 21790 909 21796 943
rect 21830 909 21836 943
rect 21790 862 21836 909
rect 21878 981 21884 1015
rect 21918 981 21924 1015
rect 21878 943 21924 981
rect 21878 909 21884 943
rect 21918 909 21924 943
rect 21878 862 21924 909
rect 23032 1015 23078 1036
rect 23032 981 23038 1015
rect 23072 981 23078 1015
rect 23032 943 23078 981
rect 23032 909 23038 943
rect 23072 909 23078 943
rect 23032 862 23078 909
rect 23120 1042 23166 1062
rect 23300 1057 23329 1091
rect 23363 1057 23390 1091
rect 23120 1036 23188 1042
rect 23300 1036 23390 1057
rect 23120 1015 23128 1036
rect 23120 981 23126 1015
rect 23180 984 23188 1036
rect 23160 981 23188 984
rect 23120 976 23188 981
rect 23386 1000 23444 1002
rect 23592 1000 23626 1146
rect 23712 1143 23778 1154
rect 23712 1109 23728 1143
rect 23762 1109 23778 1143
rect 23712 1098 23778 1109
rect 23886 1144 24510 1176
rect 24598 1164 24676 2122
rect 25190 2113 25219 2122
rect 25253 2122 27107 2147
rect 25253 2113 25280 2122
rect 25190 2092 25280 2113
rect 25276 2056 25334 2058
rect 25276 2039 25338 2056
rect 25276 2005 25288 2039
rect 25322 2005 25338 2039
rect 25276 1996 25338 2005
rect 24776 1958 25142 1962
rect 25224 1958 25290 1966
rect 24776 1930 25184 1958
rect 24776 1892 24804 1930
rect 25098 1911 25184 1930
rect 24776 1884 24842 1892
rect 24776 1850 24791 1884
rect 24825 1850 24842 1884
rect 24776 1838 24842 1850
rect 24948 1888 25016 1894
rect 24948 1836 24958 1888
rect 25010 1836 25016 1888
rect 24948 1830 25016 1836
rect 25098 1877 25144 1911
rect 25178 1877 25184 1911
rect 25224 1906 25230 1958
rect 25282 1906 25290 1958
rect 25224 1898 25240 1906
rect 25098 1839 25184 1877
rect 25098 1805 25144 1839
rect 25178 1805 25184 1839
rect 24858 1776 24926 1782
rect 24858 1724 24866 1776
rect 24918 1724 24926 1776
rect 24858 1714 24926 1724
rect 25098 1758 25184 1805
rect 25234 1877 25240 1898
rect 25274 1898 25290 1906
rect 25330 1926 25658 1958
rect 25330 1911 25426 1926
rect 25274 1877 25280 1898
rect 25234 1839 25280 1877
rect 25234 1805 25240 1839
rect 25274 1805 25280 1839
rect 25234 1758 25280 1805
rect 25330 1877 25336 1911
rect 25370 1877 25426 1911
rect 25630 1890 25658 1926
rect 25330 1839 25426 1877
rect 25330 1805 25336 1839
rect 25370 1805 25426 1839
rect 25588 1882 25658 1890
rect 25588 1848 25603 1882
rect 25637 1848 25658 1882
rect 25588 1830 25658 1848
rect 25764 1890 25828 1896
rect 25764 1838 25770 1890
rect 25822 1838 25828 1890
rect 25764 1832 25828 1838
rect 25330 1758 25426 1805
rect 24756 1643 25032 1674
rect 24756 1609 24785 1643
rect 24819 1609 24877 1643
rect 24911 1609 24969 1643
rect 25003 1609 25032 1643
rect 24756 1578 25032 1609
rect 25098 1558 25148 1758
rect 25180 1711 25238 1726
rect 25180 1677 25192 1711
rect 25226 1677 25238 1711
rect 25180 1660 25238 1677
rect 25292 1630 25350 1648
rect 25292 1596 25304 1630
rect 25338 1596 25350 1630
rect 25292 1586 25350 1596
rect 25380 1558 25426 1758
rect 25676 1774 25740 1780
rect 25676 1722 25682 1774
rect 25734 1722 25740 1774
rect 25676 1716 25740 1722
rect 25570 1643 25846 1674
rect 25570 1609 25599 1643
rect 25633 1609 25691 1643
rect 25725 1609 25783 1643
rect 25817 1609 25846 1643
rect 25570 1606 25846 1609
rect 24738 1541 24802 1548
rect 24738 1508 24744 1541
rect 24796 1508 24802 1541
rect 24914 1541 24978 1548
rect 24914 1508 24920 1541
rect 24796 1489 24920 1508
rect 24972 1489 24978 1541
rect 24744 1480 24978 1489
rect 25098 1546 25200 1558
rect 25098 1512 25160 1546
rect 25194 1512 25200 1546
rect 25098 1474 25200 1512
rect 25250 1546 25296 1558
rect 25250 1512 25256 1546
rect 25290 1512 25296 1546
rect 25250 1492 25296 1512
rect 25346 1546 25426 1558
rect 25346 1512 25352 1546
rect 25386 1512 25426 1546
rect 25098 1442 25160 1474
rect 24894 1440 25160 1442
rect 25194 1440 25200 1474
rect 24894 1428 25200 1440
rect 25240 1486 25306 1492
rect 25240 1434 25248 1486
rect 25300 1434 25306 1486
rect 25240 1428 25306 1434
rect 25346 1474 25426 1512
rect 25346 1440 25352 1474
rect 25386 1440 25426 1474
rect 25542 1578 25846 1606
rect 25346 1428 25392 1440
rect 24894 1414 25148 1428
rect 24738 1408 24804 1414
rect 24738 1356 24746 1408
rect 24798 1356 24804 1408
rect 24738 1350 24804 1356
rect 23886 1141 23916 1144
rect 23968 1141 24510 1144
rect 23886 1107 23915 1141
rect 23968 1107 24007 1141
rect 24041 1107 24099 1141
rect 24133 1139 24510 1141
rect 24133 1107 24261 1139
rect 23886 1092 23916 1107
rect 23968 1105 24261 1107
rect 24295 1105 24353 1139
rect 24387 1105 24445 1139
rect 24479 1105 24510 1139
rect 23968 1092 24510 1105
rect 23886 1074 24510 1092
rect 24578 1150 24854 1164
rect 24578 1133 24770 1150
rect 24822 1133 24854 1150
rect 24578 1099 24607 1133
rect 24641 1099 24699 1133
rect 24733 1099 24770 1133
rect 24825 1099 24854 1133
rect 24578 1098 24770 1099
rect 24822 1098 24854 1099
rect 24578 1068 24854 1098
rect 24894 1064 24922 1414
rect 25194 1390 25258 1400
rect 25194 1356 25208 1390
rect 25242 1356 25514 1390
rect 25194 1338 25258 1356
rect 25110 1292 25182 1304
rect 25110 1240 25120 1292
rect 25172 1240 25182 1292
rect 25110 1228 25182 1240
rect 25480 1174 25514 1356
rect 25542 1274 25570 1578
rect 25542 1264 25610 1274
rect 25542 1230 25558 1264
rect 25592 1230 25610 1264
rect 25542 1216 25610 1230
rect 24954 1146 25514 1174
rect 24954 1143 25020 1146
rect 24954 1109 24970 1143
rect 25004 1109 25020 1143
rect 24954 1100 25020 1109
rect 25188 1091 25278 1112
rect 23386 983 23626 1000
rect 23670 1056 23736 1062
rect 23670 1004 23678 1056
rect 23730 1004 23736 1056
rect 23670 998 23684 1004
rect 23120 943 23166 976
rect 23120 909 23126 943
rect 23160 909 23166 943
rect 23386 949 23398 983
rect 23432 972 23626 983
rect 23678 981 23684 998
rect 23718 998 23736 1004
rect 23766 1015 23812 1062
rect 24894 1036 24966 1064
rect 23718 981 23724 998
rect 23432 949 23624 972
rect 23386 940 23624 949
rect 23120 862 23166 909
rect 23334 902 23400 910
rect 23248 898 23294 902
rect 22364 840 22436 844
rect 21824 815 21890 828
rect 21824 781 21840 815
rect 21874 781 21890 815
rect 21824 772 21890 781
rect 22364 788 22373 840
rect 22425 788 22436 840
rect 22364 776 22436 788
rect 22560 838 22634 858
rect 23208 855 23294 898
rect 22560 804 22572 838
rect 22606 804 22634 838
rect 22560 780 22634 804
rect 22670 844 22738 850
rect 22670 792 22677 844
rect 22729 838 22738 844
rect 22729 832 22822 838
rect 22729 798 22768 832
rect 22802 798 22822 832
rect 22729 792 22822 798
rect 22670 788 22822 792
rect 23066 815 23132 826
rect 22670 786 22738 788
rect 23066 781 23082 815
rect 23116 781 23132 815
rect 23066 768 23132 781
rect 23208 821 23254 855
rect 23288 821 23294 855
rect 23334 850 23340 902
rect 23392 850 23400 902
rect 23334 842 23350 850
rect 23208 783 23294 821
rect 23208 749 23254 783
rect 23288 749 23294 783
rect 22146 728 22204 742
rect 22146 708 22158 728
rect 21676 694 22158 708
rect 22192 694 22204 728
rect 21676 674 22204 694
rect 23208 702 23294 749
rect 23344 821 23350 842
rect 23384 842 23400 850
rect 23440 855 23536 902
rect 23384 821 23390 842
rect 23344 783 23390 821
rect 23344 749 23350 783
rect 23384 749 23390 783
rect 23344 702 23390 749
rect 23440 821 23446 855
rect 23480 821 23536 855
rect 23440 783 23536 821
rect 23440 749 23446 783
rect 23480 749 23536 783
rect 23440 702 23536 749
rect 21568 372 21614 384
rect 21676 344 21736 674
rect 23208 648 23258 702
rect 21782 624 21858 630
rect 21782 572 21790 624
rect 21842 572 21858 624
rect 21782 566 21858 572
rect 21998 597 22620 628
rect 21416 334 21736 344
rect 21416 300 21430 334
rect 21464 300 21736 334
rect 21416 282 21736 300
rect 21998 563 22027 597
rect 22061 563 22119 597
rect 22153 563 22211 597
rect 22245 595 22620 597
rect 22245 563 22373 595
rect 21998 561 22373 563
rect 22407 561 22465 595
rect 22499 561 22557 595
rect 22591 561 22620 595
rect 21998 530 22620 561
rect 22690 602 22966 620
rect 22690 589 22813 602
rect 22865 589 22966 602
rect 23042 598 23100 606
rect 22690 555 22719 589
rect 22753 555 22811 589
rect 22865 555 22903 589
rect 22937 555 22966 589
rect 22690 550 22813 555
rect 22865 550 22966 555
rect 21998 254 22096 530
rect 22690 524 22966 550
rect 23034 592 23108 598
rect 23034 540 23045 592
rect 23097 540 23108 592
rect 23188 582 23258 648
rect 23290 655 23348 670
rect 23290 621 23302 655
rect 23336 621 23348 655
rect 23290 604 23348 621
rect 23034 534 23108 540
rect 23042 528 23100 534
rect 22758 254 22842 524
rect 23208 502 23258 582
rect 23402 574 23460 592
rect 23402 540 23414 574
rect 23448 540 23460 574
rect 23402 530 23460 540
rect 23490 502 23536 702
rect 23208 490 23310 502
rect 23208 456 23270 490
rect 23304 456 23310 490
rect 23208 418 23310 456
rect 23360 490 23406 502
rect 23360 456 23366 490
rect 23400 456 23406 490
rect 23360 436 23406 456
rect 23456 490 23536 502
rect 23456 456 23462 490
rect 23496 456 23536 490
rect 23208 384 23270 418
rect 23304 384 23310 418
rect 23208 372 23310 384
rect 23350 430 23416 436
rect 23350 378 23358 430
rect 23410 378 23416 430
rect 23350 372 23416 378
rect 23456 418 23536 456
rect 23456 384 23462 418
rect 23496 384 23536 418
rect 23564 708 23624 940
rect 23678 943 23724 981
rect 23678 909 23684 943
rect 23718 909 23724 943
rect 23678 862 23724 909
rect 23766 981 23772 1015
rect 23806 981 23812 1015
rect 23766 943 23812 981
rect 23766 909 23772 943
rect 23806 909 23812 943
rect 23766 862 23812 909
rect 24920 1015 24966 1036
rect 24920 981 24926 1015
rect 24960 981 24966 1015
rect 24920 943 24966 981
rect 24920 909 24926 943
rect 24960 909 24966 943
rect 24920 862 24966 909
rect 25008 1042 25054 1062
rect 25188 1057 25217 1091
rect 25251 1057 25278 1091
rect 25008 1036 25076 1042
rect 25188 1036 25278 1057
rect 25008 1015 25016 1036
rect 25008 981 25014 1015
rect 25068 984 25076 1036
rect 25048 981 25076 984
rect 25008 976 25076 981
rect 25274 1000 25332 1002
rect 25480 1000 25514 1146
rect 25600 1143 25666 1154
rect 25600 1109 25616 1143
rect 25650 1109 25666 1143
rect 25600 1098 25666 1109
rect 25774 1144 26398 1176
rect 26486 1164 26564 2122
rect 27078 2113 27107 2122
rect 27141 2122 28995 2147
rect 27141 2113 27168 2122
rect 27078 2092 27168 2113
rect 27164 2056 27222 2058
rect 27164 2039 27226 2056
rect 27164 2005 27176 2039
rect 27210 2005 27226 2039
rect 27164 1996 27226 2005
rect 26664 1958 27030 1962
rect 27112 1958 27178 1966
rect 26664 1930 27072 1958
rect 26664 1892 26692 1930
rect 26986 1911 27072 1930
rect 26664 1884 26730 1892
rect 26664 1850 26679 1884
rect 26713 1850 26730 1884
rect 26664 1838 26730 1850
rect 26836 1888 26904 1894
rect 26836 1836 26846 1888
rect 26898 1836 26904 1888
rect 26836 1830 26904 1836
rect 26986 1877 27032 1911
rect 27066 1877 27072 1911
rect 27112 1906 27118 1958
rect 27170 1906 27178 1958
rect 27112 1898 27128 1906
rect 26986 1839 27072 1877
rect 26986 1805 27032 1839
rect 27066 1805 27072 1839
rect 26746 1776 26814 1782
rect 26746 1724 26754 1776
rect 26806 1724 26814 1776
rect 26746 1714 26814 1724
rect 26986 1758 27072 1805
rect 27122 1877 27128 1898
rect 27162 1898 27178 1906
rect 27218 1926 27546 1958
rect 27218 1911 27314 1926
rect 27162 1877 27168 1898
rect 27122 1839 27168 1877
rect 27122 1805 27128 1839
rect 27162 1805 27168 1839
rect 27122 1758 27168 1805
rect 27218 1877 27224 1911
rect 27258 1877 27314 1911
rect 27518 1890 27546 1926
rect 27218 1839 27314 1877
rect 27218 1805 27224 1839
rect 27258 1805 27314 1839
rect 27476 1882 27546 1890
rect 27476 1848 27491 1882
rect 27525 1848 27546 1882
rect 27476 1830 27546 1848
rect 27652 1890 27716 1896
rect 27652 1838 27658 1890
rect 27710 1838 27716 1890
rect 27652 1832 27716 1838
rect 27218 1758 27314 1805
rect 26644 1643 26920 1674
rect 26644 1609 26673 1643
rect 26707 1609 26765 1643
rect 26799 1609 26857 1643
rect 26891 1609 26920 1643
rect 26644 1578 26920 1609
rect 26986 1558 27036 1758
rect 27068 1711 27126 1726
rect 27068 1677 27080 1711
rect 27114 1677 27126 1711
rect 27068 1660 27126 1677
rect 27180 1630 27238 1648
rect 27180 1596 27192 1630
rect 27226 1596 27238 1630
rect 27180 1586 27238 1596
rect 27268 1558 27314 1758
rect 27564 1774 27628 1780
rect 27564 1722 27570 1774
rect 27622 1722 27628 1774
rect 27564 1716 27628 1722
rect 27458 1643 27734 1674
rect 27458 1609 27487 1643
rect 27521 1609 27579 1643
rect 27613 1609 27671 1643
rect 27705 1609 27734 1643
rect 27458 1606 27734 1609
rect 26626 1541 26690 1548
rect 26626 1508 26632 1541
rect 26684 1508 26690 1541
rect 26802 1541 26866 1548
rect 26802 1508 26808 1541
rect 26684 1489 26808 1508
rect 26860 1489 26866 1541
rect 26632 1480 26866 1489
rect 26986 1546 27088 1558
rect 26986 1512 27048 1546
rect 27082 1512 27088 1546
rect 26986 1474 27088 1512
rect 27138 1546 27184 1558
rect 27138 1512 27144 1546
rect 27178 1512 27184 1546
rect 27138 1492 27184 1512
rect 27234 1546 27314 1558
rect 27234 1512 27240 1546
rect 27274 1512 27314 1546
rect 26986 1442 27048 1474
rect 26782 1440 27048 1442
rect 27082 1440 27088 1474
rect 26782 1428 27088 1440
rect 27128 1486 27194 1492
rect 27128 1434 27136 1486
rect 27188 1434 27194 1486
rect 27128 1428 27194 1434
rect 27234 1474 27314 1512
rect 27234 1440 27240 1474
rect 27274 1440 27314 1474
rect 27430 1578 27734 1606
rect 27234 1428 27280 1440
rect 26782 1414 27036 1428
rect 26626 1408 26692 1414
rect 26626 1356 26634 1408
rect 26686 1356 26692 1408
rect 26626 1350 26692 1356
rect 25774 1141 25804 1144
rect 25856 1141 26398 1144
rect 25774 1107 25803 1141
rect 25856 1107 25895 1141
rect 25929 1107 25987 1141
rect 26021 1139 26398 1141
rect 26021 1107 26149 1139
rect 25774 1092 25804 1107
rect 25856 1105 26149 1107
rect 26183 1105 26241 1139
rect 26275 1105 26333 1139
rect 26367 1105 26398 1139
rect 25856 1092 26398 1105
rect 25774 1074 26398 1092
rect 26466 1150 26742 1164
rect 26466 1133 26658 1150
rect 26710 1133 26742 1150
rect 26466 1099 26495 1133
rect 26529 1099 26587 1133
rect 26621 1099 26658 1133
rect 26713 1099 26742 1133
rect 26466 1098 26658 1099
rect 26710 1098 26742 1099
rect 26466 1068 26742 1098
rect 26782 1064 26810 1414
rect 27082 1390 27146 1400
rect 27082 1356 27096 1390
rect 27130 1356 27402 1390
rect 27082 1338 27146 1356
rect 26998 1292 27070 1304
rect 26998 1240 27008 1292
rect 27060 1240 27070 1292
rect 26998 1228 27070 1240
rect 27368 1174 27402 1356
rect 27430 1274 27458 1578
rect 27430 1264 27498 1274
rect 27430 1230 27446 1264
rect 27480 1230 27498 1264
rect 27430 1216 27498 1230
rect 26842 1146 27402 1174
rect 26842 1143 26908 1146
rect 26842 1109 26858 1143
rect 26892 1109 26908 1143
rect 26842 1100 26908 1109
rect 27076 1091 27166 1112
rect 25274 983 25514 1000
rect 25558 1056 25624 1062
rect 25558 1004 25566 1056
rect 25618 1004 25624 1056
rect 25558 998 25572 1004
rect 25008 943 25054 976
rect 25008 909 25014 943
rect 25048 909 25054 943
rect 25274 949 25286 983
rect 25320 972 25514 983
rect 25566 981 25572 998
rect 25606 998 25624 1004
rect 25654 1015 25700 1062
rect 26782 1036 26854 1064
rect 25606 981 25612 998
rect 25320 949 25512 972
rect 25274 940 25512 949
rect 25008 862 25054 909
rect 25222 902 25288 910
rect 25136 898 25182 902
rect 24252 840 24324 844
rect 23712 815 23778 828
rect 23712 781 23728 815
rect 23762 781 23778 815
rect 23712 772 23778 781
rect 24252 788 24261 840
rect 24313 788 24324 840
rect 24252 776 24324 788
rect 24448 838 24522 858
rect 25096 855 25182 898
rect 24448 804 24460 838
rect 24494 804 24522 838
rect 24448 780 24522 804
rect 24558 844 24626 850
rect 24558 792 24565 844
rect 24617 838 24626 844
rect 24617 832 24710 838
rect 24617 798 24656 832
rect 24690 798 24710 832
rect 24617 792 24710 798
rect 24558 788 24710 792
rect 24954 815 25020 826
rect 24558 786 24626 788
rect 24954 781 24970 815
rect 25004 781 25020 815
rect 24954 768 25020 781
rect 25096 821 25142 855
rect 25176 821 25182 855
rect 25222 850 25228 902
rect 25280 850 25288 902
rect 25222 842 25238 850
rect 25096 783 25182 821
rect 25096 749 25142 783
rect 25176 749 25182 783
rect 24034 728 24092 742
rect 24034 708 24046 728
rect 23564 694 24046 708
rect 24080 694 24092 728
rect 23564 674 24092 694
rect 25096 702 25182 749
rect 25232 821 25238 842
rect 25272 842 25288 850
rect 25328 855 25424 902
rect 25272 821 25278 842
rect 25232 783 25278 821
rect 25232 749 25238 783
rect 25272 749 25278 783
rect 25232 702 25278 749
rect 25328 821 25334 855
rect 25368 821 25424 855
rect 25328 783 25424 821
rect 25328 749 25334 783
rect 25368 749 25424 783
rect 25328 702 25424 749
rect 23456 372 23502 384
rect 23564 344 23624 674
rect 25096 648 25146 702
rect 23670 624 23746 630
rect 23670 572 23678 624
rect 23730 572 23746 624
rect 23670 566 23746 572
rect 23886 597 24508 628
rect 23304 334 23624 344
rect 23304 300 23318 334
rect 23352 300 23624 334
rect 23304 282 23624 300
rect 23886 563 23915 597
rect 23949 563 24007 597
rect 24041 563 24099 597
rect 24133 595 24508 597
rect 24133 563 24261 595
rect 23886 561 24261 563
rect 24295 561 24353 595
rect 24387 561 24445 595
rect 24479 561 24508 595
rect 23886 530 24508 561
rect 24578 602 24854 620
rect 24578 589 24701 602
rect 24753 589 24854 602
rect 24930 598 24988 606
rect 24578 555 24607 589
rect 24641 555 24699 589
rect 24753 555 24791 589
rect 24825 555 24854 589
rect 24578 550 24701 555
rect 24753 550 24854 555
rect 23886 254 23984 530
rect 24578 524 24854 550
rect 24922 592 24996 598
rect 24922 540 24933 592
rect 24985 540 24996 592
rect 25076 582 25146 648
rect 25178 655 25236 670
rect 25178 621 25190 655
rect 25224 621 25236 655
rect 25178 604 25236 621
rect 24922 534 24996 540
rect 24930 528 24988 534
rect 24646 254 24730 524
rect 25096 502 25146 582
rect 25290 574 25348 592
rect 25290 540 25302 574
rect 25336 540 25348 574
rect 25290 530 25348 540
rect 25378 502 25424 702
rect 25096 490 25198 502
rect 25096 456 25158 490
rect 25192 456 25198 490
rect 25096 418 25198 456
rect 25248 490 25294 502
rect 25248 456 25254 490
rect 25288 456 25294 490
rect 25248 436 25294 456
rect 25344 490 25424 502
rect 25344 456 25350 490
rect 25384 456 25424 490
rect 25096 384 25158 418
rect 25192 384 25198 418
rect 25096 372 25198 384
rect 25238 430 25304 436
rect 25238 378 25246 430
rect 25298 378 25304 430
rect 25238 372 25304 378
rect 25344 418 25424 456
rect 25344 384 25350 418
rect 25384 384 25424 418
rect 25452 708 25512 940
rect 25566 943 25612 981
rect 25566 909 25572 943
rect 25606 909 25612 943
rect 25566 862 25612 909
rect 25654 981 25660 1015
rect 25694 981 25700 1015
rect 25654 943 25700 981
rect 25654 909 25660 943
rect 25694 909 25700 943
rect 25654 862 25700 909
rect 26808 1015 26854 1036
rect 26808 981 26814 1015
rect 26848 981 26854 1015
rect 26808 943 26854 981
rect 26808 909 26814 943
rect 26848 909 26854 943
rect 26808 862 26854 909
rect 26896 1042 26942 1062
rect 27076 1057 27105 1091
rect 27139 1057 27166 1091
rect 26896 1036 26964 1042
rect 27076 1036 27166 1057
rect 26896 1015 26904 1036
rect 26896 981 26902 1015
rect 26956 984 26964 1036
rect 26936 981 26964 984
rect 26896 976 26964 981
rect 27162 1000 27220 1002
rect 27368 1000 27402 1146
rect 27488 1143 27554 1154
rect 27488 1109 27504 1143
rect 27538 1109 27554 1143
rect 27488 1098 27554 1109
rect 27662 1144 28286 1176
rect 28374 1164 28452 2122
rect 28966 2113 28995 2122
rect 29029 2122 30883 2147
rect 29029 2113 29056 2122
rect 28966 2092 29056 2113
rect 29052 2056 29110 2058
rect 29052 2039 29114 2056
rect 29052 2005 29064 2039
rect 29098 2005 29114 2039
rect 29052 1996 29114 2005
rect 28552 1958 28918 1962
rect 29000 1958 29066 1966
rect 28552 1930 28960 1958
rect 28552 1892 28580 1930
rect 28874 1911 28960 1930
rect 28552 1884 28618 1892
rect 28552 1850 28567 1884
rect 28601 1850 28618 1884
rect 28552 1838 28618 1850
rect 28724 1888 28792 1894
rect 28724 1836 28734 1888
rect 28786 1836 28792 1888
rect 28724 1830 28792 1836
rect 28874 1877 28920 1911
rect 28954 1877 28960 1911
rect 29000 1906 29006 1958
rect 29058 1906 29066 1958
rect 29000 1898 29016 1906
rect 28874 1839 28960 1877
rect 28874 1805 28920 1839
rect 28954 1805 28960 1839
rect 28634 1776 28702 1782
rect 28634 1724 28642 1776
rect 28694 1724 28702 1776
rect 28634 1714 28702 1724
rect 28874 1758 28960 1805
rect 29010 1877 29016 1898
rect 29050 1898 29066 1906
rect 29106 1926 29434 1958
rect 29106 1911 29202 1926
rect 29050 1877 29056 1898
rect 29010 1839 29056 1877
rect 29010 1805 29016 1839
rect 29050 1805 29056 1839
rect 29010 1758 29056 1805
rect 29106 1877 29112 1911
rect 29146 1877 29202 1911
rect 29406 1890 29434 1926
rect 29106 1839 29202 1877
rect 29106 1805 29112 1839
rect 29146 1805 29202 1839
rect 29364 1882 29434 1890
rect 29364 1848 29379 1882
rect 29413 1848 29434 1882
rect 29364 1830 29434 1848
rect 29540 1890 29604 1896
rect 29540 1838 29546 1890
rect 29598 1838 29604 1890
rect 29540 1832 29604 1838
rect 29106 1758 29202 1805
rect 28532 1643 28808 1674
rect 28532 1609 28561 1643
rect 28595 1609 28653 1643
rect 28687 1609 28745 1643
rect 28779 1609 28808 1643
rect 28532 1578 28808 1609
rect 28874 1558 28924 1758
rect 28956 1711 29014 1726
rect 28956 1677 28968 1711
rect 29002 1677 29014 1711
rect 28956 1660 29014 1677
rect 29068 1630 29126 1648
rect 29068 1596 29080 1630
rect 29114 1596 29126 1630
rect 29068 1586 29126 1596
rect 29156 1558 29202 1758
rect 29452 1774 29516 1780
rect 29452 1722 29458 1774
rect 29510 1722 29516 1774
rect 29452 1716 29516 1722
rect 29346 1643 29622 1674
rect 29346 1609 29375 1643
rect 29409 1609 29467 1643
rect 29501 1609 29559 1643
rect 29593 1609 29622 1643
rect 29346 1606 29622 1609
rect 28514 1541 28578 1548
rect 28514 1508 28520 1541
rect 28572 1508 28578 1541
rect 28690 1541 28754 1548
rect 28690 1508 28696 1541
rect 28572 1489 28696 1508
rect 28748 1489 28754 1541
rect 28520 1480 28754 1489
rect 28874 1546 28976 1558
rect 28874 1512 28936 1546
rect 28970 1512 28976 1546
rect 28874 1474 28976 1512
rect 29026 1546 29072 1558
rect 29026 1512 29032 1546
rect 29066 1512 29072 1546
rect 29026 1492 29072 1512
rect 29122 1546 29202 1558
rect 29122 1512 29128 1546
rect 29162 1512 29202 1546
rect 28874 1442 28936 1474
rect 28670 1440 28936 1442
rect 28970 1440 28976 1474
rect 28670 1428 28976 1440
rect 29016 1486 29082 1492
rect 29016 1434 29024 1486
rect 29076 1434 29082 1486
rect 29016 1428 29082 1434
rect 29122 1474 29202 1512
rect 29122 1440 29128 1474
rect 29162 1440 29202 1474
rect 29318 1578 29622 1606
rect 29122 1428 29168 1440
rect 28670 1414 28924 1428
rect 28514 1408 28580 1414
rect 28514 1356 28522 1408
rect 28574 1356 28580 1408
rect 28514 1350 28580 1356
rect 27662 1141 27692 1144
rect 27744 1141 28286 1144
rect 27662 1107 27691 1141
rect 27744 1107 27783 1141
rect 27817 1107 27875 1141
rect 27909 1139 28286 1141
rect 27909 1107 28037 1139
rect 27662 1092 27692 1107
rect 27744 1105 28037 1107
rect 28071 1105 28129 1139
rect 28163 1105 28221 1139
rect 28255 1105 28286 1139
rect 27744 1092 28286 1105
rect 27662 1074 28286 1092
rect 28354 1150 28630 1164
rect 28354 1133 28546 1150
rect 28598 1133 28630 1150
rect 28354 1099 28383 1133
rect 28417 1099 28475 1133
rect 28509 1099 28546 1133
rect 28601 1099 28630 1133
rect 28354 1098 28546 1099
rect 28598 1098 28630 1099
rect 28354 1068 28630 1098
rect 28670 1064 28698 1414
rect 28970 1390 29034 1400
rect 28970 1356 28984 1390
rect 29018 1356 29290 1390
rect 28970 1338 29034 1356
rect 28886 1292 28958 1304
rect 28886 1240 28896 1292
rect 28948 1240 28958 1292
rect 28886 1228 28958 1240
rect 29256 1174 29290 1356
rect 29318 1274 29346 1578
rect 29318 1264 29386 1274
rect 29318 1230 29334 1264
rect 29368 1230 29386 1264
rect 29318 1216 29386 1230
rect 28730 1146 29290 1174
rect 28730 1143 28796 1146
rect 28730 1109 28746 1143
rect 28780 1109 28796 1143
rect 28730 1100 28796 1109
rect 28964 1091 29054 1112
rect 27162 983 27402 1000
rect 27446 1056 27512 1062
rect 27446 1004 27454 1056
rect 27506 1004 27512 1056
rect 27446 998 27460 1004
rect 26896 943 26942 976
rect 26896 909 26902 943
rect 26936 909 26942 943
rect 27162 949 27174 983
rect 27208 972 27402 983
rect 27454 981 27460 998
rect 27494 998 27512 1004
rect 27542 1015 27588 1062
rect 28670 1036 28742 1064
rect 27494 981 27500 998
rect 27208 949 27400 972
rect 27162 940 27400 949
rect 26896 862 26942 909
rect 27110 902 27176 910
rect 27024 898 27070 902
rect 26140 840 26212 844
rect 25600 815 25666 828
rect 25600 781 25616 815
rect 25650 781 25666 815
rect 25600 772 25666 781
rect 26140 788 26149 840
rect 26201 788 26212 840
rect 26140 776 26212 788
rect 26336 838 26410 858
rect 26984 855 27070 898
rect 26336 804 26348 838
rect 26382 804 26410 838
rect 26336 780 26410 804
rect 26446 844 26514 850
rect 26446 792 26453 844
rect 26505 838 26514 844
rect 26505 832 26598 838
rect 26505 798 26544 832
rect 26578 798 26598 832
rect 26505 792 26598 798
rect 26446 788 26598 792
rect 26842 815 26908 826
rect 26446 786 26514 788
rect 26842 781 26858 815
rect 26892 781 26908 815
rect 26842 768 26908 781
rect 26984 821 27030 855
rect 27064 821 27070 855
rect 27110 850 27116 902
rect 27168 850 27176 902
rect 27110 842 27126 850
rect 26984 783 27070 821
rect 26984 749 27030 783
rect 27064 749 27070 783
rect 25922 728 25980 742
rect 25922 708 25934 728
rect 25452 694 25934 708
rect 25968 694 25980 728
rect 25452 674 25980 694
rect 26984 702 27070 749
rect 27120 821 27126 842
rect 27160 842 27176 850
rect 27216 855 27312 902
rect 27160 821 27166 842
rect 27120 783 27166 821
rect 27120 749 27126 783
rect 27160 749 27166 783
rect 27120 702 27166 749
rect 27216 821 27222 855
rect 27256 821 27312 855
rect 27216 783 27312 821
rect 27216 749 27222 783
rect 27256 749 27312 783
rect 27216 702 27312 749
rect 25344 372 25390 384
rect 25452 344 25512 674
rect 26984 648 27034 702
rect 25558 624 25634 630
rect 25558 572 25566 624
rect 25618 572 25634 624
rect 25558 566 25634 572
rect 25774 597 26396 628
rect 25192 334 25512 344
rect 25192 300 25206 334
rect 25240 300 25512 334
rect 25192 282 25512 300
rect 25774 563 25803 597
rect 25837 563 25895 597
rect 25929 563 25987 597
rect 26021 595 26396 597
rect 26021 563 26149 595
rect 25774 561 26149 563
rect 26183 561 26241 595
rect 26275 561 26333 595
rect 26367 561 26396 595
rect 25774 530 26396 561
rect 26466 602 26742 620
rect 26466 589 26589 602
rect 26641 589 26742 602
rect 26818 598 26876 606
rect 26466 555 26495 589
rect 26529 555 26587 589
rect 26641 555 26679 589
rect 26713 555 26742 589
rect 26466 550 26589 555
rect 26641 550 26742 555
rect 25774 254 25872 530
rect 26466 524 26742 550
rect 26810 592 26884 598
rect 26810 540 26821 592
rect 26873 540 26884 592
rect 26964 582 27034 648
rect 27066 655 27124 670
rect 27066 621 27078 655
rect 27112 621 27124 655
rect 27066 604 27124 621
rect 26810 534 26884 540
rect 26818 528 26876 534
rect 26534 254 26618 524
rect 26984 502 27034 582
rect 27178 574 27236 592
rect 27178 540 27190 574
rect 27224 540 27236 574
rect 27178 530 27236 540
rect 27266 502 27312 702
rect 26984 490 27086 502
rect 26984 456 27046 490
rect 27080 456 27086 490
rect 26984 418 27086 456
rect 27136 490 27182 502
rect 27136 456 27142 490
rect 27176 456 27182 490
rect 27136 436 27182 456
rect 27232 490 27312 502
rect 27232 456 27238 490
rect 27272 456 27312 490
rect 26984 384 27046 418
rect 27080 384 27086 418
rect 26984 372 27086 384
rect 27126 430 27192 436
rect 27126 378 27134 430
rect 27186 378 27192 430
rect 27126 372 27192 378
rect 27232 418 27312 456
rect 27232 384 27238 418
rect 27272 384 27312 418
rect 27340 708 27400 940
rect 27454 943 27500 981
rect 27454 909 27460 943
rect 27494 909 27500 943
rect 27454 862 27500 909
rect 27542 981 27548 1015
rect 27582 981 27588 1015
rect 27542 943 27588 981
rect 27542 909 27548 943
rect 27582 909 27588 943
rect 27542 862 27588 909
rect 28696 1015 28742 1036
rect 28696 981 28702 1015
rect 28736 981 28742 1015
rect 28696 943 28742 981
rect 28696 909 28702 943
rect 28736 909 28742 943
rect 28696 862 28742 909
rect 28784 1042 28830 1062
rect 28964 1057 28993 1091
rect 29027 1057 29054 1091
rect 28784 1036 28852 1042
rect 28964 1036 29054 1057
rect 28784 1015 28792 1036
rect 28784 981 28790 1015
rect 28844 984 28852 1036
rect 28824 981 28852 984
rect 28784 976 28852 981
rect 29050 1000 29108 1002
rect 29256 1000 29290 1146
rect 29376 1143 29442 1154
rect 29376 1109 29392 1143
rect 29426 1109 29442 1143
rect 29376 1098 29442 1109
rect 29550 1144 30174 1176
rect 30262 1164 30340 2122
rect 30854 2113 30883 2122
rect 30917 2122 32771 2147
rect 30917 2113 30944 2122
rect 30854 2092 30944 2113
rect 30940 2056 30998 2058
rect 30940 2039 31002 2056
rect 30940 2005 30952 2039
rect 30986 2005 31002 2039
rect 30940 1996 31002 2005
rect 30440 1958 30806 1962
rect 30888 1958 30954 1966
rect 30440 1930 30848 1958
rect 30440 1892 30468 1930
rect 30762 1911 30848 1930
rect 30440 1884 30506 1892
rect 30440 1850 30455 1884
rect 30489 1850 30506 1884
rect 30440 1838 30506 1850
rect 30612 1888 30680 1894
rect 30612 1836 30622 1888
rect 30674 1836 30680 1888
rect 30612 1830 30680 1836
rect 30762 1877 30808 1911
rect 30842 1877 30848 1911
rect 30888 1906 30894 1958
rect 30946 1906 30954 1958
rect 30888 1898 30904 1906
rect 30762 1839 30848 1877
rect 30762 1805 30808 1839
rect 30842 1805 30848 1839
rect 30522 1776 30590 1782
rect 30522 1724 30530 1776
rect 30582 1724 30590 1776
rect 30522 1714 30590 1724
rect 30762 1758 30848 1805
rect 30898 1877 30904 1898
rect 30938 1898 30954 1906
rect 30994 1926 31322 1958
rect 30994 1911 31090 1926
rect 30938 1877 30944 1898
rect 30898 1839 30944 1877
rect 30898 1805 30904 1839
rect 30938 1805 30944 1839
rect 30898 1758 30944 1805
rect 30994 1877 31000 1911
rect 31034 1877 31090 1911
rect 31294 1890 31322 1926
rect 30994 1839 31090 1877
rect 30994 1805 31000 1839
rect 31034 1805 31090 1839
rect 31252 1882 31322 1890
rect 31252 1848 31267 1882
rect 31301 1848 31322 1882
rect 31252 1830 31322 1848
rect 31428 1890 31492 1896
rect 31428 1838 31434 1890
rect 31486 1838 31492 1890
rect 31428 1832 31492 1838
rect 30994 1758 31090 1805
rect 30420 1643 30696 1674
rect 30420 1609 30449 1643
rect 30483 1609 30541 1643
rect 30575 1609 30633 1643
rect 30667 1609 30696 1643
rect 30420 1578 30696 1609
rect 30762 1558 30812 1758
rect 30844 1711 30902 1726
rect 30844 1677 30856 1711
rect 30890 1677 30902 1711
rect 30844 1660 30902 1677
rect 30956 1630 31014 1648
rect 30956 1596 30968 1630
rect 31002 1596 31014 1630
rect 30956 1586 31014 1596
rect 31044 1558 31090 1758
rect 31340 1774 31404 1780
rect 31340 1722 31346 1774
rect 31398 1722 31404 1774
rect 31340 1716 31404 1722
rect 31234 1643 31510 1674
rect 31234 1609 31263 1643
rect 31297 1609 31355 1643
rect 31389 1609 31447 1643
rect 31481 1609 31510 1643
rect 31234 1606 31510 1609
rect 30402 1541 30466 1548
rect 30402 1508 30408 1541
rect 30460 1508 30466 1541
rect 30578 1541 30642 1548
rect 30578 1508 30584 1541
rect 30460 1489 30584 1508
rect 30636 1489 30642 1541
rect 30408 1480 30642 1489
rect 30762 1546 30864 1558
rect 30762 1512 30824 1546
rect 30858 1512 30864 1546
rect 30762 1474 30864 1512
rect 30914 1546 30960 1558
rect 30914 1512 30920 1546
rect 30954 1512 30960 1546
rect 30914 1492 30960 1512
rect 31010 1546 31090 1558
rect 31010 1512 31016 1546
rect 31050 1512 31090 1546
rect 30762 1442 30824 1474
rect 30558 1440 30824 1442
rect 30858 1440 30864 1474
rect 30558 1428 30864 1440
rect 30904 1486 30970 1492
rect 30904 1434 30912 1486
rect 30964 1434 30970 1486
rect 30904 1428 30970 1434
rect 31010 1474 31090 1512
rect 31010 1440 31016 1474
rect 31050 1440 31090 1474
rect 31206 1578 31510 1606
rect 31010 1428 31056 1440
rect 30558 1414 30812 1428
rect 30402 1408 30468 1414
rect 30402 1356 30410 1408
rect 30462 1356 30468 1408
rect 30402 1350 30468 1356
rect 29550 1141 29580 1144
rect 29632 1141 30174 1144
rect 29550 1107 29579 1141
rect 29632 1107 29671 1141
rect 29705 1107 29763 1141
rect 29797 1139 30174 1141
rect 29797 1107 29925 1139
rect 29550 1092 29580 1107
rect 29632 1105 29925 1107
rect 29959 1105 30017 1139
rect 30051 1105 30109 1139
rect 30143 1105 30174 1139
rect 29632 1092 30174 1105
rect 29550 1074 30174 1092
rect 30242 1150 30518 1164
rect 30242 1133 30434 1150
rect 30486 1133 30518 1150
rect 30242 1099 30271 1133
rect 30305 1099 30363 1133
rect 30397 1099 30434 1133
rect 30489 1099 30518 1133
rect 30242 1098 30434 1099
rect 30486 1098 30518 1099
rect 30242 1068 30518 1098
rect 30558 1064 30586 1414
rect 30858 1390 30922 1400
rect 30858 1356 30872 1390
rect 30906 1356 31178 1390
rect 30858 1338 30922 1356
rect 30774 1292 30846 1304
rect 30774 1240 30784 1292
rect 30836 1240 30846 1292
rect 30774 1228 30846 1240
rect 31144 1174 31178 1356
rect 31206 1274 31234 1578
rect 31206 1264 31274 1274
rect 31206 1230 31222 1264
rect 31256 1230 31274 1264
rect 31206 1216 31274 1230
rect 30618 1146 31178 1174
rect 30618 1143 30684 1146
rect 30618 1109 30634 1143
rect 30668 1109 30684 1143
rect 30618 1100 30684 1109
rect 30852 1091 30942 1112
rect 29050 983 29290 1000
rect 29334 1056 29400 1062
rect 29334 1004 29342 1056
rect 29394 1004 29400 1056
rect 29334 998 29348 1004
rect 28784 943 28830 976
rect 28784 909 28790 943
rect 28824 909 28830 943
rect 29050 949 29062 983
rect 29096 972 29290 983
rect 29342 981 29348 998
rect 29382 998 29400 1004
rect 29430 1015 29476 1062
rect 30558 1036 30630 1064
rect 29382 981 29388 998
rect 29096 949 29288 972
rect 29050 940 29288 949
rect 28784 862 28830 909
rect 28998 902 29064 910
rect 28912 898 28958 902
rect 28028 840 28100 844
rect 27488 815 27554 828
rect 27488 781 27504 815
rect 27538 781 27554 815
rect 27488 772 27554 781
rect 28028 788 28037 840
rect 28089 788 28100 840
rect 28028 776 28100 788
rect 28224 838 28298 858
rect 28872 855 28958 898
rect 28224 804 28236 838
rect 28270 804 28298 838
rect 28224 780 28298 804
rect 28334 844 28402 850
rect 28334 792 28341 844
rect 28393 838 28402 844
rect 28393 832 28486 838
rect 28393 798 28432 832
rect 28466 798 28486 832
rect 28393 792 28486 798
rect 28334 788 28486 792
rect 28730 815 28796 826
rect 28334 786 28402 788
rect 28730 781 28746 815
rect 28780 781 28796 815
rect 28730 768 28796 781
rect 28872 821 28918 855
rect 28952 821 28958 855
rect 28998 850 29004 902
rect 29056 850 29064 902
rect 28998 842 29014 850
rect 28872 783 28958 821
rect 28872 749 28918 783
rect 28952 749 28958 783
rect 27810 728 27868 742
rect 27810 708 27822 728
rect 27340 694 27822 708
rect 27856 694 27868 728
rect 27340 674 27868 694
rect 28872 702 28958 749
rect 29008 821 29014 842
rect 29048 842 29064 850
rect 29104 855 29200 902
rect 29048 821 29054 842
rect 29008 783 29054 821
rect 29008 749 29014 783
rect 29048 749 29054 783
rect 29008 702 29054 749
rect 29104 821 29110 855
rect 29144 821 29200 855
rect 29104 783 29200 821
rect 29104 749 29110 783
rect 29144 749 29200 783
rect 29104 702 29200 749
rect 27232 372 27278 384
rect 27340 344 27400 674
rect 28872 648 28922 702
rect 27446 624 27522 630
rect 27446 572 27454 624
rect 27506 572 27522 624
rect 27446 566 27522 572
rect 27662 597 28284 628
rect 27080 334 27400 344
rect 27080 300 27094 334
rect 27128 300 27400 334
rect 27080 282 27400 300
rect 27662 563 27691 597
rect 27725 563 27783 597
rect 27817 563 27875 597
rect 27909 595 28284 597
rect 27909 563 28037 595
rect 27662 561 28037 563
rect 28071 561 28129 595
rect 28163 561 28221 595
rect 28255 561 28284 595
rect 27662 530 28284 561
rect 28354 602 28630 620
rect 28354 589 28477 602
rect 28529 589 28630 602
rect 28706 598 28764 606
rect 28354 555 28383 589
rect 28417 555 28475 589
rect 28529 555 28567 589
rect 28601 555 28630 589
rect 28354 550 28477 555
rect 28529 550 28630 555
rect 27662 254 27760 530
rect 28354 524 28630 550
rect 28698 592 28772 598
rect 28698 540 28709 592
rect 28761 540 28772 592
rect 28852 582 28922 648
rect 28954 655 29012 670
rect 28954 621 28966 655
rect 29000 621 29012 655
rect 28954 604 29012 621
rect 28698 534 28772 540
rect 28706 528 28764 534
rect 28422 254 28506 524
rect 28872 502 28922 582
rect 29066 574 29124 592
rect 29066 540 29078 574
rect 29112 540 29124 574
rect 29066 530 29124 540
rect 29154 502 29200 702
rect 28872 490 28974 502
rect 28872 456 28934 490
rect 28968 456 28974 490
rect 28872 418 28974 456
rect 29024 490 29070 502
rect 29024 456 29030 490
rect 29064 456 29070 490
rect 29024 436 29070 456
rect 29120 490 29200 502
rect 29120 456 29126 490
rect 29160 456 29200 490
rect 28872 384 28934 418
rect 28968 384 28974 418
rect 28872 372 28974 384
rect 29014 430 29080 436
rect 29014 378 29022 430
rect 29074 378 29080 430
rect 29014 372 29080 378
rect 29120 418 29200 456
rect 29120 384 29126 418
rect 29160 384 29200 418
rect 29228 708 29288 940
rect 29342 943 29388 981
rect 29342 909 29348 943
rect 29382 909 29388 943
rect 29342 862 29388 909
rect 29430 981 29436 1015
rect 29470 981 29476 1015
rect 29430 943 29476 981
rect 29430 909 29436 943
rect 29470 909 29476 943
rect 29430 862 29476 909
rect 30584 1015 30630 1036
rect 30584 981 30590 1015
rect 30624 981 30630 1015
rect 30584 943 30630 981
rect 30584 909 30590 943
rect 30624 909 30630 943
rect 30584 862 30630 909
rect 30672 1042 30718 1062
rect 30852 1057 30881 1091
rect 30915 1057 30942 1091
rect 30672 1036 30740 1042
rect 30852 1036 30942 1057
rect 30672 1015 30680 1036
rect 30672 981 30678 1015
rect 30732 984 30740 1036
rect 30712 981 30740 984
rect 30672 976 30740 981
rect 30938 1000 30996 1002
rect 31144 1000 31178 1146
rect 31264 1143 31330 1154
rect 31264 1109 31280 1143
rect 31314 1109 31330 1143
rect 31264 1098 31330 1109
rect 31438 1144 32062 1176
rect 32150 1164 32228 2122
rect 32742 2113 32771 2122
rect 32805 2122 34659 2147
rect 32805 2113 32832 2122
rect 32742 2092 32832 2113
rect 32828 2056 32886 2058
rect 32828 2039 32890 2056
rect 32828 2005 32840 2039
rect 32874 2005 32890 2039
rect 32828 1996 32890 2005
rect 32328 1958 32694 1962
rect 32776 1958 32842 1966
rect 32328 1930 32736 1958
rect 32328 1892 32356 1930
rect 32650 1911 32736 1930
rect 32328 1884 32394 1892
rect 32328 1850 32343 1884
rect 32377 1850 32394 1884
rect 32328 1838 32394 1850
rect 32500 1888 32568 1894
rect 32500 1836 32510 1888
rect 32562 1836 32568 1888
rect 32500 1830 32568 1836
rect 32650 1877 32696 1911
rect 32730 1877 32736 1911
rect 32776 1906 32782 1958
rect 32834 1906 32842 1958
rect 32776 1898 32792 1906
rect 32650 1839 32736 1877
rect 32650 1805 32696 1839
rect 32730 1805 32736 1839
rect 32410 1776 32478 1782
rect 32410 1724 32418 1776
rect 32470 1724 32478 1776
rect 32410 1714 32478 1724
rect 32650 1758 32736 1805
rect 32786 1877 32792 1898
rect 32826 1898 32842 1906
rect 32882 1926 33210 1958
rect 32882 1911 32978 1926
rect 32826 1877 32832 1898
rect 32786 1839 32832 1877
rect 32786 1805 32792 1839
rect 32826 1805 32832 1839
rect 32786 1758 32832 1805
rect 32882 1877 32888 1911
rect 32922 1877 32978 1911
rect 33182 1890 33210 1926
rect 32882 1839 32978 1877
rect 32882 1805 32888 1839
rect 32922 1805 32978 1839
rect 33140 1882 33210 1890
rect 33140 1848 33155 1882
rect 33189 1848 33210 1882
rect 33140 1830 33210 1848
rect 33316 1890 33380 1896
rect 33316 1838 33322 1890
rect 33374 1838 33380 1890
rect 33316 1832 33380 1838
rect 32882 1758 32978 1805
rect 32308 1643 32584 1674
rect 32308 1609 32337 1643
rect 32371 1609 32429 1643
rect 32463 1609 32521 1643
rect 32555 1609 32584 1643
rect 32308 1578 32584 1609
rect 32650 1558 32700 1758
rect 32732 1711 32790 1726
rect 32732 1677 32744 1711
rect 32778 1677 32790 1711
rect 32732 1660 32790 1677
rect 32844 1630 32902 1648
rect 32844 1596 32856 1630
rect 32890 1596 32902 1630
rect 32844 1586 32902 1596
rect 32932 1558 32978 1758
rect 33228 1774 33292 1780
rect 33228 1722 33234 1774
rect 33286 1722 33292 1774
rect 33228 1716 33292 1722
rect 33122 1643 33398 1674
rect 33122 1609 33151 1643
rect 33185 1609 33243 1643
rect 33277 1609 33335 1643
rect 33369 1609 33398 1643
rect 33122 1606 33398 1609
rect 32290 1541 32354 1548
rect 32290 1508 32296 1541
rect 32348 1508 32354 1541
rect 32466 1541 32530 1548
rect 32466 1508 32472 1541
rect 32348 1489 32472 1508
rect 32524 1489 32530 1541
rect 32296 1480 32530 1489
rect 32650 1546 32752 1558
rect 32650 1512 32712 1546
rect 32746 1512 32752 1546
rect 32650 1474 32752 1512
rect 32802 1546 32848 1558
rect 32802 1512 32808 1546
rect 32842 1512 32848 1546
rect 32802 1492 32848 1512
rect 32898 1546 32978 1558
rect 32898 1512 32904 1546
rect 32938 1512 32978 1546
rect 32650 1442 32712 1474
rect 32446 1440 32712 1442
rect 32746 1440 32752 1474
rect 32446 1428 32752 1440
rect 32792 1486 32858 1492
rect 32792 1434 32800 1486
rect 32852 1434 32858 1486
rect 32792 1428 32858 1434
rect 32898 1474 32978 1512
rect 32898 1440 32904 1474
rect 32938 1440 32978 1474
rect 33094 1578 33398 1606
rect 32898 1428 32944 1440
rect 32446 1414 32700 1428
rect 32290 1408 32356 1414
rect 32290 1356 32298 1408
rect 32350 1356 32356 1408
rect 32290 1350 32356 1356
rect 31438 1141 31468 1144
rect 31520 1141 32062 1144
rect 31438 1107 31467 1141
rect 31520 1107 31559 1141
rect 31593 1107 31651 1141
rect 31685 1139 32062 1141
rect 31685 1107 31813 1139
rect 31438 1092 31468 1107
rect 31520 1105 31813 1107
rect 31847 1105 31905 1139
rect 31939 1105 31997 1139
rect 32031 1105 32062 1139
rect 31520 1092 32062 1105
rect 31438 1074 32062 1092
rect 32130 1150 32406 1164
rect 32130 1133 32322 1150
rect 32374 1133 32406 1150
rect 32130 1099 32159 1133
rect 32193 1099 32251 1133
rect 32285 1099 32322 1133
rect 32377 1099 32406 1133
rect 32130 1098 32322 1099
rect 32374 1098 32406 1099
rect 32130 1068 32406 1098
rect 32446 1064 32474 1414
rect 32746 1390 32810 1400
rect 32746 1356 32760 1390
rect 32794 1356 33066 1390
rect 32746 1338 32810 1356
rect 32662 1292 32734 1304
rect 32662 1240 32672 1292
rect 32724 1240 32734 1292
rect 32662 1228 32734 1240
rect 33032 1174 33066 1356
rect 33094 1274 33122 1578
rect 33094 1264 33162 1274
rect 33094 1230 33110 1264
rect 33144 1230 33162 1264
rect 33094 1216 33162 1230
rect 32506 1146 33066 1174
rect 32506 1143 32572 1146
rect 32506 1109 32522 1143
rect 32556 1109 32572 1143
rect 32506 1100 32572 1109
rect 32740 1091 32830 1112
rect 30938 983 31178 1000
rect 31222 1056 31288 1062
rect 31222 1004 31230 1056
rect 31282 1004 31288 1056
rect 31222 998 31236 1004
rect 30672 943 30718 976
rect 30672 909 30678 943
rect 30712 909 30718 943
rect 30938 949 30950 983
rect 30984 972 31178 983
rect 31230 981 31236 998
rect 31270 998 31288 1004
rect 31318 1015 31364 1062
rect 32446 1036 32518 1064
rect 31270 981 31276 998
rect 30984 949 31176 972
rect 30938 940 31176 949
rect 30672 862 30718 909
rect 30886 902 30952 910
rect 30800 898 30846 902
rect 29916 840 29988 844
rect 29376 815 29442 828
rect 29376 781 29392 815
rect 29426 781 29442 815
rect 29376 772 29442 781
rect 29916 788 29925 840
rect 29977 788 29988 840
rect 29916 776 29988 788
rect 30112 838 30186 858
rect 30760 855 30846 898
rect 30112 804 30124 838
rect 30158 804 30186 838
rect 30112 780 30186 804
rect 30222 844 30290 850
rect 30222 792 30229 844
rect 30281 838 30290 844
rect 30281 832 30374 838
rect 30281 798 30320 832
rect 30354 798 30374 832
rect 30281 792 30374 798
rect 30222 788 30374 792
rect 30618 815 30684 826
rect 30222 786 30290 788
rect 30618 781 30634 815
rect 30668 781 30684 815
rect 30618 768 30684 781
rect 30760 821 30806 855
rect 30840 821 30846 855
rect 30886 850 30892 902
rect 30944 850 30952 902
rect 30886 842 30902 850
rect 30760 783 30846 821
rect 30760 749 30806 783
rect 30840 749 30846 783
rect 29698 728 29756 742
rect 29698 708 29710 728
rect 29228 694 29710 708
rect 29744 694 29756 728
rect 29228 674 29756 694
rect 30760 702 30846 749
rect 30896 821 30902 842
rect 30936 842 30952 850
rect 30992 855 31088 902
rect 30936 821 30942 842
rect 30896 783 30942 821
rect 30896 749 30902 783
rect 30936 749 30942 783
rect 30896 702 30942 749
rect 30992 821 30998 855
rect 31032 821 31088 855
rect 30992 783 31088 821
rect 30992 749 30998 783
rect 31032 749 31088 783
rect 30992 702 31088 749
rect 29120 372 29166 384
rect 29228 344 29288 674
rect 30760 648 30810 702
rect 29334 624 29410 630
rect 29334 572 29342 624
rect 29394 572 29410 624
rect 29334 566 29410 572
rect 29550 597 30172 628
rect 28968 334 29288 344
rect 28968 300 28982 334
rect 29016 300 29288 334
rect 28968 282 29288 300
rect 29550 563 29579 597
rect 29613 563 29671 597
rect 29705 563 29763 597
rect 29797 595 30172 597
rect 29797 563 29925 595
rect 29550 561 29925 563
rect 29959 561 30017 595
rect 30051 561 30109 595
rect 30143 561 30172 595
rect 29550 530 30172 561
rect 30242 602 30518 620
rect 30242 589 30365 602
rect 30417 589 30518 602
rect 30594 598 30652 606
rect 30242 555 30271 589
rect 30305 555 30363 589
rect 30417 555 30455 589
rect 30489 555 30518 589
rect 30242 550 30365 555
rect 30417 550 30518 555
rect 29550 254 29648 530
rect 30242 524 30518 550
rect 30586 592 30660 598
rect 30586 540 30597 592
rect 30649 540 30660 592
rect 30740 582 30810 648
rect 30842 655 30900 670
rect 30842 621 30854 655
rect 30888 621 30900 655
rect 30842 604 30900 621
rect 30586 534 30660 540
rect 30594 528 30652 534
rect 30310 254 30394 524
rect 30760 502 30810 582
rect 30954 574 31012 592
rect 30954 540 30966 574
rect 31000 540 31012 574
rect 30954 530 31012 540
rect 31042 502 31088 702
rect 30760 490 30862 502
rect 30760 456 30822 490
rect 30856 456 30862 490
rect 30760 418 30862 456
rect 30912 490 30958 502
rect 30912 456 30918 490
rect 30952 456 30958 490
rect 30912 436 30958 456
rect 31008 490 31088 502
rect 31008 456 31014 490
rect 31048 456 31088 490
rect 30760 384 30822 418
rect 30856 384 30862 418
rect 30760 372 30862 384
rect 30902 430 30968 436
rect 30902 378 30910 430
rect 30962 378 30968 430
rect 30902 372 30968 378
rect 31008 418 31088 456
rect 31008 384 31014 418
rect 31048 384 31088 418
rect 31116 708 31176 940
rect 31230 943 31276 981
rect 31230 909 31236 943
rect 31270 909 31276 943
rect 31230 862 31276 909
rect 31318 981 31324 1015
rect 31358 981 31364 1015
rect 31318 943 31364 981
rect 31318 909 31324 943
rect 31358 909 31364 943
rect 31318 862 31364 909
rect 32472 1015 32518 1036
rect 32472 981 32478 1015
rect 32512 981 32518 1015
rect 32472 943 32518 981
rect 32472 909 32478 943
rect 32512 909 32518 943
rect 32472 862 32518 909
rect 32560 1042 32606 1062
rect 32740 1057 32769 1091
rect 32803 1057 32830 1091
rect 32560 1036 32628 1042
rect 32740 1036 32830 1057
rect 32560 1015 32568 1036
rect 32560 981 32566 1015
rect 32620 984 32628 1036
rect 32600 981 32628 984
rect 32560 976 32628 981
rect 32826 1000 32884 1002
rect 33032 1000 33066 1146
rect 33152 1143 33218 1154
rect 33152 1109 33168 1143
rect 33202 1109 33218 1143
rect 33152 1098 33218 1109
rect 33326 1144 33950 1176
rect 34038 1164 34116 2122
rect 34630 2113 34659 2122
rect 34693 2122 36547 2147
rect 34693 2113 34720 2122
rect 34630 2092 34720 2113
rect 34716 2056 34774 2058
rect 34716 2039 34778 2056
rect 34716 2005 34728 2039
rect 34762 2005 34778 2039
rect 34716 1996 34778 2005
rect 34216 1958 34582 1962
rect 34664 1958 34730 1966
rect 34216 1930 34624 1958
rect 34216 1892 34244 1930
rect 34538 1911 34624 1930
rect 34216 1884 34282 1892
rect 34216 1850 34231 1884
rect 34265 1850 34282 1884
rect 34216 1838 34282 1850
rect 34388 1888 34456 1894
rect 34388 1836 34398 1888
rect 34450 1836 34456 1888
rect 34388 1830 34456 1836
rect 34538 1877 34584 1911
rect 34618 1877 34624 1911
rect 34664 1906 34670 1958
rect 34722 1906 34730 1958
rect 34664 1898 34680 1906
rect 34538 1839 34624 1877
rect 34538 1805 34584 1839
rect 34618 1805 34624 1839
rect 34298 1776 34366 1782
rect 34298 1724 34306 1776
rect 34358 1724 34366 1776
rect 34298 1714 34366 1724
rect 34538 1758 34624 1805
rect 34674 1877 34680 1898
rect 34714 1898 34730 1906
rect 34770 1926 35098 1958
rect 34770 1911 34866 1926
rect 34714 1877 34720 1898
rect 34674 1839 34720 1877
rect 34674 1805 34680 1839
rect 34714 1805 34720 1839
rect 34674 1758 34720 1805
rect 34770 1877 34776 1911
rect 34810 1877 34866 1911
rect 35070 1890 35098 1926
rect 34770 1839 34866 1877
rect 34770 1805 34776 1839
rect 34810 1805 34866 1839
rect 35028 1882 35098 1890
rect 35028 1848 35043 1882
rect 35077 1848 35098 1882
rect 35028 1830 35098 1848
rect 35204 1890 35268 1896
rect 35204 1838 35210 1890
rect 35262 1838 35268 1890
rect 35204 1832 35268 1838
rect 34770 1758 34866 1805
rect 34196 1643 34472 1674
rect 34196 1609 34225 1643
rect 34259 1609 34317 1643
rect 34351 1609 34409 1643
rect 34443 1609 34472 1643
rect 34196 1578 34472 1609
rect 34538 1558 34588 1758
rect 34620 1711 34678 1726
rect 34620 1677 34632 1711
rect 34666 1677 34678 1711
rect 34620 1660 34678 1677
rect 34732 1630 34790 1648
rect 34732 1596 34744 1630
rect 34778 1596 34790 1630
rect 34732 1586 34790 1596
rect 34820 1558 34866 1758
rect 35116 1774 35180 1780
rect 35116 1722 35122 1774
rect 35174 1722 35180 1774
rect 35116 1716 35180 1722
rect 35010 1643 35286 1674
rect 35010 1609 35039 1643
rect 35073 1609 35131 1643
rect 35165 1609 35223 1643
rect 35257 1609 35286 1643
rect 35010 1606 35286 1609
rect 34178 1541 34242 1548
rect 34178 1508 34184 1541
rect 34236 1508 34242 1541
rect 34354 1541 34418 1548
rect 34354 1508 34360 1541
rect 34236 1489 34360 1508
rect 34412 1489 34418 1541
rect 34184 1480 34418 1489
rect 34538 1546 34640 1558
rect 34538 1512 34600 1546
rect 34634 1512 34640 1546
rect 34538 1474 34640 1512
rect 34690 1546 34736 1558
rect 34690 1512 34696 1546
rect 34730 1512 34736 1546
rect 34690 1492 34736 1512
rect 34786 1546 34866 1558
rect 34786 1512 34792 1546
rect 34826 1512 34866 1546
rect 34538 1442 34600 1474
rect 34334 1440 34600 1442
rect 34634 1440 34640 1474
rect 34334 1428 34640 1440
rect 34680 1486 34746 1492
rect 34680 1434 34688 1486
rect 34740 1434 34746 1486
rect 34680 1428 34746 1434
rect 34786 1474 34866 1512
rect 34786 1440 34792 1474
rect 34826 1440 34866 1474
rect 34982 1578 35286 1606
rect 34786 1428 34832 1440
rect 34334 1414 34588 1428
rect 34178 1408 34244 1414
rect 34178 1356 34186 1408
rect 34238 1356 34244 1408
rect 34178 1350 34244 1356
rect 33326 1141 33356 1144
rect 33408 1141 33950 1144
rect 33326 1107 33355 1141
rect 33408 1107 33447 1141
rect 33481 1107 33539 1141
rect 33573 1139 33950 1141
rect 33573 1107 33701 1139
rect 33326 1092 33356 1107
rect 33408 1105 33701 1107
rect 33735 1105 33793 1139
rect 33827 1105 33885 1139
rect 33919 1105 33950 1139
rect 33408 1092 33950 1105
rect 33326 1074 33950 1092
rect 34018 1150 34294 1164
rect 34018 1133 34210 1150
rect 34262 1133 34294 1150
rect 34018 1099 34047 1133
rect 34081 1099 34139 1133
rect 34173 1099 34210 1133
rect 34265 1099 34294 1133
rect 34018 1098 34210 1099
rect 34262 1098 34294 1099
rect 34018 1068 34294 1098
rect 34334 1064 34362 1414
rect 34634 1390 34698 1400
rect 34634 1356 34648 1390
rect 34682 1356 34954 1390
rect 34634 1338 34698 1356
rect 34550 1292 34622 1304
rect 34550 1240 34560 1292
rect 34612 1240 34622 1292
rect 34550 1228 34622 1240
rect 34920 1174 34954 1356
rect 34982 1274 35010 1578
rect 34982 1264 35050 1274
rect 34982 1230 34998 1264
rect 35032 1230 35050 1264
rect 34982 1216 35050 1230
rect 34394 1146 34954 1174
rect 34394 1143 34460 1146
rect 34394 1109 34410 1143
rect 34444 1109 34460 1143
rect 34394 1100 34460 1109
rect 34628 1091 34718 1112
rect 32826 983 33066 1000
rect 33110 1056 33176 1062
rect 33110 1004 33118 1056
rect 33170 1004 33176 1056
rect 33110 998 33124 1004
rect 32560 943 32606 976
rect 32560 909 32566 943
rect 32600 909 32606 943
rect 32826 949 32838 983
rect 32872 972 33066 983
rect 33118 981 33124 998
rect 33158 998 33176 1004
rect 33206 1015 33252 1062
rect 34334 1036 34406 1064
rect 33158 981 33164 998
rect 32872 949 33064 972
rect 32826 940 33064 949
rect 32560 862 32606 909
rect 32774 902 32840 910
rect 32688 898 32734 902
rect 31804 840 31876 844
rect 31264 815 31330 828
rect 31264 781 31280 815
rect 31314 781 31330 815
rect 31264 772 31330 781
rect 31804 788 31813 840
rect 31865 788 31876 840
rect 31804 776 31876 788
rect 32000 838 32074 858
rect 32648 855 32734 898
rect 32000 804 32012 838
rect 32046 804 32074 838
rect 32000 780 32074 804
rect 32110 844 32178 850
rect 32110 792 32117 844
rect 32169 838 32178 844
rect 32169 832 32262 838
rect 32169 798 32208 832
rect 32242 798 32262 832
rect 32169 792 32262 798
rect 32110 788 32262 792
rect 32506 815 32572 826
rect 32110 786 32178 788
rect 32506 781 32522 815
rect 32556 781 32572 815
rect 32506 768 32572 781
rect 32648 821 32694 855
rect 32728 821 32734 855
rect 32774 850 32780 902
rect 32832 850 32840 902
rect 32774 842 32790 850
rect 32648 783 32734 821
rect 32648 749 32694 783
rect 32728 749 32734 783
rect 31586 728 31644 742
rect 31586 708 31598 728
rect 31116 694 31598 708
rect 31632 694 31644 728
rect 31116 674 31644 694
rect 32648 702 32734 749
rect 32784 821 32790 842
rect 32824 842 32840 850
rect 32880 855 32976 902
rect 32824 821 32830 842
rect 32784 783 32830 821
rect 32784 749 32790 783
rect 32824 749 32830 783
rect 32784 702 32830 749
rect 32880 821 32886 855
rect 32920 821 32976 855
rect 32880 783 32976 821
rect 32880 749 32886 783
rect 32920 749 32976 783
rect 32880 702 32976 749
rect 31008 372 31054 384
rect 31116 344 31176 674
rect 32648 648 32698 702
rect 31222 624 31298 630
rect 31222 572 31230 624
rect 31282 572 31298 624
rect 31222 566 31298 572
rect 31438 597 32060 628
rect 30856 334 31176 344
rect 30856 300 30870 334
rect 30904 300 31176 334
rect 30856 282 31176 300
rect 31438 563 31467 597
rect 31501 563 31559 597
rect 31593 563 31651 597
rect 31685 595 32060 597
rect 31685 563 31813 595
rect 31438 561 31813 563
rect 31847 561 31905 595
rect 31939 561 31997 595
rect 32031 561 32060 595
rect 31438 530 32060 561
rect 32130 602 32406 620
rect 32130 589 32253 602
rect 32305 589 32406 602
rect 32482 598 32540 606
rect 32130 555 32159 589
rect 32193 555 32251 589
rect 32305 555 32343 589
rect 32377 555 32406 589
rect 32130 550 32253 555
rect 32305 550 32406 555
rect 31438 254 31536 530
rect 32130 524 32406 550
rect 32474 592 32548 598
rect 32474 540 32485 592
rect 32537 540 32548 592
rect 32628 582 32698 648
rect 32730 655 32788 670
rect 32730 621 32742 655
rect 32776 621 32788 655
rect 32730 604 32788 621
rect 32474 534 32548 540
rect 32482 528 32540 534
rect 32198 254 32282 524
rect 32648 502 32698 582
rect 32842 574 32900 592
rect 32842 540 32854 574
rect 32888 540 32900 574
rect 32842 530 32900 540
rect 32930 502 32976 702
rect 32648 490 32750 502
rect 32648 456 32710 490
rect 32744 456 32750 490
rect 32648 418 32750 456
rect 32800 490 32846 502
rect 32800 456 32806 490
rect 32840 456 32846 490
rect 32800 436 32846 456
rect 32896 490 32976 502
rect 32896 456 32902 490
rect 32936 456 32976 490
rect 32648 384 32710 418
rect 32744 384 32750 418
rect 32648 372 32750 384
rect 32790 430 32856 436
rect 32790 378 32798 430
rect 32850 378 32856 430
rect 32790 372 32856 378
rect 32896 418 32976 456
rect 32896 384 32902 418
rect 32936 384 32976 418
rect 33004 708 33064 940
rect 33118 943 33164 981
rect 33118 909 33124 943
rect 33158 909 33164 943
rect 33118 862 33164 909
rect 33206 981 33212 1015
rect 33246 981 33252 1015
rect 33206 943 33252 981
rect 33206 909 33212 943
rect 33246 909 33252 943
rect 33206 862 33252 909
rect 34360 1015 34406 1036
rect 34360 981 34366 1015
rect 34400 981 34406 1015
rect 34360 943 34406 981
rect 34360 909 34366 943
rect 34400 909 34406 943
rect 34360 862 34406 909
rect 34448 1042 34494 1062
rect 34628 1057 34657 1091
rect 34691 1057 34718 1091
rect 34448 1036 34516 1042
rect 34628 1036 34718 1057
rect 34448 1015 34456 1036
rect 34448 981 34454 1015
rect 34508 984 34516 1036
rect 34488 981 34516 984
rect 34448 976 34516 981
rect 34714 1000 34772 1002
rect 34920 1000 34954 1146
rect 35040 1143 35106 1154
rect 35040 1109 35056 1143
rect 35090 1109 35106 1143
rect 35040 1098 35106 1109
rect 35214 1144 35838 1176
rect 35926 1164 36004 2122
rect 36518 2113 36547 2122
rect 36581 2122 38435 2147
rect 36581 2113 36608 2122
rect 36518 2092 36608 2113
rect 36604 2056 36662 2058
rect 36604 2039 36666 2056
rect 36604 2005 36616 2039
rect 36650 2005 36666 2039
rect 36604 1996 36666 2005
rect 36104 1958 36470 1962
rect 36552 1958 36618 1966
rect 36104 1930 36512 1958
rect 36104 1892 36132 1930
rect 36426 1911 36512 1930
rect 36104 1884 36170 1892
rect 36104 1850 36119 1884
rect 36153 1850 36170 1884
rect 36104 1838 36170 1850
rect 36276 1888 36344 1894
rect 36276 1836 36286 1888
rect 36338 1836 36344 1888
rect 36276 1830 36344 1836
rect 36426 1877 36472 1911
rect 36506 1877 36512 1911
rect 36552 1906 36558 1958
rect 36610 1906 36618 1958
rect 36552 1898 36568 1906
rect 36426 1839 36512 1877
rect 36426 1805 36472 1839
rect 36506 1805 36512 1839
rect 36186 1776 36254 1782
rect 36186 1724 36194 1776
rect 36246 1724 36254 1776
rect 36186 1714 36254 1724
rect 36426 1758 36512 1805
rect 36562 1877 36568 1898
rect 36602 1898 36618 1906
rect 36658 1926 36986 1958
rect 36658 1911 36754 1926
rect 36602 1877 36608 1898
rect 36562 1839 36608 1877
rect 36562 1805 36568 1839
rect 36602 1805 36608 1839
rect 36562 1758 36608 1805
rect 36658 1877 36664 1911
rect 36698 1877 36754 1911
rect 36958 1890 36986 1926
rect 36658 1839 36754 1877
rect 36658 1805 36664 1839
rect 36698 1805 36754 1839
rect 36916 1882 36986 1890
rect 36916 1848 36931 1882
rect 36965 1848 36986 1882
rect 36916 1830 36986 1848
rect 37092 1890 37156 1896
rect 37092 1838 37098 1890
rect 37150 1838 37156 1890
rect 37092 1832 37156 1838
rect 36658 1758 36754 1805
rect 36084 1643 36360 1674
rect 36084 1609 36113 1643
rect 36147 1609 36205 1643
rect 36239 1609 36297 1643
rect 36331 1609 36360 1643
rect 36084 1578 36360 1609
rect 36426 1558 36476 1758
rect 36508 1711 36566 1726
rect 36508 1677 36520 1711
rect 36554 1677 36566 1711
rect 36508 1660 36566 1677
rect 36620 1630 36678 1648
rect 36620 1596 36632 1630
rect 36666 1596 36678 1630
rect 36620 1586 36678 1596
rect 36708 1558 36754 1758
rect 37004 1774 37068 1780
rect 37004 1722 37010 1774
rect 37062 1722 37068 1774
rect 37004 1716 37068 1722
rect 36898 1643 37174 1674
rect 36898 1609 36927 1643
rect 36961 1609 37019 1643
rect 37053 1609 37111 1643
rect 37145 1609 37174 1643
rect 36898 1606 37174 1609
rect 36066 1541 36130 1548
rect 36066 1508 36072 1541
rect 36124 1508 36130 1541
rect 36242 1541 36306 1548
rect 36242 1508 36248 1541
rect 36124 1489 36248 1508
rect 36300 1489 36306 1541
rect 36072 1480 36306 1489
rect 36426 1546 36528 1558
rect 36426 1512 36488 1546
rect 36522 1512 36528 1546
rect 36426 1474 36528 1512
rect 36578 1546 36624 1558
rect 36578 1512 36584 1546
rect 36618 1512 36624 1546
rect 36578 1492 36624 1512
rect 36674 1546 36754 1558
rect 36674 1512 36680 1546
rect 36714 1512 36754 1546
rect 36426 1442 36488 1474
rect 36222 1440 36488 1442
rect 36522 1440 36528 1474
rect 36222 1428 36528 1440
rect 36568 1486 36634 1492
rect 36568 1434 36576 1486
rect 36628 1434 36634 1486
rect 36568 1428 36634 1434
rect 36674 1474 36754 1512
rect 36674 1440 36680 1474
rect 36714 1440 36754 1474
rect 36870 1578 37174 1606
rect 36674 1428 36720 1440
rect 36222 1414 36476 1428
rect 36066 1408 36132 1414
rect 36066 1356 36074 1408
rect 36126 1356 36132 1408
rect 36066 1350 36132 1356
rect 35214 1141 35244 1144
rect 35296 1141 35838 1144
rect 35214 1107 35243 1141
rect 35296 1107 35335 1141
rect 35369 1107 35427 1141
rect 35461 1139 35838 1141
rect 35461 1107 35589 1139
rect 35214 1092 35244 1107
rect 35296 1105 35589 1107
rect 35623 1105 35681 1139
rect 35715 1105 35773 1139
rect 35807 1105 35838 1139
rect 35296 1092 35838 1105
rect 35214 1074 35838 1092
rect 35906 1150 36182 1164
rect 35906 1133 36098 1150
rect 36150 1133 36182 1150
rect 35906 1099 35935 1133
rect 35969 1099 36027 1133
rect 36061 1099 36098 1133
rect 36153 1099 36182 1133
rect 35906 1098 36098 1099
rect 36150 1098 36182 1099
rect 35906 1068 36182 1098
rect 36222 1064 36250 1414
rect 36522 1390 36586 1400
rect 36522 1356 36536 1390
rect 36570 1356 36842 1390
rect 36522 1338 36586 1356
rect 36438 1292 36510 1304
rect 36438 1240 36448 1292
rect 36500 1240 36510 1292
rect 36438 1228 36510 1240
rect 36808 1174 36842 1356
rect 36870 1274 36898 1578
rect 36870 1264 36938 1274
rect 36870 1230 36886 1264
rect 36920 1230 36938 1264
rect 36870 1216 36938 1230
rect 36282 1146 36842 1174
rect 36282 1143 36348 1146
rect 36282 1109 36298 1143
rect 36332 1109 36348 1143
rect 36282 1100 36348 1109
rect 36516 1091 36606 1112
rect 34714 983 34954 1000
rect 34998 1056 35064 1062
rect 34998 1004 35006 1056
rect 35058 1004 35064 1056
rect 34998 998 35012 1004
rect 34448 943 34494 976
rect 34448 909 34454 943
rect 34488 909 34494 943
rect 34714 949 34726 983
rect 34760 972 34954 983
rect 35006 981 35012 998
rect 35046 998 35064 1004
rect 35094 1015 35140 1062
rect 36222 1036 36294 1064
rect 35046 981 35052 998
rect 34760 949 34952 972
rect 34714 940 34952 949
rect 34448 862 34494 909
rect 34662 902 34728 910
rect 34576 898 34622 902
rect 33692 840 33764 844
rect 33152 815 33218 828
rect 33152 781 33168 815
rect 33202 781 33218 815
rect 33152 772 33218 781
rect 33692 788 33701 840
rect 33753 788 33764 840
rect 33692 776 33764 788
rect 33888 838 33962 858
rect 34536 855 34622 898
rect 33888 804 33900 838
rect 33934 804 33962 838
rect 33888 780 33962 804
rect 33998 844 34066 850
rect 33998 792 34005 844
rect 34057 838 34066 844
rect 34057 832 34150 838
rect 34057 798 34096 832
rect 34130 798 34150 832
rect 34057 792 34150 798
rect 33998 788 34150 792
rect 34394 815 34460 826
rect 33998 786 34066 788
rect 34394 781 34410 815
rect 34444 781 34460 815
rect 34394 768 34460 781
rect 34536 821 34582 855
rect 34616 821 34622 855
rect 34662 850 34668 902
rect 34720 850 34728 902
rect 34662 842 34678 850
rect 34536 783 34622 821
rect 34536 749 34582 783
rect 34616 749 34622 783
rect 33474 728 33532 742
rect 33474 708 33486 728
rect 33004 694 33486 708
rect 33520 694 33532 728
rect 33004 674 33532 694
rect 34536 702 34622 749
rect 34672 821 34678 842
rect 34712 842 34728 850
rect 34768 855 34864 902
rect 34712 821 34718 842
rect 34672 783 34718 821
rect 34672 749 34678 783
rect 34712 749 34718 783
rect 34672 702 34718 749
rect 34768 821 34774 855
rect 34808 821 34864 855
rect 34768 783 34864 821
rect 34768 749 34774 783
rect 34808 749 34864 783
rect 34768 702 34864 749
rect 32896 372 32942 384
rect 33004 344 33064 674
rect 34536 648 34586 702
rect 33110 624 33186 630
rect 33110 572 33118 624
rect 33170 572 33186 624
rect 33110 566 33186 572
rect 33326 597 33948 628
rect 32744 334 33064 344
rect 32744 300 32758 334
rect 32792 300 33064 334
rect 32744 282 33064 300
rect 33326 563 33355 597
rect 33389 563 33447 597
rect 33481 563 33539 597
rect 33573 595 33948 597
rect 33573 563 33701 595
rect 33326 561 33701 563
rect 33735 561 33793 595
rect 33827 561 33885 595
rect 33919 561 33948 595
rect 33326 530 33948 561
rect 34018 602 34294 620
rect 34018 589 34141 602
rect 34193 589 34294 602
rect 34370 598 34428 606
rect 34018 555 34047 589
rect 34081 555 34139 589
rect 34193 555 34231 589
rect 34265 555 34294 589
rect 34018 550 34141 555
rect 34193 550 34294 555
rect 33326 254 33424 530
rect 34018 524 34294 550
rect 34362 592 34436 598
rect 34362 540 34373 592
rect 34425 540 34436 592
rect 34516 582 34586 648
rect 34618 655 34676 670
rect 34618 621 34630 655
rect 34664 621 34676 655
rect 34618 604 34676 621
rect 34362 534 34436 540
rect 34370 528 34428 534
rect 34086 254 34170 524
rect 34536 502 34586 582
rect 34730 574 34788 592
rect 34730 540 34742 574
rect 34776 540 34788 574
rect 34730 530 34788 540
rect 34818 502 34864 702
rect 34536 490 34638 502
rect 34536 456 34598 490
rect 34632 456 34638 490
rect 34536 418 34638 456
rect 34688 490 34734 502
rect 34688 456 34694 490
rect 34728 456 34734 490
rect 34688 436 34734 456
rect 34784 490 34864 502
rect 34784 456 34790 490
rect 34824 456 34864 490
rect 34536 384 34598 418
rect 34632 384 34638 418
rect 34536 372 34638 384
rect 34678 430 34744 436
rect 34678 378 34686 430
rect 34738 378 34744 430
rect 34678 372 34744 378
rect 34784 418 34864 456
rect 34784 384 34790 418
rect 34824 384 34864 418
rect 34892 708 34952 940
rect 35006 943 35052 981
rect 35006 909 35012 943
rect 35046 909 35052 943
rect 35006 862 35052 909
rect 35094 981 35100 1015
rect 35134 981 35140 1015
rect 35094 943 35140 981
rect 35094 909 35100 943
rect 35134 909 35140 943
rect 35094 862 35140 909
rect 36248 1015 36294 1036
rect 36248 981 36254 1015
rect 36288 981 36294 1015
rect 36248 943 36294 981
rect 36248 909 36254 943
rect 36288 909 36294 943
rect 36248 862 36294 909
rect 36336 1042 36382 1062
rect 36516 1057 36545 1091
rect 36579 1057 36606 1091
rect 36336 1036 36404 1042
rect 36516 1036 36606 1057
rect 36336 1015 36344 1036
rect 36336 981 36342 1015
rect 36396 984 36404 1036
rect 36376 981 36404 984
rect 36336 976 36404 981
rect 36602 1000 36660 1002
rect 36808 1000 36842 1146
rect 36928 1143 36994 1154
rect 36928 1109 36944 1143
rect 36978 1109 36994 1143
rect 36928 1098 36994 1109
rect 37102 1144 37726 1176
rect 37814 1164 37892 2122
rect 38406 2113 38435 2122
rect 38469 2122 40323 2147
rect 38469 2113 38496 2122
rect 38406 2092 38496 2113
rect 38492 2056 38550 2058
rect 38492 2039 38554 2056
rect 38492 2005 38504 2039
rect 38538 2005 38554 2039
rect 38492 1996 38554 2005
rect 37992 1958 38358 1962
rect 38440 1958 38506 1966
rect 37992 1930 38400 1958
rect 37992 1892 38020 1930
rect 38314 1911 38400 1930
rect 37992 1884 38058 1892
rect 37992 1850 38007 1884
rect 38041 1850 38058 1884
rect 37992 1838 38058 1850
rect 38164 1888 38232 1894
rect 38164 1836 38174 1888
rect 38226 1836 38232 1888
rect 38164 1830 38232 1836
rect 38314 1877 38360 1911
rect 38394 1877 38400 1911
rect 38440 1906 38446 1958
rect 38498 1906 38506 1958
rect 38440 1898 38456 1906
rect 38314 1839 38400 1877
rect 38314 1805 38360 1839
rect 38394 1805 38400 1839
rect 38074 1776 38142 1782
rect 38074 1724 38082 1776
rect 38134 1724 38142 1776
rect 38074 1714 38142 1724
rect 38314 1758 38400 1805
rect 38450 1877 38456 1898
rect 38490 1898 38506 1906
rect 38546 1926 38874 1958
rect 38546 1911 38642 1926
rect 38490 1877 38496 1898
rect 38450 1839 38496 1877
rect 38450 1805 38456 1839
rect 38490 1805 38496 1839
rect 38450 1758 38496 1805
rect 38546 1877 38552 1911
rect 38586 1877 38642 1911
rect 38846 1890 38874 1926
rect 38546 1839 38642 1877
rect 38546 1805 38552 1839
rect 38586 1805 38642 1839
rect 38804 1882 38874 1890
rect 38804 1848 38819 1882
rect 38853 1848 38874 1882
rect 38804 1830 38874 1848
rect 38980 1890 39044 1896
rect 38980 1838 38986 1890
rect 39038 1838 39044 1890
rect 38980 1832 39044 1838
rect 38546 1758 38642 1805
rect 37972 1643 38248 1674
rect 37972 1609 38001 1643
rect 38035 1609 38093 1643
rect 38127 1609 38185 1643
rect 38219 1609 38248 1643
rect 37972 1578 38248 1609
rect 38314 1558 38364 1758
rect 38396 1711 38454 1726
rect 38396 1677 38408 1711
rect 38442 1677 38454 1711
rect 38396 1660 38454 1677
rect 38508 1630 38566 1648
rect 38508 1596 38520 1630
rect 38554 1596 38566 1630
rect 38508 1586 38566 1596
rect 38596 1558 38642 1758
rect 38892 1774 38956 1780
rect 38892 1722 38898 1774
rect 38950 1722 38956 1774
rect 38892 1716 38956 1722
rect 38786 1643 39062 1674
rect 38786 1609 38815 1643
rect 38849 1609 38907 1643
rect 38941 1609 38999 1643
rect 39033 1609 39062 1643
rect 38786 1606 39062 1609
rect 37954 1541 38018 1548
rect 37954 1508 37960 1541
rect 38012 1508 38018 1541
rect 38130 1541 38194 1548
rect 38130 1508 38136 1541
rect 38012 1489 38136 1508
rect 38188 1489 38194 1541
rect 37960 1480 38194 1489
rect 38314 1546 38416 1558
rect 38314 1512 38376 1546
rect 38410 1512 38416 1546
rect 38314 1474 38416 1512
rect 38466 1546 38512 1558
rect 38466 1512 38472 1546
rect 38506 1512 38512 1546
rect 38466 1492 38512 1512
rect 38562 1546 38642 1558
rect 38562 1512 38568 1546
rect 38602 1512 38642 1546
rect 38314 1442 38376 1474
rect 38110 1440 38376 1442
rect 38410 1440 38416 1474
rect 38110 1428 38416 1440
rect 38456 1486 38522 1492
rect 38456 1434 38464 1486
rect 38516 1434 38522 1486
rect 38456 1428 38522 1434
rect 38562 1474 38642 1512
rect 38562 1440 38568 1474
rect 38602 1440 38642 1474
rect 38758 1578 39062 1606
rect 38562 1428 38608 1440
rect 38110 1414 38364 1428
rect 37954 1408 38020 1414
rect 37954 1356 37962 1408
rect 38014 1356 38020 1408
rect 37954 1350 38020 1356
rect 37102 1141 37132 1144
rect 37184 1141 37726 1144
rect 37102 1107 37131 1141
rect 37184 1107 37223 1141
rect 37257 1107 37315 1141
rect 37349 1139 37726 1141
rect 37349 1107 37477 1139
rect 37102 1092 37132 1107
rect 37184 1105 37477 1107
rect 37511 1105 37569 1139
rect 37603 1105 37661 1139
rect 37695 1105 37726 1139
rect 37184 1092 37726 1105
rect 37102 1074 37726 1092
rect 37794 1150 38070 1164
rect 37794 1133 37986 1150
rect 38038 1133 38070 1150
rect 37794 1099 37823 1133
rect 37857 1099 37915 1133
rect 37949 1099 37986 1133
rect 38041 1099 38070 1133
rect 37794 1098 37986 1099
rect 38038 1098 38070 1099
rect 37794 1068 38070 1098
rect 38110 1064 38138 1414
rect 38410 1390 38474 1400
rect 38410 1356 38424 1390
rect 38458 1356 38730 1390
rect 38410 1338 38474 1356
rect 38326 1292 38398 1304
rect 38326 1240 38336 1292
rect 38388 1240 38398 1292
rect 38326 1228 38398 1240
rect 38696 1174 38730 1356
rect 38758 1274 38786 1578
rect 38758 1264 38826 1274
rect 38758 1230 38774 1264
rect 38808 1230 38826 1264
rect 38758 1216 38826 1230
rect 38170 1146 38730 1174
rect 38170 1143 38236 1146
rect 38170 1109 38186 1143
rect 38220 1109 38236 1143
rect 38170 1100 38236 1109
rect 38404 1091 38494 1112
rect 36602 983 36842 1000
rect 36886 1056 36952 1062
rect 36886 1004 36894 1056
rect 36946 1004 36952 1056
rect 36886 998 36900 1004
rect 36336 943 36382 976
rect 36336 909 36342 943
rect 36376 909 36382 943
rect 36602 949 36614 983
rect 36648 972 36842 983
rect 36894 981 36900 998
rect 36934 998 36952 1004
rect 36982 1015 37028 1062
rect 38110 1036 38182 1064
rect 36934 981 36940 998
rect 36648 949 36840 972
rect 36602 940 36840 949
rect 36336 862 36382 909
rect 36550 902 36616 910
rect 36464 898 36510 902
rect 35580 840 35652 844
rect 35040 815 35106 828
rect 35040 781 35056 815
rect 35090 781 35106 815
rect 35040 772 35106 781
rect 35580 788 35589 840
rect 35641 788 35652 840
rect 35580 776 35652 788
rect 35776 838 35850 858
rect 36424 855 36510 898
rect 35776 804 35788 838
rect 35822 804 35850 838
rect 35776 780 35850 804
rect 35886 844 35954 850
rect 35886 792 35893 844
rect 35945 838 35954 844
rect 35945 832 36038 838
rect 35945 798 35984 832
rect 36018 798 36038 832
rect 35945 792 36038 798
rect 35886 788 36038 792
rect 36282 815 36348 826
rect 35886 786 35954 788
rect 36282 781 36298 815
rect 36332 781 36348 815
rect 36282 768 36348 781
rect 36424 821 36470 855
rect 36504 821 36510 855
rect 36550 850 36556 902
rect 36608 850 36616 902
rect 36550 842 36566 850
rect 36424 783 36510 821
rect 36424 749 36470 783
rect 36504 749 36510 783
rect 35362 728 35420 742
rect 35362 708 35374 728
rect 34892 694 35374 708
rect 35408 694 35420 728
rect 34892 674 35420 694
rect 36424 702 36510 749
rect 36560 821 36566 842
rect 36600 842 36616 850
rect 36656 855 36752 902
rect 36600 821 36606 842
rect 36560 783 36606 821
rect 36560 749 36566 783
rect 36600 749 36606 783
rect 36560 702 36606 749
rect 36656 821 36662 855
rect 36696 821 36752 855
rect 36656 783 36752 821
rect 36656 749 36662 783
rect 36696 749 36752 783
rect 36656 702 36752 749
rect 34784 372 34830 384
rect 34892 344 34952 674
rect 36424 648 36474 702
rect 34998 624 35074 630
rect 34998 572 35006 624
rect 35058 572 35074 624
rect 34998 566 35074 572
rect 35214 597 35836 628
rect 34632 334 34952 344
rect 34632 300 34646 334
rect 34680 300 34952 334
rect 34632 282 34952 300
rect 35214 563 35243 597
rect 35277 563 35335 597
rect 35369 563 35427 597
rect 35461 595 35836 597
rect 35461 563 35589 595
rect 35214 561 35589 563
rect 35623 561 35681 595
rect 35715 561 35773 595
rect 35807 561 35836 595
rect 35214 530 35836 561
rect 35906 602 36182 620
rect 35906 589 36029 602
rect 36081 589 36182 602
rect 36258 598 36316 606
rect 35906 555 35935 589
rect 35969 555 36027 589
rect 36081 555 36119 589
rect 36153 555 36182 589
rect 35906 550 36029 555
rect 36081 550 36182 555
rect 35214 254 35312 530
rect 35906 524 36182 550
rect 36250 592 36324 598
rect 36250 540 36261 592
rect 36313 540 36324 592
rect 36404 582 36474 648
rect 36506 655 36564 670
rect 36506 621 36518 655
rect 36552 621 36564 655
rect 36506 604 36564 621
rect 36250 534 36324 540
rect 36258 528 36316 534
rect 35974 254 36058 524
rect 36424 502 36474 582
rect 36618 574 36676 592
rect 36618 540 36630 574
rect 36664 540 36676 574
rect 36618 530 36676 540
rect 36706 502 36752 702
rect 36424 490 36526 502
rect 36424 456 36486 490
rect 36520 456 36526 490
rect 36424 418 36526 456
rect 36576 490 36622 502
rect 36576 456 36582 490
rect 36616 456 36622 490
rect 36576 436 36622 456
rect 36672 490 36752 502
rect 36672 456 36678 490
rect 36712 456 36752 490
rect 36424 384 36486 418
rect 36520 384 36526 418
rect 36424 372 36526 384
rect 36566 430 36632 436
rect 36566 378 36574 430
rect 36626 378 36632 430
rect 36566 372 36632 378
rect 36672 418 36752 456
rect 36672 384 36678 418
rect 36712 384 36752 418
rect 36780 708 36840 940
rect 36894 943 36940 981
rect 36894 909 36900 943
rect 36934 909 36940 943
rect 36894 862 36940 909
rect 36982 981 36988 1015
rect 37022 981 37028 1015
rect 36982 943 37028 981
rect 36982 909 36988 943
rect 37022 909 37028 943
rect 36982 862 37028 909
rect 38136 1015 38182 1036
rect 38136 981 38142 1015
rect 38176 981 38182 1015
rect 38136 943 38182 981
rect 38136 909 38142 943
rect 38176 909 38182 943
rect 38136 862 38182 909
rect 38224 1042 38270 1062
rect 38404 1057 38433 1091
rect 38467 1057 38494 1091
rect 38224 1036 38292 1042
rect 38404 1036 38494 1057
rect 38224 1015 38232 1036
rect 38224 981 38230 1015
rect 38284 984 38292 1036
rect 38264 981 38292 984
rect 38224 976 38292 981
rect 38490 1000 38548 1002
rect 38696 1000 38730 1146
rect 38816 1143 38882 1154
rect 38816 1109 38832 1143
rect 38866 1109 38882 1143
rect 38816 1098 38882 1109
rect 38990 1144 39614 1176
rect 39702 1164 39780 2122
rect 40294 2113 40323 2122
rect 40357 2122 42211 2147
rect 40357 2113 40384 2122
rect 40294 2092 40384 2113
rect 40380 2056 40438 2058
rect 40380 2039 40442 2056
rect 40380 2005 40392 2039
rect 40426 2005 40442 2039
rect 40380 1996 40442 2005
rect 39880 1958 40246 1962
rect 40328 1958 40394 1966
rect 39880 1930 40288 1958
rect 39880 1892 39908 1930
rect 40202 1911 40288 1930
rect 39880 1884 39946 1892
rect 39880 1850 39895 1884
rect 39929 1850 39946 1884
rect 39880 1838 39946 1850
rect 40052 1888 40120 1894
rect 40052 1836 40062 1888
rect 40114 1836 40120 1888
rect 40052 1830 40120 1836
rect 40202 1877 40248 1911
rect 40282 1877 40288 1911
rect 40328 1906 40334 1958
rect 40386 1906 40394 1958
rect 40328 1898 40344 1906
rect 40202 1839 40288 1877
rect 40202 1805 40248 1839
rect 40282 1805 40288 1839
rect 39962 1776 40030 1782
rect 39962 1724 39970 1776
rect 40022 1724 40030 1776
rect 39962 1714 40030 1724
rect 40202 1758 40288 1805
rect 40338 1877 40344 1898
rect 40378 1898 40394 1906
rect 40434 1926 40762 1958
rect 40434 1911 40530 1926
rect 40378 1877 40384 1898
rect 40338 1839 40384 1877
rect 40338 1805 40344 1839
rect 40378 1805 40384 1839
rect 40338 1758 40384 1805
rect 40434 1877 40440 1911
rect 40474 1877 40530 1911
rect 40734 1890 40762 1926
rect 40434 1839 40530 1877
rect 40434 1805 40440 1839
rect 40474 1805 40530 1839
rect 40692 1882 40762 1890
rect 40692 1848 40707 1882
rect 40741 1848 40762 1882
rect 40692 1830 40762 1848
rect 40868 1890 40932 1896
rect 40868 1838 40874 1890
rect 40926 1838 40932 1890
rect 40868 1832 40932 1838
rect 40434 1758 40530 1805
rect 39860 1643 40136 1674
rect 39860 1609 39889 1643
rect 39923 1609 39981 1643
rect 40015 1609 40073 1643
rect 40107 1609 40136 1643
rect 39860 1578 40136 1609
rect 40202 1558 40252 1758
rect 40284 1711 40342 1726
rect 40284 1677 40296 1711
rect 40330 1677 40342 1711
rect 40284 1660 40342 1677
rect 40396 1630 40454 1648
rect 40396 1596 40408 1630
rect 40442 1596 40454 1630
rect 40396 1586 40454 1596
rect 40484 1558 40530 1758
rect 40780 1774 40844 1780
rect 40780 1722 40786 1774
rect 40838 1722 40844 1774
rect 40780 1716 40844 1722
rect 40674 1643 40950 1674
rect 40674 1609 40703 1643
rect 40737 1609 40795 1643
rect 40829 1609 40887 1643
rect 40921 1609 40950 1643
rect 40674 1606 40950 1609
rect 39842 1541 39906 1548
rect 39842 1508 39848 1541
rect 39900 1508 39906 1541
rect 40018 1541 40082 1548
rect 40018 1508 40024 1541
rect 39900 1489 40024 1508
rect 40076 1489 40082 1541
rect 39848 1480 40082 1489
rect 40202 1546 40304 1558
rect 40202 1512 40264 1546
rect 40298 1512 40304 1546
rect 40202 1474 40304 1512
rect 40354 1546 40400 1558
rect 40354 1512 40360 1546
rect 40394 1512 40400 1546
rect 40354 1492 40400 1512
rect 40450 1546 40530 1558
rect 40450 1512 40456 1546
rect 40490 1512 40530 1546
rect 40202 1442 40264 1474
rect 39998 1440 40264 1442
rect 40298 1440 40304 1474
rect 39998 1428 40304 1440
rect 40344 1486 40410 1492
rect 40344 1434 40352 1486
rect 40404 1434 40410 1486
rect 40344 1428 40410 1434
rect 40450 1474 40530 1512
rect 40450 1440 40456 1474
rect 40490 1440 40530 1474
rect 40646 1578 40950 1606
rect 40450 1428 40496 1440
rect 39998 1414 40252 1428
rect 39842 1408 39908 1414
rect 39842 1356 39850 1408
rect 39902 1356 39908 1408
rect 39842 1350 39908 1356
rect 38990 1141 39020 1144
rect 39072 1141 39614 1144
rect 38990 1107 39019 1141
rect 39072 1107 39111 1141
rect 39145 1107 39203 1141
rect 39237 1139 39614 1141
rect 39237 1107 39365 1139
rect 38990 1092 39020 1107
rect 39072 1105 39365 1107
rect 39399 1105 39457 1139
rect 39491 1105 39549 1139
rect 39583 1105 39614 1139
rect 39072 1092 39614 1105
rect 38990 1074 39614 1092
rect 39682 1150 39958 1164
rect 39682 1133 39874 1150
rect 39926 1133 39958 1150
rect 39682 1099 39711 1133
rect 39745 1099 39803 1133
rect 39837 1099 39874 1133
rect 39929 1099 39958 1133
rect 39682 1098 39874 1099
rect 39926 1098 39958 1099
rect 39682 1068 39958 1098
rect 39998 1064 40026 1414
rect 40298 1390 40362 1400
rect 40298 1356 40312 1390
rect 40346 1356 40618 1390
rect 40298 1338 40362 1356
rect 40214 1292 40286 1304
rect 40214 1240 40224 1292
rect 40276 1240 40286 1292
rect 40214 1228 40286 1240
rect 40584 1174 40618 1356
rect 40646 1274 40674 1578
rect 40646 1264 40714 1274
rect 40646 1230 40662 1264
rect 40696 1230 40714 1264
rect 40646 1216 40714 1230
rect 40058 1146 40618 1174
rect 40058 1143 40124 1146
rect 40058 1109 40074 1143
rect 40108 1109 40124 1143
rect 40058 1100 40124 1109
rect 40292 1091 40382 1112
rect 38490 983 38730 1000
rect 38774 1056 38840 1062
rect 38774 1004 38782 1056
rect 38834 1004 38840 1056
rect 38774 998 38788 1004
rect 38224 943 38270 976
rect 38224 909 38230 943
rect 38264 909 38270 943
rect 38490 949 38502 983
rect 38536 972 38730 983
rect 38782 981 38788 998
rect 38822 998 38840 1004
rect 38870 1015 38916 1062
rect 39998 1036 40070 1064
rect 38822 981 38828 998
rect 38536 949 38728 972
rect 38490 940 38728 949
rect 38224 862 38270 909
rect 38438 902 38504 910
rect 38352 898 38398 902
rect 37468 840 37540 844
rect 36928 815 36994 828
rect 36928 781 36944 815
rect 36978 781 36994 815
rect 36928 772 36994 781
rect 37468 788 37477 840
rect 37529 788 37540 840
rect 37468 776 37540 788
rect 37664 838 37738 858
rect 38312 855 38398 898
rect 37664 804 37676 838
rect 37710 804 37738 838
rect 37664 780 37738 804
rect 37774 844 37842 850
rect 37774 792 37781 844
rect 37833 838 37842 844
rect 37833 832 37926 838
rect 37833 798 37872 832
rect 37906 798 37926 832
rect 37833 792 37926 798
rect 37774 788 37926 792
rect 38170 815 38236 826
rect 37774 786 37842 788
rect 38170 781 38186 815
rect 38220 781 38236 815
rect 38170 768 38236 781
rect 38312 821 38358 855
rect 38392 821 38398 855
rect 38438 850 38444 902
rect 38496 850 38504 902
rect 38438 842 38454 850
rect 38312 783 38398 821
rect 38312 749 38358 783
rect 38392 749 38398 783
rect 37250 728 37308 742
rect 37250 708 37262 728
rect 36780 694 37262 708
rect 37296 694 37308 728
rect 36780 674 37308 694
rect 38312 702 38398 749
rect 38448 821 38454 842
rect 38488 842 38504 850
rect 38544 855 38640 902
rect 38488 821 38494 842
rect 38448 783 38494 821
rect 38448 749 38454 783
rect 38488 749 38494 783
rect 38448 702 38494 749
rect 38544 821 38550 855
rect 38584 821 38640 855
rect 38544 783 38640 821
rect 38544 749 38550 783
rect 38584 749 38640 783
rect 38544 702 38640 749
rect 36672 372 36718 384
rect 36780 344 36840 674
rect 38312 648 38362 702
rect 36886 624 36962 630
rect 36886 572 36894 624
rect 36946 572 36962 624
rect 36886 566 36962 572
rect 37102 597 37724 628
rect 36520 334 36840 344
rect 36520 300 36534 334
rect 36568 300 36840 334
rect 36520 282 36840 300
rect 37102 563 37131 597
rect 37165 563 37223 597
rect 37257 563 37315 597
rect 37349 595 37724 597
rect 37349 563 37477 595
rect 37102 561 37477 563
rect 37511 561 37569 595
rect 37603 561 37661 595
rect 37695 561 37724 595
rect 37102 530 37724 561
rect 37794 602 38070 620
rect 37794 589 37917 602
rect 37969 589 38070 602
rect 38146 598 38204 606
rect 37794 555 37823 589
rect 37857 555 37915 589
rect 37969 555 38007 589
rect 38041 555 38070 589
rect 37794 550 37917 555
rect 37969 550 38070 555
rect 37102 254 37200 530
rect 37794 524 38070 550
rect 38138 592 38212 598
rect 38138 540 38149 592
rect 38201 540 38212 592
rect 38292 582 38362 648
rect 38394 655 38452 670
rect 38394 621 38406 655
rect 38440 621 38452 655
rect 38394 604 38452 621
rect 38138 534 38212 540
rect 38146 528 38204 534
rect 37862 254 37946 524
rect 38312 502 38362 582
rect 38506 574 38564 592
rect 38506 540 38518 574
rect 38552 540 38564 574
rect 38506 530 38564 540
rect 38594 502 38640 702
rect 38312 490 38414 502
rect 38312 456 38374 490
rect 38408 456 38414 490
rect 38312 418 38414 456
rect 38464 490 38510 502
rect 38464 456 38470 490
rect 38504 456 38510 490
rect 38464 436 38510 456
rect 38560 490 38640 502
rect 38560 456 38566 490
rect 38600 456 38640 490
rect 38312 384 38374 418
rect 38408 384 38414 418
rect 38312 372 38414 384
rect 38454 430 38520 436
rect 38454 378 38462 430
rect 38514 378 38520 430
rect 38454 372 38520 378
rect 38560 418 38640 456
rect 38560 384 38566 418
rect 38600 384 38640 418
rect 38668 708 38728 940
rect 38782 943 38828 981
rect 38782 909 38788 943
rect 38822 909 38828 943
rect 38782 862 38828 909
rect 38870 981 38876 1015
rect 38910 981 38916 1015
rect 38870 943 38916 981
rect 38870 909 38876 943
rect 38910 909 38916 943
rect 38870 862 38916 909
rect 40024 1015 40070 1036
rect 40024 981 40030 1015
rect 40064 981 40070 1015
rect 40024 943 40070 981
rect 40024 909 40030 943
rect 40064 909 40070 943
rect 40024 862 40070 909
rect 40112 1042 40158 1062
rect 40292 1057 40321 1091
rect 40355 1057 40382 1091
rect 40112 1036 40180 1042
rect 40292 1036 40382 1057
rect 40112 1015 40120 1036
rect 40112 981 40118 1015
rect 40172 984 40180 1036
rect 40152 981 40180 984
rect 40112 976 40180 981
rect 40378 1000 40436 1002
rect 40584 1000 40618 1146
rect 40704 1143 40770 1154
rect 40704 1109 40720 1143
rect 40754 1109 40770 1143
rect 40704 1098 40770 1109
rect 40878 1144 41502 1176
rect 41590 1164 41668 2122
rect 42182 2113 42211 2122
rect 42245 2122 44099 2147
rect 42245 2113 42272 2122
rect 42182 2092 42272 2113
rect 42268 2056 42326 2058
rect 42268 2039 42330 2056
rect 42268 2005 42280 2039
rect 42314 2005 42330 2039
rect 42268 1996 42330 2005
rect 41768 1958 42134 1962
rect 42216 1958 42282 1966
rect 41768 1930 42176 1958
rect 41768 1892 41796 1930
rect 42090 1911 42176 1930
rect 41768 1884 41834 1892
rect 41768 1850 41783 1884
rect 41817 1850 41834 1884
rect 41768 1838 41834 1850
rect 41940 1888 42008 1894
rect 41940 1836 41950 1888
rect 42002 1836 42008 1888
rect 41940 1830 42008 1836
rect 42090 1877 42136 1911
rect 42170 1877 42176 1911
rect 42216 1906 42222 1958
rect 42274 1906 42282 1958
rect 42216 1898 42232 1906
rect 42090 1839 42176 1877
rect 42090 1805 42136 1839
rect 42170 1805 42176 1839
rect 41850 1776 41918 1782
rect 41850 1724 41858 1776
rect 41910 1724 41918 1776
rect 41850 1714 41918 1724
rect 42090 1758 42176 1805
rect 42226 1877 42232 1898
rect 42266 1898 42282 1906
rect 42322 1926 42650 1958
rect 42322 1911 42418 1926
rect 42266 1877 42272 1898
rect 42226 1839 42272 1877
rect 42226 1805 42232 1839
rect 42266 1805 42272 1839
rect 42226 1758 42272 1805
rect 42322 1877 42328 1911
rect 42362 1877 42418 1911
rect 42622 1890 42650 1926
rect 42322 1839 42418 1877
rect 42322 1805 42328 1839
rect 42362 1805 42418 1839
rect 42580 1882 42650 1890
rect 42580 1848 42595 1882
rect 42629 1848 42650 1882
rect 42580 1830 42650 1848
rect 42756 1890 42820 1896
rect 42756 1838 42762 1890
rect 42814 1838 42820 1890
rect 42756 1832 42820 1838
rect 42322 1758 42418 1805
rect 41748 1643 42024 1674
rect 41748 1609 41777 1643
rect 41811 1609 41869 1643
rect 41903 1609 41961 1643
rect 41995 1609 42024 1643
rect 41748 1578 42024 1609
rect 42090 1558 42140 1758
rect 42172 1711 42230 1726
rect 42172 1677 42184 1711
rect 42218 1677 42230 1711
rect 42172 1660 42230 1677
rect 42284 1630 42342 1648
rect 42284 1596 42296 1630
rect 42330 1596 42342 1630
rect 42284 1586 42342 1596
rect 42372 1558 42418 1758
rect 42668 1774 42732 1780
rect 42668 1722 42674 1774
rect 42726 1722 42732 1774
rect 42668 1716 42732 1722
rect 42562 1643 42838 1674
rect 42562 1609 42591 1643
rect 42625 1609 42683 1643
rect 42717 1609 42775 1643
rect 42809 1609 42838 1643
rect 42562 1606 42838 1609
rect 41730 1541 41794 1548
rect 41730 1508 41736 1541
rect 41788 1508 41794 1541
rect 41906 1541 41970 1548
rect 41906 1508 41912 1541
rect 41788 1489 41912 1508
rect 41964 1489 41970 1541
rect 41736 1480 41970 1489
rect 42090 1546 42192 1558
rect 42090 1512 42152 1546
rect 42186 1512 42192 1546
rect 42090 1474 42192 1512
rect 42242 1546 42288 1558
rect 42242 1512 42248 1546
rect 42282 1512 42288 1546
rect 42242 1492 42288 1512
rect 42338 1546 42418 1558
rect 42338 1512 42344 1546
rect 42378 1512 42418 1546
rect 42090 1442 42152 1474
rect 41886 1440 42152 1442
rect 42186 1440 42192 1474
rect 41886 1428 42192 1440
rect 42232 1486 42298 1492
rect 42232 1434 42240 1486
rect 42292 1434 42298 1486
rect 42232 1428 42298 1434
rect 42338 1474 42418 1512
rect 42338 1440 42344 1474
rect 42378 1440 42418 1474
rect 42534 1578 42838 1606
rect 42338 1428 42384 1440
rect 41886 1414 42140 1428
rect 41730 1408 41796 1414
rect 41730 1356 41738 1408
rect 41790 1356 41796 1408
rect 41730 1350 41796 1356
rect 40878 1141 40908 1144
rect 40960 1141 41502 1144
rect 40878 1107 40907 1141
rect 40960 1107 40999 1141
rect 41033 1107 41091 1141
rect 41125 1139 41502 1141
rect 41125 1107 41253 1139
rect 40878 1092 40908 1107
rect 40960 1105 41253 1107
rect 41287 1105 41345 1139
rect 41379 1105 41437 1139
rect 41471 1105 41502 1139
rect 40960 1092 41502 1105
rect 40878 1074 41502 1092
rect 41570 1150 41846 1164
rect 41570 1133 41762 1150
rect 41814 1133 41846 1150
rect 41570 1099 41599 1133
rect 41633 1099 41691 1133
rect 41725 1099 41762 1133
rect 41817 1099 41846 1133
rect 41570 1098 41762 1099
rect 41814 1098 41846 1099
rect 41570 1068 41846 1098
rect 41886 1064 41914 1414
rect 42186 1390 42250 1400
rect 42186 1356 42200 1390
rect 42234 1356 42506 1390
rect 42186 1338 42250 1356
rect 42102 1292 42174 1304
rect 42102 1240 42112 1292
rect 42164 1240 42174 1292
rect 42102 1228 42174 1240
rect 42472 1174 42506 1356
rect 42534 1274 42562 1578
rect 42534 1264 42602 1274
rect 42534 1230 42550 1264
rect 42584 1230 42602 1264
rect 42534 1216 42602 1230
rect 41946 1146 42506 1174
rect 41946 1143 42012 1146
rect 41946 1109 41962 1143
rect 41996 1109 42012 1143
rect 41946 1100 42012 1109
rect 42180 1091 42270 1112
rect 40378 983 40618 1000
rect 40662 1056 40728 1062
rect 40662 1004 40670 1056
rect 40722 1004 40728 1056
rect 40662 998 40676 1004
rect 40112 943 40158 976
rect 40112 909 40118 943
rect 40152 909 40158 943
rect 40378 949 40390 983
rect 40424 972 40618 983
rect 40670 981 40676 998
rect 40710 998 40728 1004
rect 40758 1015 40804 1062
rect 41886 1036 41958 1064
rect 40710 981 40716 998
rect 40424 949 40616 972
rect 40378 940 40616 949
rect 40112 862 40158 909
rect 40326 902 40392 910
rect 40240 898 40286 902
rect 39356 840 39428 844
rect 38816 815 38882 828
rect 38816 781 38832 815
rect 38866 781 38882 815
rect 38816 772 38882 781
rect 39356 788 39365 840
rect 39417 788 39428 840
rect 39356 776 39428 788
rect 39552 838 39626 858
rect 40200 855 40286 898
rect 39552 804 39564 838
rect 39598 804 39626 838
rect 39552 780 39626 804
rect 39662 844 39730 850
rect 39662 792 39669 844
rect 39721 838 39730 844
rect 39721 832 39814 838
rect 39721 798 39760 832
rect 39794 798 39814 832
rect 39721 792 39814 798
rect 39662 788 39814 792
rect 40058 815 40124 826
rect 39662 786 39730 788
rect 40058 781 40074 815
rect 40108 781 40124 815
rect 40058 768 40124 781
rect 40200 821 40246 855
rect 40280 821 40286 855
rect 40326 850 40332 902
rect 40384 850 40392 902
rect 40326 842 40342 850
rect 40200 783 40286 821
rect 40200 749 40246 783
rect 40280 749 40286 783
rect 39138 728 39196 742
rect 39138 708 39150 728
rect 38668 694 39150 708
rect 39184 694 39196 728
rect 38668 674 39196 694
rect 40200 702 40286 749
rect 40336 821 40342 842
rect 40376 842 40392 850
rect 40432 855 40528 902
rect 40376 821 40382 842
rect 40336 783 40382 821
rect 40336 749 40342 783
rect 40376 749 40382 783
rect 40336 702 40382 749
rect 40432 821 40438 855
rect 40472 821 40528 855
rect 40432 783 40528 821
rect 40432 749 40438 783
rect 40472 749 40528 783
rect 40432 702 40528 749
rect 38560 372 38606 384
rect 38668 344 38728 674
rect 40200 648 40250 702
rect 38774 624 38850 630
rect 38774 572 38782 624
rect 38834 572 38850 624
rect 38774 566 38850 572
rect 38990 597 39612 628
rect 38408 334 38728 344
rect 38408 300 38422 334
rect 38456 300 38728 334
rect 38408 282 38728 300
rect 38990 563 39019 597
rect 39053 563 39111 597
rect 39145 563 39203 597
rect 39237 595 39612 597
rect 39237 563 39365 595
rect 38990 561 39365 563
rect 39399 561 39457 595
rect 39491 561 39549 595
rect 39583 561 39612 595
rect 38990 530 39612 561
rect 39682 602 39958 620
rect 39682 589 39805 602
rect 39857 589 39958 602
rect 40034 598 40092 606
rect 39682 555 39711 589
rect 39745 555 39803 589
rect 39857 555 39895 589
rect 39929 555 39958 589
rect 39682 550 39805 555
rect 39857 550 39958 555
rect 38990 254 39088 530
rect 39682 524 39958 550
rect 40026 592 40100 598
rect 40026 540 40037 592
rect 40089 540 40100 592
rect 40180 582 40250 648
rect 40282 655 40340 670
rect 40282 621 40294 655
rect 40328 621 40340 655
rect 40282 604 40340 621
rect 40026 534 40100 540
rect 40034 528 40092 534
rect 39750 254 39834 524
rect 40200 502 40250 582
rect 40394 574 40452 592
rect 40394 540 40406 574
rect 40440 540 40452 574
rect 40394 530 40452 540
rect 40482 502 40528 702
rect 40200 490 40302 502
rect 40200 456 40262 490
rect 40296 456 40302 490
rect 40200 418 40302 456
rect 40352 490 40398 502
rect 40352 456 40358 490
rect 40392 456 40398 490
rect 40352 436 40398 456
rect 40448 490 40528 502
rect 40448 456 40454 490
rect 40488 456 40528 490
rect 40200 384 40262 418
rect 40296 384 40302 418
rect 40200 372 40302 384
rect 40342 430 40408 436
rect 40342 378 40350 430
rect 40402 378 40408 430
rect 40342 372 40408 378
rect 40448 418 40528 456
rect 40448 384 40454 418
rect 40488 384 40528 418
rect 40556 708 40616 940
rect 40670 943 40716 981
rect 40670 909 40676 943
rect 40710 909 40716 943
rect 40670 862 40716 909
rect 40758 981 40764 1015
rect 40798 981 40804 1015
rect 40758 943 40804 981
rect 40758 909 40764 943
rect 40798 909 40804 943
rect 40758 862 40804 909
rect 41912 1015 41958 1036
rect 41912 981 41918 1015
rect 41952 981 41958 1015
rect 41912 943 41958 981
rect 41912 909 41918 943
rect 41952 909 41958 943
rect 41912 862 41958 909
rect 42000 1042 42046 1062
rect 42180 1057 42209 1091
rect 42243 1057 42270 1091
rect 42000 1036 42068 1042
rect 42180 1036 42270 1057
rect 42000 1015 42008 1036
rect 42000 981 42006 1015
rect 42060 984 42068 1036
rect 42040 981 42068 984
rect 42000 976 42068 981
rect 42266 1000 42324 1002
rect 42472 1000 42506 1146
rect 42592 1143 42658 1154
rect 42592 1109 42608 1143
rect 42642 1109 42658 1143
rect 42592 1098 42658 1109
rect 42766 1144 43390 1176
rect 43478 1164 43556 2122
rect 44070 2113 44099 2122
rect 44133 2122 45981 2147
rect 44133 2113 44160 2122
rect 44070 2092 44160 2113
rect 44156 2056 44214 2058
rect 44156 2039 44218 2056
rect 44156 2005 44168 2039
rect 44202 2005 44218 2039
rect 44156 1996 44218 2005
rect 43656 1958 44022 1962
rect 44104 1958 44170 1966
rect 43656 1930 44064 1958
rect 43656 1892 43684 1930
rect 43978 1911 44064 1930
rect 43656 1884 43722 1892
rect 43656 1850 43671 1884
rect 43705 1850 43722 1884
rect 43656 1838 43722 1850
rect 43828 1888 43896 1894
rect 43828 1836 43838 1888
rect 43890 1836 43896 1888
rect 43828 1830 43896 1836
rect 43978 1877 44024 1911
rect 44058 1877 44064 1911
rect 44104 1906 44110 1958
rect 44162 1906 44170 1958
rect 44104 1898 44120 1906
rect 43978 1839 44064 1877
rect 43978 1805 44024 1839
rect 44058 1805 44064 1839
rect 43738 1776 43806 1782
rect 43738 1724 43746 1776
rect 43798 1724 43806 1776
rect 43738 1714 43806 1724
rect 43978 1758 44064 1805
rect 44114 1877 44120 1898
rect 44154 1898 44170 1906
rect 44210 1926 44538 1958
rect 44210 1911 44306 1926
rect 44154 1877 44160 1898
rect 44114 1839 44160 1877
rect 44114 1805 44120 1839
rect 44154 1805 44160 1839
rect 44114 1758 44160 1805
rect 44210 1877 44216 1911
rect 44250 1877 44306 1911
rect 44510 1890 44538 1926
rect 44210 1839 44306 1877
rect 44210 1805 44216 1839
rect 44250 1805 44306 1839
rect 44468 1882 44538 1890
rect 44468 1848 44483 1882
rect 44517 1848 44538 1882
rect 44468 1830 44538 1848
rect 44644 1890 44708 1896
rect 44644 1838 44650 1890
rect 44702 1838 44708 1890
rect 44644 1832 44708 1838
rect 44210 1758 44306 1805
rect 43636 1643 43912 1674
rect 43636 1609 43665 1643
rect 43699 1609 43757 1643
rect 43791 1609 43849 1643
rect 43883 1609 43912 1643
rect 43636 1578 43912 1609
rect 43978 1558 44028 1758
rect 44060 1711 44118 1726
rect 44060 1677 44072 1711
rect 44106 1677 44118 1711
rect 44060 1660 44118 1677
rect 44172 1630 44230 1648
rect 44172 1596 44184 1630
rect 44218 1596 44230 1630
rect 44172 1586 44230 1596
rect 44260 1558 44306 1758
rect 44556 1774 44620 1780
rect 44556 1722 44562 1774
rect 44614 1722 44620 1774
rect 44556 1716 44620 1722
rect 44450 1643 44726 1674
rect 44450 1609 44479 1643
rect 44513 1609 44571 1643
rect 44605 1609 44663 1643
rect 44697 1609 44726 1643
rect 44450 1606 44726 1609
rect 43618 1541 43682 1548
rect 43618 1508 43624 1541
rect 43676 1508 43682 1541
rect 43794 1541 43858 1548
rect 43794 1508 43800 1541
rect 43676 1489 43800 1508
rect 43852 1489 43858 1541
rect 43624 1480 43858 1489
rect 43978 1546 44080 1558
rect 43978 1512 44040 1546
rect 44074 1512 44080 1546
rect 43978 1474 44080 1512
rect 44130 1546 44176 1558
rect 44130 1512 44136 1546
rect 44170 1512 44176 1546
rect 44130 1492 44176 1512
rect 44226 1546 44306 1558
rect 44226 1512 44232 1546
rect 44266 1512 44306 1546
rect 43978 1442 44040 1474
rect 43774 1440 44040 1442
rect 44074 1440 44080 1474
rect 43774 1428 44080 1440
rect 44120 1486 44186 1492
rect 44120 1434 44128 1486
rect 44180 1434 44186 1486
rect 44120 1428 44186 1434
rect 44226 1474 44306 1512
rect 44226 1440 44232 1474
rect 44266 1440 44306 1474
rect 44422 1578 44726 1606
rect 44226 1428 44272 1440
rect 43774 1414 44028 1428
rect 43618 1408 43684 1414
rect 43618 1356 43626 1408
rect 43678 1356 43684 1408
rect 43618 1350 43684 1356
rect 42766 1141 42796 1144
rect 42848 1141 43390 1144
rect 42766 1107 42795 1141
rect 42848 1107 42887 1141
rect 42921 1107 42979 1141
rect 43013 1139 43390 1141
rect 43013 1107 43141 1139
rect 42766 1092 42796 1107
rect 42848 1105 43141 1107
rect 43175 1105 43233 1139
rect 43267 1105 43325 1139
rect 43359 1105 43390 1139
rect 42848 1092 43390 1105
rect 42766 1074 43390 1092
rect 43458 1150 43734 1164
rect 43458 1133 43650 1150
rect 43702 1133 43734 1150
rect 43458 1099 43487 1133
rect 43521 1099 43579 1133
rect 43613 1099 43650 1133
rect 43705 1099 43734 1133
rect 43458 1098 43650 1099
rect 43702 1098 43734 1099
rect 43458 1068 43734 1098
rect 43774 1064 43802 1414
rect 44074 1390 44138 1400
rect 44074 1356 44088 1390
rect 44122 1356 44394 1390
rect 44074 1338 44138 1356
rect 43990 1292 44062 1304
rect 43990 1240 44000 1292
rect 44052 1240 44062 1292
rect 43990 1228 44062 1240
rect 44360 1174 44394 1356
rect 44422 1274 44450 1578
rect 44422 1264 44490 1274
rect 44422 1230 44438 1264
rect 44472 1230 44490 1264
rect 44422 1216 44490 1230
rect 43834 1146 44394 1174
rect 43834 1143 43900 1146
rect 43834 1109 43850 1143
rect 43884 1109 43900 1143
rect 43834 1100 43900 1109
rect 44068 1091 44158 1112
rect 42266 983 42506 1000
rect 42550 1056 42616 1062
rect 42550 1004 42558 1056
rect 42610 1004 42616 1056
rect 42550 998 42564 1004
rect 42000 943 42046 976
rect 42000 909 42006 943
rect 42040 909 42046 943
rect 42266 949 42278 983
rect 42312 972 42506 983
rect 42558 981 42564 998
rect 42598 998 42616 1004
rect 42646 1015 42692 1062
rect 43774 1036 43846 1064
rect 42598 981 42604 998
rect 42312 949 42504 972
rect 42266 940 42504 949
rect 42000 862 42046 909
rect 42214 902 42280 910
rect 42128 898 42174 902
rect 41244 840 41316 844
rect 40704 815 40770 828
rect 40704 781 40720 815
rect 40754 781 40770 815
rect 40704 772 40770 781
rect 41244 788 41253 840
rect 41305 788 41316 840
rect 41244 776 41316 788
rect 41440 838 41514 858
rect 42088 855 42174 898
rect 41440 804 41452 838
rect 41486 804 41514 838
rect 41440 780 41514 804
rect 41550 844 41618 850
rect 41550 792 41557 844
rect 41609 838 41618 844
rect 41609 832 41702 838
rect 41609 798 41648 832
rect 41682 798 41702 832
rect 41609 792 41702 798
rect 41550 788 41702 792
rect 41946 815 42012 826
rect 41550 786 41618 788
rect 41946 781 41962 815
rect 41996 781 42012 815
rect 41946 768 42012 781
rect 42088 821 42134 855
rect 42168 821 42174 855
rect 42214 850 42220 902
rect 42272 850 42280 902
rect 42214 842 42230 850
rect 42088 783 42174 821
rect 42088 749 42134 783
rect 42168 749 42174 783
rect 41026 728 41084 742
rect 41026 708 41038 728
rect 40556 694 41038 708
rect 41072 694 41084 728
rect 40556 674 41084 694
rect 42088 702 42174 749
rect 42224 821 42230 842
rect 42264 842 42280 850
rect 42320 855 42416 902
rect 42264 821 42270 842
rect 42224 783 42270 821
rect 42224 749 42230 783
rect 42264 749 42270 783
rect 42224 702 42270 749
rect 42320 821 42326 855
rect 42360 821 42416 855
rect 42320 783 42416 821
rect 42320 749 42326 783
rect 42360 749 42416 783
rect 42320 702 42416 749
rect 40448 372 40494 384
rect 40556 344 40616 674
rect 42088 648 42138 702
rect 40662 624 40738 630
rect 40662 572 40670 624
rect 40722 572 40738 624
rect 40662 566 40738 572
rect 40878 597 41500 628
rect 40296 334 40616 344
rect 40296 300 40310 334
rect 40344 300 40616 334
rect 40296 282 40616 300
rect 40878 563 40907 597
rect 40941 563 40999 597
rect 41033 563 41091 597
rect 41125 595 41500 597
rect 41125 563 41253 595
rect 40878 561 41253 563
rect 41287 561 41345 595
rect 41379 561 41437 595
rect 41471 561 41500 595
rect 40878 530 41500 561
rect 41570 602 41846 620
rect 41570 589 41693 602
rect 41745 589 41846 602
rect 41922 598 41980 606
rect 41570 555 41599 589
rect 41633 555 41691 589
rect 41745 555 41783 589
rect 41817 555 41846 589
rect 41570 550 41693 555
rect 41745 550 41846 555
rect 40878 254 40976 530
rect 41570 524 41846 550
rect 41914 592 41988 598
rect 41914 540 41925 592
rect 41977 540 41988 592
rect 42068 582 42138 648
rect 42170 655 42228 670
rect 42170 621 42182 655
rect 42216 621 42228 655
rect 42170 604 42228 621
rect 41914 534 41988 540
rect 41922 528 41980 534
rect 41638 254 41722 524
rect 42088 502 42138 582
rect 42282 574 42340 592
rect 42282 540 42294 574
rect 42328 540 42340 574
rect 42282 530 42340 540
rect 42370 502 42416 702
rect 42088 490 42190 502
rect 42088 456 42150 490
rect 42184 456 42190 490
rect 42088 418 42190 456
rect 42240 490 42286 502
rect 42240 456 42246 490
rect 42280 456 42286 490
rect 42240 436 42286 456
rect 42336 490 42416 502
rect 42336 456 42342 490
rect 42376 456 42416 490
rect 42088 384 42150 418
rect 42184 384 42190 418
rect 42088 372 42190 384
rect 42230 430 42296 436
rect 42230 378 42238 430
rect 42290 378 42296 430
rect 42230 372 42296 378
rect 42336 418 42416 456
rect 42336 384 42342 418
rect 42376 384 42416 418
rect 42444 708 42504 940
rect 42558 943 42604 981
rect 42558 909 42564 943
rect 42598 909 42604 943
rect 42558 862 42604 909
rect 42646 981 42652 1015
rect 42686 981 42692 1015
rect 42646 943 42692 981
rect 42646 909 42652 943
rect 42686 909 42692 943
rect 42646 862 42692 909
rect 43800 1015 43846 1036
rect 43800 981 43806 1015
rect 43840 981 43846 1015
rect 43800 943 43846 981
rect 43800 909 43806 943
rect 43840 909 43846 943
rect 43800 862 43846 909
rect 43888 1042 43934 1062
rect 44068 1057 44097 1091
rect 44131 1057 44158 1091
rect 43888 1036 43956 1042
rect 44068 1036 44158 1057
rect 43888 1015 43896 1036
rect 43888 981 43894 1015
rect 43948 984 43956 1036
rect 43928 981 43956 984
rect 43888 976 43956 981
rect 44154 1000 44212 1002
rect 44360 1000 44394 1146
rect 44480 1143 44546 1154
rect 44480 1109 44496 1143
rect 44530 1109 44546 1143
rect 44480 1098 44546 1109
rect 44654 1144 45278 1176
rect 45360 1164 45438 2122
rect 45952 2113 45981 2122
rect 46015 2122 47869 2147
rect 46015 2113 46042 2122
rect 45952 2092 46042 2113
rect 46038 2056 46096 2058
rect 46038 2039 46100 2056
rect 46038 2005 46050 2039
rect 46084 2005 46100 2039
rect 46038 1996 46100 2005
rect 45538 1958 45904 1962
rect 45986 1958 46052 1966
rect 45538 1930 45946 1958
rect 45538 1892 45566 1930
rect 45860 1911 45946 1930
rect 45538 1884 45604 1892
rect 45538 1850 45553 1884
rect 45587 1850 45604 1884
rect 45538 1838 45604 1850
rect 45710 1888 45778 1894
rect 45710 1836 45720 1888
rect 45772 1836 45778 1888
rect 45710 1830 45778 1836
rect 45860 1877 45906 1911
rect 45940 1877 45946 1911
rect 45986 1906 45992 1958
rect 46044 1906 46052 1958
rect 45986 1898 46002 1906
rect 45860 1839 45946 1877
rect 45860 1805 45906 1839
rect 45940 1805 45946 1839
rect 45620 1776 45688 1782
rect 45620 1724 45628 1776
rect 45680 1724 45688 1776
rect 45620 1714 45688 1724
rect 45860 1758 45946 1805
rect 45996 1877 46002 1898
rect 46036 1898 46052 1906
rect 46092 1926 46420 1958
rect 46092 1911 46188 1926
rect 46036 1877 46042 1898
rect 45996 1839 46042 1877
rect 45996 1805 46002 1839
rect 46036 1805 46042 1839
rect 45996 1758 46042 1805
rect 46092 1877 46098 1911
rect 46132 1877 46188 1911
rect 46392 1890 46420 1926
rect 46092 1839 46188 1877
rect 46092 1805 46098 1839
rect 46132 1805 46188 1839
rect 46350 1882 46420 1890
rect 46350 1848 46365 1882
rect 46399 1848 46420 1882
rect 46350 1830 46420 1848
rect 46526 1890 46590 1896
rect 46526 1838 46532 1890
rect 46584 1838 46590 1890
rect 46526 1832 46590 1838
rect 46092 1758 46188 1805
rect 45518 1643 45794 1674
rect 45518 1609 45547 1643
rect 45581 1609 45639 1643
rect 45673 1609 45731 1643
rect 45765 1609 45794 1643
rect 45518 1578 45794 1609
rect 45860 1558 45910 1758
rect 45942 1711 46000 1726
rect 45942 1677 45954 1711
rect 45988 1677 46000 1711
rect 45942 1660 46000 1677
rect 46054 1630 46112 1648
rect 46054 1596 46066 1630
rect 46100 1596 46112 1630
rect 46054 1586 46112 1596
rect 46142 1558 46188 1758
rect 46438 1774 46502 1780
rect 46438 1722 46444 1774
rect 46496 1722 46502 1774
rect 46438 1716 46502 1722
rect 46332 1643 46608 1674
rect 46332 1609 46361 1643
rect 46395 1609 46453 1643
rect 46487 1609 46545 1643
rect 46579 1609 46608 1643
rect 46332 1606 46608 1609
rect 45500 1541 45564 1548
rect 45500 1508 45506 1541
rect 45558 1508 45564 1541
rect 45676 1541 45740 1548
rect 45676 1508 45682 1541
rect 45558 1489 45682 1508
rect 45734 1489 45740 1541
rect 45506 1480 45740 1489
rect 45860 1546 45962 1558
rect 45860 1512 45922 1546
rect 45956 1512 45962 1546
rect 45860 1474 45962 1512
rect 46012 1546 46058 1558
rect 46012 1512 46018 1546
rect 46052 1512 46058 1546
rect 46012 1492 46058 1512
rect 46108 1546 46188 1558
rect 46108 1512 46114 1546
rect 46148 1512 46188 1546
rect 45860 1442 45922 1474
rect 45656 1440 45922 1442
rect 45956 1440 45962 1474
rect 45656 1428 45962 1440
rect 46002 1486 46068 1492
rect 46002 1434 46010 1486
rect 46062 1434 46068 1486
rect 46002 1428 46068 1434
rect 46108 1474 46188 1512
rect 46108 1440 46114 1474
rect 46148 1440 46188 1474
rect 46304 1578 46608 1606
rect 46108 1428 46154 1440
rect 45656 1414 45910 1428
rect 45500 1408 45566 1414
rect 45500 1356 45508 1408
rect 45560 1356 45566 1408
rect 45500 1350 45566 1356
rect 44654 1141 44684 1144
rect 44736 1141 45278 1144
rect 44654 1107 44683 1141
rect 44736 1107 44775 1141
rect 44809 1107 44867 1141
rect 44901 1139 45278 1141
rect 44901 1107 45029 1139
rect 44654 1092 44684 1107
rect 44736 1105 45029 1107
rect 45063 1105 45121 1139
rect 45155 1105 45213 1139
rect 45247 1105 45278 1139
rect 44736 1092 45278 1105
rect 44654 1074 45278 1092
rect 45340 1150 45616 1164
rect 45340 1133 45532 1150
rect 45584 1133 45616 1150
rect 45340 1099 45369 1133
rect 45403 1099 45461 1133
rect 45495 1099 45532 1133
rect 45587 1099 45616 1133
rect 45340 1098 45532 1099
rect 45584 1098 45616 1099
rect 45340 1068 45616 1098
rect 45656 1064 45684 1414
rect 45956 1390 46020 1400
rect 45956 1356 45970 1390
rect 46004 1356 46276 1390
rect 45956 1338 46020 1356
rect 45872 1292 45944 1304
rect 45872 1240 45882 1292
rect 45934 1240 45944 1292
rect 45872 1228 45944 1240
rect 46242 1174 46276 1356
rect 46304 1274 46332 1578
rect 46304 1264 46372 1274
rect 46304 1230 46320 1264
rect 46354 1230 46372 1264
rect 46304 1216 46372 1230
rect 45716 1146 46276 1174
rect 45716 1143 45782 1146
rect 45716 1109 45732 1143
rect 45766 1109 45782 1143
rect 45716 1100 45782 1109
rect 45950 1091 46040 1112
rect 44154 983 44394 1000
rect 44438 1056 44504 1062
rect 44438 1004 44446 1056
rect 44498 1004 44504 1056
rect 44438 998 44452 1004
rect 43888 943 43934 976
rect 43888 909 43894 943
rect 43928 909 43934 943
rect 44154 949 44166 983
rect 44200 972 44394 983
rect 44446 981 44452 998
rect 44486 998 44504 1004
rect 44534 1015 44580 1062
rect 45656 1036 45728 1064
rect 44486 981 44492 998
rect 44200 949 44392 972
rect 44154 940 44392 949
rect 43888 862 43934 909
rect 44102 902 44168 910
rect 44016 898 44062 902
rect 43132 840 43204 844
rect 42592 815 42658 828
rect 42592 781 42608 815
rect 42642 781 42658 815
rect 42592 772 42658 781
rect 43132 788 43141 840
rect 43193 788 43204 840
rect 43132 776 43204 788
rect 43328 838 43402 858
rect 43976 855 44062 898
rect 43328 804 43340 838
rect 43374 804 43402 838
rect 43328 780 43402 804
rect 43438 844 43506 850
rect 43438 792 43445 844
rect 43497 838 43506 844
rect 43497 832 43590 838
rect 43497 798 43536 832
rect 43570 798 43590 832
rect 43497 792 43590 798
rect 43438 788 43590 792
rect 43834 815 43900 826
rect 43438 786 43506 788
rect 43834 781 43850 815
rect 43884 781 43900 815
rect 43834 768 43900 781
rect 43976 821 44022 855
rect 44056 821 44062 855
rect 44102 850 44108 902
rect 44160 850 44168 902
rect 44102 842 44118 850
rect 43976 783 44062 821
rect 43976 749 44022 783
rect 44056 749 44062 783
rect 42914 728 42972 742
rect 42914 708 42926 728
rect 42444 694 42926 708
rect 42960 694 42972 728
rect 42444 674 42972 694
rect 43976 702 44062 749
rect 44112 821 44118 842
rect 44152 842 44168 850
rect 44208 855 44304 902
rect 44152 821 44158 842
rect 44112 783 44158 821
rect 44112 749 44118 783
rect 44152 749 44158 783
rect 44112 702 44158 749
rect 44208 821 44214 855
rect 44248 821 44304 855
rect 44208 783 44304 821
rect 44208 749 44214 783
rect 44248 749 44304 783
rect 44208 702 44304 749
rect 42336 372 42382 384
rect 42444 344 42504 674
rect 43976 648 44026 702
rect 42550 624 42626 630
rect 42550 572 42558 624
rect 42610 572 42626 624
rect 42550 566 42626 572
rect 42766 597 43388 628
rect 42184 334 42504 344
rect 42184 300 42198 334
rect 42232 300 42504 334
rect 42184 282 42504 300
rect 42766 563 42795 597
rect 42829 563 42887 597
rect 42921 563 42979 597
rect 43013 595 43388 597
rect 43013 563 43141 595
rect 42766 561 43141 563
rect 43175 561 43233 595
rect 43267 561 43325 595
rect 43359 561 43388 595
rect 42766 530 43388 561
rect 43458 602 43734 620
rect 43458 589 43581 602
rect 43633 589 43734 602
rect 43810 598 43868 606
rect 43458 555 43487 589
rect 43521 555 43579 589
rect 43633 555 43671 589
rect 43705 555 43734 589
rect 43458 550 43581 555
rect 43633 550 43734 555
rect 42766 254 42864 530
rect 43458 524 43734 550
rect 43802 592 43876 598
rect 43802 540 43813 592
rect 43865 540 43876 592
rect 43956 582 44026 648
rect 44058 655 44116 670
rect 44058 621 44070 655
rect 44104 621 44116 655
rect 44058 604 44116 621
rect 43802 534 43876 540
rect 43810 528 43868 534
rect 43526 254 43610 524
rect 43976 502 44026 582
rect 44170 574 44228 592
rect 44170 540 44182 574
rect 44216 540 44228 574
rect 44170 530 44228 540
rect 44258 502 44304 702
rect 43976 490 44078 502
rect 43976 456 44038 490
rect 44072 456 44078 490
rect 43976 418 44078 456
rect 44128 490 44174 502
rect 44128 456 44134 490
rect 44168 456 44174 490
rect 44128 436 44174 456
rect 44224 490 44304 502
rect 44224 456 44230 490
rect 44264 456 44304 490
rect 43976 384 44038 418
rect 44072 384 44078 418
rect 43976 372 44078 384
rect 44118 430 44184 436
rect 44118 378 44126 430
rect 44178 378 44184 430
rect 44118 372 44184 378
rect 44224 418 44304 456
rect 44224 384 44230 418
rect 44264 384 44304 418
rect 44332 708 44392 940
rect 44446 943 44492 981
rect 44446 909 44452 943
rect 44486 909 44492 943
rect 44446 862 44492 909
rect 44534 981 44540 1015
rect 44574 981 44580 1015
rect 44534 943 44580 981
rect 44534 909 44540 943
rect 44574 909 44580 943
rect 44534 862 44580 909
rect 45682 1015 45728 1036
rect 45682 981 45688 1015
rect 45722 981 45728 1015
rect 45682 943 45728 981
rect 45682 909 45688 943
rect 45722 909 45728 943
rect 45682 862 45728 909
rect 45770 1042 45816 1062
rect 45950 1057 45979 1091
rect 46013 1057 46040 1091
rect 45770 1036 45838 1042
rect 45950 1036 46040 1057
rect 45770 1015 45778 1036
rect 45770 981 45776 1015
rect 45830 984 45838 1036
rect 45810 981 45838 984
rect 45770 976 45838 981
rect 46036 1000 46094 1002
rect 46242 1000 46276 1146
rect 46362 1143 46428 1154
rect 46362 1109 46378 1143
rect 46412 1109 46428 1143
rect 46362 1098 46428 1109
rect 46536 1144 47160 1176
rect 47248 1164 47326 2122
rect 47840 2113 47869 2122
rect 47903 2122 49757 2147
rect 47903 2113 47930 2122
rect 47840 2092 47930 2113
rect 47926 2056 47984 2058
rect 47926 2039 47988 2056
rect 47926 2005 47938 2039
rect 47972 2005 47988 2039
rect 47926 1996 47988 2005
rect 47426 1958 47792 1962
rect 47874 1958 47940 1966
rect 47426 1930 47834 1958
rect 47426 1892 47454 1930
rect 47748 1911 47834 1930
rect 47426 1884 47492 1892
rect 47426 1850 47441 1884
rect 47475 1850 47492 1884
rect 47426 1838 47492 1850
rect 47598 1888 47666 1894
rect 47598 1836 47608 1888
rect 47660 1836 47666 1888
rect 47598 1830 47666 1836
rect 47748 1877 47794 1911
rect 47828 1877 47834 1911
rect 47874 1906 47880 1958
rect 47932 1906 47940 1958
rect 47874 1898 47890 1906
rect 47748 1839 47834 1877
rect 47748 1805 47794 1839
rect 47828 1805 47834 1839
rect 47508 1776 47576 1782
rect 47508 1724 47516 1776
rect 47568 1724 47576 1776
rect 47508 1714 47576 1724
rect 47748 1758 47834 1805
rect 47884 1877 47890 1898
rect 47924 1898 47940 1906
rect 47980 1926 48308 1958
rect 47980 1911 48076 1926
rect 47924 1877 47930 1898
rect 47884 1839 47930 1877
rect 47884 1805 47890 1839
rect 47924 1805 47930 1839
rect 47884 1758 47930 1805
rect 47980 1877 47986 1911
rect 48020 1877 48076 1911
rect 48280 1890 48308 1926
rect 47980 1839 48076 1877
rect 47980 1805 47986 1839
rect 48020 1805 48076 1839
rect 48238 1882 48308 1890
rect 48238 1848 48253 1882
rect 48287 1848 48308 1882
rect 48238 1830 48308 1848
rect 48414 1890 48478 1896
rect 48414 1838 48420 1890
rect 48472 1838 48478 1890
rect 48414 1832 48478 1838
rect 47980 1758 48076 1805
rect 47406 1643 47682 1674
rect 47406 1609 47435 1643
rect 47469 1609 47527 1643
rect 47561 1609 47619 1643
rect 47653 1609 47682 1643
rect 47406 1578 47682 1609
rect 47748 1558 47798 1758
rect 47830 1711 47888 1726
rect 47830 1677 47842 1711
rect 47876 1677 47888 1711
rect 47830 1660 47888 1677
rect 47942 1630 48000 1648
rect 47942 1596 47954 1630
rect 47988 1596 48000 1630
rect 47942 1586 48000 1596
rect 48030 1558 48076 1758
rect 48326 1774 48390 1780
rect 48326 1722 48332 1774
rect 48384 1722 48390 1774
rect 48326 1716 48390 1722
rect 48220 1643 48496 1674
rect 48220 1609 48249 1643
rect 48283 1609 48341 1643
rect 48375 1609 48433 1643
rect 48467 1609 48496 1643
rect 48220 1606 48496 1609
rect 47388 1541 47452 1548
rect 47388 1508 47394 1541
rect 47446 1508 47452 1541
rect 47564 1541 47628 1548
rect 47564 1508 47570 1541
rect 47446 1489 47570 1508
rect 47622 1489 47628 1541
rect 47394 1480 47628 1489
rect 47748 1546 47850 1558
rect 47748 1512 47810 1546
rect 47844 1512 47850 1546
rect 47748 1474 47850 1512
rect 47900 1546 47946 1558
rect 47900 1512 47906 1546
rect 47940 1512 47946 1546
rect 47900 1492 47946 1512
rect 47996 1546 48076 1558
rect 47996 1512 48002 1546
rect 48036 1512 48076 1546
rect 47748 1442 47810 1474
rect 47544 1440 47810 1442
rect 47844 1440 47850 1474
rect 47544 1428 47850 1440
rect 47890 1486 47956 1492
rect 47890 1434 47898 1486
rect 47950 1434 47956 1486
rect 47890 1428 47956 1434
rect 47996 1474 48076 1512
rect 47996 1440 48002 1474
rect 48036 1440 48076 1474
rect 48192 1578 48496 1606
rect 47996 1428 48042 1440
rect 47544 1414 47798 1428
rect 47388 1408 47454 1414
rect 47388 1356 47396 1408
rect 47448 1356 47454 1408
rect 47388 1350 47454 1356
rect 46536 1141 46566 1144
rect 46618 1141 47160 1144
rect 46536 1107 46565 1141
rect 46618 1107 46657 1141
rect 46691 1107 46749 1141
rect 46783 1139 47160 1141
rect 46783 1107 46911 1139
rect 46536 1092 46566 1107
rect 46618 1105 46911 1107
rect 46945 1105 47003 1139
rect 47037 1105 47095 1139
rect 47129 1105 47160 1139
rect 46618 1092 47160 1105
rect 46536 1074 47160 1092
rect 47228 1150 47504 1164
rect 47228 1133 47420 1150
rect 47472 1133 47504 1150
rect 47228 1099 47257 1133
rect 47291 1099 47349 1133
rect 47383 1099 47420 1133
rect 47475 1099 47504 1133
rect 47228 1098 47420 1099
rect 47472 1098 47504 1099
rect 47228 1068 47504 1098
rect 47544 1064 47572 1414
rect 47844 1390 47908 1400
rect 47844 1356 47858 1390
rect 47892 1356 48164 1390
rect 47844 1338 47908 1356
rect 47760 1292 47832 1304
rect 47760 1240 47770 1292
rect 47822 1240 47832 1292
rect 47760 1228 47832 1240
rect 48130 1174 48164 1356
rect 48192 1274 48220 1578
rect 48192 1264 48260 1274
rect 48192 1230 48208 1264
rect 48242 1230 48260 1264
rect 48192 1216 48260 1230
rect 47604 1146 48164 1174
rect 47604 1143 47670 1146
rect 47604 1109 47620 1143
rect 47654 1109 47670 1143
rect 47604 1100 47670 1109
rect 47838 1091 47928 1112
rect 46036 983 46276 1000
rect 46320 1056 46386 1062
rect 46320 1004 46328 1056
rect 46380 1004 46386 1056
rect 46320 998 46334 1004
rect 45770 943 45816 976
rect 45770 909 45776 943
rect 45810 909 45816 943
rect 46036 949 46048 983
rect 46082 972 46276 983
rect 46328 981 46334 998
rect 46368 998 46386 1004
rect 46416 1015 46462 1062
rect 47544 1036 47616 1064
rect 46368 981 46374 998
rect 46082 949 46274 972
rect 46036 940 46274 949
rect 45770 862 45816 909
rect 45984 902 46050 910
rect 45898 898 45944 902
rect 45020 840 45092 844
rect 44480 815 44546 828
rect 44480 781 44496 815
rect 44530 781 44546 815
rect 44480 772 44546 781
rect 45020 788 45029 840
rect 45081 788 45092 840
rect 45020 776 45092 788
rect 45216 838 45290 858
rect 45858 855 45944 898
rect 45216 804 45228 838
rect 45262 804 45290 838
rect 45216 780 45290 804
rect 45320 844 45388 850
rect 45320 792 45327 844
rect 45379 838 45388 844
rect 45379 832 45472 838
rect 45379 798 45418 832
rect 45452 798 45472 832
rect 45379 792 45472 798
rect 45320 788 45472 792
rect 45716 815 45782 826
rect 45320 786 45388 788
rect 45716 781 45732 815
rect 45766 781 45782 815
rect 45716 768 45782 781
rect 45858 821 45904 855
rect 45938 821 45944 855
rect 45984 850 45990 902
rect 46042 850 46050 902
rect 45984 842 46000 850
rect 45858 783 45944 821
rect 45858 749 45904 783
rect 45938 749 45944 783
rect 44802 728 44860 742
rect 44802 708 44814 728
rect 44332 694 44814 708
rect 44848 694 44860 728
rect 44332 674 44860 694
rect 45858 702 45944 749
rect 45994 821 46000 842
rect 46034 842 46050 850
rect 46090 855 46186 902
rect 46034 821 46040 842
rect 45994 783 46040 821
rect 45994 749 46000 783
rect 46034 749 46040 783
rect 45994 702 46040 749
rect 46090 821 46096 855
rect 46130 821 46186 855
rect 46090 783 46186 821
rect 46090 749 46096 783
rect 46130 749 46186 783
rect 46090 702 46186 749
rect 44224 372 44270 384
rect 44332 344 44392 674
rect 45858 648 45908 702
rect 44438 624 44514 630
rect 44438 572 44446 624
rect 44498 572 44514 624
rect 44438 566 44514 572
rect 44654 597 45276 628
rect 44072 334 44392 344
rect 44072 300 44086 334
rect 44120 300 44392 334
rect 44072 282 44392 300
rect 44654 563 44683 597
rect 44717 563 44775 597
rect 44809 563 44867 597
rect 44901 595 45276 597
rect 44901 563 45029 595
rect 44654 561 45029 563
rect 45063 561 45121 595
rect 45155 561 45213 595
rect 45247 561 45276 595
rect 44654 530 45276 561
rect 45340 602 45616 620
rect 45340 589 45463 602
rect 45515 589 45616 602
rect 45692 598 45750 606
rect 45340 555 45369 589
rect 45403 555 45461 589
rect 45515 555 45553 589
rect 45587 555 45616 589
rect 45340 550 45463 555
rect 45515 550 45616 555
rect 44654 254 44752 530
rect 45340 524 45616 550
rect 45684 592 45758 598
rect 45684 540 45695 592
rect 45747 540 45758 592
rect 45838 582 45908 648
rect 45940 655 45998 670
rect 45940 621 45952 655
rect 45986 621 45998 655
rect 45940 604 45998 621
rect 45684 534 45758 540
rect 45692 528 45750 534
rect 45408 254 45492 524
rect 45858 502 45908 582
rect 46052 574 46110 592
rect 46052 540 46064 574
rect 46098 540 46110 574
rect 46052 530 46110 540
rect 46140 502 46186 702
rect 45858 490 45960 502
rect 45858 456 45920 490
rect 45954 456 45960 490
rect 45858 418 45960 456
rect 46010 490 46056 502
rect 46010 456 46016 490
rect 46050 456 46056 490
rect 46010 436 46056 456
rect 46106 490 46186 502
rect 46106 456 46112 490
rect 46146 456 46186 490
rect 45858 384 45920 418
rect 45954 384 45960 418
rect 45858 372 45960 384
rect 46000 430 46066 436
rect 46000 378 46008 430
rect 46060 378 46066 430
rect 46000 372 46066 378
rect 46106 418 46186 456
rect 46106 384 46112 418
rect 46146 384 46186 418
rect 46214 708 46274 940
rect 46328 943 46374 981
rect 46328 909 46334 943
rect 46368 909 46374 943
rect 46328 862 46374 909
rect 46416 981 46422 1015
rect 46456 981 46462 1015
rect 46416 943 46462 981
rect 46416 909 46422 943
rect 46456 909 46462 943
rect 46416 862 46462 909
rect 47570 1015 47616 1036
rect 47570 981 47576 1015
rect 47610 981 47616 1015
rect 47570 943 47616 981
rect 47570 909 47576 943
rect 47610 909 47616 943
rect 47570 862 47616 909
rect 47658 1042 47704 1062
rect 47838 1057 47867 1091
rect 47901 1057 47928 1091
rect 47658 1036 47726 1042
rect 47838 1036 47928 1057
rect 47658 1015 47666 1036
rect 47658 981 47664 1015
rect 47718 984 47726 1036
rect 47698 981 47726 984
rect 47658 976 47726 981
rect 47924 1000 47982 1002
rect 48130 1000 48164 1146
rect 48250 1143 48316 1154
rect 48250 1109 48266 1143
rect 48300 1109 48316 1143
rect 48250 1098 48316 1109
rect 48424 1144 49048 1176
rect 49136 1164 49214 2122
rect 49728 2113 49757 2122
rect 49791 2122 51645 2147
rect 49791 2113 49818 2122
rect 49728 2092 49818 2113
rect 49814 2056 49872 2058
rect 49814 2039 49876 2056
rect 49814 2005 49826 2039
rect 49860 2005 49876 2039
rect 49814 1996 49876 2005
rect 49314 1958 49680 1962
rect 49762 1958 49828 1966
rect 49314 1930 49722 1958
rect 49314 1892 49342 1930
rect 49636 1911 49722 1930
rect 49314 1884 49380 1892
rect 49314 1850 49329 1884
rect 49363 1850 49380 1884
rect 49314 1838 49380 1850
rect 49486 1888 49554 1894
rect 49486 1836 49496 1888
rect 49548 1836 49554 1888
rect 49486 1830 49554 1836
rect 49636 1877 49682 1911
rect 49716 1877 49722 1911
rect 49762 1906 49768 1958
rect 49820 1906 49828 1958
rect 49762 1898 49778 1906
rect 49636 1839 49722 1877
rect 49636 1805 49682 1839
rect 49716 1805 49722 1839
rect 49396 1776 49464 1782
rect 49396 1724 49404 1776
rect 49456 1724 49464 1776
rect 49396 1714 49464 1724
rect 49636 1758 49722 1805
rect 49772 1877 49778 1898
rect 49812 1898 49828 1906
rect 49868 1926 50196 1958
rect 49868 1911 49964 1926
rect 49812 1877 49818 1898
rect 49772 1839 49818 1877
rect 49772 1805 49778 1839
rect 49812 1805 49818 1839
rect 49772 1758 49818 1805
rect 49868 1877 49874 1911
rect 49908 1877 49964 1911
rect 50168 1890 50196 1926
rect 49868 1839 49964 1877
rect 49868 1805 49874 1839
rect 49908 1805 49964 1839
rect 50126 1882 50196 1890
rect 50126 1848 50141 1882
rect 50175 1848 50196 1882
rect 50126 1830 50196 1848
rect 50302 1890 50366 1896
rect 50302 1838 50308 1890
rect 50360 1838 50366 1890
rect 50302 1832 50366 1838
rect 49868 1758 49964 1805
rect 49294 1643 49570 1674
rect 49294 1609 49323 1643
rect 49357 1609 49415 1643
rect 49449 1609 49507 1643
rect 49541 1609 49570 1643
rect 49294 1578 49570 1609
rect 49636 1558 49686 1758
rect 49718 1711 49776 1726
rect 49718 1677 49730 1711
rect 49764 1677 49776 1711
rect 49718 1660 49776 1677
rect 49830 1630 49888 1648
rect 49830 1596 49842 1630
rect 49876 1596 49888 1630
rect 49830 1586 49888 1596
rect 49918 1558 49964 1758
rect 50214 1774 50278 1780
rect 50214 1722 50220 1774
rect 50272 1722 50278 1774
rect 50214 1716 50278 1722
rect 50108 1643 50384 1674
rect 50108 1609 50137 1643
rect 50171 1609 50229 1643
rect 50263 1609 50321 1643
rect 50355 1609 50384 1643
rect 50108 1606 50384 1609
rect 49276 1541 49340 1548
rect 49276 1508 49282 1541
rect 49334 1508 49340 1541
rect 49452 1541 49516 1548
rect 49452 1508 49458 1541
rect 49334 1489 49458 1508
rect 49510 1489 49516 1541
rect 49282 1480 49516 1489
rect 49636 1546 49738 1558
rect 49636 1512 49698 1546
rect 49732 1512 49738 1546
rect 49636 1474 49738 1512
rect 49788 1546 49834 1558
rect 49788 1512 49794 1546
rect 49828 1512 49834 1546
rect 49788 1492 49834 1512
rect 49884 1546 49964 1558
rect 49884 1512 49890 1546
rect 49924 1512 49964 1546
rect 49636 1442 49698 1474
rect 49432 1440 49698 1442
rect 49732 1440 49738 1474
rect 49432 1428 49738 1440
rect 49778 1486 49844 1492
rect 49778 1434 49786 1486
rect 49838 1434 49844 1486
rect 49778 1428 49844 1434
rect 49884 1474 49964 1512
rect 49884 1440 49890 1474
rect 49924 1440 49964 1474
rect 50080 1578 50384 1606
rect 49884 1428 49930 1440
rect 49432 1414 49686 1428
rect 49276 1408 49342 1414
rect 49276 1356 49284 1408
rect 49336 1356 49342 1408
rect 49276 1350 49342 1356
rect 48424 1141 48454 1144
rect 48506 1141 49048 1144
rect 48424 1107 48453 1141
rect 48506 1107 48545 1141
rect 48579 1107 48637 1141
rect 48671 1139 49048 1141
rect 48671 1107 48799 1139
rect 48424 1092 48454 1107
rect 48506 1105 48799 1107
rect 48833 1105 48891 1139
rect 48925 1105 48983 1139
rect 49017 1105 49048 1139
rect 48506 1092 49048 1105
rect 48424 1074 49048 1092
rect 49116 1150 49392 1164
rect 49116 1133 49308 1150
rect 49360 1133 49392 1150
rect 49116 1099 49145 1133
rect 49179 1099 49237 1133
rect 49271 1099 49308 1133
rect 49363 1099 49392 1133
rect 49116 1098 49308 1099
rect 49360 1098 49392 1099
rect 49116 1068 49392 1098
rect 49432 1064 49460 1414
rect 49732 1390 49796 1400
rect 49732 1356 49746 1390
rect 49780 1356 50052 1390
rect 49732 1338 49796 1356
rect 49648 1292 49720 1304
rect 49648 1240 49658 1292
rect 49710 1240 49720 1292
rect 49648 1228 49720 1240
rect 50018 1174 50052 1356
rect 50080 1274 50108 1578
rect 50080 1264 50148 1274
rect 50080 1230 50096 1264
rect 50130 1230 50148 1264
rect 50080 1216 50148 1230
rect 49492 1146 50052 1174
rect 49492 1143 49558 1146
rect 49492 1109 49508 1143
rect 49542 1109 49558 1143
rect 49492 1100 49558 1109
rect 49726 1091 49816 1112
rect 47924 983 48164 1000
rect 48208 1056 48274 1062
rect 48208 1004 48216 1056
rect 48268 1004 48274 1056
rect 48208 998 48222 1004
rect 47658 943 47704 976
rect 47658 909 47664 943
rect 47698 909 47704 943
rect 47924 949 47936 983
rect 47970 972 48164 983
rect 48216 981 48222 998
rect 48256 998 48274 1004
rect 48304 1015 48350 1062
rect 49432 1036 49504 1064
rect 48256 981 48262 998
rect 47970 949 48162 972
rect 47924 940 48162 949
rect 47658 862 47704 909
rect 47872 902 47938 910
rect 47786 898 47832 902
rect 46902 840 46974 844
rect 46362 815 46428 828
rect 46362 781 46378 815
rect 46412 781 46428 815
rect 46362 772 46428 781
rect 46902 788 46911 840
rect 46963 788 46974 840
rect 46902 776 46974 788
rect 47098 838 47172 858
rect 47746 855 47832 898
rect 47098 804 47110 838
rect 47144 804 47172 838
rect 47098 780 47172 804
rect 47208 844 47276 850
rect 47208 792 47215 844
rect 47267 838 47276 844
rect 47267 832 47360 838
rect 47267 798 47306 832
rect 47340 798 47360 832
rect 47267 792 47360 798
rect 47208 788 47360 792
rect 47604 815 47670 826
rect 47208 786 47276 788
rect 47604 781 47620 815
rect 47654 781 47670 815
rect 47604 768 47670 781
rect 47746 821 47792 855
rect 47826 821 47832 855
rect 47872 850 47878 902
rect 47930 850 47938 902
rect 47872 842 47888 850
rect 47746 783 47832 821
rect 47746 749 47792 783
rect 47826 749 47832 783
rect 46684 728 46742 742
rect 46684 708 46696 728
rect 46214 694 46696 708
rect 46730 694 46742 728
rect 46214 674 46742 694
rect 47746 702 47832 749
rect 47882 821 47888 842
rect 47922 842 47938 850
rect 47978 855 48074 902
rect 47922 821 47928 842
rect 47882 783 47928 821
rect 47882 749 47888 783
rect 47922 749 47928 783
rect 47882 702 47928 749
rect 47978 821 47984 855
rect 48018 821 48074 855
rect 47978 783 48074 821
rect 47978 749 47984 783
rect 48018 749 48074 783
rect 47978 702 48074 749
rect 46106 372 46152 384
rect 46214 344 46274 674
rect 47746 648 47796 702
rect 46320 624 46396 630
rect 46320 572 46328 624
rect 46380 572 46396 624
rect 46320 566 46396 572
rect 46536 597 47158 628
rect 45954 334 46274 344
rect 45954 300 45968 334
rect 46002 300 46274 334
rect 45954 282 46274 300
rect 46536 563 46565 597
rect 46599 563 46657 597
rect 46691 563 46749 597
rect 46783 595 47158 597
rect 46783 563 46911 595
rect 46536 561 46911 563
rect 46945 561 47003 595
rect 47037 561 47095 595
rect 47129 561 47158 595
rect 46536 530 47158 561
rect 47228 602 47504 620
rect 47228 589 47351 602
rect 47403 589 47504 602
rect 47580 598 47638 606
rect 47228 555 47257 589
rect 47291 555 47349 589
rect 47403 555 47441 589
rect 47475 555 47504 589
rect 47228 550 47351 555
rect 47403 550 47504 555
rect 46536 254 46634 530
rect 47228 524 47504 550
rect 47572 592 47646 598
rect 47572 540 47583 592
rect 47635 540 47646 592
rect 47726 582 47796 648
rect 47828 655 47886 670
rect 47828 621 47840 655
rect 47874 621 47886 655
rect 47828 604 47886 621
rect 47572 534 47646 540
rect 47580 528 47638 534
rect 47296 254 47380 524
rect 47746 502 47796 582
rect 47940 574 47998 592
rect 47940 540 47952 574
rect 47986 540 47998 574
rect 47940 530 47998 540
rect 48028 502 48074 702
rect 47746 490 47848 502
rect 47746 456 47808 490
rect 47842 456 47848 490
rect 47746 418 47848 456
rect 47898 490 47944 502
rect 47898 456 47904 490
rect 47938 456 47944 490
rect 47898 436 47944 456
rect 47994 490 48074 502
rect 47994 456 48000 490
rect 48034 456 48074 490
rect 47746 384 47808 418
rect 47842 384 47848 418
rect 47746 372 47848 384
rect 47888 430 47954 436
rect 47888 378 47896 430
rect 47948 378 47954 430
rect 47888 372 47954 378
rect 47994 418 48074 456
rect 47994 384 48000 418
rect 48034 384 48074 418
rect 48102 708 48162 940
rect 48216 943 48262 981
rect 48216 909 48222 943
rect 48256 909 48262 943
rect 48216 862 48262 909
rect 48304 981 48310 1015
rect 48344 981 48350 1015
rect 48304 943 48350 981
rect 48304 909 48310 943
rect 48344 909 48350 943
rect 48304 862 48350 909
rect 49458 1015 49504 1036
rect 49458 981 49464 1015
rect 49498 981 49504 1015
rect 49458 943 49504 981
rect 49458 909 49464 943
rect 49498 909 49504 943
rect 49458 862 49504 909
rect 49546 1042 49592 1062
rect 49726 1057 49755 1091
rect 49789 1057 49816 1091
rect 49546 1036 49614 1042
rect 49726 1036 49816 1057
rect 49546 1015 49554 1036
rect 49546 981 49552 1015
rect 49606 984 49614 1036
rect 49586 981 49614 984
rect 49546 976 49614 981
rect 49812 1000 49870 1002
rect 50018 1000 50052 1146
rect 50138 1143 50204 1154
rect 50138 1109 50154 1143
rect 50188 1109 50204 1143
rect 50138 1098 50204 1109
rect 50312 1144 50936 1176
rect 51024 1164 51102 2122
rect 51616 2113 51645 2122
rect 51679 2122 53533 2147
rect 51679 2113 51706 2122
rect 51616 2092 51706 2113
rect 51702 2056 51760 2058
rect 51702 2039 51764 2056
rect 51702 2005 51714 2039
rect 51748 2005 51764 2039
rect 51702 1996 51764 2005
rect 51202 1958 51568 1962
rect 51650 1958 51716 1966
rect 51202 1930 51610 1958
rect 51202 1892 51230 1930
rect 51524 1911 51610 1930
rect 51202 1884 51268 1892
rect 51202 1850 51217 1884
rect 51251 1850 51268 1884
rect 51202 1838 51268 1850
rect 51374 1888 51442 1894
rect 51374 1836 51384 1888
rect 51436 1836 51442 1888
rect 51374 1830 51442 1836
rect 51524 1877 51570 1911
rect 51604 1877 51610 1911
rect 51650 1906 51656 1958
rect 51708 1906 51716 1958
rect 51650 1898 51666 1906
rect 51524 1839 51610 1877
rect 51524 1805 51570 1839
rect 51604 1805 51610 1839
rect 51284 1776 51352 1782
rect 51284 1724 51292 1776
rect 51344 1724 51352 1776
rect 51284 1714 51352 1724
rect 51524 1758 51610 1805
rect 51660 1877 51666 1898
rect 51700 1898 51716 1906
rect 51756 1926 52084 1958
rect 51756 1911 51852 1926
rect 51700 1877 51706 1898
rect 51660 1839 51706 1877
rect 51660 1805 51666 1839
rect 51700 1805 51706 1839
rect 51660 1758 51706 1805
rect 51756 1877 51762 1911
rect 51796 1877 51852 1911
rect 52056 1890 52084 1926
rect 51756 1839 51852 1877
rect 51756 1805 51762 1839
rect 51796 1805 51852 1839
rect 52014 1882 52084 1890
rect 52014 1848 52029 1882
rect 52063 1848 52084 1882
rect 52014 1830 52084 1848
rect 52190 1890 52254 1896
rect 52190 1838 52196 1890
rect 52248 1838 52254 1890
rect 52190 1832 52254 1838
rect 51756 1758 51852 1805
rect 51182 1643 51458 1674
rect 51182 1609 51211 1643
rect 51245 1609 51303 1643
rect 51337 1609 51395 1643
rect 51429 1609 51458 1643
rect 51182 1578 51458 1609
rect 51524 1558 51574 1758
rect 51606 1711 51664 1726
rect 51606 1677 51618 1711
rect 51652 1677 51664 1711
rect 51606 1660 51664 1677
rect 51718 1630 51776 1648
rect 51718 1596 51730 1630
rect 51764 1596 51776 1630
rect 51718 1586 51776 1596
rect 51806 1558 51852 1758
rect 52102 1774 52166 1780
rect 52102 1722 52108 1774
rect 52160 1722 52166 1774
rect 52102 1716 52166 1722
rect 51996 1643 52272 1674
rect 51996 1609 52025 1643
rect 52059 1609 52117 1643
rect 52151 1609 52209 1643
rect 52243 1609 52272 1643
rect 51996 1606 52272 1609
rect 51164 1541 51228 1548
rect 51164 1508 51170 1541
rect 51222 1508 51228 1541
rect 51340 1541 51404 1548
rect 51340 1508 51346 1541
rect 51222 1489 51346 1508
rect 51398 1489 51404 1541
rect 51170 1480 51404 1489
rect 51524 1546 51626 1558
rect 51524 1512 51586 1546
rect 51620 1512 51626 1546
rect 51524 1474 51626 1512
rect 51676 1546 51722 1558
rect 51676 1512 51682 1546
rect 51716 1512 51722 1546
rect 51676 1492 51722 1512
rect 51772 1546 51852 1558
rect 51772 1512 51778 1546
rect 51812 1512 51852 1546
rect 51524 1442 51586 1474
rect 51320 1440 51586 1442
rect 51620 1440 51626 1474
rect 51320 1428 51626 1440
rect 51666 1486 51732 1492
rect 51666 1434 51674 1486
rect 51726 1434 51732 1486
rect 51666 1428 51732 1434
rect 51772 1474 51852 1512
rect 51772 1440 51778 1474
rect 51812 1440 51852 1474
rect 51968 1578 52272 1606
rect 51772 1428 51818 1440
rect 51320 1414 51574 1428
rect 51164 1408 51230 1414
rect 51164 1356 51172 1408
rect 51224 1356 51230 1408
rect 51164 1350 51230 1356
rect 50312 1141 50342 1144
rect 50394 1141 50936 1144
rect 50312 1107 50341 1141
rect 50394 1107 50433 1141
rect 50467 1107 50525 1141
rect 50559 1139 50936 1141
rect 50559 1107 50687 1139
rect 50312 1092 50342 1107
rect 50394 1105 50687 1107
rect 50721 1105 50779 1139
rect 50813 1105 50871 1139
rect 50905 1105 50936 1139
rect 50394 1092 50936 1105
rect 50312 1074 50936 1092
rect 51004 1150 51280 1164
rect 51004 1133 51196 1150
rect 51248 1133 51280 1150
rect 51004 1099 51033 1133
rect 51067 1099 51125 1133
rect 51159 1099 51196 1133
rect 51251 1099 51280 1133
rect 51004 1098 51196 1099
rect 51248 1098 51280 1099
rect 51004 1068 51280 1098
rect 51320 1064 51348 1414
rect 51620 1390 51684 1400
rect 51620 1356 51634 1390
rect 51668 1356 51940 1390
rect 51620 1338 51684 1356
rect 51536 1292 51608 1304
rect 51536 1240 51546 1292
rect 51598 1240 51608 1292
rect 51536 1228 51608 1240
rect 51906 1174 51940 1356
rect 51968 1274 51996 1578
rect 51968 1264 52036 1274
rect 51968 1230 51984 1264
rect 52018 1230 52036 1264
rect 51968 1216 52036 1230
rect 51380 1146 51940 1174
rect 51380 1143 51446 1146
rect 51380 1109 51396 1143
rect 51430 1109 51446 1143
rect 51380 1100 51446 1109
rect 51614 1091 51704 1112
rect 49812 983 50052 1000
rect 50096 1056 50162 1062
rect 50096 1004 50104 1056
rect 50156 1004 50162 1056
rect 50096 998 50110 1004
rect 49546 943 49592 976
rect 49546 909 49552 943
rect 49586 909 49592 943
rect 49812 949 49824 983
rect 49858 972 50052 983
rect 50104 981 50110 998
rect 50144 998 50162 1004
rect 50192 1015 50238 1062
rect 51320 1036 51392 1064
rect 50144 981 50150 998
rect 49858 949 50050 972
rect 49812 940 50050 949
rect 49546 862 49592 909
rect 49760 902 49826 910
rect 49674 898 49720 902
rect 48790 840 48862 844
rect 48250 815 48316 828
rect 48250 781 48266 815
rect 48300 781 48316 815
rect 48250 772 48316 781
rect 48790 788 48799 840
rect 48851 788 48862 840
rect 48790 776 48862 788
rect 48986 838 49060 858
rect 49634 855 49720 898
rect 48986 804 48998 838
rect 49032 804 49060 838
rect 48986 780 49060 804
rect 49096 844 49164 850
rect 49096 792 49103 844
rect 49155 838 49164 844
rect 49155 832 49248 838
rect 49155 798 49194 832
rect 49228 798 49248 832
rect 49155 792 49248 798
rect 49096 788 49248 792
rect 49492 815 49558 826
rect 49096 786 49164 788
rect 49492 781 49508 815
rect 49542 781 49558 815
rect 49492 768 49558 781
rect 49634 821 49680 855
rect 49714 821 49720 855
rect 49760 850 49766 902
rect 49818 850 49826 902
rect 49760 842 49776 850
rect 49634 783 49720 821
rect 49634 749 49680 783
rect 49714 749 49720 783
rect 48572 728 48630 742
rect 48572 708 48584 728
rect 48102 694 48584 708
rect 48618 694 48630 728
rect 48102 674 48630 694
rect 49634 702 49720 749
rect 49770 821 49776 842
rect 49810 842 49826 850
rect 49866 855 49962 902
rect 49810 821 49816 842
rect 49770 783 49816 821
rect 49770 749 49776 783
rect 49810 749 49816 783
rect 49770 702 49816 749
rect 49866 821 49872 855
rect 49906 821 49962 855
rect 49866 783 49962 821
rect 49866 749 49872 783
rect 49906 749 49962 783
rect 49866 702 49962 749
rect 47994 372 48040 384
rect 48102 344 48162 674
rect 49634 648 49684 702
rect 48208 624 48284 630
rect 48208 572 48216 624
rect 48268 572 48284 624
rect 48208 566 48284 572
rect 48424 597 49046 628
rect 47842 334 48162 344
rect 47842 300 47856 334
rect 47890 300 48162 334
rect 47842 282 48162 300
rect 48424 563 48453 597
rect 48487 563 48545 597
rect 48579 563 48637 597
rect 48671 595 49046 597
rect 48671 563 48799 595
rect 48424 561 48799 563
rect 48833 561 48891 595
rect 48925 561 48983 595
rect 49017 561 49046 595
rect 48424 530 49046 561
rect 49116 602 49392 620
rect 49116 589 49239 602
rect 49291 589 49392 602
rect 49468 598 49526 606
rect 49116 555 49145 589
rect 49179 555 49237 589
rect 49291 555 49329 589
rect 49363 555 49392 589
rect 49116 550 49239 555
rect 49291 550 49392 555
rect 48424 254 48522 530
rect 49116 524 49392 550
rect 49460 592 49534 598
rect 49460 540 49471 592
rect 49523 540 49534 592
rect 49614 582 49684 648
rect 49716 655 49774 670
rect 49716 621 49728 655
rect 49762 621 49774 655
rect 49716 604 49774 621
rect 49460 534 49534 540
rect 49468 528 49526 534
rect 49184 254 49268 524
rect 49634 502 49684 582
rect 49828 574 49886 592
rect 49828 540 49840 574
rect 49874 540 49886 574
rect 49828 530 49886 540
rect 49916 502 49962 702
rect 49634 490 49736 502
rect 49634 456 49696 490
rect 49730 456 49736 490
rect 49634 418 49736 456
rect 49786 490 49832 502
rect 49786 456 49792 490
rect 49826 456 49832 490
rect 49786 436 49832 456
rect 49882 490 49962 502
rect 49882 456 49888 490
rect 49922 456 49962 490
rect 49634 384 49696 418
rect 49730 384 49736 418
rect 49634 372 49736 384
rect 49776 430 49842 436
rect 49776 378 49784 430
rect 49836 378 49842 430
rect 49776 372 49842 378
rect 49882 418 49962 456
rect 49882 384 49888 418
rect 49922 384 49962 418
rect 49990 708 50050 940
rect 50104 943 50150 981
rect 50104 909 50110 943
rect 50144 909 50150 943
rect 50104 862 50150 909
rect 50192 981 50198 1015
rect 50232 981 50238 1015
rect 50192 943 50238 981
rect 50192 909 50198 943
rect 50232 909 50238 943
rect 50192 862 50238 909
rect 51346 1015 51392 1036
rect 51346 981 51352 1015
rect 51386 981 51392 1015
rect 51346 943 51392 981
rect 51346 909 51352 943
rect 51386 909 51392 943
rect 51346 862 51392 909
rect 51434 1042 51480 1062
rect 51614 1057 51643 1091
rect 51677 1057 51704 1091
rect 51434 1036 51502 1042
rect 51614 1036 51704 1057
rect 51434 1015 51442 1036
rect 51434 981 51440 1015
rect 51494 984 51502 1036
rect 51474 981 51502 984
rect 51434 976 51502 981
rect 51700 1000 51758 1002
rect 51906 1000 51940 1146
rect 52026 1143 52092 1154
rect 52026 1109 52042 1143
rect 52076 1109 52092 1143
rect 52026 1098 52092 1109
rect 52200 1144 52824 1176
rect 52912 1164 52990 2122
rect 53504 2113 53533 2122
rect 53567 2122 55421 2147
rect 53567 2113 53594 2122
rect 53504 2092 53594 2113
rect 53590 2056 53648 2058
rect 53590 2039 53652 2056
rect 53590 2005 53602 2039
rect 53636 2005 53652 2039
rect 53590 1996 53652 2005
rect 53090 1958 53456 1962
rect 53538 1958 53604 1966
rect 53090 1930 53498 1958
rect 53090 1892 53118 1930
rect 53412 1911 53498 1930
rect 53090 1884 53156 1892
rect 53090 1850 53105 1884
rect 53139 1850 53156 1884
rect 53090 1838 53156 1850
rect 53262 1888 53330 1894
rect 53262 1836 53272 1888
rect 53324 1836 53330 1888
rect 53262 1830 53330 1836
rect 53412 1877 53458 1911
rect 53492 1877 53498 1911
rect 53538 1906 53544 1958
rect 53596 1906 53604 1958
rect 53538 1898 53554 1906
rect 53412 1839 53498 1877
rect 53412 1805 53458 1839
rect 53492 1805 53498 1839
rect 53172 1776 53240 1782
rect 53172 1724 53180 1776
rect 53232 1724 53240 1776
rect 53172 1714 53240 1724
rect 53412 1758 53498 1805
rect 53548 1877 53554 1898
rect 53588 1898 53604 1906
rect 53644 1926 53972 1958
rect 53644 1911 53740 1926
rect 53588 1877 53594 1898
rect 53548 1839 53594 1877
rect 53548 1805 53554 1839
rect 53588 1805 53594 1839
rect 53548 1758 53594 1805
rect 53644 1877 53650 1911
rect 53684 1877 53740 1911
rect 53944 1890 53972 1926
rect 53644 1839 53740 1877
rect 53644 1805 53650 1839
rect 53684 1805 53740 1839
rect 53902 1882 53972 1890
rect 53902 1848 53917 1882
rect 53951 1848 53972 1882
rect 53902 1830 53972 1848
rect 54078 1890 54142 1896
rect 54078 1838 54084 1890
rect 54136 1838 54142 1890
rect 54078 1832 54142 1838
rect 53644 1758 53740 1805
rect 53070 1643 53346 1674
rect 53070 1609 53099 1643
rect 53133 1609 53191 1643
rect 53225 1609 53283 1643
rect 53317 1609 53346 1643
rect 53070 1578 53346 1609
rect 53412 1558 53462 1758
rect 53494 1711 53552 1726
rect 53494 1677 53506 1711
rect 53540 1677 53552 1711
rect 53494 1660 53552 1677
rect 53606 1630 53664 1648
rect 53606 1596 53618 1630
rect 53652 1596 53664 1630
rect 53606 1586 53664 1596
rect 53694 1558 53740 1758
rect 53990 1774 54054 1780
rect 53990 1722 53996 1774
rect 54048 1722 54054 1774
rect 53990 1716 54054 1722
rect 53884 1643 54160 1674
rect 53884 1609 53913 1643
rect 53947 1609 54005 1643
rect 54039 1609 54097 1643
rect 54131 1609 54160 1643
rect 53884 1606 54160 1609
rect 53052 1541 53116 1548
rect 53052 1508 53058 1541
rect 53110 1508 53116 1541
rect 53228 1541 53292 1548
rect 53228 1508 53234 1541
rect 53110 1489 53234 1508
rect 53286 1489 53292 1541
rect 53058 1480 53292 1489
rect 53412 1546 53514 1558
rect 53412 1512 53474 1546
rect 53508 1512 53514 1546
rect 53412 1474 53514 1512
rect 53564 1546 53610 1558
rect 53564 1512 53570 1546
rect 53604 1512 53610 1546
rect 53564 1492 53610 1512
rect 53660 1546 53740 1558
rect 53660 1512 53666 1546
rect 53700 1512 53740 1546
rect 53412 1442 53474 1474
rect 53208 1440 53474 1442
rect 53508 1440 53514 1474
rect 53208 1428 53514 1440
rect 53554 1486 53620 1492
rect 53554 1434 53562 1486
rect 53614 1434 53620 1486
rect 53554 1428 53620 1434
rect 53660 1474 53740 1512
rect 53660 1440 53666 1474
rect 53700 1440 53740 1474
rect 53856 1578 54160 1606
rect 53660 1428 53706 1440
rect 53208 1414 53462 1428
rect 53052 1408 53118 1414
rect 53052 1356 53060 1408
rect 53112 1356 53118 1408
rect 53052 1350 53118 1356
rect 52200 1141 52230 1144
rect 52282 1141 52824 1144
rect 52200 1107 52229 1141
rect 52282 1107 52321 1141
rect 52355 1107 52413 1141
rect 52447 1139 52824 1141
rect 52447 1107 52575 1139
rect 52200 1092 52230 1107
rect 52282 1105 52575 1107
rect 52609 1105 52667 1139
rect 52701 1105 52759 1139
rect 52793 1105 52824 1139
rect 52282 1092 52824 1105
rect 52200 1074 52824 1092
rect 52892 1150 53168 1164
rect 52892 1133 53084 1150
rect 53136 1133 53168 1150
rect 52892 1099 52921 1133
rect 52955 1099 53013 1133
rect 53047 1099 53084 1133
rect 53139 1099 53168 1133
rect 52892 1098 53084 1099
rect 53136 1098 53168 1099
rect 52892 1068 53168 1098
rect 53208 1064 53236 1414
rect 53508 1390 53572 1400
rect 53508 1356 53522 1390
rect 53556 1356 53828 1390
rect 53508 1338 53572 1356
rect 53424 1292 53496 1304
rect 53424 1240 53434 1292
rect 53486 1240 53496 1292
rect 53424 1228 53496 1240
rect 53794 1174 53828 1356
rect 53856 1274 53884 1578
rect 53856 1264 53924 1274
rect 53856 1230 53872 1264
rect 53906 1230 53924 1264
rect 53856 1216 53924 1230
rect 53268 1146 53828 1174
rect 53268 1143 53334 1146
rect 53268 1109 53284 1143
rect 53318 1109 53334 1143
rect 53268 1100 53334 1109
rect 53502 1091 53592 1112
rect 51700 983 51940 1000
rect 51984 1056 52050 1062
rect 51984 1004 51992 1056
rect 52044 1004 52050 1056
rect 51984 998 51998 1004
rect 51434 943 51480 976
rect 51434 909 51440 943
rect 51474 909 51480 943
rect 51700 949 51712 983
rect 51746 972 51940 983
rect 51992 981 51998 998
rect 52032 998 52050 1004
rect 52080 1015 52126 1062
rect 53208 1036 53280 1064
rect 52032 981 52038 998
rect 51746 949 51938 972
rect 51700 940 51938 949
rect 51434 862 51480 909
rect 51648 902 51714 910
rect 51562 898 51608 902
rect 50678 840 50750 844
rect 50138 815 50204 828
rect 50138 781 50154 815
rect 50188 781 50204 815
rect 50138 772 50204 781
rect 50678 788 50687 840
rect 50739 788 50750 840
rect 50678 776 50750 788
rect 50874 838 50948 858
rect 51522 855 51608 898
rect 50874 804 50886 838
rect 50920 804 50948 838
rect 50874 780 50948 804
rect 50984 844 51052 850
rect 50984 792 50991 844
rect 51043 838 51052 844
rect 51043 832 51136 838
rect 51043 798 51082 832
rect 51116 798 51136 832
rect 51043 792 51136 798
rect 50984 788 51136 792
rect 51380 815 51446 826
rect 50984 786 51052 788
rect 51380 781 51396 815
rect 51430 781 51446 815
rect 51380 768 51446 781
rect 51522 821 51568 855
rect 51602 821 51608 855
rect 51648 850 51654 902
rect 51706 850 51714 902
rect 51648 842 51664 850
rect 51522 783 51608 821
rect 51522 749 51568 783
rect 51602 749 51608 783
rect 50460 728 50518 742
rect 50460 708 50472 728
rect 49990 694 50472 708
rect 50506 694 50518 728
rect 49990 674 50518 694
rect 51522 702 51608 749
rect 51658 821 51664 842
rect 51698 842 51714 850
rect 51754 855 51850 902
rect 51698 821 51704 842
rect 51658 783 51704 821
rect 51658 749 51664 783
rect 51698 749 51704 783
rect 51658 702 51704 749
rect 51754 821 51760 855
rect 51794 821 51850 855
rect 51754 783 51850 821
rect 51754 749 51760 783
rect 51794 749 51850 783
rect 51754 702 51850 749
rect 49882 372 49928 384
rect 49990 344 50050 674
rect 51522 648 51572 702
rect 50096 624 50172 630
rect 50096 572 50104 624
rect 50156 572 50172 624
rect 50096 566 50172 572
rect 50312 597 50934 628
rect 49730 334 50050 344
rect 49730 300 49744 334
rect 49778 300 50050 334
rect 49730 282 50050 300
rect 50312 563 50341 597
rect 50375 563 50433 597
rect 50467 563 50525 597
rect 50559 595 50934 597
rect 50559 563 50687 595
rect 50312 561 50687 563
rect 50721 561 50779 595
rect 50813 561 50871 595
rect 50905 561 50934 595
rect 50312 530 50934 561
rect 51004 602 51280 620
rect 51004 589 51127 602
rect 51179 589 51280 602
rect 51356 598 51414 606
rect 51004 555 51033 589
rect 51067 555 51125 589
rect 51179 555 51217 589
rect 51251 555 51280 589
rect 51004 550 51127 555
rect 51179 550 51280 555
rect 50312 254 50410 530
rect 51004 524 51280 550
rect 51348 592 51422 598
rect 51348 540 51359 592
rect 51411 540 51422 592
rect 51502 582 51572 648
rect 51604 655 51662 670
rect 51604 621 51616 655
rect 51650 621 51662 655
rect 51604 604 51662 621
rect 51348 534 51422 540
rect 51356 528 51414 534
rect 51072 254 51156 524
rect 51522 502 51572 582
rect 51716 574 51774 592
rect 51716 540 51728 574
rect 51762 540 51774 574
rect 51716 530 51774 540
rect 51804 502 51850 702
rect 51522 490 51624 502
rect 51522 456 51584 490
rect 51618 456 51624 490
rect 51522 418 51624 456
rect 51674 490 51720 502
rect 51674 456 51680 490
rect 51714 456 51720 490
rect 51674 436 51720 456
rect 51770 490 51850 502
rect 51770 456 51776 490
rect 51810 456 51850 490
rect 51522 384 51584 418
rect 51618 384 51624 418
rect 51522 372 51624 384
rect 51664 430 51730 436
rect 51664 378 51672 430
rect 51724 378 51730 430
rect 51664 372 51730 378
rect 51770 418 51850 456
rect 51770 384 51776 418
rect 51810 384 51850 418
rect 51878 708 51938 940
rect 51992 943 52038 981
rect 51992 909 51998 943
rect 52032 909 52038 943
rect 51992 862 52038 909
rect 52080 981 52086 1015
rect 52120 981 52126 1015
rect 52080 943 52126 981
rect 52080 909 52086 943
rect 52120 909 52126 943
rect 52080 862 52126 909
rect 53234 1015 53280 1036
rect 53234 981 53240 1015
rect 53274 981 53280 1015
rect 53234 943 53280 981
rect 53234 909 53240 943
rect 53274 909 53280 943
rect 53234 862 53280 909
rect 53322 1042 53368 1062
rect 53502 1057 53531 1091
rect 53565 1057 53592 1091
rect 53322 1036 53390 1042
rect 53502 1036 53592 1057
rect 53322 1015 53330 1036
rect 53322 981 53328 1015
rect 53382 984 53390 1036
rect 53362 981 53390 984
rect 53322 976 53390 981
rect 53588 1000 53646 1002
rect 53794 1000 53828 1146
rect 53914 1143 53980 1154
rect 53914 1109 53930 1143
rect 53964 1109 53980 1143
rect 53914 1098 53980 1109
rect 54088 1144 54712 1176
rect 54800 1164 54878 2122
rect 55392 2113 55421 2122
rect 55455 2122 57309 2147
rect 55455 2113 55482 2122
rect 55392 2092 55482 2113
rect 55478 2056 55536 2058
rect 55478 2039 55540 2056
rect 55478 2005 55490 2039
rect 55524 2005 55540 2039
rect 55478 1996 55540 2005
rect 54978 1958 55344 1962
rect 55426 1958 55492 1966
rect 54978 1930 55386 1958
rect 54978 1892 55006 1930
rect 55300 1911 55386 1930
rect 54978 1884 55044 1892
rect 54978 1850 54993 1884
rect 55027 1850 55044 1884
rect 54978 1838 55044 1850
rect 55150 1888 55218 1894
rect 55150 1836 55160 1888
rect 55212 1836 55218 1888
rect 55150 1830 55218 1836
rect 55300 1877 55346 1911
rect 55380 1877 55386 1911
rect 55426 1906 55432 1958
rect 55484 1906 55492 1958
rect 55426 1898 55442 1906
rect 55300 1839 55386 1877
rect 55300 1805 55346 1839
rect 55380 1805 55386 1839
rect 55060 1776 55128 1782
rect 55060 1724 55068 1776
rect 55120 1724 55128 1776
rect 55060 1714 55128 1724
rect 55300 1758 55386 1805
rect 55436 1877 55442 1898
rect 55476 1898 55492 1906
rect 55532 1926 55860 1958
rect 55532 1911 55628 1926
rect 55476 1877 55482 1898
rect 55436 1839 55482 1877
rect 55436 1805 55442 1839
rect 55476 1805 55482 1839
rect 55436 1758 55482 1805
rect 55532 1877 55538 1911
rect 55572 1877 55628 1911
rect 55832 1890 55860 1926
rect 55532 1839 55628 1877
rect 55532 1805 55538 1839
rect 55572 1805 55628 1839
rect 55790 1882 55860 1890
rect 55790 1848 55805 1882
rect 55839 1848 55860 1882
rect 55790 1830 55860 1848
rect 55966 1890 56030 1896
rect 55966 1838 55972 1890
rect 56024 1838 56030 1890
rect 55966 1832 56030 1838
rect 55532 1758 55628 1805
rect 54958 1643 55234 1674
rect 54958 1609 54987 1643
rect 55021 1609 55079 1643
rect 55113 1609 55171 1643
rect 55205 1609 55234 1643
rect 54958 1578 55234 1609
rect 55300 1558 55350 1758
rect 55382 1711 55440 1726
rect 55382 1677 55394 1711
rect 55428 1677 55440 1711
rect 55382 1660 55440 1677
rect 55494 1630 55552 1648
rect 55494 1596 55506 1630
rect 55540 1596 55552 1630
rect 55494 1586 55552 1596
rect 55582 1558 55628 1758
rect 55878 1774 55942 1780
rect 55878 1722 55884 1774
rect 55936 1722 55942 1774
rect 55878 1716 55942 1722
rect 55772 1643 56048 1674
rect 55772 1609 55801 1643
rect 55835 1609 55893 1643
rect 55927 1609 55985 1643
rect 56019 1609 56048 1643
rect 55772 1606 56048 1609
rect 54940 1541 55004 1548
rect 54940 1508 54946 1541
rect 54998 1508 55004 1541
rect 55116 1541 55180 1548
rect 55116 1508 55122 1541
rect 54998 1489 55122 1508
rect 55174 1489 55180 1541
rect 54946 1480 55180 1489
rect 55300 1546 55402 1558
rect 55300 1512 55362 1546
rect 55396 1512 55402 1546
rect 55300 1474 55402 1512
rect 55452 1546 55498 1558
rect 55452 1512 55458 1546
rect 55492 1512 55498 1546
rect 55452 1492 55498 1512
rect 55548 1546 55628 1558
rect 55548 1512 55554 1546
rect 55588 1512 55628 1546
rect 55300 1442 55362 1474
rect 55096 1440 55362 1442
rect 55396 1440 55402 1474
rect 55096 1428 55402 1440
rect 55442 1486 55508 1492
rect 55442 1434 55450 1486
rect 55502 1434 55508 1486
rect 55442 1428 55508 1434
rect 55548 1474 55628 1512
rect 55548 1440 55554 1474
rect 55588 1440 55628 1474
rect 55744 1578 56048 1606
rect 55548 1428 55594 1440
rect 55096 1414 55350 1428
rect 54940 1408 55006 1414
rect 54940 1356 54948 1408
rect 55000 1356 55006 1408
rect 54940 1350 55006 1356
rect 54088 1141 54118 1144
rect 54170 1141 54712 1144
rect 54088 1107 54117 1141
rect 54170 1107 54209 1141
rect 54243 1107 54301 1141
rect 54335 1139 54712 1141
rect 54335 1107 54463 1139
rect 54088 1092 54118 1107
rect 54170 1105 54463 1107
rect 54497 1105 54555 1139
rect 54589 1105 54647 1139
rect 54681 1105 54712 1139
rect 54170 1092 54712 1105
rect 54088 1074 54712 1092
rect 54780 1150 55056 1164
rect 54780 1133 54972 1150
rect 55024 1133 55056 1150
rect 54780 1099 54809 1133
rect 54843 1099 54901 1133
rect 54935 1099 54972 1133
rect 55027 1099 55056 1133
rect 54780 1098 54972 1099
rect 55024 1098 55056 1099
rect 54780 1068 55056 1098
rect 55096 1064 55124 1414
rect 55396 1390 55460 1400
rect 55396 1356 55410 1390
rect 55444 1356 55716 1390
rect 55396 1338 55460 1356
rect 55312 1292 55384 1304
rect 55312 1240 55322 1292
rect 55374 1240 55384 1292
rect 55312 1228 55384 1240
rect 55682 1174 55716 1356
rect 55744 1274 55772 1578
rect 55744 1264 55812 1274
rect 55744 1230 55760 1264
rect 55794 1230 55812 1264
rect 55744 1216 55812 1230
rect 55156 1146 55716 1174
rect 55156 1143 55222 1146
rect 55156 1109 55172 1143
rect 55206 1109 55222 1143
rect 55156 1100 55222 1109
rect 55390 1091 55480 1112
rect 53588 983 53828 1000
rect 53872 1056 53938 1062
rect 53872 1004 53880 1056
rect 53932 1004 53938 1056
rect 53872 998 53886 1004
rect 53322 943 53368 976
rect 53322 909 53328 943
rect 53362 909 53368 943
rect 53588 949 53600 983
rect 53634 972 53828 983
rect 53880 981 53886 998
rect 53920 998 53938 1004
rect 53968 1015 54014 1062
rect 55096 1036 55168 1064
rect 53920 981 53926 998
rect 53634 949 53826 972
rect 53588 940 53826 949
rect 53322 862 53368 909
rect 53536 902 53602 910
rect 53450 898 53496 902
rect 52566 840 52638 844
rect 52026 815 52092 828
rect 52026 781 52042 815
rect 52076 781 52092 815
rect 52026 772 52092 781
rect 52566 788 52575 840
rect 52627 788 52638 840
rect 52566 776 52638 788
rect 52762 838 52836 858
rect 53410 855 53496 898
rect 52762 804 52774 838
rect 52808 804 52836 838
rect 52762 780 52836 804
rect 52872 844 52940 850
rect 52872 792 52879 844
rect 52931 838 52940 844
rect 52931 832 53024 838
rect 52931 798 52970 832
rect 53004 798 53024 832
rect 52931 792 53024 798
rect 52872 788 53024 792
rect 53268 815 53334 826
rect 52872 786 52940 788
rect 53268 781 53284 815
rect 53318 781 53334 815
rect 53268 768 53334 781
rect 53410 821 53456 855
rect 53490 821 53496 855
rect 53536 850 53542 902
rect 53594 850 53602 902
rect 53536 842 53552 850
rect 53410 783 53496 821
rect 53410 749 53456 783
rect 53490 749 53496 783
rect 52348 728 52406 742
rect 52348 708 52360 728
rect 51878 694 52360 708
rect 52394 694 52406 728
rect 51878 674 52406 694
rect 53410 702 53496 749
rect 53546 821 53552 842
rect 53586 842 53602 850
rect 53642 855 53738 902
rect 53586 821 53592 842
rect 53546 783 53592 821
rect 53546 749 53552 783
rect 53586 749 53592 783
rect 53546 702 53592 749
rect 53642 821 53648 855
rect 53682 821 53738 855
rect 53642 783 53738 821
rect 53642 749 53648 783
rect 53682 749 53738 783
rect 53642 702 53738 749
rect 51770 372 51816 384
rect 51878 344 51938 674
rect 53410 648 53460 702
rect 51984 624 52060 630
rect 51984 572 51992 624
rect 52044 572 52060 624
rect 51984 566 52060 572
rect 52200 597 52822 628
rect 51618 334 51938 344
rect 51618 300 51632 334
rect 51666 300 51938 334
rect 51618 282 51938 300
rect 52200 563 52229 597
rect 52263 563 52321 597
rect 52355 563 52413 597
rect 52447 595 52822 597
rect 52447 563 52575 595
rect 52200 561 52575 563
rect 52609 561 52667 595
rect 52701 561 52759 595
rect 52793 561 52822 595
rect 52200 530 52822 561
rect 52892 602 53168 620
rect 52892 589 53015 602
rect 53067 589 53168 602
rect 53244 598 53302 606
rect 52892 555 52921 589
rect 52955 555 53013 589
rect 53067 555 53105 589
rect 53139 555 53168 589
rect 52892 550 53015 555
rect 53067 550 53168 555
rect 52200 254 52298 530
rect 52892 524 53168 550
rect 53236 592 53310 598
rect 53236 540 53247 592
rect 53299 540 53310 592
rect 53390 582 53460 648
rect 53492 655 53550 670
rect 53492 621 53504 655
rect 53538 621 53550 655
rect 53492 604 53550 621
rect 53236 534 53310 540
rect 53244 528 53302 534
rect 52960 254 53044 524
rect 53410 502 53460 582
rect 53604 574 53662 592
rect 53604 540 53616 574
rect 53650 540 53662 574
rect 53604 530 53662 540
rect 53692 502 53738 702
rect 53410 490 53512 502
rect 53410 456 53472 490
rect 53506 456 53512 490
rect 53410 418 53512 456
rect 53562 490 53608 502
rect 53562 456 53568 490
rect 53602 456 53608 490
rect 53562 436 53608 456
rect 53658 490 53738 502
rect 53658 456 53664 490
rect 53698 456 53738 490
rect 53410 384 53472 418
rect 53506 384 53512 418
rect 53410 372 53512 384
rect 53552 430 53618 436
rect 53552 378 53560 430
rect 53612 378 53618 430
rect 53552 372 53618 378
rect 53658 418 53738 456
rect 53658 384 53664 418
rect 53698 384 53738 418
rect 53766 708 53826 940
rect 53880 943 53926 981
rect 53880 909 53886 943
rect 53920 909 53926 943
rect 53880 862 53926 909
rect 53968 981 53974 1015
rect 54008 981 54014 1015
rect 53968 943 54014 981
rect 53968 909 53974 943
rect 54008 909 54014 943
rect 53968 862 54014 909
rect 55122 1015 55168 1036
rect 55122 981 55128 1015
rect 55162 981 55168 1015
rect 55122 943 55168 981
rect 55122 909 55128 943
rect 55162 909 55168 943
rect 55122 862 55168 909
rect 55210 1042 55256 1062
rect 55390 1057 55419 1091
rect 55453 1057 55480 1091
rect 55210 1036 55278 1042
rect 55390 1036 55480 1057
rect 55210 1015 55218 1036
rect 55210 981 55216 1015
rect 55270 984 55278 1036
rect 55250 981 55278 984
rect 55210 976 55278 981
rect 55476 1000 55534 1002
rect 55682 1000 55716 1146
rect 55802 1143 55868 1154
rect 55802 1109 55818 1143
rect 55852 1109 55868 1143
rect 55802 1098 55868 1109
rect 55976 1144 56600 1176
rect 56688 1164 56766 2122
rect 57280 2113 57309 2122
rect 57343 2122 59197 2147
rect 57343 2113 57370 2122
rect 57280 2092 57370 2113
rect 57366 2056 57424 2058
rect 57366 2039 57428 2056
rect 57366 2005 57378 2039
rect 57412 2005 57428 2039
rect 57366 1996 57428 2005
rect 56866 1958 57232 1962
rect 57314 1958 57380 1966
rect 56866 1930 57274 1958
rect 56866 1892 56894 1930
rect 57188 1911 57274 1930
rect 56866 1884 56932 1892
rect 56866 1850 56881 1884
rect 56915 1850 56932 1884
rect 56866 1838 56932 1850
rect 57038 1888 57106 1894
rect 57038 1836 57048 1888
rect 57100 1836 57106 1888
rect 57038 1830 57106 1836
rect 57188 1877 57234 1911
rect 57268 1877 57274 1911
rect 57314 1906 57320 1958
rect 57372 1906 57380 1958
rect 57314 1898 57330 1906
rect 57188 1839 57274 1877
rect 57188 1805 57234 1839
rect 57268 1805 57274 1839
rect 56948 1776 57016 1782
rect 56948 1724 56956 1776
rect 57008 1724 57016 1776
rect 56948 1714 57016 1724
rect 57188 1758 57274 1805
rect 57324 1877 57330 1898
rect 57364 1898 57380 1906
rect 57420 1926 57748 1958
rect 57420 1911 57516 1926
rect 57364 1877 57370 1898
rect 57324 1839 57370 1877
rect 57324 1805 57330 1839
rect 57364 1805 57370 1839
rect 57324 1758 57370 1805
rect 57420 1877 57426 1911
rect 57460 1877 57516 1911
rect 57720 1890 57748 1926
rect 57420 1839 57516 1877
rect 57420 1805 57426 1839
rect 57460 1805 57516 1839
rect 57678 1882 57748 1890
rect 57678 1848 57693 1882
rect 57727 1848 57748 1882
rect 57678 1830 57748 1848
rect 57854 1890 57918 1896
rect 57854 1838 57860 1890
rect 57912 1838 57918 1890
rect 57854 1832 57918 1838
rect 57420 1758 57516 1805
rect 56846 1643 57122 1674
rect 56846 1609 56875 1643
rect 56909 1609 56967 1643
rect 57001 1609 57059 1643
rect 57093 1609 57122 1643
rect 56846 1578 57122 1609
rect 57188 1558 57238 1758
rect 57270 1711 57328 1726
rect 57270 1677 57282 1711
rect 57316 1677 57328 1711
rect 57270 1660 57328 1677
rect 57382 1630 57440 1648
rect 57382 1596 57394 1630
rect 57428 1596 57440 1630
rect 57382 1586 57440 1596
rect 57470 1558 57516 1758
rect 57766 1774 57830 1780
rect 57766 1722 57772 1774
rect 57824 1722 57830 1774
rect 57766 1716 57830 1722
rect 57660 1643 57936 1674
rect 57660 1609 57689 1643
rect 57723 1609 57781 1643
rect 57815 1609 57873 1643
rect 57907 1609 57936 1643
rect 57660 1606 57936 1609
rect 56828 1541 56892 1548
rect 56828 1508 56834 1541
rect 56886 1508 56892 1541
rect 57004 1541 57068 1548
rect 57004 1508 57010 1541
rect 56886 1489 57010 1508
rect 57062 1489 57068 1541
rect 56834 1480 57068 1489
rect 57188 1546 57290 1558
rect 57188 1512 57250 1546
rect 57284 1512 57290 1546
rect 57188 1474 57290 1512
rect 57340 1546 57386 1558
rect 57340 1512 57346 1546
rect 57380 1512 57386 1546
rect 57340 1492 57386 1512
rect 57436 1546 57516 1558
rect 57436 1512 57442 1546
rect 57476 1512 57516 1546
rect 57188 1442 57250 1474
rect 56984 1440 57250 1442
rect 57284 1440 57290 1474
rect 56984 1428 57290 1440
rect 57330 1486 57396 1492
rect 57330 1434 57338 1486
rect 57390 1434 57396 1486
rect 57330 1428 57396 1434
rect 57436 1474 57516 1512
rect 57436 1440 57442 1474
rect 57476 1440 57516 1474
rect 57632 1578 57936 1606
rect 57436 1428 57482 1440
rect 56984 1414 57238 1428
rect 56828 1408 56894 1414
rect 56828 1356 56836 1408
rect 56888 1356 56894 1408
rect 56828 1350 56894 1356
rect 55976 1141 56006 1144
rect 56058 1141 56600 1144
rect 55976 1107 56005 1141
rect 56058 1107 56097 1141
rect 56131 1107 56189 1141
rect 56223 1139 56600 1141
rect 56223 1107 56351 1139
rect 55976 1092 56006 1107
rect 56058 1105 56351 1107
rect 56385 1105 56443 1139
rect 56477 1105 56535 1139
rect 56569 1105 56600 1139
rect 56058 1092 56600 1105
rect 55976 1074 56600 1092
rect 56668 1150 56944 1164
rect 56668 1133 56860 1150
rect 56912 1133 56944 1150
rect 56668 1099 56697 1133
rect 56731 1099 56789 1133
rect 56823 1099 56860 1133
rect 56915 1099 56944 1133
rect 56668 1098 56860 1099
rect 56912 1098 56944 1099
rect 56668 1068 56944 1098
rect 56984 1064 57012 1414
rect 57284 1390 57348 1400
rect 57284 1356 57298 1390
rect 57332 1356 57604 1390
rect 57284 1338 57348 1356
rect 57200 1292 57272 1304
rect 57200 1240 57210 1292
rect 57262 1240 57272 1292
rect 57200 1228 57272 1240
rect 57570 1174 57604 1356
rect 57632 1274 57660 1578
rect 57632 1264 57700 1274
rect 57632 1230 57648 1264
rect 57682 1230 57700 1264
rect 57632 1216 57700 1230
rect 57044 1146 57604 1174
rect 57044 1143 57110 1146
rect 57044 1109 57060 1143
rect 57094 1109 57110 1143
rect 57044 1100 57110 1109
rect 57278 1091 57368 1112
rect 55476 983 55716 1000
rect 55760 1056 55826 1062
rect 55760 1004 55768 1056
rect 55820 1004 55826 1056
rect 55760 998 55774 1004
rect 55210 943 55256 976
rect 55210 909 55216 943
rect 55250 909 55256 943
rect 55476 949 55488 983
rect 55522 972 55716 983
rect 55768 981 55774 998
rect 55808 998 55826 1004
rect 55856 1015 55902 1062
rect 56984 1036 57056 1064
rect 55808 981 55814 998
rect 55522 949 55714 972
rect 55476 940 55714 949
rect 55210 862 55256 909
rect 55424 902 55490 910
rect 55338 898 55384 902
rect 54454 840 54526 844
rect 53914 815 53980 828
rect 53914 781 53930 815
rect 53964 781 53980 815
rect 53914 772 53980 781
rect 54454 788 54463 840
rect 54515 788 54526 840
rect 54454 776 54526 788
rect 54650 838 54724 858
rect 55298 855 55384 898
rect 54650 804 54662 838
rect 54696 804 54724 838
rect 54650 780 54724 804
rect 54760 844 54828 850
rect 54760 792 54767 844
rect 54819 838 54828 844
rect 54819 832 54912 838
rect 54819 798 54858 832
rect 54892 798 54912 832
rect 54819 792 54912 798
rect 54760 788 54912 792
rect 55156 815 55222 826
rect 54760 786 54828 788
rect 55156 781 55172 815
rect 55206 781 55222 815
rect 55156 768 55222 781
rect 55298 821 55344 855
rect 55378 821 55384 855
rect 55424 850 55430 902
rect 55482 850 55490 902
rect 55424 842 55440 850
rect 55298 783 55384 821
rect 55298 749 55344 783
rect 55378 749 55384 783
rect 54236 728 54294 742
rect 54236 708 54248 728
rect 53766 694 54248 708
rect 54282 694 54294 728
rect 53766 674 54294 694
rect 55298 702 55384 749
rect 55434 821 55440 842
rect 55474 842 55490 850
rect 55530 855 55626 902
rect 55474 821 55480 842
rect 55434 783 55480 821
rect 55434 749 55440 783
rect 55474 749 55480 783
rect 55434 702 55480 749
rect 55530 821 55536 855
rect 55570 821 55626 855
rect 55530 783 55626 821
rect 55530 749 55536 783
rect 55570 749 55626 783
rect 55530 702 55626 749
rect 53658 372 53704 384
rect 53766 344 53826 674
rect 55298 648 55348 702
rect 53872 624 53948 630
rect 53872 572 53880 624
rect 53932 572 53948 624
rect 53872 566 53948 572
rect 54088 597 54710 628
rect 53506 334 53826 344
rect 53506 300 53520 334
rect 53554 300 53826 334
rect 53506 282 53826 300
rect 54088 563 54117 597
rect 54151 563 54209 597
rect 54243 563 54301 597
rect 54335 595 54710 597
rect 54335 563 54463 595
rect 54088 561 54463 563
rect 54497 561 54555 595
rect 54589 561 54647 595
rect 54681 561 54710 595
rect 54088 530 54710 561
rect 54780 602 55056 620
rect 54780 589 54903 602
rect 54955 589 55056 602
rect 55132 598 55190 606
rect 54780 555 54809 589
rect 54843 555 54901 589
rect 54955 555 54993 589
rect 55027 555 55056 589
rect 54780 550 54903 555
rect 54955 550 55056 555
rect 54088 254 54186 530
rect 54780 524 55056 550
rect 55124 592 55198 598
rect 55124 540 55135 592
rect 55187 540 55198 592
rect 55278 582 55348 648
rect 55380 655 55438 670
rect 55380 621 55392 655
rect 55426 621 55438 655
rect 55380 604 55438 621
rect 55124 534 55198 540
rect 55132 528 55190 534
rect 54848 254 54932 524
rect 55298 502 55348 582
rect 55492 574 55550 592
rect 55492 540 55504 574
rect 55538 540 55550 574
rect 55492 530 55550 540
rect 55580 502 55626 702
rect 55298 490 55400 502
rect 55298 456 55360 490
rect 55394 456 55400 490
rect 55298 418 55400 456
rect 55450 490 55496 502
rect 55450 456 55456 490
rect 55490 456 55496 490
rect 55450 436 55496 456
rect 55546 490 55626 502
rect 55546 456 55552 490
rect 55586 456 55626 490
rect 55298 384 55360 418
rect 55394 384 55400 418
rect 55298 372 55400 384
rect 55440 430 55506 436
rect 55440 378 55448 430
rect 55500 378 55506 430
rect 55440 372 55506 378
rect 55546 418 55626 456
rect 55546 384 55552 418
rect 55586 384 55626 418
rect 55654 708 55714 940
rect 55768 943 55814 981
rect 55768 909 55774 943
rect 55808 909 55814 943
rect 55768 862 55814 909
rect 55856 981 55862 1015
rect 55896 981 55902 1015
rect 55856 943 55902 981
rect 55856 909 55862 943
rect 55896 909 55902 943
rect 55856 862 55902 909
rect 57010 1015 57056 1036
rect 57010 981 57016 1015
rect 57050 981 57056 1015
rect 57010 943 57056 981
rect 57010 909 57016 943
rect 57050 909 57056 943
rect 57010 862 57056 909
rect 57098 1042 57144 1062
rect 57278 1057 57307 1091
rect 57341 1057 57368 1091
rect 57098 1036 57166 1042
rect 57278 1036 57368 1057
rect 57098 1015 57106 1036
rect 57098 981 57104 1015
rect 57158 984 57166 1036
rect 57138 981 57166 984
rect 57098 976 57166 981
rect 57364 1000 57422 1002
rect 57570 1000 57604 1146
rect 57690 1143 57756 1154
rect 57690 1109 57706 1143
rect 57740 1109 57756 1143
rect 57690 1098 57756 1109
rect 57864 1144 58488 1176
rect 58576 1164 58654 2122
rect 59168 2113 59197 2122
rect 59231 2122 60412 2147
rect 59231 2113 59258 2122
rect 59168 2092 59258 2113
rect 59254 2056 59312 2058
rect 59254 2039 59316 2056
rect 59254 2005 59266 2039
rect 59300 2005 59316 2039
rect 59254 1996 59316 2005
rect 58754 1958 59120 1962
rect 59202 1958 59268 1966
rect 58754 1930 59162 1958
rect 58754 1892 58782 1930
rect 59076 1911 59162 1930
rect 58754 1884 58820 1892
rect 58754 1850 58769 1884
rect 58803 1850 58820 1884
rect 58754 1838 58820 1850
rect 58926 1888 58994 1894
rect 58926 1836 58936 1888
rect 58988 1836 58994 1888
rect 58926 1830 58994 1836
rect 59076 1877 59122 1911
rect 59156 1877 59162 1911
rect 59202 1906 59208 1958
rect 59260 1906 59268 1958
rect 59202 1898 59218 1906
rect 59076 1839 59162 1877
rect 59076 1805 59122 1839
rect 59156 1805 59162 1839
rect 58836 1776 58904 1782
rect 58836 1724 58844 1776
rect 58896 1724 58904 1776
rect 58836 1714 58904 1724
rect 59076 1758 59162 1805
rect 59212 1877 59218 1898
rect 59252 1898 59268 1906
rect 59308 1926 59636 1958
rect 59308 1911 59404 1926
rect 59252 1877 59258 1898
rect 59212 1839 59258 1877
rect 59212 1805 59218 1839
rect 59252 1805 59258 1839
rect 59212 1758 59258 1805
rect 59308 1877 59314 1911
rect 59348 1877 59404 1911
rect 59608 1890 59636 1926
rect 59308 1839 59404 1877
rect 59308 1805 59314 1839
rect 59348 1805 59404 1839
rect 59566 1882 59636 1890
rect 59566 1848 59581 1882
rect 59615 1848 59636 1882
rect 59566 1830 59636 1848
rect 59742 1890 59806 1896
rect 59742 1838 59748 1890
rect 59800 1838 59806 1890
rect 59742 1832 59806 1838
rect 59308 1758 59404 1805
rect 58734 1643 59010 1674
rect 58734 1609 58763 1643
rect 58797 1609 58855 1643
rect 58889 1609 58947 1643
rect 58981 1609 59010 1643
rect 58734 1578 59010 1609
rect 59076 1558 59126 1758
rect 59158 1711 59216 1726
rect 59158 1677 59170 1711
rect 59204 1677 59216 1711
rect 59158 1660 59216 1677
rect 59270 1630 59328 1648
rect 59270 1596 59282 1630
rect 59316 1596 59328 1630
rect 59270 1586 59328 1596
rect 59358 1558 59404 1758
rect 59654 1774 59718 1780
rect 59654 1722 59660 1774
rect 59712 1722 59718 1774
rect 59654 1716 59718 1722
rect 59548 1643 59824 1674
rect 59548 1609 59577 1643
rect 59611 1609 59669 1643
rect 59703 1609 59761 1643
rect 59795 1609 59824 1643
rect 59548 1606 59824 1609
rect 58716 1541 58780 1548
rect 58716 1508 58722 1541
rect 58774 1508 58780 1541
rect 58892 1541 58956 1548
rect 58892 1508 58898 1541
rect 58774 1489 58898 1508
rect 58950 1489 58956 1541
rect 58722 1480 58956 1489
rect 59076 1546 59178 1558
rect 59076 1512 59138 1546
rect 59172 1512 59178 1546
rect 59076 1474 59178 1512
rect 59228 1546 59274 1558
rect 59228 1512 59234 1546
rect 59268 1512 59274 1546
rect 59228 1492 59274 1512
rect 59324 1546 59404 1558
rect 59324 1512 59330 1546
rect 59364 1512 59404 1546
rect 59076 1442 59138 1474
rect 58872 1440 59138 1442
rect 59172 1440 59178 1474
rect 58872 1428 59178 1440
rect 59218 1486 59284 1492
rect 59218 1434 59226 1486
rect 59278 1434 59284 1486
rect 59218 1428 59284 1434
rect 59324 1474 59404 1512
rect 59324 1440 59330 1474
rect 59364 1440 59404 1474
rect 59520 1578 59824 1606
rect 59324 1428 59370 1440
rect 58872 1414 59126 1428
rect 58716 1408 58782 1414
rect 58716 1356 58724 1408
rect 58776 1356 58782 1408
rect 58716 1350 58782 1356
rect 57864 1141 57894 1144
rect 57946 1141 58488 1144
rect 57864 1107 57893 1141
rect 57946 1107 57985 1141
rect 58019 1107 58077 1141
rect 58111 1139 58488 1141
rect 58111 1107 58239 1139
rect 57864 1092 57894 1107
rect 57946 1105 58239 1107
rect 58273 1105 58331 1139
rect 58365 1105 58423 1139
rect 58457 1105 58488 1139
rect 57946 1092 58488 1105
rect 57864 1074 58488 1092
rect 58556 1150 58832 1164
rect 58556 1133 58748 1150
rect 58800 1133 58832 1150
rect 58556 1099 58585 1133
rect 58619 1099 58677 1133
rect 58711 1099 58748 1133
rect 58803 1099 58832 1133
rect 58556 1098 58748 1099
rect 58800 1098 58832 1099
rect 58556 1068 58832 1098
rect 58872 1064 58900 1414
rect 59172 1390 59236 1400
rect 59172 1356 59186 1390
rect 59220 1356 59492 1390
rect 59172 1338 59236 1356
rect 59088 1292 59160 1304
rect 59088 1240 59098 1292
rect 59150 1240 59160 1292
rect 59088 1228 59160 1240
rect 59458 1174 59492 1356
rect 59520 1274 59548 1578
rect 59520 1264 59588 1274
rect 59520 1230 59536 1264
rect 59570 1230 59588 1264
rect 59520 1216 59588 1230
rect 58932 1146 59492 1174
rect 58932 1143 58998 1146
rect 58932 1109 58948 1143
rect 58982 1109 58998 1143
rect 58932 1100 58998 1109
rect 59166 1091 59256 1112
rect 57364 983 57604 1000
rect 57648 1056 57714 1062
rect 57648 1004 57656 1056
rect 57708 1004 57714 1056
rect 57648 998 57662 1004
rect 57098 943 57144 976
rect 57098 909 57104 943
rect 57138 909 57144 943
rect 57364 949 57376 983
rect 57410 972 57604 983
rect 57656 981 57662 998
rect 57696 998 57714 1004
rect 57744 1015 57790 1062
rect 58872 1036 58944 1064
rect 57696 981 57702 998
rect 57410 949 57602 972
rect 57364 940 57602 949
rect 57098 862 57144 909
rect 57312 902 57378 910
rect 57226 898 57272 902
rect 56342 840 56414 844
rect 55802 815 55868 828
rect 55802 781 55818 815
rect 55852 781 55868 815
rect 55802 772 55868 781
rect 56342 788 56351 840
rect 56403 788 56414 840
rect 56342 776 56414 788
rect 56538 838 56612 858
rect 57186 855 57272 898
rect 56538 804 56550 838
rect 56584 804 56612 838
rect 56538 780 56612 804
rect 56648 844 56716 850
rect 56648 792 56655 844
rect 56707 838 56716 844
rect 56707 832 56800 838
rect 56707 798 56746 832
rect 56780 798 56800 832
rect 56707 792 56800 798
rect 56648 788 56800 792
rect 57044 815 57110 826
rect 56648 786 56716 788
rect 57044 781 57060 815
rect 57094 781 57110 815
rect 57044 768 57110 781
rect 57186 821 57232 855
rect 57266 821 57272 855
rect 57312 850 57318 902
rect 57370 850 57378 902
rect 57312 842 57328 850
rect 57186 783 57272 821
rect 57186 749 57232 783
rect 57266 749 57272 783
rect 56124 728 56182 742
rect 56124 708 56136 728
rect 55654 694 56136 708
rect 56170 694 56182 728
rect 55654 674 56182 694
rect 57186 702 57272 749
rect 57322 821 57328 842
rect 57362 842 57378 850
rect 57418 855 57514 902
rect 57362 821 57368 842
rect 57322 783 57368 821
rect 57322 749 57328 783
rect 57362 749 57368 783
rect 57322 702 57368 749
rect 57418 821 57424 855
rect 57458 821 57514 855
rect 57418 783 57514 821
rect 57418 749 57424 783
rect 57458 749 57514 783
rect 57418 702 57514 749
rect 55546 372 55592 384
rect 55654 344 55714 674
rect 57186 648 57236 702
rect 55760 624 55836 630
rect 55760 572 55768 624
rect 55820 572 55836 624
rect 55760 566 55836 572
rect 55976 597 56598 628
rect 55394 334 55714 344
rect 55394 300 55408 334
rect 55442 300 55714 334
rect 55394 282 55714 300
rect 55976 563 56005 597
rect 56039 563 56097 597
rect 56131 563 56189 597
rect 56223 595 56598 597
rect 56223 563 56351 595
rect 55976 561 56351 563
rect 56385 561 56443 595
rect 56477 561 56535 595
rect 56569 561 56598 595
rect 55976 530 56598 561
rect 56668 602 56944 620
rect 56668 589 56791 602
rect 56843 589 56944 602
rect 57020 598 57078 606
rect 56668 555 56697 589
rect 56731 555 56789 589
rect 56843 555 56881 589
rect 56915 555 56944 589
rect 56668 550 56791 555
rect 56843 550 56944 555
rect 55976 254 56074 530
rect 56668 524 56944 550
rect 57012 592 57086 598
rect 57012 540 57023 592
rect 57075 540 57086 592
rect 57166 582 57236 648
rect 57268 655 57326 670
rect 57268 621 57280 655
rect 57314 621 57326 655
rect 57268 604 57326 621
rect 57012 534 57086 540
rect 57020 528 57078 534
rect 56736 254 56820 524
rect 57186 502 57236 582
rect 57380 574 57438 592
rect 57380 540 57392 574
rect 57426 540 57438 574
rect 57380 530 57438 540
rect 57468 502 57514 702
rect 57186 490 57288 502
rect 57186 456 57248 490
rect 57282 456 57288 490
rect 57186 418 57288 456
rect 57338 490 57384 502
rect 57338 456 57344 490
rect 57378 456 57384 490
rect 57338 436 57384 456
rect 57434 490 57514 502
rect 57434 456 57440 490
rect 57474 456 57514 490
rect 57186 384 57248 418
rect 57282 384 57288 418
rect 57186 372 57288 384
rect 57328 430 57394 436
rect 57328 378 57336 430
rect 57388 378 57394 430
rect 57328 372 57394 378
rect 57434 418 57514 456
rect 57434 384 57440 418
rect 57474 384 57514 418
rect 57542 708 57602 940
rect 57656 943 57702 981
rect 57656 909 57662 943
rect 57696 909 57702 943
rect 57656 862 57702 909
rect 57744 981 57750 1015
rect 57784 981 57790 1015
rect 57744 943 57790 981
rect 57744 909 57750 943
rect 57784 909 57790 943
rect 57744 862 57790 909
rect 58898 1015 58944 1036
rect 58898 981 58904 1015
rect 58938 981 58944 1015
rect 58898 943 58944 981
rect 58898 909 58904 943
rect 58938 909 58944 943
rect 58898 862 58944 909
rect 58986 1042 59032 1062
rect 59166 1057 59195 1091
rect 59229 1057 59256 1091
rect 58986 1036 59054 1042
rect 59166 1036 59256 1057
rect 58986 1015 58994 1036
rect 58986 981 58992 1015
rect 59046 984 59054 1036
rect 59026 981 59054 984
rect 58986 976 59054 981
rect 59252 1000 59310 1002
rect 59458 1000 59492 1146
rect 59578 1143 59644 1154
rect 59578 1109 59594 1143
rect 59628 1109 59644 1143
rect 59578 1098 59644 1109
rect 59752 1144 60376 1176
rect 59752 1141 59782 1144
rect 59834 1141 60376 1144
rect 59752 1107 59781 1141
rect 59834 1107 59873 1141
rect 59907 1107 59965 1141
rect 59999 1139 60376 1141
rect 59999 1107 60127 1139
rect 59752 1092 59782 1107
rect 59834 1105 60127 1107
rect 60161 1105 60219 1139
rect 60253 1105 60311 1139
rect 60345 1105 60376 1139
rect 59834 1092 60376 1105
rect 59752 1074 60376 1092
rect 59252 983 59492 1000
rect 59536 1056 59602 1062
rect 59536 1004 59544 1056
rect 59596 1004 59602 1056
rect 59536 998 59550 1004
rect 58986 943 59032 976
rect 58986 909 58992 943
rect 59026 909 59032 943
rect 59252 949 59264 983
rect 59298 972 59492 983
rect 59544 981 59550 998
rect 59584 998 59602 1004
rect 59632 1015 59678 1062
rect 59584 981 59590 998
rect 59298 949 59490 972
rect 59252 940 59490 949
rect 58986 862 59032 909
rect 59200 902 59266 910
rect 59114 898 59160 902
rect 58230 840 58302 844
rect 57690 815 57756 828
rect 57690 781 57706 815
rect 57740 781 57756 815
rect 57690 772 57756 781
rect 58230 788 58239 840
rect 58291 788 58302 840
rect 58230 776 58302 788
rect 58426 838 58500 858
rect 59074 855 59160 898
rect 58426 804 58438 838
rect 58472 804 58500 838
rect 58426 780 58500 804
rect 58536 844 58604 850
rect 58536 792 58543 844
rect 58595 838 58604 844
rect 58595 832 58688 838
rect 58595 798 58634 832
rect 58668 798 58688 832
rect 58595 792 58688 798
rect 58536 788 58688 792
rect 58932 815 58998 826
rect 58536 786 58604 788
rect 58932 781 58948 815
rect 58982 781 58998 815
rect 58932 768 58998 781
rect 59074 821 59120 855
rect 59154 821 59160 855
rect 59200 850 59206 902
rect 59258 850 59266 902
rect 59200 842 59216 850
rect 59074 783 59160 821
rect 59074 749 59120 783
rect 59154 749 59160 783
rect 58012 728 58070 742
rect 58012 708 58024 728
rect 57542 694 58024 708
rect 58058 694 58070 728
rect 57542 674 58070 694
rect 59074 702 59160 749
rect 59210 821 59216 842
rect 59250 842 59266 850
rect 59306 855 59402 902
rect 59250 821 59256 842
rect 59210 783 59256 821
rect 59210 749 59216 783
rect 59250 749 59256 783
rect 59210 702 59256 749
rect 59306 821 59312 855
rect 59346 821 59402 855
rect 59306 783 59402 821
rect 59306 749 59312 783
rect 59346 749 59402 783
rect 59306 702 59402 749
rect 57434 372 57480 384
rect 57542 344 57602 674
rect 59074 648 59124 702
rect 57648 624 57724 630
rect 57648 572 57656 624
rect 57708 572 57724 624
rect 57648 566 57724 572
rect 57864 597 58486 628
rect 57282 334 57602 344
rect 57282 300 57296 334
rect 57330 300 57602 334
rect 57282 282 57602 300
rect 57864 563 57893 597
rect 57927 563 57985 597
rect 58019 563 58077 597
rect 58111 595 58486 597
rect 58111 563 58239 595
rect 57864 561 58239 563
rect 58273 561 58331 595
rect 58365 561 58423 595
rect 58457 561 58486 595
rect 57864 530 58486 561
rect 58556 602 58832 620
rect 58556 589 58679 602
rect 58731 589 58832 602
rect 58908 598 58966 606
rect 58556 555 58585 589
rect 58619 555 58677 589
rect 58731 555 58769 589
rect 58803 555 58832 589
rect 58556 550 58679 555
rect 58731 550 58832 555
rect 57864 254 57962 530
rect 58556 524 58832 550
rect 58900 592 58974 598
rect 58900 540 58911 592
rect 58963 540 58974 592
rect 59054 582 59124 648
rect 59156 655 59214 670
rect 59156 621 59168 655
rect 59202 621 59214 655
rect 59156 604 59214 621
rect 58900 534 58974 540
rect 58908 528 58966 534
rect 58624 254 58708 524
rect 59074 502 59124 582
rect 59268 574 59326 592
rect 59268 540 59280 574
rect 59314 540 59326 574
rect 59268 530 59326 540
rect 59356 502 59402 702
rect 59074 490 59176 502
rect 59074 456 59136 490
rect 59170 456 59176 490
rect 59074 418 59176 456
rect 59226 490 59272 502
rect 59226 456 59232 490
rect 59266 456 59272 490
rect 59226 436 59272 456
rect 59322 490 59402 502
rect 59322 456 59328 490
rect 59362 456 59402 490
rect 59074 384 59136 418
rect 59170 384 59176 418
rect 59074 372 59176 384
rect 59216 430 59282 436
rect 59216 378 59224 430
rect 59276 378 59282 430
rect 59216 372 59282 378
rect 59322 418 59402 456
rect 59322 384 59328 418
rect 59362 384 59402 418
rect 59430 708 59490 940
rect 59544 943 59590 981
rect 59544 909 59550 943
rect 59584 909 59590 943
rect 59544 862 59590 909
rect 59632 981 59638 1015
rect 59672 981 59678 1015
rect 59632 943 59678 981
rect 59632 909 59638 943
rect 59672 909 59678 943
rect 59632 862 59678 909
rect 60118 840 60190 844
rect 59578 815 59644 828
rect 59578 781 59594 815
rect 59628 781 59644 815
rect 59578 772 59644 781
rect 60118 788 60127 840
rect 60179 788 60190 840
rect 60118 776 60190 788
rect 60314 838 60604 858
rect 60314 804 60326 838
rect 60360 804 60604 838
rect 60314 780 60604 804
rect 59900 728 59958 742
rect 59900 708 59912 728
rect 59430 694 59912 708
rect 59946 694 59958 728
rect 59430 674 59958 694
rect 59322 372 59368 384
rect 59430 344 59490 674
rect 59536 624 59612 630
rect 59536 572 59544 624
rect 59596 572 59612 624
rect 59536 566 59612 572
rect 59752 597 60374 628
rect 59170 334 59490 344
rect 59170 300 59184 334
rect 59218 300 59490 334
rect 59170 282 59490 300
rect 59752 563 59781 597
rect 59815 563 59873 597
rect 59907 563 59965 597
rect 59999 595 60374 597
rect 59999 563 60127 595
rect 59752 561 60127 563
rect 60161 561 60219 595
rect 60253 561 60311 595
rect 60345 561 60374 595
rect 59752 530 60374 561
rect 59752 254 59850 530
rect 8 225 60412 254
rect 8 191 588 225
rect 622 191 2476 225
rect 2510 191 4364 225
rect 4398 191 6252 225
rect 6286 191 8140 225
rect 8174 191 10028 225
rect 10062 191 11916 225
rect 11950 191 13804 225
rect 13838 191 15686 225
rect 15720 191 17574 225
rect 17608 191 19462 225
rect 19496 191 21350 225
rect 21384 191 23238 225
rect 23272 191 25126 225
rect 25160 191 27014 225
rect 27048 191 28902 225
rect 28936 191 30790 225
rect 30824 191 32678 225
rect 32712 191 34566 225
rect 34600 191 36454 225
rect 36488 191 38342 225
rect 38376 191 40230 225
rect 40264 191 42118 225
rect 42152 191 44006 225
rect 44040 191 45888 225
rect 45922 191 47776 225
rect 47810 191 49664 225
rect 49698 191 51552 225
rect 51586 191 53440 225
rect 53474 191 55328 225
rect 55362 191 57216 225
rect 57250 191 59104 225
rect 59138 191 60412 225
rect 8 180 60412 191
rect 8 64 1535 180
rect 1843 64 3423 180
rect 3731 64 5311 180
rect 5619 64 7199 180
rect 7507 64 9087 180
rect 9395 64 10975 180
rect 11283 64 12863 180
rect 13171 64 14751 180
rect 15059 64 16633 180
rect 16941 64 18521 180
rect 18829 64 20409 180
rect 20717 64 22297 180
rect 22605 64 24185 180
rect 24493 64 26073 180
rect 26381 64 27961 180
rect 28269 64 29849 180
rect 30157 64 31737 180
rect 32045 64 33625 180
rect 33933 64 35513 180
rect 35821 64 37401 180
rect 37709 64 39289 180
rect 39597 64 41177 180
rect 41485 64 43065 180
rect 43373 64 44953 180
rect 45261 64 46835 180
rect 47143 64 48723 180
rect 49031 64 50611 180
rect 50919 64 52499 180
rect 52807 64 54387 180
rect 54695 64 56275 180
rect 56583 64 58163 180
rect 58471 64 60051 180
rect 60359 64 60412 180
rect 8 0 60412 64
<< via1 >>
rect -377 7260 -69 7376
rect 1511 7260 1819 7376
rect 3399 7260 3707 7376
rect 5287 7260 5595 7376
rect 7175 7260 7483 7376
rect 9063 7260 9371 7376
rect 10951 7260 11259 7376
rect 12839 7260 13147 7376
rect 14721 7260 15029 7376
rect 16609 7260 16917 7376
rect 18497 7260 18805 7376
rect 20385 7260 20693 7376
rect 22273 7260 22581 7376
rect 24161 7260 24469 7376
rect 26049 7260 26357 7376
rect 27937 7260 28245 7376
rect 29825 7260 30133 7376
rect 31713 7260 32021 7376
rect 33601 7260 33909 7376
rect 35489 7260 35797 7376
rect 37377 7260 37685 7376
rect 39265 7260 39573 7376
rect 41153 7260 41461 7376
rect 43041 7260 43349 7376
rect 44923 7260 45231 7376
rect 46811 7260 47119 7376
rect 48699 7260 49007 7376
rect 50587 7260 50895 7376
rect 52475 7260 52783 7376
rect 54363 7260 54671 7376
rect 56251 7260 56559 7376
rect 58139 7260 58447 7376
rect 386 6862 438 6868
rect 386 6828 396 6862
rect 396 6828 430 6862
rect 430 6828 438 6862
rect 386 6816 438 6828
rect -197 6648 -145 6652
rect -197 6614 -185 6648
rect -185 6614 -151 6648
rect -151 6614 -145 6648
rect -197 6600 -145 6614
rect 706 7056 758 7062
rect 706 7022 716 7056
rect 716 7022 750 7056
rect 750 7022 758 7056
rect 706 7010 758 7022
rect 1019 6890 1071 6900
rect 1019 6856 1028 6890
rect 1028 6856 1062 6890
rect 1062 6856 1071 6890
rect 1019 6848 1071 6856
rect 1251 6885 1303 6890
rect 1251 6851 1271 6885
rect 1271 6851 1303 6885
rect 1251 6838 1303 6851
rect 2274 6862 2326 6868
rect 2274 6828 2284 6862
rect 2284 6828 2318 6862
rect 2318 6828 2326 6862
rect 2274 6816 2326 6828
rect 724 6585 732 6590
rect 732 6585 766 6590
rect 766 6585 776 6590
rect 724 6538 776 6585
rect 1387 6596 1439 6648
rect 1691 6648 1743 6652
rect 1691 6614 1703 6648
rect 1703 6614 1737 6648
rect 1737 6614 1743 6648
rect 1691 6600 1743 6614
rect 386 6425 398 6436
rect 398 6425 432 6436
rect 432 6425 438 6436
rect 386 6384 438 6425
rect 148 6333 200 6348
rect 148 6299 167 6333
rect 167 6299 200 6333
rect 148 6296 200 6299
rect 936 6425 956 6456
rect 956 6425 988 6456
rect 936 6404 988 6425
rect 2594 7056 2646 7062
rect 2594 7022 2604 7056
rect 2604 7022 2638 7056
rect 2638 7022 2646 7056
rect 2594 7010 2646 7022
rect 2907 6890 2959 6900
rect 2907 6856 2916 6890
rect 2916 6856 2950 6890
rect 2950 6856 2959 6890
rect 2907 6848 2959 6856
rect 3139 6885 3191 6890
rect 3139 6851 3159 6885
rect 3159 6851 3191 6885
rect 3139 6838 3191 6851
rect 4162 6862 4214 6868
rect 4162 6828 4172 6862
rect 4172 6828 4206 6862
rect 4206 6828 4214 6862
rect 4162 6816 4214 6828
rect 2612 6585 2620 6590
rect 2620 6585 2654 6590
rect 2654 6585 2664 6590
rect 2612 6538 2664 6585
rect 3275 6596 3327 6648
rect 3579 6648 3631 6652
rect 3579 6614 3591 6648
rect 3591 6614 3625 6648
rect 3625 6614 3631 6648
rect 3579 6600 3631 6614
rect 2274 6425 2286 6436
rect 2286 6425 2320 6436
rect 2320 6425 2326 6436
rect 2274 6384 2326 6425
rect 832 6193 884 6200
rect 832 6159 842 6193
rect 842 6159 876 6193
rect 876 6159 884 6193
rect 832 6148 884 6159
rect 1182 6341 1234 6342
rect 1182 6307 1213 6341
rect 1213 6307 1234 6341
rect 1182 6290 1234 6307
rect 2036 6333 2088 6348
rect 2036 6299 2055 6333
rect 2055 6299 2088 6333
rect 2036 6296 2088 6299
rect 1206 6076 1258 6084
rect 1206 6042 1214 6076
rect 1214 6042 1248 6076
rect 1248 6042 1258 6076
rect 1206 6032 1258 6042
rect 704 6000 756 6006
rect 704 5966 714 6000
rect 714 5966 748 6000
rect 748 5966 756 6000
rect 704 5954 756 5966
rect 1032 5899 1084 5951
rect 1208 5899 1260 5951
rect 270 5715 322 5718
rect 270 5681 279 5715
rect 279 5681 313 5715
rect 313 5681 322 5715
rect 270 5666 322 5681
rect 182 5592 234 5602
rect 182 5558 193 5592
rect 193 5558 227 5592
rect 227 5558 234 5592
rect 182 5550 234 5558
rect 1086 5710 1138 5716
rect 1086 5676 1097 5710
rect 1097 5676 1131 5710
rect 1131 5676 1138 5710
rect 1086 5664 1138 5676
rect 722 5529 730 5534
rect 730 5529 764 5534
rect 764 5529 774 5534
rect 722 5482 774 5529
rect 994 5594 1046 5604
rect 994 5560 1006 5594
rect 1006 5560 1040 5594
rect 1040 5560 1046 5594
rect 994 5552 1046 5560
rect 2824 6425 2844 6456
rect 2844 6425 2876 6456
rect 2824 6404 2876 6425
rect 4482 7056 4534 7062
rect 4482 7022 4492 7056
rect 4492 7022 4526 7056
rect 4526 7022 4534 7056
rect 4482 7010 4534 7022
rect 4795 6890 4847 6900
rect 4795 6856 4804 6890
rect 4804 6856 4838 6890
rect 4838 6856 4847 6890
rect 4795 6848 4847 6856
rect 5027 6885 5079 6890
rect 5027 6851 5047 6885
rect 5047 6851 5079 6885
rect 5027 6838 5079 6851
rect 6050 6862 6102 6868
rect 6050 6828 6060 6862
rect 6060 6828 6094 6862
rect 6094 6828 6102 6862
rect 6050 6816 6102 6828
rect 4500 6585 4508 6590
rect 4508 6585 4542 6590
rect 4542 6585 4552 6590
rect 4500 6538 4552 6585
rect 5163 6596 5215 6648
rect 5467 6648 5519 6652
rect 5467 6614 5479 6648
rect 5479 6614 5513 6648
rect 5513 6614 5519 6648
rect 5467 6600 5519 6614
rect 4162 6425 4174 6436
rect 4174 6425 4208 6436
rect 4208 6425 4214 6436
rect 4162 6384 4214 6425
rect 2720 6193 2772 6200
rect 2720 6159 2730 6193
rect 2730 6159 2764 6193
rect 2764 6159 2772 6193
rect 2720 6148 2772 6159
rect 3070 6341 3122 6342
rect 3070 6307 3101 6341
rect 3101 6307 3122 6341
rect 3070 6290 3122 6307
rect 3924 6333 3976 6348
rect 3924 6299 3943 6333
rect 3943 6299 3976 6333
rect 3924 6296 3976 6299
rect 3094 6076 3146 6084
rect 3094 6042 3102 6076
rect 3102 6042 3136 6076
rect 3136 6042 3146 6076
rect 3094 6032 3146 6042
rect 2592 6000 2644 6006
rect 2592 5966 2602 6000
rect 2602 5966 2636 6000
rect 2636 5966 2644 6000
rect 2592 5954 2644 5966
rect 2920 5899 2972 5951
rect 3096 5899 3148 5951
rect 2158 5715 2210 5718
rect 2158 5681 2167 5715
rect 2167 5681 2201 5715
rect 2201 5681 2210 5715
rect 2158 5666 2210 5681
rect 2070 5592 2122 5602
rect 2070 5558 2081 5592
rect 2081 5558 2115 5592
rect 2115 5558 2122 5592
rect 2070 5550 2122 5558
rect 2974 5710 3026 5716
rect 2974 5676 2985 5710
rect 2985 5676 3019 5710
rect 3019 5676 3026 5710
rect 2974 5664 3026 5676
rect 2610 5529 2618 5534
rect 2618 5529 2652 5534
rect 2652 5529 2662 5534
rect 2610 5482 2662 5529
rect 2882 5594 2934 5604
rect 2882 5560 2894 5594
rect 2894 5560 2928 5594
rect 2928 5560 2934 5594
rect 2882 5552 2934 5560
rect 4712 6425 4732 6456
rect 4732 6425 4764 6456
rect 4712 6404 4764 6425
rect 6370 7056 6422 7062
rect 6370 7022 6380 7056
rect 6380 7022 6414 7056
rect 6414 7022 6422 7056
rect 6370 7010 6422 7022
rect 6683 6890 6735 6900
rect 6683 6856 6692 6890
rect 6692 6856 6726 6890
rect 6726 6856 6735 6890
rect 6683 6848 6735 6856
rect 6915 6885 6967 6890
rect 6915 6851 6935 6885
rect 6935 6851 6967 6885
rect 6915 6838 6967 6851
rect 7938 6862 7990 6868
rect 7938 6828 7948 6862
rect 7948 6828 7982 6862
rect 7982 6828 7990 6862
rect 7938 6816 7990 6828
rect 6388 6585 6396 6590
rect 6396 6585 6430 6590
rect 6430 6585 6440 6590
rect 6388 6538 6440 6585
rect 7051 6596 7103 6648
rect 7355 6648 7407 6652
rect 7355 6614 7367 6648
rect 7367 6614 7401 6648
rect 7401 6614 7407 6648
rect 7355 6600 7407 6614
rect 6050 6425 6062 6436
rect 6062 6425 6096 6436
rect 6096 6425 6102 6436
rect 6050 6384 6102 6425
rect 4608 6193 4660 6200
rect 4608 6159 4618 6193
rect 4618 6159 4652 6193
rect 4652 6159 4660 6193
rect 4608 6148 4660 6159
rect 4958 6341 5010 6342
rect 4958 6307 4989 6341
rect 4989 6307 5010 6341
rect 4958 6290 5010 6307
rect 5812 6333 5864 6348
rect 5812 6299 5831 6333
rect 5831 6299 5864 6333
rect 5812 6296 5864 6299
rect 4982 6076 5034 6084
rect 4982 6042 4990 6076
rect 4990 6042 5024 6076
rect 5024 6042 5034 6076
rect 4982 6032 5034 6042
rect 4480 6000 4532 6006
rect 4480 5966 4490 6000
rect 4490 5966 4524 6000
rect 4524 5966 4532 6000
rect 4480 5954 4532 5966
rect 4808 5899 4860 5951
rect 4984 5899 5036 5951
rect 4046 5715 4098 5718
rect 4046 5681 4055 5715
rect 4055 5681 4089 5715
rect 4089 5681 4098 5715
rect 4046 5666 4098 5681
rect 3958 5592 4010 5602
rect 3958 5558 3969 5592
rect 3969 5558 4003 5592
rect 4003 5558 4010 5592
rect 3958 5550 4010 5558
rect 4862 5710 4914 5716
rect 4862 5676 4873 5710
rect 4873 5676 4907 5710
rect 4907 5676 4914 5710
rect 4862 5664 4914 5676
rect 4498 5529 4506 5534
rect 4506 5529 4540 5534
rect 4540 5529 4550 5534
rect 4498 5482 4550 5529
rect 4770 5594 4822 5604
rect 4770 5560 4782 5594
rect 4782 5560 4816 5594
rect 4816 5560 4822 5594
rect 4770 5552 4822 5560
rect 6600 6425 6620 6456
rect 6620 6425 6652 6456
rect 6600 6404 6652 6425
rect 8258 7056 8310 7062
rect 8258 7022 8268 7056
rect 8268 7022 8302 7056
rect 8302 7022 8310 7056
rect 8258 7010 8310 7022
rect 8571 6890 8623 6900
rect 8571 6856 8580 6890
rect 8580 6856 8614 6890
rect 8614 6856 8623 6890
rect 8571 6848 8623 6856
rect 8803 6885 8855 6890
rect 8803 6851 8823 6885
rect 8823 6851 8855 6885
rect 8803 6838 8855 6851
rect 9826 6862 9878 6868
rect 9826 6828 9836 6862
rect 9836 6828 9870 6862
rect 9870 6828 9878 6862
rect 9826 6816 9878 6828
rect 8276 6585 8284 6590
rect 8284 6585 8318 6590
rect 8318 6585 8328 6590
rect 8276 6538 8328 6585
rect 8939 6596 8991 6648
rect 9243 6648 9295 6652
rect 9243 6614 9255 6648
rect 9255 6614 9289 6648
rect 9289 6614 9295 6648
rect 9243 6600 9295 6614
rect 7938 6425 7950 6436
rect 7950 6425 7984 6436
rect 7984 6425 7990 6436
rect 7938 6384 7990 6425
rect 6496 6193 6548 6200
rect 6496 6159 6506 6193
rect 6506 6159 6540 6193
rect 6540 6159 6548 6193
rect 6496 6148 6548 6159
rect 6846 6341 6898 6342
rect 6846 6307 6877 6341
rect 6877 6307 6898 6341
rect 6846 6290 6898 6307
rect 7700 6333 7752 6348
rect 7700 6299 7719 6333
rect 7719 6299 7752 6333
rect 7700 6296 7752 6299
rect 6870 6076 6922 6084
rect 6870 6042 6878 6076
rect 6878 6042 6912 6076
rect 6912 6042 6922 6076
rect 6870 6032 6922 6042
rect 6368 6000 6420 6006
rect 6368 5966 6378 6000
rect 6378 5966 6412 6000
rect 6412 5966 6420 6000
rect 6368 5954 6420 5966
rect 6696 5899 6748 5951
rect 6872 5899 6924 5951
rect 5934 5715 5986 5718
rect 5934 5681 5943 5715
rect 5943 5681 5977 5715
rect 5977 5681 5986 5715
rect 5934 5666 5986 5681
rect 5846 5592 5898 5602
rect 5846 5558 5857 5592
rect 5857 5558 5891 5592
rect 5891 5558 5898 5592
rect 5846 5550 5898 5558
rect 6750 5710 6802 5716
rect 6750 5676 6761 5710
rect 6761 5676 6795 5710
rect 6795 5676 6802 5710
rect 6750 5664 6802 5676
rect 6386 5529 6394 5534
rect 6394 5529 6428 5534
rect 6428 5529 6438 5534
rect 6386 5482 6438 5529
rect 6658 5594 6710 5604
rect 6658 5560 6670 5594
rect 6670 5560 6704 5594
rect 6704 5560 6710 5594
rect 6658 5552 6710 5560
rect 8488 6425 8508 6456
rect 8508 6425 8540 6456
rect 8488 6404 8540 6425
rect 10146 7056 10198 7062
rect 10146 7022 10156 7056
rect 10156 7022 10190 7056
rect 10190 7022 10198 7056
rect 10146 7010 10198 7022
rect 10459 6890 10511 6900
rect 10459 6856 10468 6890
rect 10468 6856 10502 6890
rect 10502 6856 10511 6890
rect 10459 6848 10511 6856
rect 10691 6885 10743 6890
rect 10691 6851 10711 6885
rect 10711 6851 10743 6885
rect 10691 6838 10743 6851
rect 11714 6862 11766 6868
rect 11714 6828 11724 6862
rect 11724 6828 11758 6862
rect 11758 6828 11766 6862
rect 11714 6816 11766 6828
rect 10164 6585 10172 6590
rect 10172 6585 10206 6590
rect 10206 6585 10216 6590
rect 10164 6538 10216 6585
rect 10827 6596 10879 6648
rect 11131 6648 11183 6652
rect 11131 6614 11143 6648
rect 11143 6614 11177 6648
rect 11177 6614 11183 6648
rect 11131 6600 11183 6614
rect 9826 6425 9838 6436
rect 9838 6425 9872 6436
rect 9872 6425 9878 6436
rect 9826 6384 9878 6425
rect 8384 6193 8436 6200
rect 8384 6159 8394 6193
rect 8394 6159 8428 6193
rect 8428 6159 8436 6193
rect 8384 6148 8436 6159
rect 8734 6341 8786 6342
rect 8734 6307 8765 6341
rect 8765 6307 8786 6341
rect 8734 6290 8786 6307
rect 9588 6333 9640 6348
rect 9588 6299 9607 6333
rect 9607 6299 9640 6333
rect 9588 6296 9640 6299
rect 8758 6076 8810 6084
rect 8758 6042 8766 6076
rect 8766 6042 8800 6076
rect 8800 6042 8810 6076
rect 8758 6032 8810 6042
rect 8256 6000 8308 6006
rect 8256 5966 8266 6000
rect 8266 5966 8300 6000
rect 8300 5966 8308 6000
rect 8256 5954 8308 5966
rect 8584 5899 8636 5951
rect 8760 5899 8812 5951
rect 7822 5715 7874 5718
rect 7822 5681 7831 5715
rect 7831 5681 7865 5715
rect 7865 5681 7874 5715
rect 7822 5666 7874 5681
rect 7734 5592 7786 5602
rect 7734 5558 7745 5592
rect 7745 5558 7779 5592
rect 7779 5558 7786 5592
rect 7734 5550 7786 5558
rect 8638 5710 8690 5716
rect 8638 5676 8649 5710
rect 8649 5676 8683 5710
rect 8683 5676 8690 5710
rect 8638 5664 8690 5676
rect 8274 5529 8282 5534
rect 8282 5529 8316 5534
rect 8316 5529 8326 5534
rect 8274 5482 8326 5529
rect 8546 5594 8598 5604
rect 8546 5560 8558 5594
rect 8558 5560 8592 5594
rect 8592 5560 8598 5594
rect 8546 5552 8598 5560
rect 10376 6425 10396 6456
rect 10396 6425 10428 6456
rect 10376 6404 10428 6425
rect 12034 7056 12086 7062
rect 12034 7022 12044 7056
rect 12044 7022 12078 7056
rect 12078 7022 12086 7056
rect 12034 7010 12086 7022
rect 12347 6890 12399 6900
rect 12347 6856 12356 6890
rect 12356 6856 12390 6890
rect 12390 6856 12399 6890
rect 12347 6848 12399 6856
rect 12579 6885 12631 6890
rect 12579 6851 12599 6885
rect 12599 6851 12631 6885
rect 12579 6838 12631 6851
rect 13602 6862 13654 6868
rect 13602 6828 13612 6862
rect 13612 6828 13646 6862
rect 13646 6828 13654 6862
rect 13602 6816 13654 6828
rect 12052 6585 12060 6590
rect 12060 6585 12094 6590
rect 12094 6585 12104 6590
rect 12052 6538 12104 6585
rect 12715 6596 12767 6648
rect 13019 6648 13071 6652
rect 13019 6614 13031 6648
rect 13031 6614 13065 6648
rect 13065 6614 13071 6648
rect 13019 6600 13071 6614
rect 11714 6425 11726 6436
rect 11726 6425 11760 6436
rect 11760 6425 11766 6436
rect 11714 6384 11766 6425
rect 10272 6193 10324 6200
rect 10272 6159 10282 6193
rect 10282 6159 10316 6193
rect 10316 6159 10324 6193
rect 10272 6148 10324 6159
rect 10622 6341 10674 6342
rect 10622 6307 10653 6341
rect 10653 6307 10674 6341
rect 10622 6290 10674 6307
rect 11476 6333 11528 6348
rect 11476 6299 11495 6333
rect 11495 6299 11528 6333
rect 11476 6296 11528 6299
rect 10646 6076 10698 6084
rect 10646 6042 10654 6076
rect 10654 6042 10688 6076
rect 10688 6042 10698 6076
rect 10646 6032 10698 6042
rect 10144 6000 10196 6006
rect 10144 5966 10154 6000
rect 10154 5966 10188 6000
rect 10188 5966 10196 6000
rect 10144 5954 10196 5966
rect 10472 5899 10524 5951
rect 10648 5899 10700 5951
rect 9710 5715 9762 5718
rect 9710 5681 9719 5715
rect 9719 5681 9753 5715
rect 9753 5681 9762 5715
rect 9710 5666 9762 5681
rect 9622 5592 9674 5602
rect 9622 5558 9633 5592
rect 9633 5558 9667 5592
rect 9667 5558 9674 5592
rect 9622 5550 9674 5558
rect 10526 5710 10578 5716
rect 10526 5676 10537 5710
rect 10537 5676 10571 5710
rect 10571 5676 10578 5710
rect 10526 5664 10578 5676
rect 10162 5529 10170 5534
rect 10170 5529 10204 5534
rect 10204 5529 10214 5534
rect 10162 5482 10214 5529
rect 10434 5594 10486 5604
rect 10434 5560 10446 5594
rect 10446 5560 10480 5594
rect 10480 5560 10486 5594
rect 10434 5552 10486 5560
rect 12264 6425 12284 6456
rect 12284 6425 12316 6456
rect 12264 6404 12316 6425
rect 13922 7056 13974 7062
rect 13922 7022 13932 7056
rect 13932 7022 13966 7056
rect 13966 7022 13974 7056
rect 13922 7010 13974 7022
rect 14235 6890 14287 6900
rect 14235 6856 14244 6890
rect 14244 6856 14278 6890
rect 14278 6856 14287 6890
rect 14235 6848 14287 6856
rect 14467 6885 14519 6890
rect 14467 6851 14487 6885
rect 14487 6851 14519 6885
rect 14467 6838 14519 6851
rect 15484 6862 15536 6868
rect 15484 6828 15494 6862
rect 15494 6828 15528 6862
rect 15528 6828 15536 6862
rect 15484 6816 15536 6828
rect 13940 6585 13948 6590
rect 13948 6585 13982 6590
rect 13982 6585 13992 6590
rect 13940 6538 13992 6585
rect 14603 6596 14655 6648
rect 14901 6648 14953 6652
rect 14901 6614 14913 6648
rect 14913 6614 14947 6648
rect 14947 6614 14953 6648
rect 14901 6600 14953 6614
rect 13602 6425 13614 6436
rect 13614 6425 13648 6436
rect 13648 6425 13654 6436
rect 13602 6384 13654 6425
rect 12160 6193 12212 6200
rect 12160 6159 12170 6193
rect 12170 6159 12204 6193
rect 12204 6159 12212 6193
rect 12160 6148 12212 6159
rect 12510 6341 12562 6342
rect 12510 6307 12541 6341
rect 12541 6307 12562 6341
rect 12510 6290 12562 6307
rect 13364 6333 13416 6348
rect 13364 6299 13383 6333
rect 13383 6299 13416 6333
rect 13364 6296 13416 6299
rect 12534 6076 12586 6084
rect 12534 6042 12542 6076
rect 12542 6042 12576 6076
rect 12576 6042 12586 6076
rect 12534 6032 12586 6042
rect 12032 6000 12084 6006
rect 12032 5966 12042 6000
rect 12042 5966 12076 6000
rect 12076 5966 12084 6000
rect 12032 5954 12084 5966
rect 12360 5899 12412 5951
rect 12536 5899 12588 5951
rect 11598 5715 11650 5718
rect 11598 5681 11607 5715
rect 11607 5681 11641 5715
rect 11641 5681 11650 5715
rect 11598 5666 11650 5681
rect 11510 5592 11562 5602
rect 11510 5558 11521 5592
rect 11521 5558 11555 5592
rect 11555 5558 11562 5592
rect 11510 5550 11562 5558
rect 12414 5710 12466 5716
rect 12414 5676 12425 5710
rect 12425 5676 12459 5710
rect 12459 5676 12466 5710
rect 12414 5664 12466 5676
rect 12050 5529 12058 5534
rect 12058 5529 12092 5534
rect 12092 5529 12102 5534
rect 12050 5482 12102 5529
rect 12322 5594 12374 5604
rect 12322 5560 12334 5594
rect 12334 5560 12368 5594
rect 12368 5560 12374 5594
rect 12322 5552 12374 5560
rect 14152 6425 14172 6456
rect 14172 6425 14204 6456
rect 14152 6404 14204 6425
rect 15804 7056 15856 7062
rect 15804 7022 15814 7056
rect 15814 7022 15848 7056
rect 15848 7022 15856 7056
rect 15804 7010 15856 7022
rect 16117 6890 16169 6900
rect 16117 6856 16126 6890
rect 16126 6856 16160 6890
rect 16160 6856 16169 6890
rect 16117 6848 16169 6856
rect 16349 6885 16401 6890
rect 16349 6851 16369 6885
rect 16369 6851 16401 6885
rect 16349 6838 16401 6851
rect 17372 6862 17424 6868
rect 17372 6828 17382 6862
rect 17382 6828 17416 6862
rect 17416 6828 17424 6862
rect 17372 6816 17424 6828
rect 15822 6585 15830 6590
rect 15830 6585 15864 6590
rect 15864 6585 15874 6590
rect 15822 6538 15874 6585
rect 16485 6596 16537 6648
rect 16789 6648 16841 6652
rect 16789 6614 16801 6648
rect 16801 6614 16835 6648
rect 16835 6614 16841 6648
rect 16789 6600 16841 6614
rect 15484 6425 15496 6436
rect 15496 6425 15530 6436
rect 15530 6425 15536 6436
rect 15484 6384 15536 6425
rect 14048 6193 14100 6200
rect 14048 6159 14058 6193
rect 14058 6159 14092 6193
rect 14092 6159 14100 6193
rect 14048 6148 14100 6159
rect 14398 6341 14450 6342
rect 14398 6307 14429 6341
rect 14429 6307 14450 6341
rect 14398 6290 14450 6307
rect 15246 6333 15298 6348
rect 15246 6299 15265 6333
rect 15265 6299 15298 6333
rect 15246 6296 15298 6299
rect 14422 6076 14474 6084
rect 14422 6042 14430 6076
rect 14430 6042 14464 6076
rect 14464 6042 14474 6076
rect 14422 6032 14474 6042
rect 13920 6000 13972 6006
rect 13920 5966 13930 6000
rect 13930 5966 13964 6000
rect 13964 5966 13972 6000
rect 13920 5954 13972 5966
rect 14248 5899 14300 5951
rect 14424 5899 14476 5951
rect 13486 5715 13538 5718
rect 13486 5681 13495 5715
rect 13495 5681 13529 5715
rect 13529 5681 13538 5715
rect 13486 5666 13538 5681
rect 13398 5592 13450 5602
rect 13398 5558 13409 5592
rect 13409 5558 13443 5592
rect 13443 5558 13450 5592
rect 13398 5550 13450 5558
rect 14302 5710 14354 5716
rect 14302 5676 14313 5710
rect 14313 5676 14347 5710
rect 14347 5676 14354 5710
rect 14302 5664 14354 5676
rect 13938 5529 13946 5534
rect 13946 5529 13980 5534
rect 13980 5529 13990 5534
rect 13938 5482 13990 5529
rect 14210 5594 14262 5604
rect 14210 5560 14222 5594
rect 14222 5560 14256 5594
rect 14256 5560 14262 5594
rect 14210 5552 14262 5560
rect 16034 6425 16054 6456
rect 16054 6425 16086 6456
rect 16034 6404 16086 6425
rect 17692 7056 17744 7062
rect 17692 7022 17702 7056
rect 17702 7022 17736 7056
rect 17736 7022 17744 7056
rect 17692 7010 17744 7022
rect 18005 6890 18057 6900
rect 18005 6856 18014 6890
rect 18014 6856 18048 6890
rect 18048 6856 18057 6890
rect 18005 6848 18057 6856
rect 18237 6885 18289 6890
rect 18237 6851 18257 6885
rect 18257 6851 18289 6885
rect 18237 6838 18289 6851
rect 19260 6862 19312 6868
rect 19260 6828 19270 6862
rect 19270 6828 19304 6862
rect 19304 6828 19312 6862
rect 19260 6816 19312 6828
rect 17710 6585 17718 6590
rect 17718 6585 17752 6590
rect 17752 6585 17762 6590
rect 17710 6538 17762 6585
rect 18373 6596 18425 6648
rect 18677 6648 18729 6652
rect 18677 6614 18689 6648
rect 18689 6614 18723 6648
rect 18723 6614 18729 6648
rect 18677 6600 18729 6614
rect 17372 6425 17384 6436
rect 17384 6425 17418 6436
rect 17418 6425 17424 6436
rect 17372 6384 17424 6425
rect 15930 6193 15982 6200
rect 15930 6159 15940 6193
rect 15940 6159 15974 6193
rect 15974 6159 15982 6193
rect 15930 6148 15982 6159
rect 16280 6341 16332 6342
rect 16280 6307 16311 6341
rect 16311 6307 16332 6341
rect 16280 6290 16332 6307
rect 17134 6333 17186 6348
rect 17134 6299 17153 6333
rect 17153 6299 17186 6333
rect 17134 6296 17186 6299
rect 16304 6076 16356 6084
rect 16304 6042 16312 6076
rect 16312 6042 16346 6076
rect 16346 6042 16356 6076
rect 16304 6032 16356 6042
rect 15802 6000 15854 6006
rect 15802 5966 15812 6000
rect 15812 5966 15846 6000
rect 15846 5966 15854 6000
rect 15802 5954 15854 5966
rect 16130 5899 16182 5951
rect 16306 5899 16358 5951
rect 15368 5715 15420 5718
rect 15368 5681 15377 5715
rect 15377 5681 15411 5715
rect 15411 5681 15420 5715
rect 15368 5666 15420 5681
rect 15280 5592 15332 5602
rect 15280 5558 15291 5592
rect 15291 5558 15325 5592
rect 15325 5558 15332 5592
rect 15280 5550 15332 5558
rect 16184 5710 16236 5716
rect 16184 5676 16195 5710
rect 16195 5676 16229 5710
rect 16229 5676 16236 5710
rect 16184 5664 16236 5676
rect 15820 5529 15828 5534
rect 15828 5529 15862 5534
rect 15862 5529 15872 5534
rect 15820 5482 15872 5529
rect 16092 5594 16144 5604
rect 16092 5560 16104 5594
rect 16104 5560 16138 5594
rect 16138 5560 16144 5594
rect 16092 5552 16144 5560
rect 17922 6425 17942 6456
rect 17942 6425 17974 6456
rect 17922 6404 17974 6425
rect 19580 7056 19632 7062
rect 19580 7022 19590 7056
rect 19590 7022 19624 7056
rect 19624 7022 19632 7056
rect 19580 7010 19632 7022
rect 19893 6890 19945 6900
rect 19893 6856 19902 6890
rect 19902 6856 19936 6890
rect 19936 6856 19945 6890
rect 19893 6848 19945 6856
rect 20125 6885 20177 6890
rect 20125 6851 20145 6885
rect 20145 6851 20177 6885
rect 20125 6838 20177 6851
rect 21148 6862 21200 6868
rect 21148 6828 21158 6862
rect 21158 6828 21192 6862
rect 21192 6828 21200 6862
rect 21148 6816 21200 6828
rect 19598 6585 19606 6590
rect 19606 6585 19640 6590
rect 19640 6585 19650 6590
rect 19598 6538 19650 6585
rect 20261 6596 20313 6648
rect 20565 6648 20617 6652
rect 20565 6614 20577 6648
rect 20577 6614 20611 6648
rect 20611 6614 20617 6648
rect 20565 6600 20617 6614
rect 19260 6425 19272 6436
rect 19272 6425 19306 6436
rect 19306 6425 19312 6436
rect 19260 6384 19312 6425
rect 17818 6193 17870 6200
rect 17818 6159 17828 6193
rect 17828 6159 17862 6193
rect 17862 6159 17870 6193
rect 17818 6148 17870 6159
rect 18168 6341 18220 6342
rect 18168 6307 18199 6341
rect 18199 6307 18220 6341
rect 18168 6290 18220 6307
rect 19022 6333 19074 6348
rect 19022 6299 19041 6333
rect 19041 6299 19074 6333
rect 19022 6296 19074 6299
rect 18192 6076 18244 6084
rect 18192 6042 18200 6076
rect 18200 6042 18234 6076
rect 18234 6042 18244 6076
rect 18192 6032 18244 6042
rect 17690 6000 17742 6006
rect 17690 5966 17700 6000
rect 17700 5966 17734 6000
rect 17734 5966 17742 6000
rect 17690 5954 17742 5966
rect 18018 5899 18070 5951
rect 18194 5899 18246 5951
rect 17256 5715 17308 5718
rect 17256 5681 17265 5715
rect 17265 5681 17299 5715
rect 17299 5681 17308 5715
rect 17256 5666 17308 5681
rect 17168 5592 17220 5602
rect 17168 5558 17179 5592
rect 17179 5558 17213 5592
rect 17213 5558 17220 5592
rect 17168 5550 17220 5558
rect 18072 5710 18124 5716
rect 18072 5676 18083 5710
rect 18083 5676 18117 5710
rect 18117 5676 18124 5710
rect 18072 5664 18124 5676
rect 17708 5529 17716 5534
rect 17716 5529 17750 5534
rect 17750 5529 17760 5534
rect 17708 5482 17760 5529
rect 17980 5594 18032 5604
rect 17980 5560 17992 5594
rect 17992 5560 18026 5594
rect 18026 5560 18032 5594
rect 17980 5552 18032 5560
rect 19810 6425 19830 6456
rect 19830 6425 19862 6456
rect 19810 6404 19862 6425
rect 21468 7056 21520 7062
rect 21468 7022 21478 7056
rect 21478 7022 21512 7056
rect 21512 7022 21520 7056
rect 21468 7010 21520 7022
rect 21781 6890 21833 6900
rect 21781 6856 21790 6890
rect 21790 6856 21824 6890
rect 21824 6856 21833 6890
rect 21781 6848 21833 6856
rect 22013 6885 22065 6890
rect 22013 6851 22033 6885
rect 22033 6851 22065 6885
rect 22013 6838 22065 6851
rect 23036 6862 23088 6868
rect 23036 6828 23046 6862
rect 23046 6828 23080 6862
rect 23080 6828 23088 6862
rect 23036 6816 23088 6828
rect 21486 6585 21494 6590
rect 21494 6585 21528 6590
rect 21528 6585 21538 6590
rect 21486 6538 21538 6585
rect 22149 6596 22201 6648
rect 22453 6648 22505 6652
rect 22453 6614 22465 6648
rect 22465 6614 22499 6648
rect 22499 6614 22505 6648
rect 22453 6600 22505 6614
rect 21148 6425 21160 6436
rect 21160 6425 21194 6436
rect 21194 6425 21200 6436
rect 21148 6384 21200 6425
rect 19706 6193 19758 6200
rect 19706 6159 19716 6193
rect 19716 6159 19750 6193
rect 19750 6159 19758 6193
rect 19706 6148 19758 6159
rect 20056 6341 20108 6342
rect 20056 6307 20087 6341
rect 20087 6307 20108 6341
rect 20056 6290 20108 6307
rect 20910 6333 20962 6348
rect 20910 6299 20929 6333
rect 20929 6299 20962 6333
rect 20910 6296 20962 6299
rect 20080 6076 20132 6084
rect 20080 6042 20088 6076
rect 20088 6042 20122 6076
rect 20122 6042 20132 6076
rect 20080 6032 20132 6042
rect 19578 6000 19630 6006
rect 19578 5966 19588 6000
rect 19588 5966 19622 6000
rect 19622 5966 19630 6000
rect 19578 5954 19630 5966
rect 19906 5899 19958 5951
rect 20082 5899 20134 5951
rect 19144 5715 19196 5718
rect 19144 5681 19153 5715
rect 19153 5681 19187 5715
rect 19187 5681 19196 5715
rect 19144 5666 19196 5681
rect 19056 5592 19108 5602
rect 19056 5558 19067 5592
rect 19067 5558 19101 5592
rect 19101 5558 19108 5592
rect 19056 5550 19108 5558
rect 19960 5710 20012 5716
rect 19960 5676 19971 5710
rect 19971 5676 20005 5710
rect 20005 5676 20012 5710
rect 19960 5664 20012 5676
rect 19596 5529 19604 5534
rect 19604 5529 19638 5534
rect 19638 5529 19648 5534
rect 19596 5482 19648 5529
rect 19868 5594 19920 5604
rect 19868 5560 19880 5594
rect 19880 5560 19914 5594
rect 19914 5560 19920 5594
rect 19868 5552 19920 5560
rect 21698 6425 21718 6456
rect 21718 6425 21750 6456
rect 21698 6404 21750 6425
rect 23356 7056 23408 7062
rect 23356 7022 23366 7056
rect 23366 7022 23400 7056
rect 23400 7022 23408 7056
rect 23356 7010 23408 7022
rect 23669 6890 23721 6900
rect 23669 6856 23678 6890
rect 23678 6856 23712 6890
rect 23712 6856 23721 6890
rect 23669 6848 23721 6856
rect 23901 6885 23953 6890
rect 23901 6851 23921 6885
rect 23921 6851 23953 6885
rect 23901 6838 23953 6851
rect 24924 6862 24976 6868
rect 24924 6828 24934 6862
rect 24934 6828 24968 6862
rect 24968 6828 24976 6862
rect 24924 6816 24976 6828
rect 23374 6585 23382 6590
rect 23382 6585 23416 6590
rect 23416 6585 23426 6590
rect 23374 6538 23426 6585
rect 24037 6596 24089 6648
rect 24341 6648 24393 6652
rect 24341 6614 24353 6648
rect 24353 6614 24387 6648
rect 24387 6614 24393 6648
rect 24341 6600 24393 6614
rect 23036 6425 23048 6436
rect 23048 6425 23082 6436
rect 23082 6425 23088 6436
rect 23036 6384 23088 6425
rect 21594 6193 21646 6200
rect 21594 6159 21604 6193
rect 21604 6159 21638 6193
rect 21638 6159 21646 6193
rect 21594 6148 21646 6159
rect 21944 6341 21996 6342
rect 21944 6307 21975 6341
rect 21975 6307 21996 6341
rect 21944 6290 21996 6307
rect 22798 6333 22850 6348
rect 22798 6299 22817 6333
rect 22817 6299 22850 6333
rect 22798 6296 22850 6299
rect 21968 6076 22020 6084
rect 21968 6042 21976 6076
rect 21976 6042 22010 6076
rect 22010 6042 22020 6076
rect 21968 6032 22020 6042
rect 21466 6000 21518 6006
rect 21466 5966 21476 6000
rect 21476 5966 21510 6000
rect 21510 5966 21518 6000
rect 21466 5954 21518 5966
rect 21794 5899 21846 5951
rect 21970 5899 22022 5951
rect 21032 5715 21084 5718
rect 21032 5681 21041 5715
rect 21041 5681 21075 5715
rect 21075 5681 21084 5715
rect 21032 5666 21084 5681
rect 20944 5592 20996 5602
rect 20944 5558 20955 5592
rect 20955 5558 20989 5592
rect 20989 5558 20996 5592
rect 20944 5550 20996 5558
rect 21848 5710 21900 5716
rect 21848 5676 21859 5710
rect 21859 5676 21893 5710
rect 21893 5676 21900 5710
rect 21848 5664 21900 5676
rect 21484 5529 21492 5534
rect 21492 5529 21526 5534
rect 21526 5529 21536 5534
rect 21484 5482 21536 5529
rect 21756 5594 21808 5604
rect 21756 5560 21768 5594
rect 21768 5560 21802 5594
rect 21802 5560 21808 5594
rect 21756 5552 21808 5560
rect 23586 6425 23606 6456
rect 23606 6425 23638 6456
rect 23586 6404 23638 6425
rect 25244 7056 25296 7062
rect 25244 7022 25254 7056
rect 25254 7022 25288 7056
rect 25288 7022 25296 7056
rect 25244 7010 25296 7022
rect 25557 6890 25609 6900
rect 25557 6856 25566 6890
rect 25566 6856 25600 6890
rect 25600 6856 25609 6890
rect 25557 6848 25609 6856
rect 25789 6885 25841 6890
rect 25789 6851 25809 6885
rect 25809 6851 25841 6885
rect 25789 6838 25841 6851
rect 26812 6862 26864 6868
rect 26812 6828 26822 6862
rect 26822 6828 26856 6862
rect 26856 6828 26864 6862
rect 26812 6816 26864 6828
rect 25262 6585 25270 6590
rect 25270 6585 25304 6590
rect 25304 6585 25314 6590
rect 25262 6538 25314 6585
rect 25925 6596 25977 6648
rect 26229 6648 26281 6652
rect 26229 6614 26241 6648
rect 26241 6614 26275 6648
rect 26275 6614 26281 6648
rect 26229 6600 26281 6614
rect 24924 6425 24936 6436
rect 24936 6425 24970 6436
rect 24970 6425 24976 6436
rect 24924 6384 24976 6425
rect 23482 6193 23534 6200
rect 23482 6159 23492 6193
rect 23492 6159 23526 6193
rect 23526 6159 23534 6193
rect 23482 6148 23534 6159
rect 23832 6341 23884 6342
rect 23832 6307 23863 6341
rect 23863 6307 23884 6341
rect 23832 6290 23884 6307
rect 24686 6333 24738 6348
rect 24686 6299 24705 6333
rect 24705 6299 24738 6333
rect 24686 6296 24738 6299
rect 23856 6076 23908 6084
rect 23856 6042 23864 6076
rect 23864 6042 23898 6076
rect 23898 6042 23908 6076
rect 23856 6032 23908 6042
rect 23354 6000 23406 6006
rect 23354 5966 23364 6000
rect 23364 5966 23398 6000
rect 23398 5966 23406 6000
rect 23354 5954 23406 5966
rect 23682 5899 23734 5951
rect 23858 5899 23910 5951
rect 22920 5715 22972 5718
rect 22920 5681 22929 5715
rect 22929 5681 22963 5715
rect 22963 5681 22972 5715
rect 22920 5666 22972 5681
rect 22832 5592 22884 5602
rect 22832 5558 22843 5592
rect 22843 5558 22877 5592
rect 22877 5558 22884 5592
rect 22832 5550 22884 5558
rect 23736 5710 23788 5716
rect 23736 5676 23747 5710
rect 23747 5676 23781 5710
rect 23781 5676 23788 5710
rect 23736 5664 23788 5676
rect 23372 5529 23380 5534
rect 23380 5529 23414 5534
rect 23414 5529 23424 5534
rect 23372 5482 23424 5529
rect 23644 5594 23696 5604
rect 23644 5560 23656 5594
rect 23656 5560 23690 5594
rect 23690 5560 23696 5594
rect 23644 5552 23696 5560
rect 25474 6425 25494 6456
rect 25494 6425 25526 6456
rect 25474 6404 25526 6425
rect 27132 7056 27184 7062
rect 27132 7022 27142 7056
rect 27142 7022 27176 7056
rect 27176 7022 27184 7056
rect 27132 7010 27184 7022
rect 27445 6890 27497 6900
rect 27445 6856 27454 6890
rect 27454 6856 27488 6890
rect 27488 6856 27497 6890
rect 27445 6848 27497 6856
rect 27677 6885 27729 6890
rect 27677 6851 27697 6885
rect 27697 6851 27729 6885
rect 27677 6838 27729 6851
rect 28700 6862 28752 6868
rect 28700 6828 28710 6862
rect 28710 6828 28744 6862
rect 28744 6828 28752 6862
rect 28700 6816 28752 6828
rect 27150 6585 27158 6590
rect 27158 6585 27192 6590
rect 27192 6585 27202 6590
rect 27150 6538 27202 6585
rect 27813 6596 27865 6648
rect 28117 6648 28169 6652
rect 28117 6614 28129 6648
rect 28129 6614 28163 6648
rect 28163 6614 28169 6648
rect 28117 6600 28169 6614
rect 26812 6425 26824 6436
rect 26824 6425 26858 6436
rect 26858 6425 26864 6436
rect 26812 6384 26864 6425
rect 25370 6193 25422 6200
rect 25370 6159 25380 6193
rect 25380 6159 25414 6193
rect 25414 6159 25422 6193
rect 25370 6148 25422 6159
rect 25720 6341 25772 6342
rect 25720 6307 25751 6341
rect 25751 6307 25772 6341
rect 25720 6290 25772 6307
rect 26574 6333 26626 6348
rect 26574 6299 26593 6333
rect 26593 6299 26626 6333
rect 26574 6296 26626 6299
rect 25744 6076 25796 6084
rect 25744 6042 25752 6076
rect 25752 6042 25786 6076
rect 25786 6042 25796 6076
rect 25744 6032 25796 6042
rect 25242 6000 25294 6006
rect 25242 5966 25252 6000
rect 25252 5966 25286 6000
rect 25286 5966 25294 6000
rect 25242 5954 25294 5966
rect 25570 5899 25622 5951
rect 25746 5899 25798 5951
rect 24808 5715 24860 5718
rect 24808 5681 24817 5715
rect 24817 5681 24851 5715
rect 24851 5681 24860 5715
rect 24808 5666 24860 5681
rect 24720 5592 24772 5602
rect 24720 5558 24731 5592
rect 24731 5558 24765 5592
rect 24765 5558 24772 5592
rect 24720 5550 24772 5558
rect 25624 5710 25676 5716
rect 25624 5676 25635 5710
rect 25635 5676 25669 5710
rect 25669 5676 25676 5710
rect 25624 5664 25676 5676
rect 25260 5529 25268 5534
rect 25268 5529 25302 5534
rect 25302 5529 25312 5534
rect 25260 5482 25312 5529
rect 25532 5594 25584 5604
rect 25532 5560 25544 5594
rect 25544 5560 25578 5594
rect 25578 5560 25584 5594
rect 25532 5552 25584 5560
rect 27362 6425 27382 6456
rect 27382 6425 27414 6456
rect 27362 6404 27414 6425
rect 29020 7056 29072 7062
rect 29020 7022 29030 7056
rect 29030 7022 29064 7056
rect 29064 7022 29072 7056
rect 29020 7010 29072 7022
rect 29333 6890 29385 6900
rect 29333 6856 29342 6890
rect 29342 6856 29376 6890
rect 29376 6856 29385 6890
rect 29333 6848 29385 6856
rect 29565 6885 29617 6890
rect 29565 6851 29585 6885
rect 29585 6851 29617 6885
rect 29565 6838 29617 6851
rect 30588 6862 30640 6868
rect 30588 6828 30598 6862
rect 30598 6828 30632 6862
rect 30632 6828 30640 6862
rect 30588 6816 30640 6828
rect 29038 6585 29046 6590
rect 29046 6585 29080 6590
rect 29080 6585 29090 6590
rect 29038 6538 29090 6585
rect 29701 6596 29753 6648
rect 30005 6648 30057 6652
rect 30005 6614 30017 6648
rect 30017 6614 30051 6648
rect 30051 6614 30057 6648
rect 30005 6600 30057 6614
rect 28700 6425 28712 6436
rect 28712 6425 28746 6436
rect 28746 6425 28752 6436
rect 28700 6384 28752 6425
rect 27258 6193 27310 6200
rect 27258 6159 27268 6193
rect 27268 6159 27302 6193
rect 27302 6159 27310 6193
rect 27258 6148 27310 6159
rect 27608 6341 27660 6342
rect 27608 6307 27639 6341
rect 27639 6307 27660 6341
rect 27608 6290 27660 6307
rect 28462 6333 28514 6348
rect 28462 6299 28481 6333
rect 28481 6299 28514 6333
rect 28462 6296 28514 6299
rect 27632 6076 27684 6084
rect 27632 6042 27640 6076
rect 27640 6042 27674 6076
rect 27674 6042 27684 6076
rect 27632 6032 27684 6042
rect 27130 6000 27182 6006
rect 27130 5966 27140 6000
rect 27140 5966 27174 6000
rect 27174 5966 27182 6000
rect 27130 5954 27182 5966
rect 27458 5899 27510 5951
rect 27634 5899 27686 5951
rect 26696 5715 26748 5718
rect 26696 5681 26705 5715
rect 26705 5681 26739 5715
rect 26739 5681 26748 5715
rect 26696 5666 26748 5681
rect 26608 5592 26660 5602
rect 26608 5558 26619 5592
rect 26619 5558 26653 5592
rect 26653 5558 26660 5592
rect 26608 5550 26660 5558
rect 27512 5710 27564 5716
rect 27512 5676 27523 5710
rect 27523 5676 27557 5710
rect 27557 5676 27564 5710
rect 27512 5664 27564 5676
rect 27148 5529 27156 5534
rect 27156 5529 27190 5534
rect 27190 5529 27200 5534
rect 27148 5482 27200 5529
rect 27420 5594 27472 5604
rect 27420 5560 27432 5594
rect 27432 5560 27466 5594
rect 27466 5560 27472 5594
rect 27420 5552 27472 5560
rect 29250 6425 29270 6456
rect 29270 6425 29302 6456
rect 29250 6404 29302 6425
rect 30908 7056 30960 7062
rect 30908 7022 30918 7056
rect 30918 7022 30952 7056
rect 30952 7022 30960 7056
rect 30908 7010 30960 7022
rect 31221 6890 31273 6900
rect 31221 6856 31230 6890
rect 31230 6856 31264 6890
rect 31264 6856 31273 6890
rect 31221 6848 31273 6856
rect 31453 6885 31505 6890
rect 31453 6851 31473 6885
rect 31473 6851 31505 6885
rect 31453 6838 31505 6851
rect 32476 6862 32528 6868
rect 32476 6828 32486 6862
rect 32486 6828 32520 6862
rect 32520 6828 32528 6862
rect 32476 6816 32528 6828
rect 30926 6585 30934 6590
rect 30934 6585 30968 6590
rect 30968 6585 30978 6590
rect 30926 6538 30978 6585
rect 31589 6596 31641 6648
rect 31893 6648 31945 6652
rect 31893 6614 31905 6648
rect 31905 6614 31939 6648
rect 31939 6614 31945 6648
rect 31893 6600 31945 6614
rect 30588 6425 30600 6436
rect 30600 6425 30634 6436
rect 30634 6425 30640 6436
rect 30588 6384 30640 6425
rect 29146 6193 29198 6200
rect 29146 6159 29156 6193
rect 29156 6159 29190 6193
rect 29190 6159 29198 6193
rect 29146 6148 29198 6159
rect 29496 6341 29548 6342
rect 29496 6307 29527 6341
rect 29527 6307 29548 6341
rect 29496 6290 29548 6307
rect 30350 6333 30402 6348
rect 30350 6299 30369 6333
rect 30369 6299 30402 6333
rect 30350 6296 30402 6299
rect 29520 6076 29572 6084
rect 29520 6042 29528 6076
rect 29528 6042 29562 6076
rect 29562 6042 29572 6076
rect 29520 6032 29572 6042
rect 29018 6000 29070 6006
rect 29018 5966 29028 6000
rect 29028 5966 29062 6000
rect 29062 5966 29070 6000
rect 29018 5954 29070 5966
rect 29346 5899 29398 5951
rect 29522 5899 29574 5951
rect 28584 5715 28636 5718
rect 28584 5681 28593 5715
rect 28593 5681 28627 5715
rect 28627 5681 28636 5715
rect 28584 5666 28636 5681
rect 28496 5592 28548 5602
rect 28496 5558 28507 5592
rect 28507 5558 28541 5592
rect 28541 5558 28548 5592
rect 28496 5550 28548 5558
rect 29400 5710 29452 5716
rect 29400 5676 29411 5710
rect 29411 5676 29445 5710
rect 29445 5676 29452 5710
rect 29400 5664 29452 5676
rect 29036 5529 29044 5534
rect 29044 5529 29078 5534
rect 29078 5529 29088 5534
rect 29036 5482 29088 5529
rect 29308 5594 29360 5604
rect 29308 5560 29320 5594
rect 29320 5560 29354 5594
rect 29354 5560 29360 5594
rect 29308 5552 29360 5560
rect 31138 6425 31158 6456
rect 31158 6425 31190 6456
rect 31138 6404 31190 6425
rect 32796 7056 32848 7062
rect 32796 7022 32806 7056
rect 32806 7022 32840 7056
rect 32840 7022 32848 7056
rect 32796 7010 32848 7022
rect 33109 6890 33161 6900
rect 33109 6856 33118 6890
rect 33118 6856 33152 6890
rect 33152 6856 33161 6890
rect 33109 6848 33161 6856
rect 33341 6885 33393 6890
rect 33341 6851 33361 6885
rect 33361 6851 33393 6885
rect 33341 6838 33393 6851
rect 34364 6862 34416 6868
rect 34364 6828 34374 6862
rect 34374 6828 34408 6862
rect 34408 6828 34416 6862
rect 34364 6816 34416 6828
rect 32814 6585 32822 6590
rect 32822 6585 32856 6590
rect 32856 6585 32866 6590
rect 32814 6538 32866 6585
rect 33477 6596 33529 6648
rect 33781 6648 33833 6652
rect 33781 6614 33793 6648
rect 33793 6614 33827 6648
rect 33827 6614 33833 6648
rect 33781 6600 33833 6614
rect 32476 6425 32488 6436
rect 32488 6425 32522 6436
rect 32522 6425 32528 6436
rect 32476 6384 32528 6425
rect 31034 6193 31086 6200
rect 31034 6159 31044 6193
rect 31044 6159 31078 6193
rect 31078 6159 31086 6193
rect 31034 6148 31086 6159
rect 31384 6341 31436 6342
rect 31384 6307 31415 6341
rect 31415 6307 31436 6341
rect 31384 6290 31436 6307
rect 32238 6333 32290 6348
rect 32238 6299 32257 6333
rect 32257 6299 32290 6333
rect 32238 6296 32290 6299
rect 31408 6076 31460 6084
rect 31408 6042 31416 6076
rect 31416 6042 31450 6076
rect 31450 6042 31460 6076
rect 31408 6032 31460 6042
rect 30906 6000 30958 6006
rect 30906 5966 30916 6000
rect 30916 5966 30950 6000
rect 30950 5966 30958 6000
rect 30906 5954 30958 5966
rect 31234 5899 31286 5951
rect 31410 5899 31462 5951
rect 30472 5715 30524 5718
rect 30472 5681 30481 5715
rect 30481 5681 30515 5715
rect 30515 5681 30524 5715
rect 30472 5666 30524 5681
rect 30384 5592 30436 5602
rect 30384 5558 30395 5592
rect 30395 5558 30429 5592
rect 30429 5558 30436 5592
rect 30384 5550 30436 5558
rect 31288 5710 31340 5716
rect 31288 5676 31299 5710
rect 31299 5676 31333 5710
rect 31333 5676 31340 5710
rect 31288 5664 31340 5676
rect 30924 5529 30932 5534
rect 30932 5529 30966 5534
rect 30966 5529 30976 5534
rect 30924 5482 30976 5529
rect 31196 5594 31248 5604
rect 31196 5560 31208 5594
rect 31208 5560 31242 5594
rect 31242 5560 31248 5594
rect 31196 5552 31248 5560
rect 33026 6425 33046 6456
rect 33046 6425 33078 6456
rect 33026 6404 33078 6425
rect 34684 7056 34736 7062
rect 34684 7022 34694 7056
rect 34694 7022 34728 7056
rect 34728 7022 34736 7056
rect 34684 7010 34736 7022
rect 34997 6890 35049 6900
rect 34997 6856 35006 6890
rect 35006 6856 35040 6890
rect 35040 6856 35049 6890
rect 34997 6848 35049 6856
rect 35229 6885 35281 6890
rect 35229 6851 35249 6885
rect 35249 6851 35281 6885
rect 35229 6838 35281 6851
rect 36252 6862 36304 6868
rect 36252 6828 36262 6862
rect 36262 6828 36296 6862
rect 36296 6828 36304 6862
rect 36252 6816 36304 6828
rect 34702 6585 34710 6590
rect 34710 6585 34744 6590
rect 34744 6585 34754 6590
rect 34702 6538 34754 6585
rect 35365 6596 35417 6648
rect 35669 6648 35721 6652
rect 35669 6614 35681 6648
rect 35681 6614 35715 6648
rect 35715 6614 35721 6648
rect 35669 6600 35721 6614
rect 34364 6425 34376 6436
rect 34376 6425 34410 6436
rect 34410 6425 34416 6436
rect 34364 6384 34416 6425
rect 32922 6193 32974 6200
rect 32922 6159 32932 6193
rect 32932 6159 32966 6193
rect 32966 6159 32974 6193
rect 32922 6148 32974 6159
rect 33272 6341 33324 6342
rect 33272 6307 33303 6341
rect 33303 6307 33324 6341
rect 33272 6290 33324 6307
rect 34126 6333 34178 6348
rect 34126 6299 34145 6333
rect 34145 6299 34178 6333
rect 34126 6296 34178 6299
rect 33296 6076 33348 6084
rect 33296 6042 33304 6076
rect 33304 6042 33338 6076
rect 33338 6042 33348 6076
rect 33296 6032 33348 6042
rect 32794 6000 32846 6006
rect 32794 5966 32804 6000
rect 32804 5966 32838 6000
rect 32838 5966 32846 6000
rect 32794 5954 32846 5966
rect 33122 5899 33174 5951
rect 33298 5899 33350 5951
rect 32360 5715 32412 5718
rect 32360 5681 32369 5715
rect 32369 5681 32403 5715
rect 32403 5681 32412 5715
rect 32360 5666 32412 5681
rect 32272 5592 32324 5602
rect 32272 5558 32283 5592
rect 32283 5558 32317 5592
rect 32317 5558 32324 5592
rect 32272 5550 32324 5558
rect 33176 5710 33228 5716
rect 33176 5676 33187 5710
rect 33187 5676 33221 5710
rect 33221 5676 33228 5710
rect 33176 5664 33228 5676
rect 32812 5529 32820 5534
rect 32820 5529 32854 5534
rect 32854 5529 32864 5534
rect 32812 5482 32864 5529
rect 33084 5594 33136 5604
rect 33084 5560 33096 5594
rect 33096 5560 33130 5594
rect 33130 5560 33136 5594
rect 33084 5552 33136 5560
rect 34914 6425 34934 6456
rect 34934 6425 34966 6456
rect 34914 6404 34966 6425
rect 36572 7056 36624 7062
rect 36572 7022 36582 7056
rect 36582 7022 36616 7056
rect 36616 7022 36624 7056
rect 36572 7010 36624 7022
rect 36885 6890 36937 6900
rect 36885 6856 36894 6890
rect 36894 6856 36928 6890
rect 36928 6856 36937 6890
rect 36885 6848 36937 6856
rect 37117 6885 37169 6890
rect 37117 6851 37137 6885
rect 37137 6851 37169 6885
rect 37117 6838 37169 6851
rect 38140 6862 38192 6868
rect 38140 6828 38150 6862
rect 38150 6828 38184 6862
rect 38184 6828 38192 6862
rect 38140 6816 38192 6828
rect 36590 6585 36598 6590
rect 36598 6585 36632 6590
rect 36632 6585 36642 6590
rect 36590 6538 36642 6585
rect 37253 6596 37305 6648
rect 37557 6648 37609 6652
rect 37557 6614 37569 6648
rect 37569 6614 37603 6648
rect 37603 6614 37609 6648
rect 37557 6600 37609 6614
rect 36252 6425 36264 6436
rect 36264 6425 36298 6436
rect 36298 6425 36304 6436
rect 36252 6384 36304 6425
rect 34810 6193 34862 6200
rect 34810 6159 34820 6193
rect 34820 6159 34854 6193
rect 34854 6159 34862 6193
rect 34810 6148 34862 6159
rect 35160 6341 35212 6342
rect 35160 6307 35191 6341
rect 35191 6307 35212 6341
rect 35160 6290 35212 6307
rect 36014 6333 36066 6348
rect 36014 6299 36033 6333
rect 36033 6299 36066 6333
rect 36014 6296 36066 6299
rect 35184 6076 35236 6084
rect 35184 6042 35192 6076
rect 35192 6042 35226 6076
rect 35226 6042 35236 6076
rect 35184 6032 35236 6042
rect 34682 6000 34734 6006
rect 34682 5966 34692 6000
rect 34692 5966 34726 6000
rect 34726 5966 34734 6000
rect 34682 5954 34734 5966
rect 35010 5899 35062 5951
rect 35186 5899 35238 5951
rect 34248 5715 34300 5718
rect 34248 5681 34257 5715
rect 34257 5681 34291 5715
rect 34291 5681 34300 5715
rect 34248 5666 34300 5681
rect 34160 5592 34212 5602
rect 34160 5558 34171 5592
rect 34171 5558 34205 5592
rect 34205 5558 34212 5592
rect 34160 5550 34212 5558
rect 35064 5710 35116 5716
rect 35064 5676 35075 5710
rect 35075 5676 35109 5710
rect 35109 5676 35116 5710
rect 35064 5664 35116 5676
rect 34700 5529 34708 5534
rect 34708 5529 34742 5534
rect 34742 5529 34752 5534
rect 34700 5482 34752 5529
rect 34972 5594 35024 5604
rect 34972 5560 34984 5594
rect 34984 5560 35018 5594
rect 35018 5560 35024 5594
rect 34972 5552 35024 5560
rect 36802 6425 36822 6456
rect 36822 6425 36854 6456
rect 36802 6404 36854 6425
rect 38460 7056 38512 7062
rect 38460 7022 38470 7056
rect 38470 7022 38504 7056
rect 38504 7022 38512 7056
rect 38460 7010 38512 7022
rect 38773 6890 38825 6900
rect 38773 6856 38782 6890
rect 38782 6856 38816 6890
rect 38816 6856 38825 6890
rect 38773 6848 38825 6856
rect 39005 6885 39057 6890
rect 39005 6851 39025 6885
rect 39025 6851 39057 6885
rect 39005 6838 39057 6851
rect 40028 6862 40080 6868
rect 40028 6828 40038 6862
rect 40038 6828 40072 6862
rect 40072 6828 40080 6862
rect 40028 6816 40080 6828
rect 38478 6585 38486 6590
rect 38486 6585 38520 6590
rect 38520 6585 38530 6590
rect 38478 6538 38530 6585
rect 39141 6596 39193 6648
rect 39445 6648 39497 6652
rect 39445 6614 39457 6648
rect 39457 6614 39491 6648
rect 39491 6614 39497 6648
rect 39445 6600 39497 6614
rect 38140 6425 38152 6436
rect 38152 6425 38186 6436
rect 38186 6425 38192 6436
rect 38140 6384 38192 6425
rect 36698 6193 36750 6200
rect 36698 6159 36708 6193
rect 36708 6159 36742 6193
rect 36742 6159 36750 6193
rect 36698 6148 36750 6159
rect 37048 6341 37100 6342
rect 37048 6307 37079 6341
rect 37079 6307 37100 6341
rect 37048 6290 37100 6307
rect 37902 6333 37954 6348
rect 37902 6299 37921 6333
rect 37921 6299 37954 6333
rect 37902 6296 37954 6299
rect 37072 6076 37124 6084
rect 37072 6042 37080 6076
rect 37080 6042 37114 6076
rect 37114 6042 37124 6076
rect 37072 6032 37124 6042
rect 36570 6000 36622 6006
rect 36570 5966 36580 6000
rect 36580 5966 36614 6000
rect 36614 5966 36622 6000
rect 36570 5954 36622 5966
rect 36898 5899 36950 5951
rect 37074 5899 37126 5951
rect 36136 5715 36188 5718
rect 36136 5681 36145 5715
rect 36145 5681 36179 5715
rect 36179 5681 36188 5715
rect 36136 5666 36188 5681
rect 36048 5592 36100 5602
rect 36048 5558 36059 5592
rect 36059 5558 36093 5592
rect 36093 5558 36100 5592
rect 36048 5550 36100 5558
rect 36952 5710 37004 5716
rect 36952 5676 36963 5710
rect 36963 5676 36997 5710
rect 36997 5676 37004 5710
rect 36952 5664 37004 5676
rect 36588 5529 36596 5534
rect 36596 5529 36630 5534
rect 36630 5529 36640 5534
rect 36588 5482 36640 5529
rect 36860 5594 36912 5604
rect 36860 5560 36872 5594
rect 36872 5560 36906 5594
rect 36906 5560 36912 5594
rect 36860 5552 36912 5560
rect 38690 6425 38710 6456
rect 38710 6425 38742 6456
rect 38690 6404 38742 6425
rect 40348 7056 40400 7062
rect 40348 7022 40358 7056
rect 40358 7022 40392 7056
rect 40392 7022 40400 7056
rect 40348 7010 40400 7022
rect 40661 6890 40713 6900
rect 40661 6856 40670 6890
rect 40670 6856 40704 6890
rect 40704 6856 40713 6890
rect 40661 6848 40713 6856
rect 40893 6885 40945 6890
rect 40893 6851 40913 6885
rect 40913 6851 40945 6885
rect 40893 6838 40945 6851
rect 41916 6862 41968 6868
rect 41916 6828 41926 6862
rect 41926 6828 41960 6862
rect 41960 6828 41968 6862
rect 41916 6816 41968 6828
rect 40366 6585 40374 6590
rect 40374 6585 40408 6590
rect 40408 6585 40418 6590
rect 40366 6538 40418 6585
rect 41029 6596 41081 6648
rect 41333 6648 41385 6652
rect 41333 6614 41345 6648
rect 41345 6614 41379 6648
rect 41379 6614 41385 6648
rect 41333 6600 41385 6614
rect 40028 6425 40040 6436
rect 40040 6425 40074 6436
rect 40074 6425 40080 6436
rect 40028 6384 40080 6425
rect 38586 6193 38638 6200
rect 38586 6159 38596 6193
rect 38596 6159 38630 6193
rect 38630 6159 38638 6193
rect 38586 6148 38638 6159
rect 38936 6341 38988 6342
rect 38936 6307 38967 6341
rect 38967 6307 38988 6341
rect 38936 6290 38988 6307
rect 39790 6333 39842 6348
rect 39790 6299 39809 6333
rect 39809 6299 39842 6333
rect 39790 6296 39842 6299
rect 38960 6076 39012 6084
rect 38960 6042 38968 6076
rect 38968 6042 39002 6076
rect 39002 6042 39012 6076
rect 38960 6032 39012 6042
rect 38458 6000 38510 6006
rect 38458 5966 38468 6000
rect 38468 5966 38502 6000
rect 38502 5966 38510 6000
rect 38458 5954 38510 5966
rect 38786 5899 38838 5951
rect 38962 5899 39014 5951
rect 38024 5715 38076 5718
rect 38024 5681 38033 5715
rect 38033 5681 38067 5715
rect 38067 5681 38076 5715
rect 38024 5666 38076 5681
rect 37936 5592 37988 5602
rect 37936 5558 37947 5592
rect 37947 5558 37981 5592
rect 37981 5558 37988 5592
rect 37936 5550 37988 5558
rect 38840 5710 38892 5716
rect 38840 5676 38851 5710
rect 38851 5676 38885 5710
rect 38885 5676 38892 5710
rect 38840 5664 38892 5676
rect 38476 5529 38484 5534
rect 38484 5529 38518 5534
rect 38518 5529 38528 5534
rect 38476 5482 38528 5529
rect 38748 5594 38800 5604
rect 38748 5560 38760 5594
rect 38760 5560 38794 5594
rect 38794 5560 38800 5594
rect 38748 5552 38800 5560
rect 40578 6425 40598 6456
rect 40598 6425 40630 6456
rect 40578 6404 40630 6425
rect 42236 7056 42288 7062
rect 42236 7022 42246 7056
rect 42246 7022 42280 7056
rect 42280 7022 42288 7056
rect 42236 7010 42288 7022
rect 42549 6890 42601 6900
rect 42549 6856 42558 6890
rect 42558 6856 42592 6890
rect 42592 6856 42601 6890
rect 42549 6848 42601 6856
rect 42781 6885 42833 6890
rect 42781 6851 42801 6885
rect 42801 6851 42833 6885
rect 42781 6838 42833 6851
rect 43804 6862 43856 6868
rect 43804 6828 43814 6862
rect 43814 6828 43848 6862
rect 43848 6828 43856 6862
rect 43804 6816 43856 6828
rect 42254 6585 42262 6590
rect 42262 6585 42296 6590
rect 42296 6585 42306 6590
rect 42254 6538 42306 6585
rect 42917 6596 42969 6648
rect 43221 6648 43273 6652
rect 43221 6614 43233 6648
rect 43233 6614 43267 6648
rect 43267 6614 43273 6648
rect 43221 6600 43273 6614
rect 41916 6425 41928 6436
rect 41928 6425 41962 6436
rect 41962 6425 41968 6436
rect 41916 6384 41968 6425
rect 40474 6193 40526 6200
rect 40474 6159 40484 6193
rect 40484 6159 40518 6193
rect 40518 6159 40526 6193
rect 40474 6148 40526 6159
rect 40824 6341 40876 6342
rect 40824 6307 40855 6341
rect 40855 6307 40876 6341
rect 40824 6290 40876 6307
rect 41678 6333 41730 6348
rect 41678 6299 41697 6333
rect 41697 6299 41730 6333
rect 41678 6296 41730 6299
rect 40848 6076 40900 6084
rect 40848 6042 40856 6076
rect 40856 6042 40890 6076
rect 40890 6042 40900 6076
rect 40848 6032 40900 6042
rect 40346 6000 40398 6006
rect 40346 5966 40356 6000
rect 40356 5966 40390 6000
rect 40390 5966 40398 6000
rect 40346 5954 40398 5966
rect 40674 5899 40726 5951
rect 40850 5899 40902 5951
rect 39912 5715 39964 5718
rect 39912 5681 39921 5715
rect 39921 5681 39955 5715
rect 39955 5681 39964 5715
rect 39912 5666 39964 5681
rect 39824 5592 39876 5602
rect 39824 5558 39835 5592
rect 39835 5558 39869 5592
rect 39869 5558 39876 5592
rect 39824 5550 39876 5558
rect 40728 5710 40780 5716
rect 40728 5676 40739 5710
rect 40739 5676 40773 5710
rect 40773 5676 40780 5710
rect 40728 5664 40780 5676
rect 40364 5529 40372 5534
rect 40372 5529 40406 5534
rect 40406 5529 40416 5534
rect 40364 5482 40416 5529
rect 40636 5594 40688 5604
rect 40636 5560 40648 5594
rect 40648 5560 40682 5594
rect 40682 5560 40688 5594
rect 40636 5552 40688 5560
rect 42466 6425 42486 6456
rect 42486 6425 42518 6456
rect 42466 6404 42518 6425
rect 44124 7056 44176 7062
rect 44124 7022 44134 7056
rect 44134 7022 44168 7056
rect 44168 7022 44176 7056
rect 44124 7010 44176 7022
rect 44437 6890 44489 6900
rect 44437 6856 44446 6890
rect 44446 6856 44480 6890
rect 44480 6856 44489 6890
rect 44437 6848 44489 6856
rect 44669 6885 44721 6890
rect 44669 6851 44689 6885
rect 44689 6851 44721 6885
rect 44669 6838 44721 6851
rect 45686 6862 45738 6868
rect 45686 6828 45696 6862
rect 45696 6828 45730 6862
rect 45730 6828 45738 6862
rect 45686 6816 45738 6828
rect 44142 6585 44150 6590
rect 44150 6585 44184 6590
rect 44184 6585 44194 6590
rect 44142 6538 44194 6585
rect 44805 6596 44857 6648
rect 45103 6648 45155 6652
rect 45103 6614 45115 6648
rect 45115 6614 45149 6648
rect 45149 6614 45155 6648
rect 45103 6600 45155 6614
rect 43804 6425 43816 6436
rect 43816 6425 43850 6436
rect 43850 6425 43856 6436
rect 43804 6384 43856 6425
rect 42362 6193 42414 6200
rect 42362 6159 42372 6193
rect 42372 6159 42406 6193
rect 42406 6159 42414 6193
rect 42362 6148 42414 6159
rect 42712 6341 42764 6342
rect 42712 6307 42743 6341
rect 42743 6307 42764 6341
rect 42712 6290 42764 6307
rect 43566 6333 43618 6348
rect 43566 6299 43585 6333
rect 43585 6299 43618 6333
rect 43566 6296 43618 6299
rect 42736 6076 42788 6084
rect 42736 6042 42744 6076
rect 42744 6042 42778 6076
rect 42778 6042 42788 6076
rect 42736 6032 42788 6042
rect 42234 6000 42286 6006
rect 42234 5966 42244 6000
rect 42244 5966 42278 6000
rect 42278 5966 42286 6000
rect 42234 5954 42286 5966
rect 42562 5899 42614 5951
rect 42738 5899 42790 5951
rect 41800 5715 41852 5718
rect 41800 5681 41809 5715
rect 41809 5681 41843 5715
rect 41843 5681 41852 5715
rect 41800 5666 41852 5681
rect 41712 5592 41764 5602
rect 41712 5558 41723 5592
rect 41723 5558 41757 5592
rect 41757 5558 41764 5592
rect 41712 5550 41764 5558
rect 42616 5710 42668 5716
rect 42616 5676 42627 5710
rect 42627 5676 42661 5710
rect 42661 5676 42668 5710
rect 42616 5664 42668 5676
rect 42252 5529 42260 5534
rect 42260 5529 42294 5534
rect 42294 5529 42304 5534
rect 42252 5482 42304 5529
rect 42524 5594 42576 5604
rect 42524 5560 42536 5594
rect 42536 5560 42570 5594
rect 42570 5560 42576 5594
rect 42524 5552 42576 5560
rect 44354 6425 44374 6456
rect 44374 6425 44406 6456
rect 44354 6404 44406 6425
rect 46006 7056 46058 7062
rect 46006 7022 46016 7056
rect 46016 7022 46050 7056
rect 46050 7022 46058 7056
rect 46006 7010 46058 7022
rect 46319 6890 46371 6900
rect 46319 6856 46328 6890
rect 46328 6856 46362 6890
rect 46362 6856 46371 6890
rect 46319 6848 46371 6856
rect 46551 6885 46603 6890
rect 46551 6851 46571 6885
rect 46571 6851 46603 6885
rect 46551 6838 46603 6851
rect 47574 6862 47626 6868
rect 47574 6828 47584 6862
rect 47584 6828 47618 6862
rect 47618 6828 47626 6862
rect 47574 6816 47626 6828
rect 46024 6585 46032 6590
rect 46032 6585 46066 6590
rect 46066 6585 46076 6590
rect 46024 6538 46076 6585
rect 46687 6596 46739 6648
rect 46991 6648 47043 6652
rect 46991 6614 47003 6648
rect 47003 6614 47037 6648
rect 47037 6614 47043 6648
rect 46991 6600 47043 6614
rect 45686 6425 45698 6436
rect 45698 6425 45732 6436
rect 45732 6425 45738 6436
rect 45686 6384 45738 6425
rect 44250 6193 44302 6200
rect 44250 6159 44260 6193
rect 44260 6159 44294 6193
rect 44294 6159 44302 6193
rect 44250 6148 44302 6159
rect 44600 6341 44652 6342
rect 44600 6307 44631 6341
rect 44631 6307 44652 6341
rect 44600 6290 44652 6307
rect 45448 6333 45500 6348
rect 45448 6299 45467 6333
rect 45467 6299 45500 6333
rect 45448 6296 45500 6299
rect 44624 6076 44676 6084
rect 44624 6042 44632 6076
rect 44632 6042 44666 6076
rect 44666 6042 44676 6076
rect 44624 6032 44676 6042
rect 44122 6000 44174 6006
rect 44122 5966 44132 6000
rect 44132 5966 44166 6000
rect 44166 5966 44174 6000
rect 44122 5954 44174 5966
rect 44450 5899 44502 5951
rect 44626 5899 44678 5951
rect 43688 5715 43740 5718
rect 43688 5681 43697 5715
rect 43697 5681 43731 5715
rect 43731 5681 43740 5715
rect 43688 5666 43740 5681
rect 43600 5592 43652 5602
rect 43600 5558 43611 5592
rect 43611 5558 43645 5592
rect 43645 5558 43652 5592
rect 43600 5550 43652 5558
rect 44504 5710 44556 5716
rect 44504 5676 44515 5710
rect 44515 5676 44549 5710
rect 44549 5676 44556 5710
rect 44504 5664 44556 5676
rect 44140 5529 44148 5534
rect 44148 5529 44182 5534
rect 44182 5529 44192 5534
rect 44140 5482 44192 5529
rect 44412 5594 44464 5604
rect 44412 5560 44424 5594
rect 44424 5560 44458 5594
rect 44458 5560 44464 5594
rect 44412 5552 44464 5560
rect 46236 6425 46256 6456
rect 46256 6425 46288 6456
rect 46236 6404 46288 6425
rect 47894 7056 47946 7062
rect 47894 7022 47904 7056
rect 47904 7022 47938 7056
rect 47938 7022 47946 7056
rect 47894 7010 47946 7022
rect 48207 6890 48259 6900
rect 48207 6856 48216 6890
rect 48216 6856 48250 6890
rect 48250 6856 48259 6890
rect 48207 6848 48259 6856
rect 48439 6885 48491 6890
rect 48439 6851 48459 6885
rect 48459 6851 48491 6885
rect 48439 6838 48491 6851
rect 49462 6862 49514 6868
rect 49462 6828 49472 6862
rect 49472 6828 49506 6862
rect 49506 6828 49514 6862
rect 49462 6816 49514 6828
rect 47912 6585 47920 6590
rect 47920 6585 47954 6590
rect 47954 6585 47964 6590
rect 47912 6538 47964 6585
rect 48575 6596 48627 6648
rect 48879 6648 48931 6652
rect 48879 6614 48891 6648
rect 48891 6614 48925 6648
rect 48925 6614 48931 6648
rect 48879 6600 48931 6614
rect 47574 6425 47586 6436
rect 47586 6425 47620 6436
rect 47620 6425 47626 6436
rect 47574 6384 47626 6425
rect 46132 6193 46184 6200
rect 46132 6159 46142 6193
rect 46142 6159 46176 6193
rect 46176 6159 46184 6193
rect 46132 6148 46184 6159
rect 46482 6341 46534 6342
rect 46482 6307 46513 6341
rect 46513 6307 46534 6341
rect 46482 6290 46534 6307
rect 47336 6333 47388 6348
rect 47336 6299 47355 6333
rect 47355 6299 47388 6333
rect 47336 6296 47388 6299
rect 46506 6076 46558 6084
rect 46506 6042 46514 6076
rect 46514 6042 46548 6076
rect 46548 6042 46558 6076
rect 46506 6032 46558 6042
rect 46004 6000 46056 6006
rect 46004 5966 46014 6000
rect 46014 5966 46048 6000
rect 46048 5966 46056 6000
rect 46004 5954 46056 5966
rect 46332 5899 46384 5951
rect 46508 5899 46560 5951
rect 45570 5715 45622 5718
rect 45570 5681 45579 5715
rect 45579 5681 45613 5715
rect 45613 5681 45622 5715
rect 45570 5666 45622 5681
rect 45482 5592 45534 5602
rect 45482 5558 45493 5592
rect 45493 5558 45527 5592
rect 45527 5558 45534 5592
rect 45482 5550 45534 5558
rect 46386 5710 46438 5716
rect 46386 5676 46397 5710
rect 46397 5676 46431 5710
rect 46431 5676 46438 5710
rect 46386 5664 46438 5676
rect 46022 5529 46030 5534
rect 46030 5529 46064 5534
rect 46064 5529 46074 5534
rect 46022 5482 46074 5529
rect 46294 5594 46346 5604
rect 46294 5560 46306 5594
rect 46306 5560 46340 5594
rect 46340 5560 46346 5594
rect 46294 5552 46346 5560
rect 48124 6425 48144 6456
rect 48144 6425 48176 6456
rect 48124 6404 48176 6425
rect 49782 7056 49834 7062
rect 49782 7022 49792 7056
rect 49792 7022 49826 7056
rect 49826 7022 49834 7056
rect 49782 7010 49834 7022
rect 50095 6890 50147 6900
rect 50095 6856 50104 6890
rect 50104 6856 50138 6890
rect 50138 6856 50147 6890
rect 50095 6848 50147 6856
rect 50327 6885 50379 6890
rect 50327 6851 50347 6885
rect 50347 6851 50379 6885
rect 50327 6838 50379 6851
rect 51350 6862 51402 6868
rect 51350 6828 51360 6862
rect 51360 6828 51394 6862
rect 51394 6828 51402 6862
rect 51350 6816 51402 6828
rect 49800 6585 49808 6590
rect 49808 6585 49842 6590
rect 49842 6585 49852 6590
rect 49800 6538 49852 6585
rect 50463 6596 50515 6648
rect 50767 6648 50819 6652
rect 50767 6614 50779 6648
rect 50779 6614 50813 6648
rect 50813 6614 50819 6648
rect 50767 6600 50819 6614
rect 49462 6425 49474 6436
rect 49474 6425 49508 6436
rect 49508 6425 49514 6436
rect 49462 6384 49514 6425
rect 48020 6193 48072 6200
rect 48020 6159 48030 6193
rect 48030 6159 48064 6193
rect 48064 6159 48072 6193
rect 48020 6148 48072 6159
rect 48370 6341 48422 6342
rect 48370 6307 48401 6341
rect 48401 6307 48422 6341
rect 48370 6290 48422 6307
rect 49224 6333 49276 6348
rect 49224 6299 49243 6333
rect 49243 6299 49276 6333
rect 49224 6296 49276 6299
rect 48394 6076 48446 6084
rect 48394 6042 48402 6076
rect 48402 6042 48436 6076
rect 48436 6042 48446 6076
rect 48394 6032 48446 6042
rect 47892 6000 47944 6006
rect 47892 5966 47902 6000
rect 47902 5966 47936 6000
rect 47936 5966 47944 6000
rect 47892 5954 47944 5966
rect 48220 5899 48272 5951
rect 48396 5899 48448 5951
rect 47458 5715 47510 5718
rect 47458 5681 47467 5715
rect 47467 5681 47501 5715
rect 47501 5681 47510 5715
rect 47458 5666 47510 5681
rect 47370 5592 47422 5602
rect 47370 5558 47381 5592
rect 47381 5558 47415 5592
rect 47415 5558 47422 5592
rect 47370 5550 47422 5558
rect 48274 5710 48326 5716
rect 48274 5676 48285 5710
rect 48285 5676 48319 5710
rect 48319 5676 48326 5710
rect 48274 5664 48326 5676
rect 47910 5529 47918 5534
rect 47918 5529 47952 5534
rect 47952 5529 47962 5534
rect 47910 5482 47962 5529
rect 48182 5594 48234 5604
rect 48182 5560 48194 5594
rect 48194 5560 48228 5594
rect 48228 5560 48234 5594
rect 48182 5552 48234 5560
rect 50012 6425 50032 6456
rect 50032 6425 50064 6456
rect 50012 6404 50064 6425
rect 51670 7056 51722 7062
rect 51670 7022 51680 7056
rect 51680 7022 51714 7056
rect 51714 7022 51722 7056
rect 51670 7010 51722 7022
rect 51983 6890 52035 6900
rect 51983 6856 51992 6890
rect 51992 6856 52026 6890
rect 52026 6856 52035 6890
rect 51983 6848 52035 6856
rect 52215 6885 52267 6890
rect 52215 6851 52235 6885
rect 52235 6851 52267 6885
rect 52215 6838 52267 6851
rect 53238 6862 53290 6868
rect 53238 6828 53248 6862
rect 53248 6828 53282 6862
rect 53282 6828 53290 6862
rect 53238 6816 53290 6828
rect 51688 6585 51696 6590
rect 51696 6585 51730 6590
rect 51730 6585 51740 6590
rect 51688 6538 51740 6585
rect 52351 6596 52403 6648
rect 52655 6648 52707 6652
rect 52655 6614 52667 6648
rect 52667 6614 52701 6648
rect 52701 6614 52707 6648
rect 52655 6600 52707 6614
rect 51350 6425 51362 6436
rect 51362 6425 51396 6436
rect 51396 6425 51402 6436
rect 51350 6384 51402 6425
rect 49908 6193 49960 6200
rect 49908 6159 49918 6193
rect 49918 6159 49952 6193
rect 49952 6159 49960 6193
rect 49908 6148 49960 6159
rect 50258 6341 50310 6342
rect 50258 6307 50289 6341
rect 50289 6307 50310 6341
rect 50258 6290 50310 6307
rect 51112 6333 51164 6348
rect 51112 6299 51131 6333
rect 51131 6299 51164 6333
rect 51112 6296 51164 6299
rect 50282 6076 50334 6084
rect 50282 6042 50290 6076
rect 50290 6042 50324 6076
rect 50324 6042 50334 6076
rect 50282 6032 50334 6042
rect 49780 6000 49832 6006
rect 49780 5966 49790 6000
rect 49790 5966 49824 6000
rect 49824 5966 49832 6000
rect 49780 5954 49832 5966
rect 50108 5899 50160 5951
rect 50284 5899 50336 5951
rect 49346 5715 49398 5718
rect 49346 5681 49355 5715
rect 49355 5681 49389 5715
rect 49389 5681 49398 5715
rect 49346 5666 49398 5681
rect 49258 5592 49310 5602
rect 49258 5558 49269 5592
rect 49269 5558 49303 5592
rect 49303 5558 49310 5592
rect 49258 5550 49310 5558
rect 50162 5710 50214 5716
rect 50162 5676 50173 5710
rect 50173 5676 50207 5710
rect 50207 5676 50214 5710
rect 50162 5664 50214 5676
rect 49798 5529 49806 5534
rect 49806 5529 49840 5534
rect 49840 5529 49850 5534
rect 49798 5482 49850 5529
rect 50070 5594 50122 5604
rect 50070 5560 50082 5594
rect 50082 5560 50116 5594
rect 50116 5560 50122 5594
rect 50070 5552 50122 5560
rect 51900 6425 51920 6456
rect 51920 6425 51952 6456
rect 51900 6404 51952 6425
rect 53558 7056 53610 7062
rect 53558 7022 53568 7056
rect 53568 7022 53602 7056
rect 53602 7022 53610 7056
rect 53558 7010 53610 7022
rect 53871 6890 53923 6900
rect 53871 6856 53880 6890
rect 53880 6856 53914 6890
rect 53914 6856 53923 6890
rect 53871 6848 53923 6856
rect 54103 6885 54155 6890
rect 54103 6851 54123 6885
rect 54123 6851 54155 6885
rect 54103 6838 54155 6851
rect 55126 6862 55178 6868
rect 55126 6828 55136 6862
rect 55136 6828 55170 6862
rect 55170 6828 55178 6862
rect 55126 6816 55178 6828
rect 53576 6585 53584 6590
rect 53584 6585 53618 6590
rect 53618 6585 53628 6590
rect 53576 6538 53628 6585
rect 54239 6596 54291 6648
rect 54543 6648 54595 6652
rect 54543 6614 54555 6648
rect 54555 6614 54589 6648
rect 54589 6614 54595 6648
rect 54543 6600 54595 6614
rect 53238 6425 53250 6436
rect 53250 6425 53284 6436
rect 53284 6425 53290 6436
rect 53238 6384 53290 6425
rect 51796 6193 51848 6200
rect 51796 6159 51806 6193
rect 51806 6159 51840 6193
rect 51840 6159 51848 6193
rect 51796 6148 51848 6159
rect 52146 6341 52198 6342
rect 52146 6307 52177 6341
rect 52177 6307 52198 6341
rect 52146 6290 52198 6307
rect 53000 6333 53052 6348
rect 53000 6299 53019 6333
rect 53019 6299 53052 6333
rect 53000 6296 53052 6299
rect 52170 6076 52222 6084
rect 52170 6042 52178 6076
rect 52178 6042 52212 6076
rect 52212 6042 52222 6076
rect 52170 6032 52222 6042
rect 51668 6000 51720 6006
rect 51668 5966 51678 6000
rect 51678 5966 51712 6000
rect 51712 5966 51720 6000
rect 51668 5954 51720 5966
rect 51996 5899 52048 5951
rect 52172 5899 52224 5951
rect 51234 5715 51286 5718
rect 51234 5681 51243 5715
rect 51243 5681 51277 5715
rect 51277 5681 51286 5715
rect 51234 5666 51286 5681
rect 51146 5592 51198 5602
rect 51146 5558 51157 5592
rect 51157 5558 51191 5592
rect 51191 5558 51198 5592
rect 51146 5550 51198 5558
rect 52050 5710 52102 5716
rect 52050 5676 52061 5710
rect 52061 5676 52095 5710
rect 52095 5676 52102 5710
rect 52050 5664 52102 5676
rect 51686 5529 51694 5534
rect 51694 5529 51728 5534
rect 51728 5529 51738 5534
rect 51686 5482 51738 5529
rect 51958 5594 52010 5604
rect 51958 5560 51970 5594
rect 51970 5560 52004 5594
rect 52004 5560 52010 5594
rect 51958 5552 52010 5560
rect 53788 6425 53808 6456
rect 53808 6425 53840 6456
rect 53788 6404 53840 6425
rect 55446 7056 55498 7062
rect 55446 7022 55456 7056
rect 55456 7022 55490 7056
rect 55490 7022 55498 7056
rect 55446 7010 55498 7022
rect 55759 6890 55811 6900
rect 55759 6856 55768 6890
rect 55768 6856 55802 6890
rect 55802 6856 55811 6890
rect 55759 6848 55811 6856
rect 55991 6885 56043 6890
rect 55991 6851 56011 6885
rect 56011 6851 56043 6885
rect 55991 6838 56043 6851
rect 57014 6862 57066 6868
rect 57014 6828 57024 6862
rect 57024 6828 57058 6862
rect 57058 6828 57066 6862
rect 57014 6816 57066 6828
rect 55464 6585 55472 6590
rect 55472 6585 55506 6590
rect 55506 6585 55516 6590
rect 55464 6538 55516 6585
rect 56127 6596 56179 6648
rect 56431 6648 56483 6652
rect 56431 6614 56443 6648
rect 56443 6614 56477 6648
rect 56477 6614 56483 6648
rect 56431 6600 56483 6614
rect 55126 6425 55138 6436
rect 55138 6425 55172 6436
rect 55172 6425 55178 6436
rect 55126 6384 55178 6425
rect 53684 6193 53736 6200
rect 53684 6159 53694 6193
rect 53694 6159 53728 6193
rect 53728 6159 53736 6193
rect 53684 6148 53736 6159
rect 54034 6341 54086 6342
rect 54034 6307 54065 6341
rect 54065 6307 54086 6341
rect 54034 6290 54086 6307
rect 54888 6333 54940 6348
rect 54888 6299 54907 6333
rect 54907 6299 54940 6333
rect 54888 6296 54940 6299
rect 54058 6076 54110 6084
rect 54058 6042 54066 6076
rect 54066 6042 54100 6076
rect 54100 6042 54110 6076
rect 54058 6032 54110 6042
rect 53556 6000 53608 6006
rect 53556 5966 53566 6000
rect 53566 5966 53600 6000
rect 53600 5966 53608 6000
rect 53556 5954 53608 5966
rect 53884 5899 53936 5951
rect 54060 5899 54112 5951
rect 53122 5715 53174 5718
rect 53122 5681 53131 5715
rect 53131 5681 53165 5715
rect 53165 5681 53174 5715
rect 53122 5666 53174 5681
rect 53034 5592 53086 5602
rect 53034 5558 53045 5592
rect 53045 5558 53079 5592
rect 53079 5558 53086 5592
rect 53034 5550 53086 5558
rect 53938 5710 53990 5716
rect 53938 5676 53949 5710
rect 53949 5676 53983 5710
rect 53983 5676 53990 5710
rect 53938 5664 53990 5676
rect 53574 5529 53582 5534
rect 53582 5529 53616 5534
rect 53616 5529 53626 5534
rect 53574 5482 53626 5529
rect 53846 5594 53898 5604
rect 53846 5560 53858 5594
rect 53858 5560 53892 5594
rect 53892 5560 53898 5594
rect 53846 5552 53898 5560
rect 55676 6425 55696 6456
rect 55696 6425 55728 6456
rect 55676 6404 55728 6425
rect 57334 7056 57386 7062
rect 57334 7022 57344 7056
rect 57344 7022 57378 7056
rect 57378 7022 57386 7056
rect 57334 7010 57386 7022
rect 57647 6890 57699 6900
rect 57647 6856 57656 6890
rect 57656 6856 57690 6890
rect 57690 6856 57699 6890
rect 57647 6848 57699 6856
rect 57879 6885 57931 6890
rect 57879 6851 57899 6885
rect 57899 6851 57931 6885
rect 57879 6838 57931 6851
rect 58902 6862 58954 6868
rect 58902 6828 58912 6862
rect 58912 6828 58946 6862
rect 58946 6828 58954 6862
rect 58902 6816 58954 6828
rect 57352 6585 57360 6590
rect 57360 6585 57394 6590
rect 57394 6585 57404 6590
rect 57352 6538 57404 6585
rect 58015 6596 58067 6648
rect 58319 6648 58371 6652
rect 58319 6614 58331 6648
rect 58331 6614 58365 6648
rect 58365 6614 58371 6648
rect 58319 6600 58371 6614
rect 57014 6425 57026 6436
rect 57026 6425 57060 6436
rect 57060 6425 57066 6436
rect 57014 6384 57066 6425
rect 55572 6193 55624 6200
rect 55572 6159 55582 6193
rect 55582 6159 55616 6193
rect 55616 6159 55624 6193
rect 55572 6148 55624 6159
rect 55922 6341 55974 6342
rect 55922 6307 55953 6341
rect 55953 6307 55974 6341
rect 55922 6290 55974 6307
rect 56776 6333 56828 6348
rect 56776 6299 56795 6333
rect 56795 6299 56828 6333
rect 56776 6296 56828 6299
rect 55946 6076 55998 6084
rect 55946 6042 55954 6076
rect 55954 6042 55988 6076
rect 55988 6042 55998 6076
rect 55946 6032 55998 6042
rect 55444 6000 55496 6006
rect 55444 5966 55454 6000
rect 55454 5966 55488 6000
rect 55488 5966 55496 6000
rect 55444 5954 55496 5966
rect 55772 5899 55824 5951
rect 55948 5899 56000 5951
rect 55010 5715 55062 5718
rect 55010 5681 55019 5715
rect 55019 5681 55053 5715
rect 55053 5681 55062 5715
rect 55010 5666 55062 5681
rect 54922 5592 54974 5602
rect 54922 5558 54933 5592
rect 54933 5558 54967 5592
rect 54967 5558 54974 5592
rect 54922 5550 54974 5558
rect 55826 5710 55878 5716
rect 55826 5676 55837 5710
rect 55837 5676 55871 5710
rect 55871 5676 55878 5710
rect 55826 5664 55878 5676
rect 55462 5529 55470 5534
rect 55470 5529 55504 5534
rect 55504 5529 55514 5534
rect 55462 5482 55514 5529
rect 55734 5594 55786 5604
rect 55734 5560 55746 5594
rect 55746 5560 55780 5594
rect 55780 5560 55786 5594
rect 55734 5552 55786 5560
rect 57564 6425 57584 6456
rect 57584 6425 57616 6456
rect 57564 6404 57616 6425
rect 59222 7056 59274 7062
rect 59222 7022 59232 7056
rect 59232 7022 59266 7056
rect 59266 7022 59274 7056
rect 59222 7010 59274 7022
rect 59535 6890 59587 6900
rect 59535 6856 59544 6890
rect 59544 6856 59578 6890
rect 59578 6856 59587 6890
rect 59535 6848 59587 6856
rect 59767 6885 59819 6890
rect 59767 6851 59787 6885
rect 59787 6851 59819 6885
rect 59767 6838 59819 6851
rect 59240 6585 59248 6590
rect 59248 6585 59282 6590
rect 59282 6585 59292 6590
rect 59240 6538 59292 6585
rect 59903 6596 59955 6648
rect 58902 6425 58914 6436
rect 58914 6425 58948 6436
rect 58948 6425 58954 6436
rect 58902 6384 58954 6425
rect 57460 6193 57512 6200
rect 57460 6159 57470 6193
rect 57470 6159 57504 6193
rect 57504 6159 57512 6193
rect 57460 6148 57512 6159
rect 57810 6341 57862 6342
rect 57810 6307 57841 6341
rect 57841 6307 57862 6341
rect 57810 6290 57862 6307
rect 58664 6333 58716 6348
rect 58664 6299 58683 6333
rect 58683 6299 58716 6333
rect 58664 6296 58716 6299
rect 57834 6076 57886 6084
rect 57834 6042 57842 6076
rect 57842 6042 57876 6076
rect 57876 6042 57886 6076
rect 57834 6032 57886 6042
rect 57332 6000 57384 6006
rect 57332 5966 57342 6000
rect 57342 5966 57376 6000
rect 57376 5966 57384 6000
rect 57332 5954 57384 5966
rect 57660 5899 57712 5951
rect 57836 5899 57888 5951
rect 56898 5715 56950 5718
rect 56898 5681 56907 5715
rect 56907 5681 56941 5715
rect 56941 5681 56950 5715
rect 56898 5666 56950 5681
rect 56810 5592 56862 5602
rect 56810 5558 56821 5592
rect 56821 5558 56855 5592
rect 56855 5558 56862 5592
rect 56810 5550 56862 5558
rect 57714 5710 57766 5716
rect 57714 5676 57725 5710
rect 57725 5676 57759 5710
rect 57759 5676 57766 5710
rect 57714 5664 57766 5676
rect 57350 5529 57358 5534
rect 57358 5529 57392 5534
rect 57392 5529 57402 5534
rect 57350 5482 57402 5529
rect 57622 5594 57674 5604
rect 57622 5560 57634 5594
rect 57634 5560 57668 5594
rect 57668 5560 57674 5594
rect 57622 5552 57674 5560
rect 59452 6425 59472 6456
rect 59472 6425 59504 6456
rect 59452 6404 59504 6425
rect 59348 6193 59400 6200
rect 59348 6159 59358 6193
rect 59358 6159 59392 6193
rect 59392 6159 59400 6193
rect 59348 6148 59400 6159
rect 59698 6341 59750 6342
rect 59698 6307 59729 6341
rect 59729 6307 59750 6341
rect 59698 6290 59750 6307
rect 59722 6076 59774 6084
rect 59722 6042 59730 6076
rect 59730 6042 59764 6076
rect 59764 6042 59774 6076
rect 59722 6032 59774 6042
rect 59220 6000 59272 6006
rect 59220 5966 59230 6000
rect 59230 5966 59264 6000
rect 59264 5966 59272 6000
rect 59220 5954 59272 5966
rect 59548 5899 59600 5951
rect 59724 5899 59776 5951
rect 58786 5715 58838 5718
rect 58786 5681 58795 5715
rect 58795 5681 58829 5715
rect 58829 5681 58838 5715
rect 58786 5666 58838 5681
rect 58698 5592 58750 5602
rect 58698 5558 58709 5592
rect 58709 5558 58743 5592
rect 58743 5558 58750 5592
rect 58698 5550 58750 5558
rect 59602 5710 59654 5716
rect 59602 5676 59613 5710
rect 59613 5676 59647 5710
rect 59647 5676 59654 5710
rect 59602 5664 59654 5676
rect 59238 5529 59246 5534
rect 59246 5529 59280 5534
rect 59280 5529 59290 5534
rect 59238 5482 59290 5529
rect 59510 5594 59562 5604
rect 59510 5560 59522 5594
rect 59522 5560 59556 5594
rect 59556 5560 59562 5594
rect 59510 5552 59562 5560
rect -377 5136 -69 5252
rect 1511 5136 1819 5252
rect 3399 5136 3707 5252
rect 5287 5136 5595 5252
rect 7175 5136 7483 5252
rect 9063 5136 9371 5252
rect 10951 5136 11259 5252
rect 12839 5136 13147 5252
rect 14721 5136 15029 5252
rect 16609 5136 16917 5252
rect 18497 5136 18805 5252
rect 20385 5136 20693 5252
rect 22273 5136 22581 5252
rect 24161 5136 24469 5252
rect 26049 5136 26357 5252
rect 27937 5136 28245 5252
rect 29825 5136 30133 5252
rect 31713 5136 32021 5252
rect 33601 5136 33909 5252
rect 35489 5136 35797 5252
rect 37377 5136 37685 5252
rect 39265 5136 39573 5252
rect 41153 5136 41461 5252
rect 43041 5136 43349 5252
rect 44923 5136 45231 5252
rect 46811 5136 47119 5252
rect 48699 5136 49007 5252
rect 50587 5136 50895 5252
rect 52475 5136 52783 5252
rect 54363 5136 54671 5252
rect 56251 5136 56559 5252
rect 58139 5136 58447 5252
rect 5864 4967 5916 5019
rect 5979 5009 6031 5019
rect 5979 4975 5996 5009
rect 5996 4975 6031 5009
rect 5979 4967 6031 4975
rect 6106 5007 6158 5019
rect 6106 4973 6132 5007
rect 6132 4973 6158 5007
rect 6106 4967 6158 4973
rect 6223 4967 6275 5019
rect 6337 4967 6389 5019
rect 6456 4993 6508 5018
rect 6456 4966 6466 4993
rect 6466 4966 6500 4993
rect 6500 4966 6508 4993
rect 6554 4966 6606 5018
rect 6650 4996 6702 5018
rect 6650 4966 6671 4996
rect 6671 4966 6702 4996
rect 6758 5001 6810 5018
rect 6758 4967 6799 5001
rect 6799 4967 6810 5001
rect 6758 4966 6810 4967
rect 6857 4966 6909 5018
rect 6951 5002 7003 5018
rect 6951 4968 6972 5002
rect 6972 4968 7003 5002
rect 6951 4966 7003 4968
rect 7665 4965 7717 5017
rect 7761 4965 7813 5017
rect 7850 5003 7902 5016
rect 7850 4969 7879 5003
rect 7879 4969 7902 5003
rect 7850 4964 7902 4969
rect 7950 4964 8002 5016
rect 8047 5012 8099 5016
rect 8047 4978 8049 5012
rect 8049 4978 8099 5012
rect 8184 5010 8236 5016
rect 8047 4964 8099 4978
rect 8184 4976 8217 5010
rect 8217 4976 8236 5010
rect 8184 4964 8236 4976
rect 8338 4997 8390 5016
rect 8338 4964 8350 4997
rect 8350 4964 8384 4997
rect 8384 4964 8390 4997
rect 8464 5002 8516 5014
rect 8464 4968 8515 5002
rect 8515 4968 8516 5002
rect 8464 4962 8516 4968
rect 8566 4962 8618 5014
rect 8673 5006 8725 5014
rect 8673 4972 8688 5006
rect 8688 4972 8722 5006
rect 8722 4972 8725 5006
rect 8673 4962 8725 4972
rect 8785 4960 8837 5012
rect 7264 4761 7316 4813
rect 7345 4760 7397 4812
rect 20891 4996 20943 5020
rect 20891 4968 20901 4996
rect 20901 4968 20935 4996
rect 20935 4968 20943 4996
rect 20988 4968 21040 5020
rect 21085 4998 21137 5020
rect 21085 4968 21094 4998
rect 21094 4968 21137 4998
rect 21191 5000 21243 5020
rect 21191 4968 21230 5000
rect 21230 4968 21243 5000
rect 21296 4968 21348 5020
rect 21413 5006 21465 5020
rect 21413 4972 21434 5006
rect 21434 4972 21465 5006
rect 21413 4968 21465 4972
rect 21547 5018 21599 5019
rect 21547 4993 21606 5018
rect 21547 4967 21564 4993
rect 21554 4966 21564 4967
rect 21564 4966 21598 4993
rect 21598 4966 21606 4993
rect 21676 4969 21728 5021
rect 21792 4969 21844 5021
rect 21898 4997 21950 5021
rect 21898 4969 21900 4997
rect 21900 4969 21934 4997
rect 21934 4969 21950 4997
rect 22005 4969 22057 5021
rect 22780 4994 22832 5017
rect 22780 4965 22808 4994
rect 22808 4965 22832 4994
rect 22877 4965 22929 5017
rect 22974 4996 23026 5017
rect 22974 4965 22978 4996
rect 22978 4965 23026 4996
rect 23080 5002 23132 5017
rect 23080 4968 23110 5002
rect 23110 4968 23132 5002
rect 23080 4965 23132 4968
rect 23185 4965 23237 5017
rect 23302 5001 23354 5017
rect 23302 4967 23313 5001
rect 23313 4967 23354 5001
rect 23302 4965 23354 4967
rect 23436 4997 23488 5016
rect 23436 4964 23448 4997
rect 23448 4964 23482 4997
rect 23482 4964 23488 4997
rect 23565 4966 23617 5018
rect 23681 4966 23733 5018
rect 23787 4997 23839 5018
rect 23787 4966 23817 4997
rect 23817 4966 23839 4997
rect 23894 4966 23946 5018
rect 22380 4758 22432 4810
rect 22475 4758 22527 4810
rect 36066 4967 36118 5019
rect 36181 5009 36233 5019
rect 36181 4975 36198 5009
rect 36198 4975 36233 5009
rect 36181 4967 36233 4975
rect 36308 5007 36360 5019
rect 36308 4973 36334 5007
rect 36334 4973 36360 5007
rect 36308 4967 36360 4973
rect 36425 4967 36477 5019
rect 36539 4967 36591 5019
rect 36658 4993 36710 5018
rect 36658 4966 36668 4993
rect 36668 4966 36702 4993
rect 36702 4966 36710 4993
rect 36756 4966 36808 5018
rect 36852 4996 36904 5018
rect 36852 4966 36873 4996
rect 36873 4966 36904 4996
rect 36960 5001 37012 5018
rect 36960 4967 37001 5001
rect 37001 4967 37012 5001
rect 36960 4966 37012 4967
rect 37059 4966 37111 5018
rect 37153 5002 37205 5018
rect 37153 4968 37174 5002
rect 37174 4968 37205 5002
rect 37153 4966 37205 4968
rect 37867 4965 37919 5017
rect 37963 4965 38015 5017
rect 38052 5003 38104 5016
rect 38052 4969 38081 5003
rect 38081 4969 38104 5003
rect 38052 4964 38104 4969
rect 38152 4964 38204 5016
rect 38249 5012 38301 5016
rect 38249 4978 38251 5012
rect 38251 4978 38301 5012
rect 38386 5010 38438 5016
rect 38249 4964 38301 4978
rect 38386 4976 38419 5010
rect 38419 4976 38438 5010
rect 38386 4964 38438 4976
rect 38540 4997 38592 5016
rect 38540 4964 38552 4997
rect 38552 4964 38586 4997
rect 38586 4964 38592 4997
rect 38666 5002 38718 5014
rect 38666 4968 38717 5002
rect 38717 4968 38718 5002
rect 38666 4962 38718 4968
rect 38768 4962 38820 5014
rect 38875 5006 38927 5014
rect 38875 4972 38890 5006
rect 38890 4972 38924 5006
rect 38924 4972 38927 5006
rect 38875 4962 38927 4972
rect 38987 4960 39039 5012
rect 14443 4695 14495 4747
rect 14521 4695 14573 4747
rect 14614 4695 14666 4747
rect 30402 4718 30454 4770
rect 30515 4718 30567 4770
rect 30616 4718 30668 4770
rect 37457 4760 37509 4812
rect 37559 4760 37611 4812
rect 51093 4996 51145 5020
rect 51093 4968 51103 4996
rect 51103 4968 51137 4996
rect 51137 4968 51145 4996
rect 51190 4968 51242 5020
rect 51287 4998 51339 5020
rect 51287 4968 51296 4998
rect 51296 4968 51339 4998
rect 51393 5000 51445 5020
rect 51393 4968 51432 5000
rect 51432 4968 51445 5000
rect 51498 4968 51550 5020
rect 51615 5006 51667 5020
rect 51615 4972 51636 5006
rect 51636 4972 51667 5006
rect 51615 4968 51667 4972
rect 51749 5018 51801 5019
rect 51749 4993 51808 5018
rect 51749 4967 51766 4993
rect 51756 4966 51766 4967
rect 51766 4966 51800 4993
rect 51800 4966 51808 4993
rect 51878 4969 51930 5021
rect 51994 4969 52046 5021
rect 52100 4997 52152 5021
rect 52100 4969 52102 4997
rect 52102 4969 52136 4997
rect 52136 4969 52152 4997
rect 52207 4969 52259 5021
rect 52982 4994 53034 5017
rect 52982 4965 53010 4994
rect 53010 4965 53034 4994
rect 53079 4965 53131 5017
rect 53176 4996 53228 5017
rect 53176 4965 53180 4996
rect 53180 4965 53228 4996
rect 53282 5002 53334 5017
rect 53282 4968 53312 5002
rect 53312 4968 53334 5002
rect 53282 4965 53334 4968
rect 53387 4965 53439 5017
rect 53504 5001 53556 5017
rect 53504 4967 53515 5001
rect 53515 4967 53556 5001
rect 53504 4965 53556 4967
rect 53638 4997 53690 5016
rect 53638 4964 53650 4997
rect 53650 4964 53684 4997
rect 53684 4964 53690 4997
rect 53767 4966 53819 5018
rect 53883 4966 53935 5018
rect 53989 4997 54041 5018
rect 53989 4966 54019 4997
rect 54019 4966 54041 4997
rect 54096 4966 54148 5018
rect 6272 4665 6324 4667
rect 6379 4665 6431 4669
rect 6481 4665 6533 4669
rect 6581 4665 6633 4670
rect 44594 4695 44646 4747
rect 44677 4695 44729 4747
rect 52575 4733 52627 4785
rect 52670 4733 52722 4785
rect 21302 4665 21354 4673
rect 21405 4665 21457 4673
rect 21488 4665 21540 4673
rect 21589 4665 21641 4673
rect 21676 4665 21728 4673
rect 6272 4631 6279 4665
rect 6279 4631 6324 4665
rect 6379 4631 6429 4665
rect 6429 4631 6431 4665
rect 6481 4631 6521 4665
rect 6521 4631 6533 4665
rect 6581 4631 6613 4665
rect 6613 4631 6633 4665
rect 6272 4615 6324 4631
rect 6379 4617 6431 4631
rect 6481 4617 6533 4631
rect 6581 4618 6633 4631
rect 21302 4631 21343 4665
rect 21343 4631 21354 4665
rect 21405 4631 21435 4665
rect 21435 4631 21457 4665
rect 21488 4631 21527 4665
rect 21527 4631 21540 4665
rect 21589 4631 21619 4665
rect 21619 4631 21641 4665
rect 21676 4631 21711 4665
rect 21711 4631 21728 4665
rect 21302 4621 21354 4631
rect 21405 4621 21457 4631
rect 21488 4621 21540 4631
rect 21589 4621 21641 4631
rect 21676 4621 21728 4631
rect 36434 4665 36486 4669
rect 36434 4631 36447 4665
rect 36447 4631 36481 4665
rect 36481 4631 36486 4665
rect 36434 4617 36486 4631
rect 36522 4665 36574 4669
rect 36522 4631 36539 4665
rect 36539 4631 36573 4665
rect 36573 4631 36574 4665
rect 36522 4617 36574 4631
rect 36607 4665 36659 4674
rect 36607 4631 36631 4665
rect 36631 4631 36659 4665
rect 36607 4622 36659 4631
rect 53350 4663 53402 4666
rect 53444 4663 53496 4666
rect 53521 4663 53573 4666
rect 53350 4629 53369 4663
rect 53369 4629 53402 4663
rect 53444 4629 53461 4663
rect 53461 4629 53496 4663
rect 53521 4629 53553 4663
rect 53553 4629 53573 4663
rect 53350 4614 53402 4629
rect 53444 4614 53496 4629
rect 53521 4614 53573 4629
rect 53601 4663 53653 4665
rect 53601 4629 53611 4663
rect 53611 4629 53645 4663
rect 53645 4629 53653 4663
rect 53601 4613 53653 4629
rect 53675 4663 53727 4666
rect 53675 4629 53703 4663
rect 53703 4629 53727 4663
rect 53675 4614 53727 4629
rect 30414 4132 30466 4147
rect 30414 4098 30424 4132
rect 30424 4098 30458 4132
rect 30458 4098 30466 4132
rect 30517 4098 30569 4150
rect 30618 4098 30670 4150
rect 30414 4095 30466 4098
rect 44600 3916 44652 3922
rect 44600 3882 44606 3916
rect 44606 3882 44640 3916
rect 44640 3882 44652 3916
rect 44600 3870 44652 3882
rect 44690 3916 44742 3923
rect 44690 3882 44698 3916
rect 44698 3882 44732 3916
rect 44732 3882 44742 3916
rect 44690 3871 44742 3882
rect 14467 3756 14519 3770
rect 14467 3722 14498 3756
rect 14498 3722 14519 3756
rect 14467 3718 14519 3722
rect 14590 3718 14642 3770
rect 31195 3720 31247 3741
rect 31195 3689 31229 3720
rect 31229 3689 31247 3720
rect 31355 3726 31407 3741
rect 31355 3692 31363 3726
rect 31363 3692 31397 3726
rect 31397 3692 31407 3726
rect 31355 3689 31407 3692
rect 31488 3724 31540 3741
rect 31488 3690 31530 3724
rect 31530 3690 31540 3724
rect 31488 3689 31540 3690
rect 31601 3689 31653 3741
rect 37460 3661 37512 3713
rect 37563 3662 37615 3714
rect 52573 3657 52625 3709
rect 52664 3662 52716 3714
rect 7265 3506 7317 3558
rect 7361 3506 7413 3558
rect 22376 3497 22428 3549
rect 22475 3504 22527 3556
rect 30370 3543 30422 3595
rect 30466 3545 30518 3597
rect 30577 3588 30629 3600
rect 30577 3554 30584 3588
rect 30584 3554 30618 3588
rect 30618 3554 30629 3588
rect 30577 3548 30629 3554
rect 30669 3588 30721 3597
rect 30669 3554 30676 3588
rect 30676 3554 30710 3588
rect 30710 3554 30721 3588
rect 30669 3545 30721 3554
rect 45023 3517 45075 3569
rect 45128 3521 45180 3573
rect 14881 3357 14933 3409
rect 14986 3361 15038 3413
rect 46035 3372 46087 3382
rect 46127 3372 46179 3383
rect 46217 3372 46269 3382
rect 46305 3372 46357 3381
rect 46035 3338 46076 3372
rect 46076 3338 46087 3372
rect 46127 3338 46168 3372
rect 46168 3338 46179 3372
rect 46217 3338 46260 3372
rect 46260 3338 46269 3372
rect 46305 3338 46352 3372
rect 46352 3338 46357 3372
rect 46035 3330 46087 3338
rect 46127 3331 46179 3338
rect 46217 3330 46269 3338
rect 46305 3329 46357 3338
rect 13680 3212 13732 3221
rect 13680 3178 13728 3212
rect 13728 3178 13732 3212
rect 13680 3169 13732 3178
rect 13764 3169 13816 3221
rect 13857 3170 13909 3222
rect 31184 3121 31236 3173
rect 31328 3121 31380 3173
rect 31472 3121 31524 3173
rect 45031 3120 45083 3172
rect 45120 3123 45172 3175
rect 31183 3037 31235 3089
rect 31327 3037 31379 3089
rect 31471 3037 31523 3089
rect 45031 3044 45083 3096
rect 45124 3044 45176 3096
rect 14885 2940 14937 2992
rect 14979 2935 15031 2987
rect 14885 2860 14937 2912
rect 14979 2862 15031 2914
rect 6266 2811 6318 2817
rect 6364 2811 6416 2817
rect 6459 2811 6511 2817
rect 6564 2811 6616 2817
rect 6266 2777 6279 2811
rect 6279 2777 6318 2811
rect 6364 2777 6371 2811
rect 6371 2777 6416 2811
rect 6459 2777 6463 2811
rect 6463 2777 6511 2811
rect 6564 2777 6613 2811
rect 6613 2777 6616 2811
rect 6266 2765 6318 2777
rect 6364 2765 6416 2777
rect 6459 2765 6511 2777
rect 6564 2765 6616 2777
rect 21316 2811 21368 2822
rect 21416 2811 21468 2822
rect 21515 2811 21567 2822
rect 21316 2777 21343 2811
rect 21343 2777 21368 2811
rect 21416 2777 21435 2811
rect 21435 2777 21468 2811
rect 21515 2777 21527 2811
rect 21527 2777 21561 2811
rect 21561 2777 21567 2811
rect 21316 2770 21368 2777
rect 21416 2770 21468 2777
rect 21515 2770 21567 2777
rect 21618 2811 21670 2822
rect 21618 2777 21619 2811
rect 21619 2777 21653 2811
rect 21653 2777 21670 2811
rect 21618 2770 21670 2777
rect 36424 2811 36476 2816
rect 36512 2811 36564 2816
rect 36610 2811 36662 2812
rect 36424 2777 36447 2811
rect 36447 2777 36476 2811
rect 36512 2777 36539 2811
rect 36539 2777 36564 2811
rect 36610 2777 36631 2811
rect 36631 2777 36662 2811
rect 36424 2764 36476 2777
rect 36512 2764 36564 2777
rect 36610 2760 36662 2777
rect 53346 2809 53398 2813
rect 53434 2809 53486 2813
rect 53346 2775 53369 2809
rect 53369 2775 53398 2809
rect 53434 2775 53461 2809
rect 53461 2775 53486 2809
rect 53346 2761 53398 2775
rect 53434 2761 53486 2775
rect 53517 2809 53569 2813
rect 53517 2775 53519 2809
rect 53519 2775 53553 2809
rect 53553 2775 53569 2809
rect 53517 2761 53569 2775
rect 53604 2809 53656 2813
rect 53604 2775 53611 2809
rect 53611 2775 53645 2809
rect 53645 2775 53656 2809
rect 53604 2761 53656 2775
rect 7265 2623 7317 2675
rect 7345 2621 7397 2673
rect 22381 2638 22433 2690
rect 22464 2638 22516 2690
rect 37459 2628 37511 2680
rect 37550 2628 37602 2680
rect 52576 2613 52628 2665
rect 52659 2613 52711 2665
rect 5834 2422 5886 2474
rect 5941 2443 5963 2474
rect 5963 2443 5993 2474
rect 5941 2422 5993 2443
rect 6047 2422 6099 2474
rect 6163 2422 6215 2474
rect 6292 2443 6298 2476
rect 6298 2443 6332 2476
rect 6332 2443 6344 2476
rect 6292 2424 6344 2443
rect 6426 2473 6478 2475
rect 6426 2439 6467 2473
rect 6467 2439 6478 2473
rect 6426 2423 6478 2439
rect 6543 2423 6595 2475
rect 6648 2472 6700 2475
rect 6648 2438 6670 2472
rect 6670 2438 6700 2472
rect 6648 2423 6700 2438
rect 6754 2444 6802 2475
rect 6802 2444 6806 2475
rect 6754 2423 6806 2444
rect 6851 2423 6903 2475
rect 6948 2446 6972 2475
rect 6972 2446 7000 2475
rect 6948 2423 7000 2446
rect 7723 2419 7775 2471
rect 7830 2443 7846 2471
rect 7846 2443 7880 2471
rect 7880 2443 7882 2471
rect 7830 2419 7882 2443
rect 7936 2419 7988 2471
rect 8052 2419 8104 2471
rect 8174 2447 8182 2474
rect 8182 2447 8216 2474
rect 8216 2473 8226 2474
rect 8216 2447 8233 2473
rect 8174 2422 8233 2447
rect 8181 2421 8233 2422
rect 8315 2468 8367 2472
rect 8315 2434 8346 2468
rect 8346 2434 8367 2468
rect 8315 2420 8367 2434
rect 8432 2420 8484 2472
rect 8537 2440 8550 2472
rect 8550 2440 8589 2472
rect 8537 2420 8589 2440
rect 8643 2442 8686 2472
rect 8686 2442 8695 2472
rect 8643 2420 8695 2442
rect 8740 2420 8792 2472
rect 8837 2444 8845 2472
rect 8845 2444 8879 2472
rect 8879 2444 8889 2472
rect 8837 2420 8889 2444
rect 20943 2428 20995 2480
rect 21055 2468 21107 2478
rect 21055 2434 21058 2468
rect 21058 2434 21092 2468
rect 21092 2434 21107 2468
rect 21055 2426 21107 2434
rect 21162 2426 21214 2478
rect 21264 2472 21316 2478
rect 21264 2438 21265 2472
rect 21265 2438 21316 2472
rect 21264 2426 21316 2438
rect 21390 2443 21396 2476
rect 21396 2443 21430 2476
rect 21430 2443 21442 2476
rect 21390 2424 21442 2443
rect 21544 2464 21596 2476
rect 21544 2430 21563 2464
rect 21563 2430 21596 2464
rect 21681 2462 21733 2476
rect 21544 2424 21596 2430
rect 21681 2428 21731 2462
rect 21731 2428 21733 2462
rect 21681 2424 21733 2428
rect 21778 2424 21830 2476
rect 21878 2471 21930 2476
rect 21878 2437 21901 2471
rect 21901 2437 21930 2471
rect 21878 2424 21930 2437
rect 21967 2423 22019 2475
rect 22063 2423 22115 2475
rect 22777 2472 22829 2474
rect 22777 2438 22808 2472
rect 22808 2438 22829 2472
rect 22777 2422 22829 2438
rect 22871 2422 22923 2474
rect 22970 2473 23022 2474
rect 22970 2439 22981 2473
rect 22981 2439 23022 2473
rect 22970 2422 23022 2439
rect 23078 2444 23109 2474
rect 23109 2444 23130 2474
rect 23078 2422 23130 2444
rect 23174 2422 23226 2474
rect 23272 2447 23280 2474
rect 23280 2447 23314 2474
rect 23314 2447 23324 2474
rect 23272 2422 23324 2447
rect 23391 2421 23443 2473
rect 23505 2421 23557 2473
rect 23622 2467 23674 2473
rect 23622 2433 23648 2467
rect 23648 2433 23674 2467
rect 23622 2421 23674 2433
rect 23749 2465 23801 2473
rect 23749 2431 23784 2465
rect 23784 2431 23801 2465
rect 23749 2421 23801 2431
rect 23864 2421 23916 2473
rect 36036 2422 36088 2474
rect 36143 2443 36165 2474
rect 36165 2443 36195 2474
rect 36143 2422 36195 2443
rect 36249 2422 36301 2474
rect 36365 2422 36417 2474
rect 36494 2443 36500 2476
rect 36500 2443 36534 2476
rect 36534 2443 36546 2476
rect 36494 2424 36546 2443
rect 36628 2473 36680 2475
rect 36628 2439 36669 2473
rect 36669 2439 36680 2473
rect 36628 2423 36680 2439
rect 36745 2423 36797 2475
rect 36850 2472 36902 2475
rect 36850 2438 36872 2472
rect 36872 2438 36902 2472
rect 36850 2423 36902 2438
rect 36956 2444 37004 2475
rect 37004 2444 37008 2475
rect 36956 2423 37008 2444
rect 37053 2423 37105 2475
rect 37150 2446 37174 2475
rect 37174 2446 37202 2475
rect 37150 2423 37202 2446
rect 37925 2419 37977 2471
rect 38032 2443 38048 2471
rect 38048 2443 38082 2471
rect 38082 2443 38084 2471
rect 38032 2419 38084 2443
rect 38138 2419 38190 2471
rect 38254 2419 38306 2471
rect 38376 2447 38384 2474
rect 38384 2447 38418 2474
rect 38418 2473 38428 2474
rect 38418 2447 38435 2473
rect 38376 2422 38435 2447
rect 38383 2421 38435 2422
rect 38517 2468 38569 2472
rect 38517 2434 38548 2468
rect 38548 2434 38569 2468
rect 38517 2420 38569 2434
rect 38634 2420 38686 2472
rect 38739 2440 38752 2472
rect 38752 2440 38791 2472
rect 38739 2420 38791 2440
rect 38845 2442 38888 2472
rect 38888 2442 38897 2472
rect 38845 2420 38897 2442
rect 38942 2420 38994 2472
rect 39039 2444 39047 2472
rect 39047 2444 39081 2472
rect 39081 2444 39091 2472
rect 39039 2420 39091 2444
rect 51145 2428 51197 2480
rect 51257 2468 51309 2478
rect 51257 2434 51260 2468
rect 51260 2434 51294 2468
rect 51294 2434 51309 2468
rect 51257 2426 51309 2434
rect 51364 2426 51416 2478
rect 51466 2472 51518 2478
rect 51466 2438 51467 2472
rect 51467 2438 51518 2472
rect 51466 2426 51518 2438
rect 51592 2443 51598 2476
rect 51598 2443 51632 2476
rect 51632 2443 51644 2476
rect 51592 2424 51644 2443
rect 51746 2464 51798 2476
rect 51746 2430 51765 2464
rect 51765 2430 51798 2464
rect 51883 2462 51935 2476
rect 51746 2424 51798 2430
rect 51883 2428 51933 2462
rect 51933 2428 51935 2462
rect 51883 2424 51935 2428
rect 51980 2424 52032 2476
rect 52080 2471 52132 2476
rect 52080 2437 52103 2471
rect 52103 2437 52132 2471
rect 52080 2424 52132 2437
rect 52169 2423 52221 2475
rect 52265 2423 52317 2475
rect 52979 2472 53031 2474
rect 52979 2438 53010 2472
rect 53010 2438 53031 2472
rect 52979 2422 53031 2438
rect 53073 2422 53125 2474
rect 53172 2473 53224 2474
rect 53172 2439 53183 2473
rect 53183 2439 53224 2473
rect 53172 2422 53224 2439
rect 53280 2444 53311 2474
rect 53311 2444 53332 2474
rect 53280 2422 53332 2444
rect 53376 2422 53428 2474
rect 53474 2447 53482 2474
rect 53482 2447 53516 2474
rect 53516 2447 53526 2474
rect 53474 2422 53526 2447
rect 53593 2421 53645 2473
rect 53707 2421 53759 2473
rect 53824 2467 53876 2473
rect 53824 2433 53850 2467
rect 53850 2433 53876 2467
rect 53824 2421 53876 2433
rect 53951 2465 54003 2473
rect 53951 2431 53986 2465
rect 53986 2431 54003 2465
rect 53951 2421 54003 2431
rect 54066 2421 54118 2473
rect 1535 2188 1843 2304
rect 3423 2188 3731 2304
rect 5311 2188 5619 2304
rect 7199 2188 7507 2304
rect 9087 2188 9395 2304
rect 10975 2188 11283 2304
rect 12863 2188 13171 2304
rect 14751 2188 15059 2304
rect 16633 2188 16941 2304
rect 18521 2188 18829 2304
rect 20409 2188 20717 2304
rect 22297 2188 22605 2304
rect 24185 2188 24493 2304
rect 26073 2188 26381 2304
rect 27961 2188 28269 2304
rect 29849 2188 30157 2304
rect 31737 2188 32045 2304
rect 33625 2188 33933 2304
rect 35513 2188 35821 2304
rect 37401 2188 37709 2304
rect 39289 2188 39597 2304
rect 41177 2188 41485 2304
rect 43065 2188 43373 2304
rect 44953 2188 45261 2304
rect 46835 2188 47143 2304
rect 48723 2188 49031 2304
rect 50611 2188 50919 2304
rect 52499 2188 52807 2304
rect 54387 2188 54695 2304
rect 56275 2188 56583 2304
rect 58163 2188 58471 2304
rect 60051 2188 60359 2304
rect 420 1880 472 1888
rect 420 1846 426 1880
rect 426 1846 460 1880
rect 460 1846 472 1880
rect 420 1836 472 1846
rect 692 1911 744 1958
rect 692 1906 702 1911
rect 702 1906 736 1911
rect 736 1906 744 1911
rect 328 1764 380 1776
rect 328 1730 335 1764
rect 335 1730 369 1764
rect 369 1730 380 1764
rect 328 1724 380 1730
rect 1232 1882 1284 1890
rect 1232 1848 1239 1882
rect 1239 1848 1273 1882
rect 1273 1848 1284 1882
rect 1232 1838 1284 1848
rect 1144 1759 1196 1774
rect 1144 1725 1153 1759
rect 1153 1725 1187 1759
rect 1187 1725 1196 1759
rect 1144 1722 1196 1725
rect 206 1489 258 1541
rect 382 1489 434 1541
rect 710 1474 762 1486
rect 710 1440 718 1474
rect 718 1440 752 1474
rect 752 1440 762 1474
rect 710 1434 762 1440
rect 208 1398 260 1408
rect 208 1364 218 1398
rect 218 1364 252 1398
rect 252 1364 260 1398
rect 208 1356 260 1364
rect 232 1133 284 1150
rect 232 1099 253 1133
rect 253 1099 284 1133
rect 232 1098 284 1099
rect 582 1281 634 1292
rect 582 1247 590 1281
rect 590 1247 624 1281
rect 624 1247 634 1281
rect 582 1240 634 1247
rect 478 1015 530 1036
rect 478 984 510 1015
rect 510 984 530 1015
rect 2308 1880 2360 1888
rect 2308 1846 2314 1880
rect 2314 1846 2348 1880
rect 2348 1846 2360 1880
rect 2308 1836 2360 1846
rect 2580 1911 2632 1958
rect 2580 1906 2590 1911
rect 2590 1906 2624 1911
rect 2624 1906 2632 1911
rect 2216 1764 2268 1776
rect 2216 1730 2223 1764
rect 2223 1730 2257 1764
rect 2257 1730 2268 1764
rect 2216 1724 2268 1730
rect 3120 1882 3172 1890
rect 3120 1848 3127 1882
rect 3127 1848 3161 1882
rect 3161 1848 3172 1882
rect 3120 1838 3172 1848
rect 3032 1759 3084 1774
rect 3032 1725 3041 1759
rect 3041 1725 3075 1759
rect 3075 1725 3084 1759
rect 3032 1722 3084 1725
rect 2094 1489 2146 1541
rect 2270 1489 2322 1541
rect 2598 1474 2650 1486
rect 2598 1440 2606 1474
rect 2606 1440 2640 1474
rect 2640 1440 2650 1474
rect 2598 1434 2650 1440
rect 2096 1398 2148 1408
rect 2096 1364 2106 1398
rect 2106 1364 2140 1398
rect 2140 1364 2148 1398
rect 2096 1356 2148 1364
rect 1266 1141 1318 1144
rect 1266 1107 1299 1141
rect 1299 1107 1318 1141
rect 1266 1092 1318 1107
rect 2120 1133 2172 1150
rect 2120 1099 2141 1133
rect 2141 1099 2172 1133
rect 2120 1098 2172 1099
rect 2470 1281 2522 1292
rect 2470 1247 2478 1281
rect 2478 1247 2512 1281
rect 2512 1247 2522 1281
rect 2470 1240 2522 1247
rect 1028 1015 1080 1056
rect 1028 1004 1034 1015
rect 1034 1004 1068 1015
rect 1068 1004 1080 1015
rect 27 792 79 844
rect 690 855 742 902
rect 690 850 700 855
rect 700 850 734 855
rect 734 850 742 855
rect 163 589 215 602
rect 163 555 195 589
rect 195 555 215 589
rect 163 550 215 555
rect 395 584 447 592
rect 395 550 404 584
rect 404 550 438 584
rect 438 550 447 584
rect 395 540 447 550
rect 708 418 760 430
rect 708 384 716 418
rect 716 384 750 418
rect 750 384 760 418
rect 708 378 760 384
rect 2366 1015 2418 1036
rect 2366 984 2398 1015
rect 2398 984 2418 1015
rect 4196 1880 4248 1888
rect 4196 1846 4202 1880
rect 4202 1846 4236 1880
rect 4236 1846 4248 1880
rect 4196 1836 4248 1846
rect 4468 1911 4520 1958
rect 4468 1906 4478 1911
rect 4478 1906 4512 1911
rect 4512 1906 4520 1911
rect 4104 1764 4156 1776
rect 4104 1730 4111 1764
rect 4111 1730 4145 1764
rect 4145 1730 4156 1764
rect 4104 1724 4156 1730
rect 5008 1882 5060 1890
rect 5008 1848 5015 1882
rect 5015 1848 5049 1882
rect 5049 1848 5060 1882
rect 5008 1838 5060 1848
rect 4920 1759 4972 1774
rect 4920 1725 4929 1759
rect 4929 1725 4963 1759
rect 4963 1725 4972 1759
rect 4920 1722 4972 1725
rect 3982 1489 4034 1541
rect 4158 1489 4210 1541
rect 4486 1474 4538 1486
rect 4486 1440 4494 1474
rect 4494 1440 4528 1474
rect 4528 1440 4538 1474
rect 4486 1434 4538 1440
rect 3984 1398 4036 1408
rect 3984 1364 3994 1398
rect 3994 1364 4028 1398
rect 4028 1364 4036 1398
rect 3984 1356 4036 1364
rect 3154 1141 3206 1144
rect 3154 1107 3187 1141
rect 3187 1107 3206 1141
rect 3154 1092 3206 1107
rect 4008 1133 4060 1150
rect 4008 1099 4029 1133
rect 4029 1099 4060 1133
rect 4008 1098 4060 1099
rect 4358 1281 4410 1292
rect 4358 1247 4366 1281
rect 4366 1247 4400 1281
rect 4400 1247 4410 1281
rect 4358 1240 4410 1247
rect 2916 1015 2968 1056
rect 2916 1004 2922 1015
rect 2922 1004 2956 1015
rect 2956 1004 2968 1015
rect 1611 826 1663 840
rect 1611 792 1617 826
rect 1617 792 1651 826
rect 1651 792 1663 826
rect 1611 788 1663 792
rect 1915 792 1967 844
rect 2578 855 2630 902
rect 2578 850 2588 855
rect 2588 850 2622 855
rect 2622 850 2630 855
rect 1028 612 1080 624
rect 1028 578 1036 612
rect 1036 578 1070 612
rect 1070 578 1080 612
rect 1028 572 1080 578
rect 2051 589 2103 602
rect 2051 555 2083 589
rect 2083 555 2103 589
rect 2051 550 2103 555
rect 2283 584 2335 592
rect 2283 550 2292 584
rect 2292 550 2326 584
rect 2326 550 2335 584
rect 2283 540 2335 550
rect 2596 418 2648 430
rect 2596 384 2604 418
rect 2604 384 2638 418
rect 2638 384 2648 418
rect 2596 378 2648 384
rect 4254 1015 4306 1036
rect 4254 984 4286 1015
rect 4286 984 4306 1015
rect 6084 1880 6136 1888
rect 6084 1846 6090 1880
rect 6090 1846 6124 1880
rect 6124 1846 6136 1880
rect 6084 1836 6136 1846
rect 6356 1911 6408 1958
rect 6356 1906 6366 1911
rect 6366 1906 6400 1911
rect 6400 1906 6408 1911
rect 5992 1764 6044 1776
rect 5992 1730 5999 1764
rect 5999 1730 6033 1764
rect 6033 1730 6044 1764
rect 5992 1724 6044 1730
rect 6896 1882 6948 1890
rect 6896 1848 6903 1882
rect 6903 1848 6937 1882
rect 6937 1848 6948 1882
rect 6896 1838 6948 1848
rect 6808 1759 6860 1774
rect 6808 1725 6817 1759
rect 6817 1725 6851 1759
rect 6851 1725 6860 1759
rect 6808 1722 6860 1725
rect 5870 1489 5922 1541
rect 6046 1489 6098 1541
rect 6374 1474 6426 1486
rect 6374 1440 6382 1474
rect 6382 1440 6416 1474
rect 6416 1440 6426 1474
rect 6374 1434 6426 1440
rect 5872 1398 5924 1408
rect 5872 1364 5882 1398
rect 5882 1364 5916 1398
rect 5916 1364 5924 1398
rect 5872 1356 5924 1364
rect 5042 1141 5094 1144
rect 5042 1107 5075 1141
rect 5075 1107 5094 1141
rect 5042 1092 5094 1107
rect 5896 1133 5948 1150
rect 5896 1099 5917 1133
rect 5917 1099 5948 1133
rect 5896 1098 5948 1099
rect 6246 1281 6298 1292
rect 6246 1247 6254 1281
rect 6254 1247 6288 1281
rect 6288 1247 6298 1281
rect 6246 1240 6298 1247
rect 4804 1015 4856 1056
rect 4804 1004 4810 1015
rect 4810 1004 4844 1015
rect 4844 1004 4856 1015
rect 3499 826 3551 840
rect 3499 792 3505 826
rect 3505 792 3539 826
rect 3539 792 3551 826
rect 3499 788 3551 792
rect 3803 792 3855 844
rect 4466 855 4518 902
rect 4466 850 4476 855
rect 4476 850 4510 855
rect 4510 850 4518 855
rect 2916 612 2968 624
rect 2916 578 2924 612
rect 2924 578 2958 612
rect 2958 578 2968 612
rect 2916 572 2968 578
rect 3939 589 3991 602
rect 3939 555 3971 589
rect 3971 555 3991 589
rect 3939 550 3991 555
rect 4171 584 4223 592
rect 4171 550 4180 584
rect 4180 550 4214 584
rect 4214 550 4223 584
rect 4171 540 4223 550
rect 4484 418 4536 430
rect 4484 384 4492 418
rect 4492 384 4526 418
rect 4526 384 4536 418
rect 4484 378 4536 384
rect 6142 1015 6194 1036
rect 6142 984 6174 1015
rect 6174 984 6194 1015
rect 7972 1880 8024 1888
rect 7972 1846 7978 1880
rect 7978 1846 8012 1880
rect 8012 1846 8024 1880
rect 7972 1836 8024 1846
rect 8244 1911 8296 1958
rect 8244 1906 8254 1911
rect 8254 1906 8288 1911
rect 8288 1906 8296 1911
rect 7880 1764 7932 1776
rect 7880 1730 7887 1764
rect 7887 1730 7921 1764
rect 7921 1730 7932 1764
rect 7880 1724 7932 1730
rect 8784 1882 8836 1890
rect 8784 1848 8791 1882
rect 8791 1848 8825 1882
rect 8825 1848 8836 1882
rect 8784 1838 8836 1848
rect 8696 1759 8748 1774
rect 8696 1725 8705 1759
rect 8705 1725 8739 1759
rect 8739 1725 8748 1759
rect 8696 1722 8748 1725
rect 7758 1489 7810 1541
rect 7934 1489 7986 1541
rect 8262 1474 8314 1486
rect 8262 1440 8270 1474
rect 8270 1440 8304 1474
rect 8304 1440 8314 1474
rect 8262 1434 8314 1440
rect 7760 1398 7812 1408
rect 7760 1364 7770 1398
rect 7770 1364 7804 1398
rect 7804 1364 7812 1398
rect 7760 1356 7812 1364
rect 6930 1141 6982 1144
rect 6930 1107 6963 1141
rect 6963 1107 6982 1141
rect 6930 1092 6982 1107
rect 7784 1133 7836 1150
rect 7784 1099 7805 1133
rect 7805 1099 7836 1133
rect 7784 1098 7836 1099
rect 8134 1281 8186 1292
rect 8134 1247 8142 1281
rect 8142 1247 8176 1281
rect 8176 1247 8186 1281
rect 8134 1240 8186 1247
rect 6692 1015 6744 1056
rect 6692 1004 6698 1015
rect 6698 1004 6732 1015
rect 6732 1004 6744 1015
rect 5387 826 5439 840
rect 5387 792 5393 826
rect 5393 792 5427 826
rect 5427 792 5439 826
rect 5387 788 5439 792
rect 5691 792 5743 844
rect 6354 855 6406 902
rect 6354 850 6364 855
rect 6364 850 6398 855
rect 6398 850 6406 855
rect 4804 612 4856 624
rect 4804 578 4812 612
rect 4812 578 4846 612
rect 4846 578 4856 612
rect 4804 572 4856 578
rect 5827 589 5879 602
rect 5827 555 5859 589
rect 5859 555 5879 589
rect 5827 550 5879 555
rect 6059 584 6111 592
rect 6059 550 6068 584
rect 6068 550 6102 584
rect 6102 550 6111 584
rect 6059 540 6111 550
rect 6372 418 6424 430
rect 6372 384 6380 418
rect 6380 384 6414 418
rect 6414 384 6424 418
rect 6372 378 6424 384
rect 8030 1015 8082 1036
rect 8030 984 8062 1015
rect 8062 984 8082 1015
rect 9860 1880 9912 1888
rect 9860 1846 9866 1880
rect 9866 1846 9900 1880
rect 9900 1846 9912 1880
rect 9860 1836 9912 1846
rect 10132 1911 10184 1958
rect 10132 1906 10142 1911
rect 10142 1906 10176 1911
rect 10176 1906 10184 1911
rect 9768 1764 9820 1776
rect 9768 1730 9775 1764
rect 9775 1730 9809 1764
rect 9809 1730 9820 1764
rect 9768 1724 9820 1730
rect 10672 1882 10724 1890
rect 10672 1848 10679 1882
rect 10679 1848 10713 1882
rect 10713 1848 10724 1882
rect 10672 1838 10724 1848
rect 10584 1759 10636 1774
rect 10584 1725 10593 1759
rect 10593 1725 10627 1759
rect 10627 1725 10636 1759
rect 10584 1722 10636 1725
rect 9646 1489 9698 1541
rect 9822 1489 9874 1541
rect 10150 1474 10202 1486
rect 10150 1440 10158 1474
rect 10158 1440 10192 1474
rect 10192 1440 10202 1474
rect 10150 1434 10202 1440
rect 9648 1398 9700 1408
rect 9648 1364 9658 1398
rect 9658 1364 9692 1398
rect 9692 1364 9700 1398
rect 9648 1356 9700 1364
rect 8818 1141 8870 1144
rect 8818 1107 8851 1141
rect 8851 1107 8870 1141
rect 8818 1092 8870 1107
rect 9672 1133 9724 1150
rect 9672 1099 9693 1133
rect 9693 1099 9724 1133
rect 9672 1098 9724 1099
rect 10022 1281 10074 1292
rect 10022 1247 10030 1281
rect 10030 1247 10064 1281
rect 10064 1247 10074 1281
rect 10022 1240 10074 1247
rect 8580 1015 8632 1056
rect 8580 1004 8586 1015
rect 8586 1004 8620 1015
rect 8620 1004 8632 1015
rect 7275 826 7327 840
rect 7275 792 7281 826
rect 7281 792 7315 826
rect 7315 792 7327 826
rect 7275 788 7327 792
rect 7579 792 7631 844
rect 8242 855 8294 902
rect 8242 850 8252 855
rect 8252 850 8286 855
rect 8286 850 8294 855
rect 6692 612 6744 624
rect 6692 578 6700 612
rect 6700 578 6734 612
rect 6734 578 6744 612
rect 6692 572 6744 578
rect 7715 589 7767 602
rect 7715 555 7747 589
rect 7747 555 7767 589
rect 7715 550 7767 555
rect 7947 584 7999 592
rect 7947 550 7956 584
rect 7956 550 7990 584
rect 7990 550 7999 584
rect 7947 540 7999 550
rect 8260 418 8312 430
rect 8260 384 8268 418
rect 8268 384 8302 418
rect 8302 384 8312 418
rect 8260 378 8312 384
rect 9918 1015 9970 1036
rect 9918 984 9950 1015
rect 9950 984 9970 1015
rect 11748 1880 11800 1888
rect 11748 1846 11754 1880
rect 11754 1846 11788 1880
rect 11788 1846 11800 1880
rect 11748 1836 11800 1846
rect 12020 1911 12072 1958
rect 12020 1906 12030 1911
rect 12030 1906 12064 1911
rect 12064 1906 12072 1911
rect 11656 1764 11708 1776
rect 11656 1730 11663 1764
rect 11663 1730 11697 1764
rect 11697 1730 11708 1764
rect 11656 1724 11708 1730
rect 12560 1882 12612 1890
rect 12560 1848 12567 1882
rect 12567 1848 12601 1882
rect 12601 1848 12612 1882
rect 12560 1838 12612 1848
rect 12472 1759 12524 1774
rect 12472 1725 12481 1759
rect 12481 1725 12515 1759
rect 12515 1725 12524 1759
rect 12472 1722 12524 1725
rect 11534 1489 11586 1541
rect 11710 1489 11762 1541
rect 12038 1474 12090 1486
rect 12038 1440 12046 1474
rect 12046 1440 12080 1474
rect 12080 1440 12090 1474
rect 12038 1434 12090 1440
rect 11536 1398 11588 1408
rect 11536 1364 11546 1398
rect 11546 1364 11580 1398
rect 11580 1364 11588 1398
rect 11536 1356 11588 1364
rect 10706 1141 10758 1144
rect 10706 1107 10739 1141
rect 10739 1107 10758 1141
rect 10706 1092 10758 1107
rect 11560 1133 11612 1150
rect 11560 1099 11581 1133
rect 11581 1099 11612 1133
rect 11560 1098 11612 1099
rect 11910 1281 11962 1292
rect 11910 1247 11918 1281
rect 11918 1247 11952 1281
rect 11952 1247 11962 1281
rect 11910 1240 11962 1247
rect 10468 1015 10520 1056
rect 10468 1004 10474 1015
rect 10474 1004 10508 1015
rect 10508 1004 10520 1015
rect 9163 826 9215 840
rect 9163 792 9169 826
rect 9169 792 9203 826
rect 9203 792 9215 826
rect 9163 788 9215 792
rect 9467 792 9519 844
rect 10130 855 10182 902
rect 10130 850 10140 855
rect 10140 850 10174 855
rect 10174 850 10182 855
rect 8580 612 8632 624
rect 8580 578 8588 612
rect 8588 578 8622 612
rect 8622 578 8632 612
rect 8580 572 8632 578
rect 9603 589 9655 602
rect 9603 555 9635 589
rect 9635 555 9655 589
rect 9603 550 9655 555
rect 9835 584 9887 592
rect 9835 550 9844 584
rect 9844 550 9878 584
rect 9878 550 9887 584
rect 9835 540 9887 550
rect 10148 418 10200 430
rect 10148 384 10156 418
rect 10156 384 10190 418
rect 10190 384 10200 418
rect 10148 378 10200 384
rect 11806 1015 11858 1036
rect 11806 984 11838 1015
rect 11838 984 11858 1015
rect 13636 1880 13688 1888
rect 13636 1846 13642 1880
rect 13642 1846 13676 1880
rect 13676 1846 13688 1880
rect 13636 1836 13688 1846
rect 13908 1911 13960 1958
rect 13908 1906 13918 1911
rect 13918 1906 13952 1911
rect 13952 1906 13960 1911
rect 13544 1764 13596 1776
rect 13544 1730 13551 1764
rect 13551 1730 13585 1764
rect 13585 1730 13596 1764
rect 13544 1724 13596 1730
rect 14448 1882 14500 1890
rect 14448 1848 14455 1882
rect 14455 1848 14489 1882
rect 14489 1848 14500 1882
rect 14448 1838 14500 1848
rect 14360 1759 14412 1774
rect 14360 1725 14369 1759
rect 14369 1725 14403 1759
rect 14403 1725 14412 1759
rect 14360 1722 14412 1725
rect 13422 1489 13474 1541
rect 13598 1489 13650 1541
rect 13926 1474 13978 1486
rect 13926 1440 13934 1474
rect 13934 1440 13968 1474
rect 13968 1440 13978 1474
rect 13926 1434 13978 1440
rect 13424 1398 13476 1408
rect 13424 1364 13434 1398
rect 13434 1364 13468 1398
rect 13468 1364 13476 1398
rect 13424 1356 13476 1364
rect 12594 1141 12646 1144
rect 12594 1107 12627 1141
rect 12627 1107 12646 1141
rect 12594 1092 12646 1107
rect 13448 1133 13500 1150
rect 13448 1099 13469 1133
rect 13469 1099 13500 1133
rect 13448 1098 13500 1099
rect 13798 1281 13850 1292
rect 13798 1247 13806 1281
rect 13806 1247 13840 1281
rect 13840 1247 13850 1281
rect 13798 1240 13850 1247
rect 12356 1015 12408 1056
rect 12356 1004 12362 1015
rect 12362 1004 12396 1015
rect 12396 1004 12408 1015
rect 11051 826 11103 840
rect 11051 792 11057 826
rect 11057 792 11091 826
rect 11091 792 11103 826
rect 11051 788 11103 792
rect 11355 792 11407 844
rect 12018 855 12070 902
rect 12018 850 12028 855
rect 12028 850 12062 855
rect 12062 850 12070 855
rect 10468 612 10520 624
rect 10468 578 10476 612
rect 10476 578 10510 612
rect 10510 578 10520 612
rect 10468 572 10520 578
rect 11491 589 11543 602
rect 11491 555 11523 589
rect 11523 555 11543 589
rect 11491 550 11543 555
rect 11723 584 11775 592
rect 11723 550 11732 584
rect 11732 550 11766 584
rect 11766 550 11775 584
rect 11723 540 11775 550
rect 12036 418 12088 430
rect 12036 384 12044 418
rect 12044 384 12078 418
rect 12078 384 12088 418
rect 12036 378 12088 384
rect 13694 1015 13746 1036
rect 13694 984 13726 1015
rect 13726 984 13746 1015
rect 15518 1880 15570 1888
rect 15518 1846 15524 1880
rect 15524 1846 15558 1880
rect 15558 1846 15570 1880
rect 15518 1836 15570 1846
rect 15790 1911 15842 1958
rect 15790 1906 15800 1911
rect 15800 1906 15834 1911
rect 15834 1906 15842 1911
rect 15426 1764 15478 1776
rect 15426 1730 15433 1764
rect 15433 1730 15467 1764
rect 15467 1730 15478 1764
rect 15426 1724 15478 1730
rect 16330 1882 16382 1890
rect 16330 1848 16337 1882
rect 16337 1848 16371 1882
rect 16371 1848 16382 1882
rect 16330 1838 16382 1848
rect 16242 1759 16294 1774
rect 16242 1725 16251 1759
rect 16251 1725 16285 1759
rect 16285 1725 16294 1759
rect 16242 1722 16294 1725
rect 15304 1489 15356 1541
rect 15480 1489 15532 1541
rect 15808 1474 15860 1486
rect 15808 1440 15816 1474
rect 15816 1440 15850 1474
rect 15850 1440 15860 1474
rect 15808 1434 15860 1440
rect 15306 1398 15358 1408
rect 15306 1364 15316 1398
rect 15316 1364 15350 1398
rect 15350 1364 15358 1398
rect 15306 1356 15358 1364
rect 14482 1141 14534 1144
rect 14482 1107 14515 1141
rect 14515 1107 14534 1141
rect 14482 1092 14534 1107
rect 15330 1133 15382 1150
rect 15330 1099 15351 1133
rect 15351 1099 15382 1133
rect 15330 1098 15382 1099
rect 15680 1281 15732 1292
rect 15680 1247 15688 1281
rect 15688 1247 15722 1281
rect 15722 1247 15732 1281
rect 15680 1240 15732 1247
rect 14244 1015 14296 1056
rect 14244 1004 14250 1015
rect 14250 1004 14284 1015
rect 14284 1004 14296 1015
rect 12939 826 12991 840
rect 12939 792 12945 826
rect 12945 792 12979 826
rect 12979 792 12991 826
rect 12939 788 12991 792
rect 13243 792 13295 844
rect 13906 855 13958 902
rect 13906 850 13916 855
rect 13916 850 13950 855
rect 13950 850 13958 855
rect 12356 612 12408 624
rect 12356 578 12364 612
rect 12364 578 12398 612
rect 12398 578 12408 612
rect 12356 572 12408 578
rect 13379 589 13431 602
rect 13379 555 13411 589
rect 13411 555 13431 589
rect 13379 550 13431 555
rect 13611 584 13663 592
rect 13611 550 13620 584
rect 13620 550 13654 584
rect 13654 550 13663 584
rect 13611 540 13663 550
rect 13924 418 13976 430
rect 13924 384 13932 418
rect 13932 384 13966 418
rect 13966 384 13976 418
rect 13924 378 13976 384
rect 15576 1015 15628 1036
rect 15576 984 15608 1015
rect 15608 984 15628 1015
rect 17406 1880 17458 1888
rect 17406 1846 17412 1880
rect 17412 1846 17446 1880
rect 17446 1846 17458 1880
rect 17406 1836 17458 1846
rect 17678 1911 17730 1958
rect 17678 1906 17688 1911
rect 17688 1906 17722 1911
rect 17722 1906 17730 1911
rect 17314 1764 17366 1776
rect 17314 1730 17321 1764
rect 17321 1730 17355 1764
rect 17355 1730 17366 1764
rect 17314 1724 17366 1730
rect 18218 1882 18270 1890
rect 18218 1848 18225 1882
rect 18225 1848 18259 1882
rect 18259 1848 18270 1882
rect 18218 1838 18270 1848
rect 18130 1759 18182 1774
rect 18130 1725 18139 1759
rect 18139 1725 18173 1759
rect 18173 1725 18182 1759
rect 18130 1722 18182 1725
rect 17192 1489 17244 1541
rect 17368 1489 17420 1541
rect 17696 1474 17748 1486
rect 17696 1440 17704 1474
rect 17704 1440 17738 1474
rect 17738 1440 17748 1474
rect 17696 1434 17748 1440
rect 17194 1398 17246 1408
rect 17194 1364 17204 1398
rect 17204 1364 17238 1398
rect 17238 1364 17246 1398
rect 17194 1356 17246 1364
rect 16364 1141 16416 1144
rect 16364 1107 16397 1141
rect 16397 1107 16416 1141
rect 16364 1092 16416 1107
rect 17218 1133 17270 1150
rect 17218 1099 17239 1133
rect 17239 1099 17270 1133
rect 17218 1098 17270 1099
rect 17568 1281 17620 1292
rect 17568 1247 17576 1281
rect 17576 1247 17610 1281
rect 17610 1247 17620 1281
rect 17568 1240 17620 1247
rect 16126 1015 16178 1056
rect 16126 1004 16132 1015
rect 16132 1004 16166 1015
rect 16166 1004 16178 1015
rect 14827 826 14879 840
rect 14827 792 14833 826
rect 14833 792 14867 826
rect 14867 792 14879 826
rect 14827 788 14879 792
rect 15125 792 15177 844
rect 15788 855 15840 902
rect 15788 850 15798 855
rect 15798 850 15832 855
rect 15832 850 15840 855
rect 14244 612 14296 624
rect 14244 578 14252 612
rect 14252 578 14286 612
rect 14286 578 14296 612
rect 14244 572 14296 578
rect 15261 589 15313 602
rect 15261 555 15293 589
rect 15293 555 15313 589
rect 15261 550 15313 555
rect 15493 584 15545 592
rect 15493 550 15502 584
rect 15502 550 15536 584
rect 15536 550 15545 584
rect 15493 540 15545 550
rect 15806 418 15858 430
rect 15806 384 15814 418
rect 15814 384 15848 418
rect 15848 384 15858 418
rect 15806 378 15858 384
rect 17464 1015 17516 1036
rect 17464 984 17496 1015
rect 17496 984 17516 1015
rect 19294 1880 19346 1888
rect 19294 1846 19300 1880
rect 19300 1846 19334 1880
rect 19334 1846 19346 1880
rect 19294 1836 19346 1846
rect 19566 1911 19618 1958
rect 19566 1906 19576 1911
rect 19576 1906 19610 1911
rect 19610 1906 19618 1911
rect 19202 1764 19254 1776
rect 19202 1730 19209 1764
rect 19209 1730 19243 1764
rect 19243 1730 19254 1764
rect 19202 1724 19254 1730
rect 20106 1882 20158 1890
rect 20106 1848 20113 1882
rect 20113 1848 20147 1882
rect 20147 1848 20158 1882
rect 20106 1838 20158 1848
rect 20018 1759 20070 1774
rect 20018 1725 20027 1759
rect 20027 1725 20061 1759
rect 20061 1725 20070 1759
rect 20018 1722 20070 1725
rect 19080 1489 19132 1541
rect 19256 1489 19308 1541
rect 19584 1474 19636 1486
rect 19584 1440 19592 1474
rect 19592 1440 19626 1474
rect 19626 1440 19636 1474
rect 19584 1434 19636 1440
rect 19082 1398 19134 1408
rect 19082 1364 19092 1398
rect 19092 1364 19126 1398
rect 19126 1364 19134 1398
rect 19082 1356 19134 1364
rect 18252 1141 18304 1144
rect 18252 1107 18285 1141
rect 18285 1107 18304 1141
rect 18252 1092 18304 1107
rect 19106 1133 19158 1150
rect 19106 1099 19127 1133
rect 19127 1099 19158 1133
rect 19106 1098 19158 1099
rect 19456 1281 19508 1292
rect 19456 1247 19464 1281
rect 19464 1247 19498 1281
rect 19498 1247 19508 1281
rect 19456 1240 19508 1247
rect 18014 1015 18066 1056
rect 18014 1004 18020 1015
rect 18020 1004 18054 1015
rect 18054 1004 18066 1015
rect 16709 826 16761 840
rect 16709 792 16715 826
rect 16715 792 16749 826
rect 16749 792 16761 826
rect 16709 788 16761 792
rect 17013 792 17065 844
rect 17676 855 17728 902
rect 17676 850 17686 855
rect 17686 850 17720 855
rect 17720 850 17728 855
rect 16126 612 16178 624
rect 16126 578 16134 612
rect 16134 578 16168 612
rect 16168 578 16178 612
rect 16126 572 16178 578
rect 17149 589 17201 602
rect 17149 555 17181 589
rect 17181 555 17201 589
rect 17149 550 17201 555
rect 17381 584 17433 592
rect 17381 550 17390 584
rect 17390 550 17424 584
rect 17424 550 17433 584
rect 17381 540 17433 550
rect 17694 418 17746 430
rect 17694 384 17702 418
rect 17702 384 17736 418
rect 17736 384 17746 418
rect 17694 378 17746 384
rect 19352 1015 19404 1036
rect 19352 984 19384 1015
rect 19384 984 19404 1015
rect 21182 1880 21234 1888
rect 21182 1846 21188 1880
rect 21188 1846 21222 1880
rect 21222 1846 21234 1880
rect 21182 1836 21234 1846
rect 21454 1911 21506 1958
rect 21454 1906 21464 1911
rect 21464 1906 21498 1911
rect 21498 1906 21506 1911
rect 21090 1764 21142 1776
rect 21090 1730 21097 1764
rect 21097 1730 21131 1764
rect 21131 1730 21142 1764
rect 21090 1724 21142 1730
rect 21994 1882 22046 1890
rect 21994 1848 22001 1882
rect 22001 1848 22035 1882
rect 22035 1848 22046 1882
rect 21994 1838 22046 1848
rect 21906 1759 21958 1774
rect 21906 1725 21915 1759
rect 21915 1725 21949 1759
rect 21949 1725 21958 1759
rect 21906 1722 21958 1725
rect 20968 1489 21020 1541
rect 21144 1489 21196 1541
rect 21472 1474 21524 1486
rect 21472 1440 21480 1474
rect 21480 1440 21514 1474
rect 21514 1440 21524 1474
rect 21472 1434 21524 1440
rect 20970 1398 21022 1408
rect 20970 1364 20980 1398
rect 20980 1364 21014 1398
rect 21014 1364 21022 1398
rect 20970 1356 21022 1364
rect 20140 1141 20192 1144
rect 20140 1107 20173 1141
rect 20173 1107 20192 1141
rect 20140 1092 20192 1107
rect 20994 1133 21046 1150
rect 20994 1099 21015 1133
rect 21015 1099 21046 1133
rect 20994 1098 21046 1099
rect 21344 1281 21396 1292
rect 21344 1247 21352 1281
rect 21352 1247 21386 1281
rect 21386 1247 21396 1281
rect 21344 1240 21396 1247
rect 19902 1015 19954 1056
rect 19902 1004 19908 1015
rect 19908 1004 19942 1015
rect 19942 1004 19954 1015
rect 18597 826 18649 840
rect 18597 792 18603 826
rect 18603 792 18637 826
rect 18637 792 18649 826
rect 18597 788 18649 792
rect 18901 792 18953 844
rect 19564 855 19616 902
rect 19564 850 19574 855
rect 19574 850 19608 855
rect 19608 850 19616 855
rect 18014 612 18066 624
rect 18014 578 18022 612
rect 18022 578 18056 612
rect 18056 578 18066 612
rect 18014 572 18066 578
rect 19037 589 19089 602
rect 19037 555 19069 589
rect 19069 555 19089 589
rect 19037 550 19089 555
rect 19269 584 19321 592
rect 19269 550 19278 584
rect 19278 550 19312 584
rect 19312 550 19321 584
rect 19269 540 19321 550
rect 19582 418 19634 430
rect 19582 384 19590 418
rect 19590 384 19624 418
rect 19624 384 19634 418
rect 19582 378 19634 384
rect 21240 1015 21292 1036
rect 21240 984 21272 1015
rect 21272 984 21292 1015
rect 23070 1880 23122 1888
rect 23070 1846 23076 1880
rect 23076 1846 23110 1880
rect 23110 1846 23122 1880
rect 23070 1836 23122 1846
rect 23342 1911 23394 1958
rect 23342 1906 23352 1911
rect 23352 1906 23386 1911
rect 23386 1906 23394 1911
rect 22978 1764 23030 1776
rect 22978 1730 22985 1764
rect 22985 1730 23019 1764
rect 23019 1730 23030 1764
rect 22978 1724 23030 1730
rect 23882 1882 23934 1890
rect 23882 1848 23889 1882
rect 23889 1848 23923 1882
rect 23923 1848 23934 1882
rect 23882 1838 23934 1848
rect 23794 1759 23846 1774
rect 23794 1725 23803 1759
rect 23803 1725 23837 1759
rect 23837 1725 23846 1759
rect 23794 1722 23846 1725
rect 22856 1489 22908 1541
rect 23032 1489 23084 1541
rect 23360 1474 23412 1486
rect 23360 1440 23368 1474
rect 23368 1440 23402 1474
rect 23402 1440 23412 1474
rect 23360 1434 23412 1440
rect 22858 1398 22910 1408
rect 22858 1364 22868 1398
rect 22868 1364 22902 1398
rect 22902 1364 22910 1398
rect 22858 1356 22910 1364
rect 22028 1141 22080 1144
rect 22028 1107 22061 1141
rect 22061 1107 22080 1141
rect 22028 1092 22080 1107
rect 22882 1133 22934 1150
rect 22882 1099 22903 1133
rect 22903 1099 22934 1133
rect 22882 1098 22934 1099
rect 23232 1281 23284 1292
rect 23232 1247 23240 1281
rect 23240 1247 23274 1281
rect 23274 1247 23284 1281
rect 23232 1240 23284 1247
rect 21790 1015 21842 1056
rect 21790 1004 21796 1015
rect 21796 1004 21830 1015
rect 21830 1004 21842 1015
rect 20485 826 20537 840
rect 20485 792 20491 826
rect 20491 792 20525 826
rect 20525 792 20537 826
rect 20485 788 20537 792
rect 20789 792 20841 844
rect 21452 855 21504 902
rect 21452 850 21462 855
rect 21462 850 21496 855
rect 21496 850 21504 855
rect 19902 612 19954 624
rect 19902 578 19910 612
rect 19910 578 19944 612
rect 19944 578 19954 612
rect 19902 572 19954 578
rect 20925 589 20977 602
rect 20925 555 20957 589
rect 20957 555 20977 589
rect 20925 550 20977 555
rect 21157 584 21209 592
rect 21157 550 21166 584
rect 21166 550 21200 584
rect 21200 550 21209 584
rect 21157 540 21209 550
rect 21470 418 21522 430
rect 21470 384 21478 418
rect 21478 384 21512 418
rect 21512 384 21522 418
rect 21470 378 21522 384
rect 23128 1015 23180 1036
rect 23128 984 23160 1015
rect 23160 984 23180 1015
rect 24958 1880 25010 1888
rect 24958 1846 24964 1880
rect 24964 1846 24998 1880
rect 24998 1846 25010 1880
rect 24958 1836 25010 1846
rect 25230 1911 25282 1958
rect 25230 1906 25240 1911
rect 25240 1906 25274 1911
rect 25274 1906 25282 1911
rect 24866 1764 24918 1776
rect 24866 1730 24873 1764
rect 24873 1730 24907 1764
rect 24907 1730 24918 1764
rect 24866 1724 24918 1730
rect 25770 1882 25822 1890
rect 25770 1848 25777 1882
rect 25777 1848 25811 1882
rect 25811 1848 25822 1882
rect 25770 1838 25822 1848
rect 25682 1759 25734 1774
rect 25682 1725 25691 1759
rect 25691 1725 25725 1759
rect 25725 1725 25734 1759
rect 25682 1722 25734 1725
rect 24744 1489 24796 1541
rect 24920 1489 24972 1541
rect 25248 1474 25300 1486
rect 25248 1440 25256 1474
rect 25256 1440 25290 1474
rect 25290 1440 25300 1474
rect 25248 1434 25300 1440
rect 24746 1398 24798 1408
rect 24746 1364 24756 1398
rect 24756 1364 24790 1398
rect 24790 1364 24798 1398
rect 24746 1356 24798 1364
rect 23916 1141 23968 1144
rect 23916 1107 23949 1141
rect 23949 1107 23968 1141
rect 23916 1092 23968 1107
rect 24770 1133 24822 1150
rect 24770 1099 24791 1133
rect 24791 1099 24822 1133
rect 24770 1098 24822 1099
rect 25120 1281 25172 1292
rect 25120 1247 25128 1281
rect 25128 1247 25162 1281
rect 25162 1247 25172 1281
rect 25120 1240 25172 1247
rect 23678 1015 23730 1056
rect 23678 1004 23684 1015
rect 23684 1004 23718 1015
rect 23718 1004 23730 1015
rect 22373 826 22425 840
rect 22373 792 22379 826
rect 22379 792 22413 826
rect 22413 792 22425 826
rect 22373 788 22425 792
rect 22677 792 22729 844
rect 23340 855 23392 902
rect 23340 850 23350 855
rect 23350 850 23384 855
rect 23384 850 23392 855
rect 21790 612 21842 624
rect 21790 578 21798 612
rect 21798 578 21832 612
rect 21832 578 21842 612
rect 21790 572 21842 578
rect 22813 589 22865 602
rect 22813 555 22845 589
rect 22845 555 22865 589
rect 22813 550 22865 555
rect 23045 584 23097 592
rect 23045 550 23054 584
rect 23054 550 23088 584
rect 23088 550 23097 584
rect 23045 540 23097 550
rect 23358 418 23410 430
rect 23358 384 23366 418
rect 23366 384 23400 418
rect 23400 384 23410 418
rect 23358 378 23410 384
rect 25016 1015 25068 1036
rect 25016 984 25048 1015
rect 25048 984 25068 1015
rect 26846 1880 26898 1888
rect 26846 1846 26852 1880
rect 26852 1846 26886 1880
rect 26886 1846 26898 1880
rect 26846 1836 26898 1846
rect 27118 1911 27170 1958
rect 27118 1906 27128 1911
rect 27128 1906 27162 1911
rect 27162 1906 27170 1911
rect 26754 1764 26806 1776
rect 26754 1730 26761 1764
rect 26761 1730 26795 1764
rect 26795 1730 26806 1764
rect 26754 1724 26806 1730
rect 27658 1882 27710 1890
rect 27658 1848 27665 1882
rect 27665 1848 27699 1882
rect 27699 1848 27710 1882
rect 27658 1838 27710 1848
rect 27570 1759 27622 1774
rect 27570 1725 27579 1759
rect 27579 1725 27613 1759
rect 27613 1725 27622 1759
rect 27570 1722 27622 1725
rect 26632 1489 26684 1541
rect 26808 1489 26860 1541
rect 27136 1474 27188 1486
rect 27136 1440 27144 1474
rect 27144 1440 27178 1474
rect 27178 1440 27188 1474
rect 27136 1434 27188 1440
rect 26634 1398 26686 1408
rect 26634 1364 26644 1398
rect 26644 1364 26678 1398
rect 26678 1364 26686 1398
rect 26634 1356 26686 1364
rect 25804 1141 25856 1144
rect 25804 1107 25837 1141
rect 25837 1107 25856 1141
rect 25804 1092 25856 1107
rect 26658 1133 26710 1150
rect 26658 1099 26679 1133
rect 26679 1099 26710 1133
rect 26658 1098 26710 1099
rect 27008 1281 27060 1292
rect 27008 1247 27016 1281
rect 27016 1247 27050 1281
rect 27050 1247 27060 1281
rect 27008 1240 27060 1247
rect 25566 1015 25618 1056
rect 25566 1004 25572 1015
rect 25572 1004 25606 1015
rect 25606 1004 25618 1015
rect 24261 826 24313 840
rect 24261 792 24267 826
rect 24267 792 24301 826
rect 24301 792 24313 826
rect 24261 788 24313 792
rect 24565 792 24617 844
rect 25228 855 25280 902
rect 25228 850 25238 855
rect 25238 850 25272 855
rect 25272 850 25280 855
rect 23678 612 23730 624
rect 23678 578 23686 612
rect 23686 578 23720 612
rect 23720 578 23730 612
rect 23678 572 23730 578
rect 24701 589 24753 602
rect 24701 555 24733 589
rect 24733 555 24753 589
rect 24701 550 24753 555
rect 24933 584 24985 592
rect 24933 550 24942 584
rect 24942 550 24976 584
rect 24976 550 24985 584
rect 24933 540 24985 550
rect 25246 418 25298 430
rect 25246 384 25254 418
rect 25254 384 25288 418
rect 25288 384 25298 418
rect 25246 378 25298 384
rect 26904 1015 26956 1036
rect 26904 984 26936 1015
rect 26936 984 26956 1015
rect 28734 1880 28786 1888
rect 28734 1846 28740 1880
rect 28740 1846 28774 1880
rect 28774 1846 28786 1880
rect 28734 1836 28786 1846
rect 29006 1911 29058 1958
rect 29006 1906 29016 1911
rect 29016 1906 29050 1911
rect 29050 1906 29058 1911
rect 28642 1764 28694 1776
rect 28642 1730 28649 1764
rect 28649 1730 28683 1764
rect 28683 1730 28694 1764
rect 28642 1724 28694 1730
rect 29546 1882 29598 1890
rect 29546 1848 29553 1882
rect 29553 1848 29587 1882
rect 29587 1848 29598 1882
rect 29546 1838 29598 1848
rect 29458 1759 29510 1774
rect 29458 1725 29467 1759
rect 29467 1725 29501 1759
rect 29501 1725 29510 1759
rect 29458 1722 29510 1725
rect 28520 1489 28572 1541
rect 28696 1489 28748 1541
rect 29024 1474 29076 1486
rect 29024 1440 29032 1474
rect 29032 1440 29066 1474
rect 29066 1440 29076 1474
rect 29024 1434 29076 1440
rect 28522 1398 28574 1408
rect 28522 1364 28532 1398
rect 28532 1364 28566 1398
rect 28566 1364 28574 1398
rect 28522 1356 28574 1364
rect 27692 1141 27744 1144
rect 27692 1107 27725 1141
rect 27725 1107 27744 1141
rect 27692 1092 27744 1107
rect 28546 1133 28598 1150
rect 28546 1099 28567 1133
rect 28567 1099 28598 1133
rect 28546 1098 28598 1099
rect 28896 1281 28948 1292
rect 28896 1247 28904 1281
rect 28904 1247 28938 1281
rect 28938 1247 28948 1281
rect 28896 1240 28948 1247
rect 27454 1015 27506 1056
rect 27454 1004 27460 1015
rect 27460 1004 27494 1015
rect 27494 1004 27506 1015
rect 26149 826 26201 840
rect 26149 792 26155 826
rect 26155 792 26189 826
rect 26189 792 26201 826
rect 26149 788 26201 792
rect 26453 792 26505 844
rect 27116 855 27168 902
rect 27116 850 27126 855
rect 27126 850 27160 855
rect 27160 850 27168 855
rect 25566 612 25618 624
rect 25566 578 25574 612
rect 25574 578 25608 612
rect 25608 578 25618 612
rect 25566 572 25618 578
rect 26589 589 26641 602
rect 26589 555 26621 589
rect 26621 555 26641 589
rect 26589 550 26641 555
rect 26821 584 26873 592
rect 26821 550 26830 584
rect 26830 550 26864 584
rect 26864 550 26873 584
rect 26821 540 26873 550
rect 27134 418 27186 430
rect 27134 384 27142 418
rect 27142 384 27176 418
rect 27176 384 27186 418
rect 27134 378 27186 384
rect 28792 1015 28844 1036
rect 28792 984 28824 1015
rect 28824 984 28844 1015
rect 30622 1880 30674 1888
rect 30622 1846 30628 1880
rect 30628 1846 30662 1880
rect 30662 1846 30674 1880
rect 30622 1836 30674 1846
rect 30894 1911 30946 1958
rect 30894 1906 30904 1911
rect 30904 1906 30938 1911
rect 30938 1906 30946 1911
rect 30530 1764 30582 1776
rect 30530 1730 30537 1764
rect 30537 1730 30571 1764
rect 30571 1730 30582 1764
rect 30530 1724 30582 1730
rect 31434 1882 31486 1890
rect 31434 1848 31441 1882
rect 31441 1848 31475 1882
rect 31475 1848 31486 1882
rect 31434 1838 31486 1848
rect 31346 1759 31398 1774
rect 31346 1725 31355 1759
rect 31355 1725 31389 1759
rect 31389 1725 31398 1759
rect 31346 1722 31398 1725
rect 30408 1489 30460 1541
rect 30584 1489 30636 1541
rect 30912 1474 30964 1486
rect 30912 1440 30920 1474
rect 30920 1440 30954 1474
rect 30954 1440 30964 1474
rect 30912 1434 30964 1440
rect 30410 1398 30462 1408
rect 30410 1364 30420 1398
rect 30420 1364 30454 1398
rect 30454 1364 30462 1398
rect 30410 1356 30462 1364
rect 29580 1141 29632 1144
rect 29580 1107 29613 1141
rect 29613 1107 29632 1141
rect 29580 1092 29632 1107
rect 30434 1133 30486 1150
rect 30434 1099 30455 1133
rect 30455 1099 30486 1133
rect 30434 1098 30486 1099
rect 30784 1281 30836 1292
rect 30784 1247 30792 1281
rect 30792 1247 30826 1281
rect 30826 1247 30836 1281
rect 30784 1240 30836 1247
rect 29342 1015 29394 1056
rect 29342 1004 29348 1015
rect 29348 1004 29382 1015
rect 29382 1004 29394 1015
rect 28037 826 28089 840
rect 28037 792 28043 826
rect 28043 792 28077 826
rect 28077 792 28089 826
rect 28037 788 28089 792
rect 28341 792 28393 844
rect 29004 855 29056 902
rect 29004 850 29014 855
rect 29014 850 29048 855
rect 29048 850 29056 855
rect 27454 612 27506 624
rect 27454 578 27462 612
rect 27462 578 27496 612
rect 27496 578 27506 612
rect 27454 572 27506 578
rect 28477 589 28529 602
rect 28477 555 28509 589
rect 28509 555 28529 589
rect 28477 550 28529 555
rect 28709 584 28761 592
rect 28709 550 28718 584
rect 28718 550 28752 584
rect 28752 550 28761 584
rect 28709 540 28761 550
rect 29022 418 29074 430
rect 29022 384 29030 418
rect 29030 384 29064 418
rect 29064 384 29074 418
rect 29022 378 29074 384
rect 30680 1015 30732 1036
rect 30680 984 30712 1015
rect 30712 984 30732 1015
rect 32510 1880 32562 1888
rect 32510 1846 32516 1880
rect 32516 1846 32550 1880
rect 32550 1846 32562 1880
rect 32510 1836 32562 1846
rect 32782 1911 32834 1958
rect 32782 1906 32792 1911
rect 32792 1906 32826 1911
rect 32826 1906 32834 1911
rect 32418 1764 32470 1776
rect 32418 1730 32425 1764
rect 32425 1730 32459 1764
rect 32459 1730 32470 1764
rect 32418 1724 32470 1730
rect 33322 1882 33374 1890
rect 33322 1848 33329 1882
rect 33329 1848 33363 1882
rect 33363 1848 33374 1882
rect 33322 1838 33374 1848
rect 33234 1759 33286 1774
rect 33234 1725 33243 1759
rect 33243 1725 33277 1759
rect 33277 1725 33286 1759
rect 33234 1722 33286 1725
rect 32296 1489 32348 1541
rect 32472 1489 32524 1541
rect 32800 1474 32852 1486
rect 32800 1440 32808 1474
rect 32808 1440 32842 1474
rect 32842 1440 32852 1474
rect 32800 1434 32852 1440
rect 32298 1398 32350 1408
rect 32298 1364 32308 1398
rect 32308 1364 32342 1398
rect 32342 1364 32350 1398
rect 32298 1356 32350 1364
rect 31468 1141 31520 1144
rect 31468 1107 31501 1141
rect 31501 1107 31520 1141
rect 31468 1092 31520 1107
rect 32322 1133 32374 1150
rect 32322 1099 32343 1133
rect 32343 1099 32374 1133
rect 32322 1098 32374 1099
rect 32672 1281 32724 1292
rect 32672 1247 32680 1281
rect 32680 1247 32714 1281
rect 32714 1247 32724 1281
rect 32672 1240 32724 1247
rect 31230 1015 31282 1056
rect 31230 1004 31236 1015
rect 31236 1004 31270 1015
rect 31270 1004 31282 1015
rect 29925 826 29977 840
rect 29925 792 29931 826
rect 29931 792 29965 826
rect 29965 792 29977 826
rect 29925 788 29977 792
rect 30229 792 30281 844
rect 30892 855 30944 902
rect 30892 850 30902 855
rect 30902 850 30936 855
rect 30936 850 30944 855
rect 29342 612 29394 624
rect 29342 578 29350 612
rect 29350 578 29384 612
rect 29384 578 29394 612
rect 29342 572 29394 578
rect 30365 589 30417 602
rect 30365 555 30397 589
rect 30397 555 30417 589
rect 30365 550 30417 555
rect 30597 584 30649 592
rect 30597 550 30606 584
rect 30606 550 30640 584
rect 30640 550 30649 584
rect 30597 540 30649 550
rect 30910 418 30962 430
rect 30910 384 30918 418
rect 30918 384 30952 418
rect 30952 384 30962 418
rect 30910 378 30962 384
rect 32568 1015 32620 1036
rect 32568 984 32600 1015
rect 32600 984 32620 1015
rect 34398 1880 34450 1888
rect 34398 1846 34404 1880
rect 34404 1846 34438 1880
rect 34438 1846 34450 1880
rect 34398 1836 34450 1846
rect 34670 1911 34722 1958
rect 34670 1906 34680 1911
rect 34680 1906 34714 1911
rect 34714 1906 34722 1911
rect 34306 1764 34358 1776
rect 34306 1730 34313 1764
rect 34313 1730 34347 1764
rect 34347 1730 34358 1764
rect 34306 1724 34358 1730
rect 35210 1882 35262 1890
rect 35210 1848 35217 1882
rect 35217 1848 35251 1882
rect 35251 1848 35262 1882
rect 35210 1838 35262 1848
rect 35122 1759 35174 1774
rect 35122 1725 35131 1759
rect 35131 1725 35165 1759
rect 35165 1725 35174 1759
rect 35122 1722 35174 1725
rect 34184 1489 34236 1541
rect 34360 1489 34412 1541
rect 34688 1474 34740 1486
rect 34688 1440 34696 1474
rect 34696 1440 34730 1474
rect 34730 1440 34740 1474
rect 34688 1434 34740 1440
rect 34186 1398 34238 1408
rect 34186 1364 34196 1398
rect 34196 1364 34230 1398
rect 34230 1364 34238 1398
rect 34186 1356 34238 1364
rect 33356 1141 33408 1144
rect 33356 1107 33389 1141
rect 33389 1107 33408 1141
rect 33356 1092 33408 1107
rect 34210 1133 34262 1150
rect 34210 1099 34231 1133
rect 34231 1099 34262 1133
rect 34210 1098 34262 1099
rect 34560 1281 34612 1292
rect 34560 1247 34568 1281
rect 34568 1247 34602 1281
rect 34602 1247 34612 1281
rect 34560 1240 34612 1247
rect 33118 1015 33170 1056
rect 33118 1004 33124 1015
rect 33124 1004 33158 1015
rect 33158 1004 33170 1015
rect 31813 826 31865 840
rect 31813 792 31819 826
rect 31819 792 31853 826
rect 31853 792 31865 826
rect 31813 788 31865 792
rect 32117 792 32169 844
rect 32780 855 32832 902
rect 32780 850 32790 855
rect 32790 850 32824 855
rect 32824 850 32832 855
rect 31230 612 31282 624
rect 31230 578 31238 612
rect 31238 578 31272 612
rect 31272 578 31282 612
rect 31230 572 31282 578
rect 32253 589 32305 602
rect 32253 555 32285 589
rect 32285 555 32305 589
rect 32253 550 32305 555
rect 32485 584 32537 592
rect 32485 550 32494 584
rect 32494 550 32528 584
rect 32528 550 32537 584
rect 32485 540 32537 550
rect 32798 418 32850 430
rect 32798 384 32806 418
rect 32806 384 32840 418
rect 32840 384 32850 418
rect 32798 378 32850 384
rect 34456 1015 34508 1036
rect 34456 984 34488 1015
rect 34488 984 34508 1015
rect 36286 1880 36338 1888
rect 36286 1846 36292 1880
rect 36292 1846 36326 1880
rect 36326 1846 36338 1880
rect 36286 1836 36338 1846
rect 36558 1911 36610 1958
rect 36558 1906 36568 1911
rect 36568 1906 36602 1911
rect 36602 1906 36610 1911
rect 36194 1764 36246 1776
rect 36194 1730 36201 1764
rect 36201 1730 36235 1764
rect 36235 1730 36246 1764
rect 36194 1724 36246 1730
rect 37098 1882 37150 1890
rect 37098 1848 37105 1882
rect 37105 1848 37139 1882
rect 37139 1848 37150 1882
rect 37098 1838 37150 1848
rect 37010 1759 37062 1774
rect 37010 1725 37019 1759
rect 37019 1725 37053 1759
rect 37053 1725 37062 1759
rect 37010 1722 37062 1725
rect 36072 1489 36124 1541
rect 36248 1489 36300 1541
rect 36576 1474 36628 1486
rect 36576 1440 36584 1474
rect 36584 1440 36618 1474
rect 36618 1440 36628 1474
rect 36576 1434 36628 1440
rect 36074 1398 36126 1408
rect 36074 1364 36084 1398
rect 36084 1364 36118 1398
rect 36118 1364 36126 1398
rect 36074 1356 36126 1364
rect 35244 1141 35296 1144
rect 35244 1107 35277 1141
rect 35277 1107 35296 1141
rect 35244 1092 35296 1107
rect 36098 1133 36150 1150
rect 36098 1099 36119 1133
rect 36119 1099 36150 1133
rect 36098 1098 36150 1099
rect 36448 1281 36500 1292
rect 36448 1247 36456 1281
rect 36456 1247 36490 1281
rect 36490 1247 36500 1281
rect 36448 1240 36500 1247
rect 35006 1015 35058 1056
rect 35006 1004 35012 1015
rect 35012 1004 35046 1015
rect 35046 1004 35058 1015
rect 33701 826 33753 840
rect 33701 792 33707 826
rect 33707 792 33741 826
rect 33741 792 33753 826
rect 33701 788 33753 792
rect 34005 792 34057 844
rect 34668 855 34720 902
rect 34668 850 34678 855
rect 34678 850 34712 855
rect 34712 850 34720 855
rect 33118 612 33170 624
rect 33118 578 33126 612
rect 33126 578 33160 612
rect 33160 578 33170 612
rect 33118 572 33170 578
rect 34141 589 34193 602
rect 34141 555 34173 589
rect 34173 555 34193 589
rect 34141 550 34193 555
rect 34373 584 34425 592
rect 34373 550 34382 584
rect 34382 550 34416 584
rect 34416 550 34425 584
rect 34373 540 34425 550
rect 34686 418 34738 430
rect 34686 384 34694 418
rect 34694 384 34728 418
rect 34728 384 34738 418
rect 34686 378 34738 384
rect 36344 1015 36396 1036
rect 36344 984 36376 1015
rect 36376 984 36396 1015
rect 38174 1880 38226 1888
rect 38174 1846 38180 1880
rect 38180 1846 38214 1880
rect 38214 1846 38226 1880
rect 38174 1836 38226 1846
rect 38446 1911 38498 1958
rect 38446 1906 38456 1911
rect 38456 1906 38490 1911
rect 38490 1906 38498 1911
rect 38082 1764 38134 1776
rect 38082 1730 38089 1764
rect 38089 1730 38123 1764
rect 38123 1730 38134 1764
rect 38082 1724 38134 1730
rect 38986 1882 39038 1890
rect 38986 1848 38993 1882
rect 38993 1848 39027 1882
rect 39027 1848 39038 1882
rect 38986 1838 39038 1848
rect 38898 1759 38950 1774
rect 38898 1725 38907 1759
rect 38907 1725 38941 1759
rect 38941 1725 38950 1759
rect 38898 1722 38950 1725
rect 37960 1489 38012 1541
rect 38136 1489 38188 1541
rect 38464 1474 38516 1486
rect 38464 1440 38472 1474
rect 38472 1440 38506 1474
rect 38506 1440 38516 1474
rect 38464 1434 38516 1440
rect 37962 1398 38014 1408
rect 37962 1364 37972 1398
rect 37972 1364 38006 1398
rect 38006 1364 38014 1398
rect 37962 1356 38014 1364
rect 37132 1141 37184 1144
rect 37132 1107 37165 1141
rect 37165 1107 37184 1141
rect 37132 1092 37184 1107
rect 37986 1133 38038 1150
rect 37986 1099 38007 1133
rect 38007 1099 38038 1133
rect 37986 1098 38038 1099
rect 38336 1281 38388 1292
rect 38336 1247 38344 1281
rect 38344 1247 38378 1281
rect 38378 1247 38388 1281
rect 38336 1240 38388 1247
rect 36894 1015 36946 1056
rect 36894 1004 36900 1015
rect 36900 1004 36934 1015
rect 36934 1004 36946 1015
rect 35589 826 35641 840
rect 35589 792 35595 826
rect 35595 792 35629 826
rect 35629 792 35641 826
rect 35589 788 35641 792
rect 35893 792 35945 844
rect 36556 855 36608 902
rect 36556 850 36566 855
rect 36566 850 36600 855
rect 36600 850 36608 855
rect 35006 612 35058 624
rect 35006 578 35014 612
rect 35014 578 35048 612
rect 35048 578 35058 612
rect 35006 572 35058 578
rect 36029 589 36081 602
rect 36029 555 36061 589
rect 36061 555 36081 589
rect 36029 550 36081 555
rect 36261 584 36313 592
rect 36261 550 36270 584
rect 36270 550 36304 584
rect 36304 550 36313 584
rect 36261 540 36313 550
rect 36574 418 36626 430
rect 36574 384 36582 418
rect 36582 384 36616 418
rect 36616 384 36626 418
rect 36574 378 36626 384
rect 38232 1015 38284 1036
rect 38232 984 38264 1015
rect 38264 984 38284 1015
rect 40062 1880 40114 1888
rect 40062 1846 40068 1880
rect 40068 1846 40102 1880
rect 40102 1846 40114 1880
rect 40062 1836 40114 1846
rect 40334 1911 40386 1958
rect 40334 1906 40344 1911
rect 40344 1906 40378 1911
rect 40378 1906 40386 1911
rect 39970 1764 40022 1776
rect 39970 1730 39977 1764
rect 39977 1730 40011 1764
rect 40011 1730 40022 1764
rect 39970 1724 40022 1730
rect 40874 1882 40926 1890
rect 40874 1848 40881 1882
rect 40881 1848 40915 1882
rect 40915 1848 40926 1882
rect 40874 1838 40926 1848
rect 40786 1759 40838 1774
rect 40786 1725 40795 1759
rect 40795 1725 40829 1759
rect 40829 1725 40838 1759
rect 40786 1722 40838 1725
rect 39848 1489 39900 1541
rect 40024 1489 40076 1541
rect 40352 1474 40404 1486
rect 40352 1440 40360 1474
rect 40360 1440 40394 1474
rect 40394 1440 40404 1474
rect 40352 1434 40404 1440
rect 39850 1398 39902 1408
rect 39850 1364 39860 1398
rect 39860 1364 39894 1398
rect 39894 1364 39902 1398
rect 39850 1356 39902 1364
rect 39020 1141 39072 1144
rect 39020 1107 39053 1141
rect 39053 1107 39072 1141
rect 39020 1092 39072 1107
rect 39874 1133 39926 1150
rect 39874 1099 39895 1133
rect 39895 1099 39926 1133
rect 39874 1098 39926 1099
rect 40224 1281 40276 1292
rect 40224 1247 40232 1281
rect 40232 1247 40266 1281
rect 40266 1247 40276 1281
rect 40224 1240 40276 1247
rect 38782 1015 38834 1056
rect 38782 1004 38788 1015
rect 38788 1004 38822 1015
rect 38822 1004 38834 1015
rect 37477 826 37529 840
rect 37477 792 37483 826
rect 37483 792 37517 826
rect 37517 792 37529 826
rect 37477 788 37529 792
rect 37781 792 37833 844
rect 38444 855 38496 902
rect 38444 850 38454 855
rect 38454 850 38488 855
rect 38488 850 38496 855
rect 36894 612 36946 624
rect 36894 578 36902 612
rect 36902 578 36936 612
rect 36936 578 36946 612
rect 36894 572 36946 578
rect 37917 589 37969 602
rect 37917 555 37949 589
rect 37949 555 37969 589
rect 37917 550 37969 555
rect 38149 584 38201 592
rect 38149 550 38158 584
rect 38158 550 38192 584
rect 38192 550 38201 584
rect 38149 540 38201 550
rect 38462 418 38514 430
rect 38462 384 38470 418
rect 38470 384 38504 418
rect 38504 384 38514 418
rect 38462 378 38514 384
rect 40120 1015 40172 1036
rect 40120 984 40152 1015
rect 40152 984 40172 1015
rect 41950 1880 42002 1888
rect 41950 1846 41956 1880
rect 41956 1846 41990 1880
rect 41990 1846 42002 1880
rect 41950 1836 42002 1846
rect 42222 1911 42274 1958
rect 42222 1906 42232 1911
rect 42232 1906 42266 1911
rect 42266 1906 42274 1911
rect 41858 1764 41910 1776
rect 41858 1730 41865 1764
rect 41865 1730 41899 1764
rect 41899 1730 41910 1764
rect 41858 1724 41910 1730
rect 42762 1882 42814 1890
rect 42762 1848 42769 1882
rect 42769 1848 42803 1882
rect 42803 1848 42814 1882
rect 42762 1838 42814 1848
rect 42674 1759 42726 1774
rect 42674 1725 42683 1759
rect 42683 1725 42717 1759
rect 42717 1725 42726 1759
rect 42674 1722 42726 1725
rect 41736 1489 41788 1541
rect 41912 1489 41964 1541
rect 42240 1474 42292 1486
rect 42240 1440 42248 1474
rect 42248 1440 42282 1474
rect 42282 1440 42292 1474
rect 42240 1434 42292 1440
rect 41738 1398 41790 1408
rect 41738 1364 41748 1398
rect 41748 1364 41782 1398
rect 41782 1364 41790 1398
rect 41738 1356 41790 1364
rect 40908 1141 40960 1144
rect 40908 1107 40941 1141
rect 40941 1107 40960 1141
rect 40908 1092 40960 1107
rect 41762 1133 41814 1150
rect 41762 1099 41783 1133
rect 41783 1099 41814 1133
rect 41762 1098 41814 1099
rect 42112 1281 42164 1292
rect 42112 1247 42120 1281
rect 42120 1247 42154 1281
rect 42154 1247 42164 1281
rect 42112 1240 42164 1247
rect 40670 1015 40722 1056
rect 40670 1004 40676 1015
rect 40676 1004 40710 1015
rect 40710 1004 40722 1015
rect 39365 826 39417 840
rect 39365 792 39371 826
rect 39371 792 39405 826
rect 39405 792 39417 826
rect 39365 788 39417 792
rect 39669 792 39721 844
rect 40332 855 40384 902
rect 40332 850 40342 855
rect 40342 850 40376 855
rect 40376 850 40384 855
rect 38782 612 38834 624
rect 38782 578 38790 612
rect 38790 578 38824 612
rect 38824 578 38834 612
rect 38782 572 38834 578
rect 39805 589 39857 602
rect 39805 555 39837 589
rect 39837 555 39857 589
rect 39805 550 39857 555
rect 40037 584 40089 592
rect 40037 550 40046 584
rect 40046 550 40080 584
rect 40080 550 40089 584
rect 40037 540 40089 550
rect 40350 418 40402 430
rect 40350 384 40358 418
rect 40358 384 40392 418
rect 40392 384 40402 418
rect 40350 378 40402 384
rect 42008 1015 42060 1036
rect 42008 984 42040 1015
rect 42040 984 42060 1015
rect 43838 1880 43890 1888
rect 43838 1846 43844 1880
rect 43844 1846 43878 1880
rect 43878 1846 43890 1880
rect 43838 1836 43890 1846
rect 44110 1911 44162 1958
rect 44110 1906 44120 1911
rect 44120 1906 44154 1911
rect 44154 1906 44162 1911
rect 43746 1764 43798 1776
rect 43746 1730 43753 1764
rect 43753 1730 43787 1764
rect 43787 1730 43798 1764
rect 43746 1724 43798 1730
rect 44650 1882 44702 1890
rect 44650 1848 44657 1882
rect 44657 1848 44691 1882
rect 44691 1848 44702 1882
rect 44650 1838 44702 1848
rect 44562 1759 44614 1774
rect 44562 1725 44571 1759
rect 44571 1725 44605 1759
rect 44605 1725 44614 1759
rect 44562 1722 44614 1725
rect 43624 1489 43676 1541
rect 43800 1489 43852 1541
rect 44128 1474 44180 1486
rect 44128 1440 44136 1474
rect 44136 1440 44170 1474
rect 44170 1440 44180 1474
rect 44128 1434 44180 1440
rect 43626 1398 43678 1408
rect 43626 1364 43636 1398
rect 43636 1364 43670 1398
rect 43670 1364 43678 1398
rect 43626 1356 43678 1364
rect 42796 1141 42848 1144
rect 42796 1107 42829 1141
rect 42829 1107 42848 1141
rect 42796 1092 42848 1107
rect 43650 1133 43702 1150
rect 43650 1099 43671 1133
rect 43671 1099 43702 1133
rect 43650 1098 43702 1099
rect 44000 1281 44052 1292
rect 44000 1247 44008 1281
rect 44008 1247 44042 1281
rect 44042 1247 44052 1281
rect 44000 1240 44052 1247
rect 42558 1015 42610 1056
rect 42558 1004 42564 1015
rect 42564 1004 42598 1015
rect 42598 1004 42610 1015
rect 41253 826 41305 840
rect 41253 792 41259 826
rect 41259 792 41293 826
rect 41293 792 41305 826
rect 41253 788 41305 792
rect 41557 792 41609 844
rect 42220 855 42272 902
rect 42220 850 42230 855
rect 42230 850 42264 855
rect 42264 850 42272 855
rect 40670 612 40722 624
rect 40670 578 40678 612
rect 40678 578 40712 612
rect 40712 578 40722 612
rect 40670 572 40722 578
rect 41693 589 41745 602
rect 41693 555 41725 589
rect 41725 555 41745 589
rect 41693 550 41745 555
rect 41925 584 41977 592
rect 41925 550 41934 584
rect 41934 550 41968 584
rect 41968 550 41977 584
rect 41925 540 41977 550
rect 42238 418 42290 430
rect 42238 384 42246 418
rect 42246 384 42280 418
rect 42280 384 42290 418
rect 42238 378 42290 384
rect 43896 1015 43948 1036
rect 43896 984 43928 1015
rect 43928 984 43948 1015
rect 45720 1880 45772 1888
rect 45720 1846 45726 1880
rect 45726 1846 45760 1880
rect 45760 1846 45772 1880
rect 45720 1836 45772 1846
rect 45992 1911 46044 1958
rect 45992 1906 46002 1911
rect 46002 1906 46036 1911
rect 46036 1906 46044 1911
rect 45628 1764 45680 1776
rect 45628 1730 45635 1764
rect 45635 1730 45669 1764
rect 45669 1730 45680 1764
rect 45628 1724 45680 1730
rect 46532 1882 46584 1890
rect 46532 1848 46539 1882
rect 46539 1848 46573 1882
rect 46573 1848 46584 1882
rect 46532 1838 46584 1848
rect 46444 1759 46496 1774
rect 46444 1725 46453 1759
rect 46453 1725 46487 1759
rect 46487 1725 46496 1759
rect 46444 1722 46496 1725
rect 45506 1489 45558 1541
rect 45682 1489 45734 1541
rect 46010 1474 46062 1486
rect 46010 1440 46018 1474
rect 46018 1440 46052 1474
rect 46052 1440 46062 1474
rect 46010 1434 46062 1440
rect 45508 1398 45560 1408
rect 45508 1364 45518 1398
rect 45518 1364 45552 1398
rect 45552 1364 45560 1398
rect 45508 1356 45560 1364
rect 44684 1141 44736 1144
rect 44684 1107 44717 1141
rect 44717 1107 44736 1141
rect 44684 1092 44736 1107
rect 45532 1133 45584 1150
rect 45532 1099 45553 1133
rect 45553 1099 45584 1133
rect 45532 1098 45584 1099
rect 45882 1281 45934 1292
rect 45882 1247 45890 1281
rect 45890 1247 45924 1281
rect 45924 1247 45934 1281
rect 45882 1240 45934 1247
rect 44446 1015 44498 1056
rect 44446 1004 44452 1015
rect 44452 1004 44486 1015
rect 44486 1004 44498 1015
rect 43141 826 43193 840
rect 43141 792 43147 826
rect 43147 792 43181 826
rect 43181 792 43193 826
rect 43141 788 43193 792
rect 43445 792 43497 844
rect 44108 855 44160 902
rect 44108 850 44118 855
rect 44118 850 44152 855
rect 44152 850 44160 855
rect 42558 612 42610 624
rect 42558 578 42566 612
rect 42566 578 42600 612
rect 42600 578 42610 612
rect 42558 572 42610 578
rect 43581 589 43633 602
rect 43581 555 43613 589
rect 43613 555 43633 589
rect 43581 550 43633 555
rect 43813 584 43865 592
rect 43813 550 43822 584
rect 43822 550 43856 584
rect 43856 550 43865 584
rect 43813 540 43865 550
rect 44126 418 44178 430
rect 44126 384 44134 418
rect 44134 384 44168 418
rect 44168 384 44178 418
rect 44126 378 44178 384
rect 45778 1015 45830 1036
rect 45778 984 45810 1015
rect 45810 984 45830 1015
rect 47608 1880 47660 1888
rect 47608 1846 47614 1880
rect 47614 1846 47648 1880
rect 47648 1846 47660 1880
rect 47608 1836 47660 1846
rect 47880 1911 47932 1958
rect 47880 1906 47890 1911
rect 47890 1906 47924 1911
rect 47924 1906 47932 1911
rect 47516 1764 47568 1776
rect 47516 1730 47523 1764
rect 47523 1730 47557 1764
rect 47557 1730 47568 1764
rect 47516 1724 47568 1730
rect 48420 1882 48472 1890
rect 48420 1848 48427 1882
rect 48427 1848 48461 1882
rect 48461 1848 48472 1882
rect 48420 1838 48472 1848
rect 48332 1759 48384 1774
rect 48332 1725 48341 1759
rect 48341 1725 48375 1759
rect 48375 1725 48384 1759
rect 48332 1722 48384 1725
rect 47394 1489 47446 1541
rect 47570 1489 47622 1541
rect 47898 1474 47950 1486
rect 47898 1440 47906 1474
rect 47906 1440 47940 1474
rect 47940 1440 47950 1474
rect 47898 1434 47950 1440
rect 47396 1398 47448 1408
rect 47396 1364 47406 1398
rect 47406 1364 47440 1398
rect 47440 1364 47448 1398
rect 47396 1356 47448 1364
rect 46566 1141 46618 1144
rect 46566 1107 46599 1141
rect 46599 1107 46618 1141
rect 46566 1092 46618 1107
rect 47420 1133 47472 1150
rect 47420 1099 47441 1133
rect 47441 1099 47472 1133
rect 47420 1098 47472 1099
rect 47770 1281 47822 1292
rect 47770 1247 47778 1281
rect 47778 1247 47812 1281
rect 47812 1247 47822 1281
rect 47770 1240 47822 1247
rect 46328 1015 46380 1056
rect 46328 1004 46334 1015
rect 46334 1004 46368 1015
rect 46368 1004 46380 1015
rect 45029 826 45081 840
rect 45029 792 45035 826
rect 45035 792 45069 826
rect 45069 792 45081 826
rect 45029 788 45081 792
rect 45327 792 45379 844
rect 45990 855 46042 902
rect 45990 850 46000 855
rect 46000 850 46034 855
rect 46034 850 46042 855
rect 44446 612 44498 624
rect 44446 578 44454 612
rect 44454 578 44488 612
rect 44488 578 44498 612
rect 44446 572 44498 578
rect 45463 589 45515 602
rect 45463 555 45495 589
rect 45495 555 45515 589
rect 45463 550 45515 555
rect 45695 584 45747 592
rect 45695 550 45704 584
rect 45704 550 45738 584
rect 45738 550 45747 584
rect 45695 540 45747 550
rect 46008 418 46060 430
rect 46008 384 46016 418
rect 46016 384 46050 418
rect 46050 384 46060 418
rect 46008 378 46060 384
rect 47666 1015 47718 1036
rect 47666 984 47698 1015
rect 47698 984 47718 1015
rect 49496 1880 49548 1888
rect 49496 1846 49502 1880
rect 49502 1846 49536 1880
rect 49536 1846 49548 1880
rect 49496 1836 49548 1846
rect 49768 1911 49820 1958
rect 49768 1906 49778 1911
rect 49778 1906 49812 1911
rect 49812 1906 49820 1911
rect 49404 1764 49456 1776
rect 49404 1730 49411 1764
rect 49411 1730 49445 1764
rect 49445 1730 49456 1764
rect 49404 1724 49456 1730
rect 50308 1882 50360 1890
rect 50308 1848 50315 1882
rect 50315 1848 50349 1882
rect 50349 1848 50360 1882
rect 50308 1838 50360 1848
rect 50220 1759 50272 1774
rect 50220 1725 50229 1759
rect 50229 1725 50263 1759
rect 50263 1725 50272 1759
rect 50220 1722 50272 1725
rect 49282 1489 49334 1541
rect 49458 1489 49510 1541
rect 49786 1474 49838 1486
rect 49786 1440 49794 1474
rect 49794 1440 49828 1474
rect 49828 1440 49838 1474
rect 49786 1434 49838 1440
rect 49284 1398 49336 1408
rect 49284 1364 49294 1398
rect 49294 1364 49328 1398
rect 49328 1364 49336 1398
rect 49284 1356 49336 1364
rect 48454 1141 48506 1144
rect 48454 1107 48487 1141
rect 48487 1107 48506 1141
rect 48454 1092 48506 1107
rect 49308 1133 49360 1150
rect 49308 1099 49329 1133
rect 49329 1099 49360 1133
rect 49308 1098 49360 1099
rect 49658 1281 49710 1292
rect 49658 1247 49666 1281
rect 49666 1247 49700 1281
rect 49700 1247 49710 1281
rect 49658 1240 49710 1247
rect 48216 1015 48268 1056
rect 48216 1004 48222 1015
rect 48222 1004 48256 1015
rect 48256 1004 48268 1015
rect 46911 826 46963 840
rect 46911 792 46917 826
rect 46917 792 46951 826
rect 46951 792 46963 826
rect 46911 788 46963 792
rect 47215 792 47267 844
rect 47878 855 47930 902
rect 47878 850 47888 855
rect 47888 850 47922 855
rect 47922 850 47930 855
rect 46328 612 46380 624
rect 46328 578 46336 612
rect 46336 578 46370 612
rect 46370 578 46380 612
rect 46328 572 46380 578
rect 47351 589 47403 602
rect 47351 555 47383 589
rect 47383 555 47403 589
rect 47351 550 47403 555
rect 47583 584 47635 592
rect 47583 550 47592 584
rect 47592 550 47626 584
rect 47626 550 47635 584
rect 47583 540 47635 550
rect 47896 418 47948 430
rect 47896 384 47904 418
rect 47904 384 47938 418
rect 47938 384 47948 418
rect 47896 378 47948 384
rect 49554 1015 49606 1036
rect 49554 984 49586 1015
rect 49586 984 49606 1015
rect 51384 1880 51436 1888
rect 51384 1846 51390 1880
rect 51390 1846 51424 1880
rect 51424 1846 51436 1880
rect 51384 1836 51436 1846
rect 51656 1911 51708 1958
rect 51656 1906 51666 1911
rect 51666 1906 51700 1911
rect 51700 1906 51708 1911
rect 51292 1764 51344 1776
rect 51292 1730 51299 1764
rect 51299 1730 51333 1764
rect 51333 1730 51344 1764
rect 51292 1724 51344 1730
rect 52196 1882 52248 1890
rect 52196 1848 52203 1882
rect 52203 1848 52237 1882
rect 52237 1848 52248 1882
rect 52196 1838 52248 1848
rect 52108 1759 52160 1774
rect 52108 1725 52117 1759
rect 52117 1725 52151 1759
rect 52151 1725 52160 1759
rect 52108 1722 52160 1725
rect 51170 1489 51222 1541
rect 51346 1489 51398 1541
rect 51674 1474 51726 1486
rect 51674 1440 51682 1474
rect 51682 1440 51716 1474
rect 51716 1440 51726 1474
rect 51674 1434 51726 1440
rect 51172 1398 51224 1408
rect 51172 1364 51182 1398
rect 51182 1364 51216 1398
rect 51216 1364 51224 1398
rect 51172 1356 51224 1364
rect 50342 1141 50394 1144
rect 50342 1107 50375 1141
rect 50375 1107 50394 1141
rect 50342 1092 50394 1107
rect 51196 1133 51248 1150
rect 51196 1099 51217 1133
rect 51217 1099 51248 1133
rect 51196 1098 51248 1099
rect 51546 1281 51598 1292
rect 51546 1247 51554 1281
rect 51554 1247 51588 1281
rect 51588 1247 51598 1281
rect 51546 1240 51598 1247
rect 50104 1015 50156 1056
rect 50104 1004 50110 1015
rect 50110 1004 50144 1015
rect 50144 1004 50156 1015
rect 48799 826 48851 840
rect 48799 792 48805 826
rect 48805 792 48839 826
rect 48839 792 48851 826
rect 48799 788 48851 792
rect 49103 792 49155 844
rect 49766 855 49818 902
rect 49766 850 49776 855
rect 49776 850 49810 855
rect 49810 850 49818 855
rect 48216 612 48268 624
rect 48216 578 48224 612
rect 48224 578 48258 612
rect 48258 578 48268 612
rect 48216 572 48268 578
rect 49239 589 49291 602
rect 49239 555 49271 589
rect 49271 555 49291 589
rect 49239 550 49291 555
rect 49471 584 49523 592
rect 49471 550 49480 584
rect 49480 550 49514 584
rect 49514 550 49523 584
rect 49471 540 49523 550
rect 49784 418 49836 430
rect 49784 384 49792 418
rect 49792 384 49826 418
rect 49826 384 49836 418
rect 49784 378 49836 384
rect 51442 1015 51494 1036
rect 51442 984 51474 1015
rect 51474 984 51494 1015
rect 53272 1880 53324 1888
rect 53272 1846 53278 1880
rect 53278 1846 53312 1880
rect 53312 1846 53324 1880
rect 53272 1836 53324 1846
rect 53544 1911 53596 1958
rect 53544 1906 53554 1911
rect 53554 1906 53588 1911
rect 53588 1906 53596 1911
rect 53180 1764 53232 1776
rect 53180 1730 53187 1764
rect 53187 1730 53221 1764
rect 53221 1730 53232 1764
rect 53180 1724 53232 1730
rect 54084 1882 54136 1890
rect 54084 1848 54091 1882
rect 54091 1848 54125 1882
rect 54125 1848 54136 1882
rect 54084 1838 54136 1848
rect 53996 1759 54048 1774
rect 53996 1725 54005 1759
rect 54005 1725 54039 1759
rect 54039 1725 54048 1759
rect 53996 1722 54048 1725
rect 53058 1489 53110 1541
rect 53234 1489 53286 1541
rect 53562 1474 53614 1486
rect 53562 1440 53570 1474
rect 53570 1440 53604 1474
rect 53604 1440 53614 1474
rect 53562 1434 53614 1440
rect 53060 1398 53112 1408
rect 53060 1364 53070 1398
rect 53070 1364 53104 1398
rect 53104 1364 53112 1398
rect 53060 1356 53112 1364
rect 52230 1141 52282 1144
rect 52230 1107 52263 1141
rect 52263 1107 52282 1141
rect 52230 1092 52282 1107
rect 53084 1133 53136 1150
rect 53084 1099 53105 1133
rect 53105 1099 53136 1133
rect 53084 1098 53136 1099
rect 53434 1281 53486 1292
rect 53434 1247 53442 1281
rect 53442 1247 53476 1281
rect 53476 1247 53486 1281
rect 53434 1240 53486 1247
rect 51992 1015 52044 1056
rect 51992 1004 51998 1015
rect 51998 1004 52032 1015
rect 52032 1004 52044 1015
rect 50687 826 50739 840
rect 50687 792 50693 826
rect 50693 792 50727 826
rect 50727 792 50739 826
rect 50687 788 50739 792
rect 50991 792 51043 844
rect 51654 855 51706 902
rect 51654 850 51664 855
rect 51664 850 51698 855
rect 51698 850 51706 855
rect 50104 612 50156 624
rect 50104 578 50112 612
rect 50112 578 50146 612
rect 50146 578 50156 612
rect 50104 572 50156 578
rect 51127 589 51179 602
rect 51127 555 51159 589
rect 51159 555 51179 589
rect 51127 550 51179 555
rect 51359 584 51411 592
rect 51359 550 51368 584
rect 51368 550 51402 584
rect 51402 550 51411 584
rect 51359 540 51411 550
rect 51672 418 51724 430
rect 51672 384 51680 418
rect 51680 384 51714 418
rect 51714 384 51724 418
rect 51672 378 51724 384
rect 53330 1015 53382 1036
rect 53330 984 53362 1015
rect 53362 984 53382 1015
rect 55160 1880 55212 1888
rect 55160 1846 55166 1880
rect 55166 1846 55200 1880
rect 55200 1846 55212 1880
rect 55160 1836 55212 1846
rect 55432 1911 55484 1958
rect 55432 1906 55442 1911
rect 55442 1906 55476 1911
rect 55476 1906 55484 1911
rect 55068 1764 55120 1776
rect 55068 1730 55075 1764
rect 55075 1730 55109 1764
rect 55109 1730 55120 1764
rect 55068 1724 55120 1730
rect 55972 1882 56024 1890
rect 55972 1848 55979 1882
rect 55979 1848 56013 1882
rect 56013 1848 56024 1882
rect 55972 1838 56024 1848
rect 55884 1759 55936 1774
rect 55884 1725 55893 1759
rect 55893 1725 55927 1759
rect 55927 1725 55936 1759
rect 55884 1722 55936 1725
rect 54946 1489 54998 1541
rect 55122 1489 55174 1541
rect 55450 1474 55502 1486
rect 55450 1440 55458 1474
rect 55458 1440 55492 1474
rect 55492 1440 55502 1474
rect 55450 1434 55502 1440
rect 54948 1398 55000 1408
rect 54948 1364 54958 1398
rect 54958 1364 54992 1398
rect 54992 1364 55000 1398
rect 54948 1356 55000 1364
rect 54118 1141 54170 1144
rect 54118 1107 54151 1141
rect 54151 1107 54170 1141
rect 54118 1092 54170 1107
rect 54972 1133 55024 1150
rect 54972 1099 54993 1133
rect 54993 1099 55024 1133
rect 54972 1098 55024 1099
rect 55322 1281 55374 1292
rect 55322 1247 55330 1281
rect 55330 1247 55364 1281
rect 55364 1247 55374 1281
rect 55322 1240 55374 1247
rect 53880 1015 53932 1056
rect 53880 1004 53886 1015
rect 53886 1004 53920 1015
rect 53920 1004 53932 1015
rect 52575 826 52627 840
rect 52575 792 52581 826
rect 52581 792 52615 826
rect 52615 792 52627 826
rect 52575 788 52627 792
rect 52879 792 52931 844
rect 53542 855 53594 902
rect 53542 850 53552 855
rect 53552 850 53586 855
rect 53586 850 53594 855
rect 51992 612 52044 624
rect 51992 578 52000 612
rect 52000 578 52034 612
rect 52034 578 52044 612
rect 51992 572 52044 578
rect 53015 589 53067 602
rect 53015 555 53047 589
rect 53047 555 53067 589
rect 53015 550 53067 555
rect 53247 584 53299 592
rect 53247 550 53256 584
rect 53256 550 53290 584
rect 53290 550 53299 584
rect 53247 540 53299 550
rect 53560 418 53612 430
rect 53560 384 53568 418
rect 53568 384 53602 418
rect 53602 384 53612 418
rect 53560 378 53612 384
rect 55218 1015 55270 1036
rect 55218 984 55250 1015
rect 55250 984 55270 1015
rect 57048 1880 57100 1888
rect 57048 1846 57054 1880
rect 57054 1846 57088 1880
rect 57088 1846 57100 1880
rect 57048 1836 57100 1846
rect 57320 1911 57372 1958
rect 57320 1906 57330 1911
rect 57330 1906 57364 1911
rect 57364 1906 57372 1911
rect 56956 1764 57008 1776
rect 56956 1730 56963 1764
rect 56963 1730 56997 1764
rect 56997 1730 57008 1764
rect 56956 1724 57008 1730
rect 57860 1882 57912 1890
rect 57860 1848 57867 1882
rect 57867 1848 57901 1882
rect 57901 1848 57912 1882
rect 57860 1838 57912 1848
rect 57772 1759 57824 1774
rect 57772 1725 57781 1759
rect 57781 1725 57815 1759
rect 57815 1725 57824 1759
rect 57772 1722 57824 1725
rect 56834 1489 56886 1541
rect 57010 1489 57062 1541
rect 57338 1474 57390 1486
rect 57338 1440 57346 1474
rect 57346 1440 57380 1474
rect 57380 1440 57390 1474
rect 57338 1434 57390 1440
rect 56836 1398 56888 1408
rect 56836 1364 56846 1398
rect 56846 1364 56880 1398
rect 56880 1364 56888 1398
rect 56836 1356 56888 1364
rect 56006 1141 56058 1144
rect 56006 1107 56039 1141
rect 56039 1107 56058 1141
rect 56006 1092 56058 1107
rect 56860 1133 56912 1150
rect 56860 1099 56881 1133
rect 56881 1099 56912 1133
rect 56860 1098 56912 1099
rect 57210 1281 57262 1292
rect 57210 1247 57218 1281
rect 57218 1247 57252 1281
rect 57252 1247 57262 1281
rect 57210 1240 57262 1247
rect 55768 1015 55820 1056
rect 55768 1004 55774 1015
rect 55774 1004 55808 1015
rect 55808 1004 55820 1015
rect 54463 826 54515 840
rect 54463 792 54469 826
rect 54469 792 54503 826
rect 54503 792 54515 826
rect 54463 788 54515 792
rect 54767 792 54819 844
rect 55430 855 55482 902
rect 55430 850 55440 855
rect 55440 850 55474 855
rect 55474 850 55482 855
rect 53880 612 53932 624
rect 53880 578 53888 612
rect 53888 578 53922 612
rect 53922 578 53932 612
rect 53880 572 53932 578
rect 54903 589 54955 602
rect 54903 555 54935 589
rect 54935 555 54955 589
rect 54903 550 54955 555
rect 55135 584 55187 592
rect 55135 550 55144 584
rect 55144 550 55178 584
rect 55178 550 55187 584
rect 55135 540 55187 550
rect 55448 418 55500 430
rect 55448 384 55456 418
rect 55456 384 55490 418
rect 55490 384 55500 418
rect 55448 378 55500 384
rect 57106 1015 57158 1036
rect 57106 984 57138 1015
rect 57138 984 57158 1015
rect 58936 1880 58988 1888
rect 58936 1846 58942 1880
rect 58942 1846 58976 1880
rect 58976 1846 58988 1880
rect 58936 1836 58988 1846
rect 59208 1911 59260 1958
rect 59208 1906 59218 1911
rect 59218 1906 59252 1911
rect 59252 1906 59260 1911
rect 58844 1764 58896 1776
rect 58844 1730 58851 1764
rect 58851 1730 58885 1764
rect 58885 1730 58896 1764
rect 58844 1724 58896 1730
rect 59748 1882 59800 1890
rect 59748 1848 59755 1882
rect 59755 1848 59789 1882
rect 59789 1848 59800 1882
rect 59748 1838 59800 1848
rect 59660 1759 59712 1774
rect 59660 1725 59669 1759
rect 59669 1725 59703 1759
rect 59703 1725 59712 1759
rect 59660 1722 59712 1725
rect 58722 1489 58774 1541
rect 58898 1489 58950 1541
rect 59226 1474 59278 1486
rect 59226 1440 59234 1474
rect 59234 1440 59268 1474
rect 59268 1440 59278 1474
rect 59226 1434 59278 1440
rect 58724 1398 58776 1408
rect 58724 1364 58734 1398
rect 58734 1364 58768 1398
rect 58768 1364 58776 1398
rect 58724 1356 58776 1364
rect 57894 1141 57946 1144
rect 57894 1107 57927 1141
rect 57927 1107 57946 1141
rect 57894 1092 57946 1107
rect 58748 1133 58800 1150
rect 58748 1099 58769 1133
rect 58769 1099 58800 1133
rect 58748 1098 58800 1099
rect 59098 1281 59150 1292
rect 59098 1247 59106 1281
rect 59106 1247 59140 1281
rect 59140 1247 59150 1281
rect 59098 1240 59150 1247
rect 57656 1015 57708 1056
rect 57656 1004 57662 1015
rect 57662 1004 57696 1015
rect 57696 1004 57708 1015
rect 56351 826 56403 840
rect 56351 792 56357 826
rect 56357 792 56391 826
rect 56391 792 56403 826
rect 56351 788 56403 792
rect 56655 792 56707 844
rect 57318 855 57370 902
rect 57318 850 57328 855
rect 57328 850 57362 855
rect 57362 850 57370 855
rect 55768 612 55820 624
rect 55768 578 55776 612
rect 55776 578 55810 612
rect 55810 578 55820 612
rect 55768 572 55820 578
rect 56791 589 56843 602
rect 56791 555 56823 589
rect 56823 555 56843 589
rect 56791 550 56843 555
rect 57023 584 57075 592
rect 57023 550 57032 584
rect 57032 550 57066 584
rect 57066 550 57075 584
rect 57023 540 57075 550
rect 57336 418 57388 430
rect 57336 384 57344 418
rect 57344 384 57378 418
rect 57378 384 57388 418
rect 57336 378 57388 384
rect 58994 1015 59046 1036
rect 58994 984 59026 1015
rect 59026 984 59046 1015
rect 59782 1141 59834 1144
rect 59782 1107 59815 1141
rect 59815 1107 59834 1141
rect 59782 1092 59834 1107
rect 59544 1015 59596 1056
rect 59544 1004 59550 1015
rect 59550 1004 59584 1015
rect 59584 1004 59596 1015
rect 58239 826 58291 840
rect 58239 792 58245 826
rect 58245 792 58279 826
rect 58279 792 58291 826
rect 58239 788 58291 792
rect 58543 792 58595 844
rect 59206 855 59258 902
rect 59206 850 59216 855
rect 59216 850 59250 855
rect 59250 850 59258 855
rect 57656 612 57708 624
rect 57656 578 57664 612
rect 57664 578 57698 612
rect 57698 578 57708 612
rect 57656 572 57708 578
rect 58679 589 58731 602
rect 58679 555 58711 589
rect 58711 555 58731 589
rect 58679 550 58731 555
rect 58911 584 58963 592
rect 58911 550 58920 584
rect 58920 550 58954 584
rect 58954 550 58963 584
rect 58911 540 58963 550
rect 59224 418 59276 430
rect 59224 384 59232 418
rect 59232 384 59266 418
rect 59266 384 59276 418
rect 59224 378 59276 384
rect 60127 826 60179 840
rect 60127 792 60133 826
rect 60133 792 60167 826
rect 60167 792 60179 826
rect 60127 788 60179 792
rect 59544 612 59596 624
rect 59544 578 59552 612
rect 59552 578 59586 612
rect 59586 578 59596 612
rect 59544 572 59596 578
rect 1535 64 1843 180
rect 3423 64 3731 180
rect 5311 64 5619 180
rect 7199 64 7507 180
rect 9087 64 9395 180
rect 10975 64 11283 180
rect 12863 64 13171 180
rect 14751 64 15059 180
rect 16633 64 16941 180
rect 18521 64 18829 180
rect 20409 64 20717 180
rect 22297 64 22605 180
rect 24185 64 24493 180
rect 26073 64 26381 180
rect 27961 64 28269 180
rect 29849 64 30157 180
rect 31737 64 32045 180
rect 33625 64 33933 180
rect 35513 64 35821 180
rect 37401 64 37709 180
rect 39289 64 39597 180
rect 41177 64 41485 180
rect 43065 64 43373 180
rect 44953 64 45261 180
rect 46835 64 47143 180
rect 48723 64 49031 180
rect 50611 64 50919 180
rect 52499 64 52807 180
rect 54387 64 54695 180
rect 56275 64 56583 180
rect 58163 64 58471 180
rect 60051 64 60359 180
<< metal2 >>
rect -398 7376 -48 7390
rect -398 7260 -377 7376
rect -69 7260 -48 7376
rect 1490 7376 1840 7390
rect -398 7246 -48 7260
rect 700 7062 766 7068
rect 700 7060 706 7062
rect 78 7032 706 7060
rect -206 6652 -126 6664
rect -206 6600 -197 6652
rect -145 6628 -126 6652
rect 78 6628 106 7032
rect 700 7010 706 7032
rect 758 7010 766 7062
rect 700 7004 766 7010
rect 370 6870 446 6874
rect 370 6868 538 6870
rect 370 6816 386 6868
rect 438 6842 538 6868
rect 438 6816 446 6842
rect 370 6810 446 6816
rect -145 6600 106 6628
rect -206 6592 106 6600
rect 78 5966 106 6592
rect 178 6436 446 6442
rect 178 6414 386 6436
rect 178 6356 206 6414
rect 380 6384 386 6414
rect 438 6384 446 6436
rect 380 6378 446 6384
rect 142 6348 206 6356
rect 142 6296 148 6348
rect 200 6296 206 6348
rect 142 6288 206 6296
rect -636 5930 106 5966
rect -636 5876 -520 5930
rect -629 1510 -539 5876
rect 510 5724 538 6842
rect 716 6598 766 7004
rect 1018 6900 1072 6916
rect 1018 6860 1019 6900
rect 858 6848 1019 6860
rect 1071 6848 1072 6900
rect 858 6832 1072 6848
rect 1242 6890 1306 6906
rect 1242 6838 1251 6890
rect 1303 6838 1306 6890
rect 716 6590 782 6598
rect 716 6538 724 6590
rect 776 6538 782 6590
rect 716 6530 782 6538
rect 858 6326 886 6832
rect 1242 6824 1306 6838
rect 928 6456 994 6464
rect 928 6404 936 6456
rect 988 6422 994 6456
rect 988 6404 1210 6422
rect 928 6398 1210 6404
rect 966 6394 1210 6398
rect 1182 6348 1210 6394
rect 1182 6342 1244 6348
rect 858 6298 1146 6326
rect 822 6212 858 6214
rect 822 6200 894 6212
rect 822 6148 832 6200
rect 884 6148 894 6200
rect 822 6136 894 6148
rect 698 6006 764 6012
rect 698 5954 704 6006
rect 756 5960 764 6006
rect 756 5954 1090 5960
rect 698 5951 1090 5954
rect 698 5948 1032 5951
rect 712 5932 1032 5948
rect 264 5718 538 5724
rect 264 5666 270 5718
rect 322 5696 538 5718
rect 322 5666 328 5696
rect 264 5660 328 5666
rect 176 5602 240 5608
rect 176 5550 182 5602
rect 234 5564 240 5602
rect 234 5550 242 5564
rect 176 5544 242 5550
rect 214 5440 242 5544
rect 714 5542 764 5932
rect 1026 5899 1032 5932
rect 1084 5899 1090 5951
rect 1026 5892 1090 5899
rect 1118 5726 1146 6298
rect 1234 6290 1244 6342
rect 1182 6284 1244 6290
rect 1278 6240 1306 6824
rect 1390 6654 1446 7270
rect 1490 7260 1511 7376
rect 1819 7260 1840 7376
rect 3378 7376 3728 7390
rect 1490 7246 1840 7260
rect 2588 7062 2654 7068
rect 2588 7060 2594 7062
rect 1966 7032 2594 7060
rect 1378 6648 1446 6654
rect 1378 6596 1387 6648
rect 1439 6596 1446 6648
rect 1378 6590 1446 6596
rect 1682 6652 1762 6664
rect 1682 6600 1691 6652
rect 1743 6628 1762 6652
rect 1966 6628 1994 7032
rect 2588 7010 2594 7032
rect 2646 7010 2654 7062
rect 2588 7004 2654 7010
rect 2258 6870 2334 6874
rect 2258 6868 2426 6870
rect 2258 6816 2274 6868
rect 2326 6842 2426 6868
rect 2326 6816 2334 6842
rect 2258 6810 2334 6816
rect 1743 6600 1994 6628
rect 1682 6592 1994 6600
rect 1238 6212 1306 6240
rect 1238 6090 1266 6212
rect 1200 6084 1266 6090
rect 1200 6032 1206 6084
rect 1258 6032 1266 6084
rect 1200 6026 1266 6032
rect 1966 5966 1994 6592
rect 2066 6436 2334 6442
rect 2066 6414 2274 6436
rect 2066 6356 2094 6414
rect 2268 6384 2274 6414
rect 2326 6384 2334 6436
rect 2268 6378 2334 6384
rect 2030 6348 2094 6356
rect 2030 6296 2036 6348
rect 2088 6296 2094 6348
rect 2030 6288 2094 6296
rect 1266 5960 1994 5966
rect 1260 5958 1994 5960
rect 1202 5951 1994 5958
rect 1202 5899 1208 5951
rect 1260 5930 1994 5951
rect 1260 5899 1266 5930
rect 1202 5892 1266 5899
rect 1078 5716 1146 5726
rect 2398 5724 2426 6842
rect 2604 6598 2654 7004
rect 2906 6900 2960 6916
rect 2906 6860 2907 6900
rect 2746 6848 2907 6860
rect 2959 6848 2960 6900
rect 2746 6832 2960 6848
rect 3130 6890 3194 6906
rect 3130 6838 3139 6890
rect 3191 6838 3194 6890
rect 2604 6590 2670 6598
rect 2604 6538 2612 6590
rect 2664 6538 2670 6590
rect 2604 6530 2670 6538
rect 2746 6326 2774 6832
rect 3130 6824 3194 6838
rect 2816 6456 2882 6464
rect 2816 6404 2824 6456
rect 2876 6422 2882 6456
rect 2876 6404 3098 6422
rect 2816 6398 3098 6404
rect 2854 6394 3098 6398
rect 3070 6348 3098 6394
rect 3070 6342 3132 6348
rect 2746 6298 3034 6326
rect 2710 6212 2746 6214
rect 2710 6200 2782 6212
rect 2710 6148 2720 6200
rect 2772 6148 2782 6200
rect 2710 6136 2782 6148
rect 2586 6006 2652 6012
rect 2586 5954 2592 6006
rect 2644 5960 2652 6006
rect 2644 5954 2978 5960
rect 2586 5951 2978 5954
rect 2586 5948 2920 5951
rect 2600 5932 2920 5948
rect 1078 5664 1086 5716
rect 1138 5664 1146 5716
rect 1078 5658 1146 5664
rect 2152 5718 2426 5724
rect 2152 5666 2158 5718
rect 2210 5696 2426 5718
rect 2210 5666 2216 5696
rect 2152 5660 2216 5666
rect 988 5604 1056 5610
rect 988 5552 994 5604
rect 1046 5552 1056 5604
rect 988 5546 1056 5552
rect 2064 5602 2128 5608
rect 2064 5550 2070 5602
rect 2122 5564 2128 5602
rect 2122 5550 2130 5564
rect 714 5534 780 5542
rect 714 5482 722 5534
rect 774 5482 780 5534
rect 714 5474 780 5482
rect 988 5440 1016 5546
rect 2064 5544 2130 5550
rect 2102 5440 2130 5544
rect 2602 5542 2652 5932
rect 2914 5899 2920 5932
rect 2972 5899 2978 5951
rect 2914 5892 2978 5899
rect 3006 5726 3034 6298
rect 3122 6290 3132 6342
rect 3070 6284 3132 6290
rect 3166 6240 3194 6824
rect 3278 6654 3334 7270
rect 3378 7260 3399 7376
rect 3707 7260 3728 7376
rect 5266 7376 5616 7390
rect 3378 7246 3728 7260
rect 4476 7062 4542 7068
rect 4476 7060 4482 7062
rect 3854 7032 4482 7060
rect 3266 6648 3334 6654
rect 3266 6596 3275 6648
rect 3327 6596 3334 6648
rect 3266 6590 3334 6596
rect 3570 6652 3650 6664
rect 3570 6600 3579 6652
rect 3631 6628 3650 6652
rect 3854 6628 3882 7032
rect 4476 7010 4482 7032
rect 4534 7010 4542 7062
rect 4476 7004 4542 7010
rect 4146 6870 4222 6874
rect 4146 6868 4314 6870
rect 4146 6816 4162 6868
rect 4214 6842 4314 6868
rect 4214 6816 4222 6842
rect 4146 6810 4222 6816
rect 3631 6600 3882 6628
rect 3570 6592 3882 6600
rect 3126 6212 3194 6240
rect 3126 6090 3154 6212
rect 3088 6084 3154 6090
rect 3088 6032 3094 6084
rect 3146 6032 3154 6084
rect 3088 6026 3154 6032
rect 3854 5966 3882 6592
rect 3954 6436 4222 6442
rect 3954 6414 4162 6436
rect 3954 6356 3982 6414
rect 4156 6384 4162 6414
rect 4214 6384 4222 6436
rect 4156 6378 4222 6384
rect 3918 6348 3982 6356
rect 3918 6296 3924 6348
rect 3976 6296 3982 6348
rect 3918 6288 3982 6296
rect 3154 5960 3882 5966
rect 3148 5958 3882 5960
rect 3090 5951 3882 5958
rect 3090 5899 3096 5951
rect 3148 5930 3882 5951
rect 3148 5899 3154 5930
rect 3090 5892 3154 5899
rect 2966 5716 3034 5726
rect 4286 5724 4314 6842
rect 4492 6598 4542 7004
rect 4794 6900 4848 6916
rect 4794 6860 4795 6900
rect 4634 6848 4795 6860
rect 4847 6848 4848 6900
rect 4634 6832 4848 6848
rect 5018 6890 5082 6906
rect 5018 6838 5027 6890
rect 5079 6838 5082 6890
rect 4492 6590 4558 6598
rect 4492 6538 4500 6590
rect 4552 6538 4558 6590
rect 4492 6530 4558 6538
rect 4634 6326 4662 6832
rect 5018 6824 5082 6838
rect 4704 6456 4770 6464
rect 4704 6404 4712 6456
rect 4764 6422 4770 6456
rect 4764 6404 4986 6422
rect 4704 6398 4986 6404
rect 4742 6394 4986 6398
rect 4958 6348 4986 6394
rect 4958 6342 5020 6348
rect 4634 6298 4922 6326
rect 4598 6212 4634 6214
rect 4598 6200 4670 6212
rect 4598 6148 4608 6200
rect 4660 6148 4670 6200
rect 4598 6136 4670 6148
rect 4474 6006 4540 6012
rect 4474 5954 4480 6006
rect 4532 5960 4540 6006
rect 4532 5954 4866 5960
rect 4474 5951 4866 5954
rect 4474 5948 4808 5951
rect 4488 5932 4808 5948
rect 2966 5664 2974 5716
rect 3026 5664 3034 5716
rect 2966 5658 3034 5664
rect 4040 5718 4314 5724
rect 4040 5666 4046 5718
rect 4098 5696 4314 5718
rect 4098 5666 4104 5696
rect 4040 5660 4104 5666
rect 2876 5604 2944 5610
rect 2876 5552 2882 5604
rect 2934 5552 2944 5604
rect 2876 5546 2944 5552
rect 3952 5602 4016 5608
rect 3952 5550 3958 5602
rect 4010 5564 4016 5602
rect 4010 5550 4018 5564
rect 2602 5534 2668 5542
rect 2602 5482 2610 5534
rect 2662 5482 2668 5534
rect 2602 5474 2668 5482
rect 2876 5440 2904 5546
rect 3952 5544 4018 5550
rect 3990 5440 4018 5544
rect 4490 5542 4540 5932
rect 4802 5899 4808 5932
rect 4860 5899 4866 5951
rect 4802 5892 4866 5899
rect 4894 5726 4922 6298
rect 5010 6290 5020 6342
rect 4958 6284 5020 6290
rect 5054 6240 5082 6824
rect 5166 6654 5222 7270
rect 5266 7260 5287 7376
rect 5595 7260 5616 7376
rect 7154 7376 7504 7390
rect 5266 7246 5616 7260
rect 6364 7062 6430 7068
rect 6364 7060 6370 7062
rect 5742 7032 6370 7060
rect 5154 6648 5222 6654
rect 5154 6596 5163 6648
rect 5215 6596 5222 6648
rect 5154 6590 5222 6596
rect 5458 6652 5538 6664
rect 5458 6600 5467 6652
rect 5519 6628 5538 6652
rect 5742 6628 5770 7032
rect 6364 7010 6370 7032
rect 6422 7010 6430 7062
rect 6364 7004 6430 7010
rect 6034 6870 6110 6874
rect 6034 6868 6202 6870
rect 6034 6816 6050 6868
rect 6102 6842 6202 6868
rect 6102 6816 6110 6842
rect 6034 6810 6110 6816
rect 5519 6600 5770 6628
rect 5458 6592 5770 6600
rect 5014 6212 5082 6240
rect 5014 6090 5042 6212
rect 4976 6084 5042 6090
rect 4976 6032 4982 6084
rect 5034 6032 5042 6084
rect 4976 6026 5042 6032
rect 5742 5966 5770 6592
rect 5842 6436 6110 6442
rect 5842 6414 6050 6436
rect 5842 6356 5870 6414
rect 6044 6384 6050 6414
rect 6102 6384 6110 6436
rect 6044 6378 6110 6384
rect 5806 6348 5870 6356
rect 5806 6296 5812 6348
rect 5864 6296 5870 6348
rect 5806 6288 5870 6296
rect 5042 5960 5770 5966
rect 5036 5958 5770 5960
rect 4978 5951 5770 5958
rect 4978 5899 4984 5951
rect 5036 5930 5770 5951
rect 5036 5899 5042 5930
rect 4978 5892 5042 5899
rect 4854 5716 4922 5726
rect 6174 5724 6202 6842
rect 6380 6598 6430 7004
rect 6682 6900 6736 6916
rect 6682 6860 6683 6900
rect 6522 6848 6683 6860
rect 6735 6848 6736 6900
rect 6522 6832 6736 6848
rect 6906 6890 6970 6906
rect 6906 6838 6915 6890
rect 6967 6838 6970 6890
rect 6380 6590 6446 6598
rect 6380 6538 6388 6590
rect 6440 6538 6446 6590
rect 6380 6530 6446 6538
rect 6522 6326 6550 6832
rect 6906 6824 6970 6838
rect 6592 6456 6658 6464
rect 6592 6404 6600 6456
rect 6652 6422 6658 6456
rect 6652 6404 6874 6422
rect 6592 6398 6874 6404
rect 6630 6394 6874 6398
rect 6846 6348 6874 6394
rect 6846 6342 6908 6348
rect 6522 6298 6810 6326
rect 6486 6212 6522 6214
rect 6486 6200 6558 6212
rect 6486 6148 6496 6200
rect 6548 6148 6558 6200
rect 6486 6136 6558 6148
rect 6362 6006 6428 6012
rect 6362 5954 6368 6006
rect 6420 5960 6428 6006
rect 6420 5954 6754 5960
rect 6362 5951 6754 5954
rect 6362 5948 6696 5951
rect 6376 5932 6696 5948
rect 4854 5664 4862 5716
rect 4914 5664 4922 5716
rect 4854 5658 4922 5664
rect 5928 5718 6202 5724
rect 5928 5666 5934 5718
rect 5986 5696 6202 5718
rect 5986 5666 5992 5696
rect 5928 5660 5992 5666
rect 4764 5604 4832 5610
rect 4764 5552 4770 5604
rect 4822 5552 4832 5604
rect 4764 5546 4832 5552
rect 5840 5602 5904 5608
rect 5840 5550 5846 5602
rect 5898 5564 5904 5602
rect 5898 5550 5906 5564
rect 4490 5534 4556 5542
rect 4490 5482 4498 5534
rect 4550 5482 4556 5534
rect 4490 5474 4556 5482
rect 4764 5440 4792 5546
rect 5840 5544 5906 5550
rect 5878 5444 5906 5544
rect 6378 5542 6428 5932
rect 6690 5899 6696 5932
rect 6748 5899 6754 5951
rect 6690 5892 6754 5899
rect 6782 5726 6810 6298
rect 6898 6290 6908 6342
rect 6846 6284 6908 6290
rect 6942 6240 6970 6824
rect 7054 6654 7110 7270
rect 7154 7260 7175 7376
rect 7483 7260 7504 7376
rect 9042 7376 9392 7390
rect 7154 7246 7504 7260
rect 8252 7062 8318 7068
rect 8252 7060 8258 7062
rect 7630 7032 8258 7060
rect 7042 6648 7110 6654
rect 7042 6596 7051 6648
rect 7103 6596 7110 6648
rect 7042 6590 7110 6596
rect 7346 6652 7426 6664
rect 7346 6600 7355 6652
rect 7407 6628 7426 6652
rect 7630 6628 7658 7032
rect 8252 7010 8258 7032
rect 8310 7010 8318 7062
rect 8252 7004 8318 7010
rect 7922 6870 7998 6874
rect 7922 6868 8090 6870
rect 7922 6816 7938 6868
rect 7990 6842 8090 6868
rect 7990 6816 7998 6842
rect 7922 6810 7998 6816
rect 7407 6600 7658 6628
rect 7346 6592 7658 6600
rect 6902 6212 6970 6240
rect 6902 6090 6930 6212
rect 6864 6084 6930 6090
rect 6864 6032 6870 6084
rect 6922 6032 6930 6084
rect 6864 6026 6930 6032
rect 7630 5966 7658 6592
rect 7730 6436 7998 6442
rect 7730 6414 7938 6436
rect 7730 6356 7758 6414
rect 7932 6384 7938 6414
rect 7990 6384 7998 6436
rect 7932 6378 7998 6384
rect 7694 6348 7758 6356
rect 7694 6296 7700 6348
rect 7752 6296 7758 6348
rect 7694 6288 7758 6296
rect 6930 5960 7658 5966
rect 6924 5958 7658 5960
rect 6866 5951 7658 5958
rect 6866 5899 6872 5951
rect 6924 5930 7658 5951
rect 6924 5899 6930 5930
rect 6866 5892 6930 5899
rect 6742 5716 6810 5726
rect 8062 5724 8090 6842
rect 8268 6598 8318 7004
rect 8570 6900 8624 6916
rect 8570 6860 8571 6900
rect 8410 6848 8571 6860
rect 8623 6848 8624 6900
rect 8410 6832 8624 6848
rect 8794 6890 8858 6906
rect 8794 6838 8803 6890
rect 8855 6838 8858 6890
rect 8268 6590 8334 6598
rect 8268 6538 8276 6590
rect 8328 6538 8334 6590
rect 8268 6530 8334 6538
rect 8410 6326 8438 6832
rect 8794 6824 8858 6838
rect 8480 6456 8546 6464
rect 8480 6404 8488 6456
rect 8540 6422 8546 6456
rect 8540 6404 8762 6422
rect 8480 6398 8762 6404
rect 8518 6394 8762 6398
rect 8734 6348 8762 6394
rect 8734 6342 8796 6348
rect 8410 6298 8698 6326
rect 8374 6212 8410 6214
rect 8374 6200 8446 6212
rect 8374 6148 8384 6200
rect 8436 6148 8446 6200
rect 8374 6136 8446 6148
rect 8250 6006 8316 6012
rect 8250 5954 8256 6006
rect 8308 5960 8316 6006
rect 8308 5954 8642 5960
rect 8250 5951 8642 5954
rect 8250 5948 8584 5951
rect 8264 5932 8584 5948
rect 6742 5664 6750 5716
rect 6802 5664 6810 5716
rect 6742 5658 6810 5664
rect 7816 5718 8090 5724
rect 7816 5666 7822 5718
rect 7874 5696 8090 5718
rect 7874 5666 7880 5696
rect 7816 5660 7880 5666
rect 6652 5604 6720 5610
rect 6652 5552 6658 5604
rect 6710 5552 6720 5604
rect 6652 5546 6720 5552
rect 7728 5602 7792 5608
rect 7728 5550 7734 5602
rect 7786 5564 7792 5602
rect 7786 5550 7794 5564
rect 6378 5534 6444 5542
rect 6378 5482 6386 5534
rect 6438 5482 6444 5534
rect 6378 5474 6444 5482
rect 6652 5444 6680 5546
rect 7728 5544 7794 5550
rect 7766 5444 7794 5544
rect 8266 5542 8316 5932
rect 8578 5899 8584 5932
rect 8636 5899 8642 5951
rect 8578 5892 8642 5899
rect 8670 5726 8698 6298
rect 8786 6290 8796 6342
rect 8734 6284 8796 6290
rect 8830 6240 8858 6824
rect 8942 6654 8998 7270
rect 9042 7260 9063 7376
rect 9371 7260 9392 7376
rect 10930 7376 11280 7390
rect 9042 7246 9392 7260
rect 10140 7062 10206 7068
rect 10140 7060 10146 7062
rect 9518 7032 10146 7060
rect 8930 6648 8998 6654
rect 8930 6596 8939 6648
rect 8991 6596 8998 6648
rect 8930 6590 8998 6596
rect 9234 6652 9314 6664
rect 9234 6600 9243 6652
rect 9295 6628 9314 6652
rect 9518 6628 9546 7032
rect 10140 7010 10146 7032
rect 10198 7010 10206 7062
rect 10140 7004 10206 7010
rect 9810 6870 9886 6874
rect 9810 6868 9978 6870
rect 9810 6816 9826 6868
rect 9878 6842 9978 6868
rect 9878 6816 9886 6842
rect 9810 6810 9886 6816
rect 9295 6600 9546 6628
rect 9234 6592 9546 6600
rect 8790 6212 8858 6240
rect 8790 6090 8818 6212
rect 8752 6084 8818 6090
rect 8752 6032 8758 6084
rect 8810 6032 8818 6084
rect 8752 6026 8818 6032
rect 9518 5966 9546 6592
rect 9618 6436 9886 6442
rect 9618 6414 9826 6436
rect 9618 6356 9646 6414
rect 9820 6384 9826 6414
rect 9878 6384 9886 6436
rect 9820 6378 9886 6384
rect 9582 6348 9646 6356
rect 9582 6296 9588 6348
rect 9640 6296 9646 6348
rect 9582 6288 9646 6296
rect 8818 5960 9546 5966
rect 8812 5958 9546 5960
rect 8754 5951 9546 5958
rect 8754 5899 8760 5951
rect 8812 5930 9546 5951
rect 8812 5899 8818 5930
rect 8754 5892 8818 5899
rect 8630 5716 8698 5726
rect 9950 5724 9978 6842
rect 10156 6598 10206 7004
rect 10458 6900 10512 6916
rect 10458 6860 10459 6900
rect 10298 6848 10459 6860
rect 10511 6848 10512 6900
rect 10298 6832 10512 6848
rect 10682 6890 10746 6906
rect 10682 6838 10691 6890
rect 10743 6838 10746 6890
rect 10156 6590 10222 6598
rect 10156 6538 10164 6590
rect 10216 6538 10222 6590
rect 10156 6530 10222 6538
rect 10298 6326 10326 6832
rect 10682 6824 10746 6838
rect 10368 6456 10434 6464
rect 10368 6404 10376 6456
rect 10428 6422 10434 6456
rect 10428 6404 10650 6422
rect 10368 6398 10650 6404
rect 10406 6394 10650 6398
rect 10622 6348 10650 6394
rect 10622 6342 10684 6348
rect 10298 6298 10586 6326
rect 10262 6212 10298 6214
rect 10262 6200 10334 6212
rect 10262 6148 10272 6200
rect 10324 6148 10334 6200
rect 10262 6136 10334 6148
rect 10138 6006 10204 6012
rect 10138 5954 10144 6006
rect 10196 5960 10204 6006
rect 10196 5954 10530 5960
rect 10138 5951 10530 5954
rect 10138 5948 10472 5951
rect 10152 5932 10472 5948
rect 8630 5664 8638 5716
rect 8690 5664 8698 5716
rect 8630 5658 8698 5664
rect 9704 5718 9978 5724
rect 9704 5666 9710 5718
rect 9762 5696 9978 5718
rect 9762 5666 9768 5696
rect 9704 5660 9768 5666
rect 8540 5604 8608 5610
rect 8540 5552 8546 5604
rect 8598 5552 8608 5604
rect 8540 5546 8608 5552
rect 9616 5602 9680 5608
rect 9616 5550 9622 5602
rect 9674 5564 9680 5602
rect 9674 5550 9682 5564
rect 8266 5534 8332 5542
rect 8266 5482 8274 5534
rect 8326 5482 8332 5534
rect 8266 5474 8332 5482
rect 8540 5444 8568 5546
rect 9616 5544 9682 5550
rect 5772 5440 7096 5444
rect 7660 5440 8980 5444
rect 9654 5440 9682 5544
rect 10154 5542 10204 5932
rect 10466 5899 10472 5932
rect 10524 5899 10530 5951
rect 10466 5892 10530 5899
rect 10558 5726 10586 6298
rect 10674 6290 10684 6342
rect 10622 6284 10684 6290
rect 10718 6240 10746 6824
rect 10830 6654 10886 7270
rect 10930 7260 10951 7376
rect 11259 7260 11280 7376
rect 12818 7376 13168 7390
rect 10930 7246 11280 7260
rect 12028 7062 12094 7068
rect 12028 7060 12034 7062
rect 11406 7032 12034 7060
rect 10818 6648 10886 6654
rect 10818 6596 10827 6648
rect 10879 6596 10886 6648
rect 10818 6590 10886 6596
rect 11122 6652 11202 6664
rect 11122 6600 11131 6652
rect 11183 6628 11202 6652
rect 11406 6628 11434 7032
rect 12028 7010 12034 7032
rect 12086 7010 12094 7062
rect 12028 7004 12094 7010
rect 11698 6870 11774 6874
rect 11698 6868 11866 6870
rect 11698 6816 11714 6868
rect 11766 6842 11866 6868
rect 11766 6816 11774 6842
rect 11698 6810 11774 6816
rect 11183 6600 11434 6628
rect 11122 6592 11434 6600
rect 10678 6212 10746 6240
rect 10678 6090 10706 6212
rect 10640 6084 10706 6090
rect 10640 6032 10646 6084
rect 10698 6032 10706 6084
rect 10640 6026 10706 6032
rect 11406 5966 11434 6592
rect 11506 6436 11774 6442
rect 11506 6414 11714 6436
rect 11506 6356 11534 6414
rect 11708 6384 11714 6414
rect 11766 6384 11774 6436
rect 11708 6378 11774 6384
rect 11470 6348 11534 6356
rect 11470 6296 11476 6348
rect 11528 6296 11534 6348
rect 11470 6288 11534 6296
rect 10706 5960 11434 5966
rect 10700 5958 11434 5960
rect 10642 5951 11434 5958
rect 10642 5899 10648 5951
rect 10700 5930 11434 5951
rect 10700 5899 10706 5930
rect 10642 5892 10706 5899
rect 10518 5716 10586 5726
rect 11838 5724 11866 6842
rect 12044 6598 12094 7004
rect 12346 6900 12400 6916
rect 12346 6860 12347 6900
rect 12186 6848 12347 6860
rect 12399 6848 12400 6900
rect 12186 6832 12400 6848
rect 12570 6890 12634 6906
rect 12570 6838 12579 6890
rect 12631 6838 12634 6890
rect 12044 6590 12110 6598
rect 12044 6538 12052 6590
rect 12104 6538 12110 6590
rect 12044 6530 12110 6538
rect 12186 6326 12214 6832
rect 12570 6824 12634 6838
rect 12256 6456 12322 6464
rect 12256 6404 12264 6456
rect 12316 6422 12322 6456
rect 12316 6404 12538 6422
rect 12256 6398 12538 6404
rect 12294 6394 12538 6398
rect 12510 6348 12538 6394
rect 12510 6342 12572 6348
rect 12186 6298 12474 6326
rect 12150 6212 12186 6214
rect 12150 6200 12222 6212
rect 12150 6148 12160 6200
rect 12212 6148 12222 6200
rect 12150 6136 12222 6148
rect 12026 6006 12092 6012
rect 12026 5954 12032 6006
rect 12084 5960 12092 6006
rect 12084 5954 12418 5960
rect 12026 5951 12418 5954
rect 12026 5948 12360 5951
rect 12040 5932 12360 5948
rect 10518 5664 10526 5716
rect 10578 5664 10586 5716
rect 10518 5658 10586 5664
rect 11592 5718 11866 5724
rect 11592 5666 11598 5718
rect 11650 5696 11866 5718
rect 11650 5666 11656 5696
rect 11592 5660 11656 5666
rect 10428 5604 10496 5610
rect 10428 5552 10434 5604
rect 10486 5552 10496 5604
rect 10428 5546 10496 5552
rect 11504 5602 11568 5608
rect 11504 5550 11510 5602
rect 11562 5564 11568 5602
rect 11562 5550 11570 5564
rect 10154 5534 10220 5542
rect 10154 5482 10162 5534
rect 10214 5482 10220 5534
rect 10154 5474 10220 5482
rect 10428 5440 10456 5546
rect 11504 5544 11570 5550
rect 11542 5440 11570 5544
rect 12042 5542 12092 5932
rect 12354 5899 12360 5932
rect 12412 5899 12418 5951
rect 12354 5892 12418 5899
rect 12446 5726 12474 6298
rect 12562 6290 12572 6342
rect 12510 6284 12572 6290
rect 12606 6240 12634 6824
rect 12718 6654 12774 7270
rect 12818 7260 12839 7376
rect 13147 7260 13168 7376
rect 14700 7376 15050 7390
rect 12818 7246 13168 7260
rect 13916 7062 13982 7068
rect 13916 7060 13922 7062
rect 13294 7032 13922 7060
rect 12706 6648 12774 6654
rect 12706 6596 12715 6648
rect 12767 6596 12774 6648
rect 12706 6590 12774 6596
rect 13010 6652 13090 6664
rect 13010 6600 13019 6652
rect 13071 6628 13090 6652
rect 13294 6628 13322 7032
rect 13916 7010 13922 7032
rect 13974 7010 13982 7062
rect 13916 7004 13982 7010
rect 13586 6870 13662 6874
rect 13586 6868 13754 6870
rect 13586 6816 13602 6868
rect 13654 6842 13754 6868
rect 13654 6816 13662 6842
rect 13586 6810 13662 6816
rect 13071 6600 13322 6628
rect 13010 6592 13322 6600
rect 12566 6212 12634 6240
rect 12566 6090 12594 6212
rect 12528 6084 12594 6090
rect 12528 6032 12534 6084
rect 12586 6032 12594 6084
rect 12528 6026 12594 6032
rect 13294 5966 13322 6592
rect 13394 6436 13662 6442
rect 13394 6414 13602 6436
rect 13394 6356 13422 6414
rect 13596 6384 13602 6414
rect 13654 6384 13662 6436
rect 13596 6378 13662 6384
rect 13358 6348 13422 6356
rect 13358 6296 13364 6348
rect 13416 6296 13422 6348
rect 13358 6288 13422 6296
rect 12594 5960 13322 5966
rect 12588 5958 13322 5960
rect 12530 5951 13322 5958
rect 12530 5899 12536 5951
rect 12588 5930 13322 5951
rect 12588 5899 12594 5930
rect 12530 5892 12594 5899
rect 12406 5716 12474 5726
rect 13726 5724 13754 6842
rect 13932 6598 13982 7004
rect 14234 6900 14288 6916
rect 14234 6860 14235 6900
rect 14074 6848 14235 6860
rect 14287 6848 14288 6900
rect 14074 6832 14288 6848
rect 14458 6890 14522 6906
rect 14458 6838 14467 6890
rect 14519 6838 14522 6890
rect 13932 6590 13998 6598
rect 13932 6538 13940 6590
rect 13992 6538 13998 6590
rect 13932 6530 13998 6538
rect 14074 6326 14102 6832
rect 14458 6824 14522 6838
rect 14144 6456 14210 6464
rect 14144 6404 14152 6456
rect 14204 6422 14210 6456
rect 14204 6404 14426 6422
rect 14144 6398 14426 6404
rect 14182 6394 14426 6398
rect 14398 6348 14426 6394
rect 14398 6342 14460 6348
rect 14074 6298 14362 6326
rect 14038 6212 14074 6214
rect 14038 6200 14110 6212
rect 14038 6148 14048 6200
rect 14100 6148 14110 6200
rect 14038 6136 14110 6148
rect 13914 6006 13980 6012
rect 13914 5954 13920 6006
rect 13972 5960 13980 6006
rect 13972 5954 14306 5960
rect 13914 5951 14306 5954
rect 13914 5948 14248 5951
rect 13928 5932 14248 5948
rect 12406 5664 12414 5716
rect 12466 5664 12474 5716
rect 12406 5658 12474 5664
rect 13480 5718 13754 5724
rect 13480 5666 13486 5718
rect 13538 5696 13754 5718
rect 13538 5666 13544 5696
rect 13480 5660 13544 5666
rect 12316 5604 12384 5610
rect 12316 5552 12322 5604
rect 12374 5552 12384 5604
rect 12316 5546 12384 5552
rect 13392 5602 13456 5608
rect 13392 5550 13398 5602
rect 13450 5564 13456 5602
rect 13450 5550 13458 5564
rect 12042 5534 12108 5542
rect 12042 5482 12050 5534
rect 12102 5482 12108 5534
rect 12042 5474 12108 5482
rect 12316 5440 12344 5546
rect 13392 5544 13458 5550
rect 13430 5440 13458 5544
rect 13930 5542 13980 5932
rect 14242 5899 14248 5932
rect 14300 5899 14306 5951
rect 14242 5892 14306 5899
rect 14334 5726 14362 6298
rect 14450 6290 14460 6342
rect 14398 6284 14460 6290
rect 14494 6240 14522 6824
rect 14606 6654 14662 7270
rect 14700 7260 14721 7376
rect 15029 7260 15050 7376
rect 16588 7376 16938 7390
rect 14700 7246 15050 7260
rect 15798 7062 15864 7068
rect 15798 7060 15804 7062
rect 15176 7032 15804 7060
rect 14594 6648 14662 6654
rect 14594 6596 14603 6648
rect 14655 6596 14662 6648
rect 14594 6590 14662 6596
rect 14892 6652 14972 6664
rect 14892 6600 14901 6652
rect 14953 6628 14972 6652
rect 15176 6628 15204 7032
rect 15798 7010 15804 7032
rect 15856 7010 15864 7062
rect 15798 7004 15864 7010
rect 15468 6870 15544 6874
rect 15468 6868 15636 6870
rect 15468 6816 15484 6868
rect 15536 6842 15636 6868
rect 15536 6816 15544 6842
rect 15468 6810 15544 6816
rect 14953 6600 15204 6628
rect 14892 6592 15204 6600
rect 14454 6212 14522 6240
rect 14454 6090 14482 6212
rect 14416 6084 14482 6090
rect 14416 6032 14422 6084
rect 14474 6032 14482 6084
rect 14416 6026 14482 6032
rect 15176 5966 15204 6592
rect 15276 6436 15544 6442
rect 15276 6414 15484 6436
rect 15276 6356 15304 6414
rect 15478 6384 15484 6414
rect 15536 6384 15544 6436
rect 15478 6378 15544 6384
rect 15240 6348 15304 6356
rect 15240 6296 15246 6348
rect 15298 6296 15304 6348
rect 15240 6288 15304 6296
rect 14482 5960 15204 5966
rect 14476 5958 15204 5960
rect 14418 5951 15204 5958
rect 14418 5899 14424 5951
rect 14476 5930 15204 5951
rect 14476 5899 14482 5930
rect 14418 5892 14482 5899
rect 14294 5716 14362 5726
rect 15608 5724 15636 6842
rect 15814 6598 15864 7004
rect 16116 6900 16170 6916
rect 16116 6860 16117 6900
rect 15956 6848 16117 6860
rect 16169 6848 16170 6900
rect 15956 6832 16170 6848
rect 16340 6890 16404 6906
rect 16340 6838 16349 6890
rect 16401 6838 16404 6890
rect 15814 6590 15880 6598
rect 15814 6538 15822 6590
rect 15874 6538 15880 6590
rect 15814 6530 15880 6538
rect 15956 6326 15984 6832
rect 16340 6824 16404 6838
rect 16026 6456 16092 6464
rect 16026 6404 16034 6456
rect 16086 6422 16092 6456
rect 16086 6404 16308 6422
rect 16026 6398 16308 6404
rect 16064 6394 16308 6398
rect 16280 6348 16308 6394
rect 16280 6342 16342 6348
rect 15956 6298 16244 6326
rect 15920 6212 15956 6214
rect 15920 6200 15992 6212
rect 15920 6148 15930 6200
rect 15982 6148 15992 6200
rect 15920 6136 15992 6148
rect 15796 6006 15862 6012
rect 15796 5954 15802 6006
rect 15854 5960 15862 6006
rect 15854 5954 16188 5960
rect 15796 5951 16188 5954
rect 15796 5948 16130 5951
rect 15810 5932 16130 5948
rect 14294 5664 14302 5716
rect 14354 5664 14362 5716
rect 14294 5658 14362 5664
rect 15362 5718 15636 5724
rect 15362 5666 15368 5718
rect 15420 5696 15636 5718
rect 15420 5666 15426 5696
rect 15362 5660 15426 5666
rect 14204 5604 14272 5610
rect 14204 5552 14210 5604
rect 14262 5552 14272 5604
rect 14204 5546 14272 5552
rect 15274 5602 15338 5608
rect 15274 5550 15280 5602
rect 15332 5564 15338 5602
rect 15332 5550 15340 5564
rect 13930 5534 13996 5542
rect 13930 5482 13938 5534
rect 13990 5482 13996 5534
rect 13930 5474 13996 5482
rect 14204 5440 14232 5546
rect 15274 5544 15340 5550
rect 15312 5444 15340 5544
rect 15812 5542 15862 5932
rect 16124 5899 16130 5932
rect 16182 5899 16188 5951
rect 16124 5892 16188 5899
rect 16216 5726 16244 6298
rect 16332 6290 16342 6342
rect 16280 6284 16342 6290
rect 16376 6240 16404 6824
rect 16494 6654 16544 7270
rect 16588 7260 16609 7376
rect 16917 7260 16938 7376
rect 18476 7376 18826 7390
rect 16588 7246 16938 7260
rect 17686 7062 17752 7068
rect 17686 7060 17692 7062
rect 17064 7032 17692 7060
rect 16476 6648 16544 6654
rect 16476 6596 16485 6648
rect 16537 6596 16544 6648
rect 16476 6590 16544 6596
rect 16780 6652 16860 6664
rect 16780 6600 16789 6652
rect 16841 6628 16860 6652
rect 17064 6628 17092 7032
rect 17686 7010 17692 7032
rect 17744 7010 17752 7062
rect 17686 7004 17752 7010
rect 17356 6870 17432 6874
rect 17356 6868 17524 6870
rect 17356 6816 17372 6868
rect 17424 6842 17524 6868
rect 17424 6816 17432 6842
rect 17356 6810 17432 6816
rect 16841 6600 17092 6628
rect 16780 6592 17092 6600
rect 16336 6212 16404 6240
rect 16336 6090 16364 6212
rect 16298 6084 16364 6090
rect 16298 6032 16304 6084
rect 16356 6032 16364 6084
rect 16298 6026 16364 6032
rect 17064 5966 17092 6592
rect 17164 6436 17432 6442
rect 17164 6414 17372 6436
rect 17164 6356 17192 6414
rect 17366 6384 17372 6414
rect 17424 6384 17432 6436
rect 17366 6378 17432 6384
rect 17128 6348 17192 6356
rect 17128 6296 17134 6348
rect 17186 6296 17192 6348
rect 17128 6288 17192 6296
rect 16364 5960 17092 5966
rect 16358 5958 17092 5960
rect 16300 5951 17092 5958
rect 16300 5899 16306 5951
rect 16358 5930 17092 5951
rect 16358 5899 16364 5930
rect 16300 5892 16364 5899
rect 16176 5716 16244 5726
rect 17496 5724 17524 6842
rect 17702 6598 17752 7004
rect 18004 6900 18058 6916
rect 18004 6860 18005 6900
rect 17844 6848 18005 6860
rect 18057 6848 18058 6900
rect 17844 6832 18058 6848
rect 18228 6890 18292 6906
rect 18228 6838 18237 6890
rect 18289 6838 18292 6890
rect 17702 6590 17768 6598
rect 17702 6538 17710 6590
rect 17762 6538 17768 6590
rect 17702 6530 17768 6538
rect 17844 6326 17872 6832
rect 18228 6824 18292 6838
rect 17914 6456 17980 6464
rect 17914 6404 17922 6456
rect 17974 6422 17980 6456
rect 17974 6404 18196 6422
rect 17914 6398 18196 6404
rect 17952 6394 18196 6398
rect 18168 6348 18196 6394
rect 18168 6342 18230 6348
rect 17844 6298 18132 6326
rect 17808 6212 17844 6214
rect 17808 6200 17880 6212
rect 17808 6148 17818 6200
rect 17870 6148 17880 6200
rect 17808 6136 17880 6148
rect 17684 6006 17750 6012
rect 17684 5954 17690 6006
rect 17742 5960 17750 6006
rect 17742 5954 18076 5960
rect 17684 5951 18076 5954
rect 17684 5948 18018 5951
rect 17698 5932 18018 5948
rect 16176 5664 16184 5716
rect 16236 5664 16244 5716
rect 16176 5658 16244 5664
rect 17250 5718 17524 5724
rect 17250 5666 17256 5718
rect 17308 5696 17524 5718
rect 17308 5666 17314 5696
rect 17250 5660 17314 5666
rect 16086 5604 16154 5610
rect 16086 5552 16092 5604
rect 16144 5552 16154 5604
rect 16086 5546 16154 5552
rect 17162 5602 17226 5608
rect 17162 5550 17168 5602
rect 17220 5564 17226 5602
rect 17220 5550 17228 5564
rect 15812 5534 15878 5542
rect 15812 5482 15820 5534
rect 15872 5482 15878 5534
rect 15812 5474 15878 5482
rect 16086 5444 16114 5546
rect 17162 5544 17228 5550
rect 17200 5444 17228 5544
rect 17700 5542 17750 5932
rect 18012 5899 18018 5932
rect 18070 5899 18076 5951
rect 18012 5892 18076 5899
rect 18104 5726 18132 6298
rect 18220 6290 18230 6342
rect 18168 6284 18230 6290
rect 18264 6240 18292 6824
rect 18382 6654 18432 7270
rect 18476 7260 18497 7376
rect 18805 7260 18826 7376
rect 20364 7376 20714 7390
rect 18476 7246 18826 7260
rect 19574 7062 19640 7068
rect 19574 7060 19580 7062
rect 18952 7032 19580 7060
rect 18364 6648 18432 6654
rect 18364 6596 18373 6648
rect 18425 6596 18432 6648
rect 18364 6590 18432 6596
rect 18668 6652 18748 6664
rect 18668 6600 18677 6652
rect 18729 6628 18748 6652
rect 18952 6628 18980 7032
rect 19574 7010 19580 7032
rect 19632 7010 19640 7062
rect 19574 7004 19640 7010
rect 19244 6870 19320 6874
rect 19244 6868 19412 6870
rect 19244 6816 19260 6868
rect 19312 6842 19412 6868
rect 19312 6816 19320 6842
rect 19244 6810 19320 6816
rect 18729 6600 18980 6628
rect 18668 6592 18980 6600
rect 18224 6212 18292 6240
rect 18224 6090 18252 6212
rect 18186 6084 18252 6090
rect 18186 6032 18192 6084
rect 18244 6032 18252 6084
rect 18186 6026 18252 6032
rect 18952 5966 18980 6592
rect 19052 6436 19320 6442
rect 19052 6414 19260 6436
rect 19052 6356 19080 6414
rect 19254 6384 19260 6414
rect 19312 6384 19320 6436
rect 19254 6378 19320 6384
rect 19016 6348 19080 6356
rect 19016 6296 19022 6348
rect 19074 6296 19080 6348
rect 19016 6288 19080 6296
rect 18252 5960 18980 5966
rect 18246 5958 18980 5960
rect 18188 5951 18980 5958
rect 18188 5899 18194 5951
rect 18246 5930 18980 5951
rect 18246 5899 18252 5930
rect 18188 5892 18252 5899
rect 18064 5716 18132 5726
rect 19384 5724 19412 6842
rect 19590 6598 19640 7004
rect 19892 6900 19946 6916
rect 19892 6860 19893 6900
rect 19732 6848 19893 6860
rect 19945 6848 19946 6900
rect 19732 6832 19946 6848
rect 20116 6890 20180 6906
rect 20116 6838 20125 6890
rect 20177 6838 20180 6890
rect 19590 6590 19656 6598
rect 19590 6538 19598 6590
rect 19650 6538 19656 6590
rect 19590 6530 19656 6538
rect 19732 6326 19760 6832
rect 20116 6824 20180 6838
rect 19802 6456 19868 6464
rect 19802 6404 19810 6456
rect 19862 6422 19868 6456
rect 19862 6404 20084 6422
rect 19802 6398 20084 6404
rect 19840 6394 20084 6398
rect 20056 6348 20084 6394
rect 20056 6342 20118 6348
rect 19732 6298 20020 6326
rect 19696 6212 19732 6214
rect 19696 6200 19768 6212
rect 19696 6148 19706 6200
rect 19758 6148 19768 6200
rect 19696 6136 19768 6148
rect 19572 6006 19638 6012
rect 19572 5954 19578 6006
rect 19630 5960 19638 6006
rect 19630 5954 19964 5960
rect 19572 5951 19964 5954
rect 19572 5948 19906 5951
rect 19586 5932 19906 5948
rect 18064 5664 18072 5716
rect 18124 5664 18132 5716
rect 18064 5658 18132 5664
rect 19138 5718 19412 5724
rect 19138 5666 19144 5718
rect 19196 5696 19412 5718
rect 19196 5666 19202 5696
rect 19138 5660 19202 5666
rect 17974 5604 18042 5610
rect 17974 5552 17980 5604
rect 18032 5552 18042 5604
rect 17974 5546 18042 5552
rect 19050 5602 19114 5608
rect 19050 5550 19056 5602
rect 19108 5564 19114 5602
rect 19108 5550 19116 5564
rect 17700 5534 17766 5542
rect 17700 5482 17708 5534
rect 17760 5482 17766 5534
rect 17700 5474 17766 5482
rect 17974 5444 18002 5546
rect 19050 5544 19116 5550
rect 19088 5444 19116 5544
rect 19588 5542 19638 5932
rect 19900 5899 19906 5932
rect 19958 5899 19964 5951
rect 19900 5892 19964 5899
rect 19992 5726 20020 6298
rect 20108 6290 20118 6342
rect 20056 6284 20118 6290
rect 20152 6240 20180 6824
rect 20270 6654 20320 7270
rect 20364 7260 20385 7376
rect 20693 7260 20714 7376
rect 22252 7376 22602 7390
rect 20364 7246 20714 7260
rect 21462 7062 21528 7068
rect 21462 7060 21468 7062
rect 20840 7032 21468 7060
rect 20252 6648 20320 6654
rect 20252 6596 20261 6648
rect 20313 6596 20320 6648
rect 20252 6590 20320 6596
rect 20556 6652 20636 6664
rect 20556 6600 20565 6652
rect 20617 6628 20636 6652
rect 20840 6628 20868 7032
rect 21462 7010 21468 7032
rect 21520 7010 21528 7062
rect 21462 7004 21528 7010
rect 21132 6870 21208 6874
rect 21132 6868 21300 6870
rect 21132 6816 21148 6868
rect 21200 6842 21300 6868
rect 21200 6816 21208 6842
rect 21132 6810 21208 6816
rect 20617 6600 20868 6628
rect 20556 6592 20868 6600
rect 20112 6212 20180 6240
rect 20112 6090 20140 6212
rect 20074 6084 20140 6090
rect 20074 6032 20080 6084
rect 20132 6032 20140 6084
rect 20074 6026 20140 6032
rect 20840 5966 20868 6592
rect 20940 6436 21208 6442
rect 20940 6414 21148 6436
rect 20940 6356 20968 6414
rect 21142 6384 21148 6414
rect 21200 6384 21208 6436
rect 21142 6378 21208 6384
rect 20904 6348 20968 6356
rect 20904 6296 20910 6348
rect 20962 6296 20968 6348
rect 20904 6288 20968 6296
rect 20140 5960 20868 5966
rect 20134 5958 20868 5960
rect 20076 5951 20868 5958
rect 20076 5899 20082 5951
rect 20134 5930 20868 5951
rect 20134 5899 20140 5930
rect 20076 5892 20140 5899
rect 19952 5716 20020 5726
rect 21272 5724 21300 6842
rect 21478 6598 21528 7004
rect 21780 6900 21834 6916
rect 21780 6860 21781 6900
rect 21620 6848 21781 6860
rect 21833 6848 21834 6900
rect 21620 6832 21834 6848
rect 22004 6890 22068 6906
rect 22004 6838 22013 6890
rect 22065 6838 22068 6890
rect 21478 6590 21544 6598
rect 21478 6538 21486 6590
rect 21538 6538 21544 6590
rect 21478 6530 21544 6538
rect 21620 6326 21648 6832
rect 22004 6824 22068 6838
rect 21690 6456 21756 6464
rect 21690 6404 21698 6456
rect 21750 6422 21756 6456
rect 21750 6404 21972 6422
rect 21690 6398 21972 6404
rect 21728 6394 21972 6398
rect 21944 6348 21972 6394
rect 21944 6342 22006 6348
rect 21620 6298 21908 6326
rect 21584 6212 21620 6214
rect 21584 6200 21656 6212
rect 21584 6148 21594 6200
rect 21646 6148 21656 6200
rect 21584 6136 21656 6148
rect 21460 6006 21526 6012
rect 21460 5954 21466 6006
rect 21518 5960 21526 6006
rect 21518 5954 21852 5960
rect 21460 5951 21852 5954
rect 21460 5948 21794 5951
rect 21474 5932 21794 5948
rect 19952 5664 19960 5716
rect 20012 5664 20020 5716
rect 19952 5658 20020 5664
rect 21026 5718 21300 5724
rect 21026 5666 21032 5718
rect 21084 5696 21300 5718
rect 21084 5666 21090 5696
rect 21026 5660 21090 5666
rect 19862 5604 19930 5610
rect 19862 5552 19868 5604
rect 19920 5552 19930 5604
rect 19862 5546 19930 5552
rect 20938 5602 21002 5608
rect 20938 5550 20944 5602
rect 20996 5564 21002 5602
rect 20996 5550 21004 5564
rect 19588 5534 19654 5542
rect 19588 5482 19596 5534
rect 19648 5482 19654 5534
rect 19588 5474 19654 5482
rect 19862 5444 19890 5546
rect 20938 5544 21004 5550
rect 20976 5444 21004 5544
rect 21476 5542 21526 5932
rect 21788 5899 21794 5932
rect 21846 5899 21852 5951
rect 21788 5892 21852 5899
rect 21880 5726 21908 6298
rect 21996 6290 22006 6342
rect 21944 6284 22006 6290
rect 22040 6240 22068 6824
rect 22158 6654 22208 7270
rect 22252 7260 22273 7376
rect 22581 7260 22602 7376
rect 24140 7376 24490 7390
rect 22252 7246 22602 7260
rect 23350 7062 23416 7068
rect 23350 7060 23356 7062
rect 22728 7032 23356 7060
rect 22140 6648 22208 6654
rect 22140 6596 22149 6648
rect 22201 6596 22208 6648
rect 22140 6590 22208 6596
rect 22444 6652 22524 6664
rect 22444 6600 22453 6652
rect 22505 6628 22524 6652
rect 22728 6628 22756 7032
rect 23350 7010 23356 7032
rect 23408 7010 23416 7062
rect 23350 7004 23416 7010
rect 23020 6870 23096 6874
rect 23020 6868 23188 6870
rect 23020 6816 23036 6868
rect 23088 6842 23188 6868
rect 23088 6816 23096 6842
rect 23020 6810 23096 6816
rect 22505 6600 22756 6628
rect 22444 6592 22756 6600
rect 22000 6212 22068 6240
rect 22000 6090 22028 6212
rect 21962 6084 22028 6090
rect 21962 6032 21968 6084
rect 22020 6032 22028 6084
rect 21962 6026 22028 6032
rect 22728 5966 22756 6592
rect 22828 6436 23096 6442
rect 22828 6414 23036 6436
rect 22828 6356 22856 6414
rect 23030 6384 23036 6414
rect 23088 6384 23096 6436
rect 23030 6378 23096 6384
rect 22792 6348 22856 6356
rect 22792 6296 22798 6348
rect 22850 6296 22856 6348
rect 22792 6288 22856 6296
rect 22028 5960 22756 5966
rect 22022 5958 22756 5960
rect 21964 5951 22756 5958
rect 21964 5899 21970 5951
rect 22022 5930 22756 5951
rect 22022 5899 22028 5930
rect 21964 5892 22028 5899
rect 21840 5716 21908 5726
rect 23160 5724 23188 6842
rect 23366 6598 23416 7004
rect 23668 6900 23722 6916
rect 23668 6860 23669 6900
rect 23508 6848 23669 6860
rect 23721 6848 23722 6900
rect 23508 6832 23722 6848
rect 23892 6890 23956 6906
rect 23892 6838 23901 6890
rect 23953 6838 23956 6890
rect 23366 6590 23432 6598
rect 23366 6538 23374 6590
rect 23426 6538 23432 6590
rect 23366 6530 23432 6538
rect 23508 6326 23536 6832
rect 23892 6824 23956 6838
rect 23578 6456 23644 6464
rect 23578 6404 23586 6456
rect 23638 6422 23644 6456
rect 23638 6404 23860 6422
rect 23578 6398 23860 6404
rect 23616 6394 23860 6398
rect 23832 6348 23860 6394
rect 23832 6342 23894 6348
rect 23508 6298 23796 6326
rect 23472 6212 23508 6214
rect 23472 6200 23544 6212
rect 23472 6148 23482 6200
rect 23534 6148 23544 6200
rect 23472 6136 23544 6148
rect 23348 6006 23414 6012
rect 23348 5954 23354 6006
rect 23406 5960 23414 6006
rect 23406 5954 23740 5960
rect 23348 5951 23740 5954
rect 23348 5948 23682 5951
rect 23362 5932 23682 5948
rect 21840 5664 21848 5716
rect 21900 5664 21908 5716
rect 21840 5658 21908 5664
rect 22914 5718 23188 5724
rect 22914 5666 22920 5718
rect 22972 5696 23188 5718
rect 22972 5666 22978 5696
rect 22914 5660 22978 5666
rect 21750 5604 21818 5610
rect 21750 5552 21756 5604
rect 21808 5552 21818 5604
rect 21750 5546 21818 5552
rect 22826 5602 22890 5608
rect 22826 5550 22832 5602
rect 22884 5564 22890 5602
rect 22884 5550 22892 5564
rect 21476 5534 21542 5542
rect 21476 5482 21484 5534
rect 21536 5482 21542 5534
rect 21476 5474 21542 5482
rect 21750 5444 21778 5546
rect 22826 5544 22892 5550
rect 22864 5444 22892 5544
rect 23364 5542 23414 5932
rect 23676 5899 23682 5932
rect 23734 5899 23740 5951
rect 23676 5892 23740 5899
rect 23768 5726 23796 6298
rect 23884 6290 23894 6342
rect 23832 6284 23894 6290
rect 23928 6240 23956 6824
rect 24046 6654 24096 7270
rect 24140 7260 24161 7376
rect 24469 7260 24490 7376
rect 26028 7376 26378 7390
rect 24140 7246 24490 7260
rect 25238 7062 25304 7068
rect 25238 7060 25244 7062
rect 24616 7032 25244 7060
rect 24028 6648 24096 6654
rect 24028 6596 24037 6648
rect 24089 6596 24096 6648
rect 24028 6590 24096 6596
rect 24332 6652 24412 6664
rect 24332 6600 24341 6652
rect 24393 6628 24412 6652
rect 24616 6628 24644 7032
rect 25238 7010 25244 7032
rect 25296 7010 25304 7062
rect 25238 7004 25304 7010
rect 24908 6870 24984 6874
rect 24908 6868 25076 6870
rect 24908 6816 24924 6868
rect 24976 6842 25076 6868
rect 24976 6816 24984 6842
rect 24908 6810 24984 6816
rect 24393 6600 24644 6628
rect 24332 6592 24644 6600
rect 23888 6212 23956 6240
rect 23888 6090 23916 6212
rect 23850 6084 23916 6090
rect 23850 6032 23856 6084
rect 23908 6032 23916 6084
rect 23850 6026 23916 6032
rect 24616 5966 24644 6592
rect 24716 6436 24984 6442
rect 24716 6414 24924 6436
rect 24716 6356 24744 6414
rect 24918 6384 24924 6414
rect 24976 6384 24984 6436
rect 24918 6378 24984 6384
rect 24680 6348 24744 6356
rect 24680 6296 24686 6348
rect 24738 6296 24744 6348
rect 24680 6288 24744 6296
rect 23916 5960 24644 5966
rect 23910 5958 24644 5960
rect 23852 5951 24644 5958
rect 23852 5899 23858 5951
rect 23910 5930 24644 5951
rect 23910 5899 23916 5930
rect 23852 5892 23916 5899
rect 23728 5716 23796 5726
rect 25048 5724 25076 6842
rect 25254 6598 25304 7004
rect 25556 6900 25610 6916
rect 25556 6860 25557 6900
rect 25396 6848 25557 6860
rect 25609 6848 25610 6900
rect 25396 6832 25610 6848
rect 25780 6890 25844 6906
rect 25780 6838 25789 6890
rect 25841 6838 25844 6890
rect 25254 6590 25320 6598
rect 25254 6538 25262 6590
rect 25314 6538 25320 6590
rect 25254 6530 25320 6538
rect 25396 6326 25424 6832
rect 25780 6824 25844 6838
rect 25466 6456 25532 6464
rect 25466 6404 25474 6456
rect 25526 6422 25532 6456
rect 25526 6404 25748 6422
rect 25466 6398 25748 6404
rect 25504 6394 25748 6398
rect 25720 6348 25748 6394
rect 25720 6342 25782 6348
rect 25396 6298 25684 6326
rect 25360 6212 25396 6214
rect 25360 6200 25432 6212
rect 25360 6148 25370 6200
rect 25422 6148 25432 6200
rect 25360 6136 25432 6148
rect 25236 6006 25302 6012
rect 25236 5954 25242 6006
rect 25294 5960 25302 6006
rect 25294 5954 25628 5960
rect 25236 5951 25628 5954
rect 25236 5948 25570 5951
rect 25250 5932 25570 5948
rect 23728 5664 23736 5716
rect 23788 5664 23796 5716
rect 23728 5658 23796 5664
rect 24802 5718 25076 5724
rect 24802 5666 24808 5718
rect 24860 5696 25076 5718
rect 24860 5666 24866 5696
rect 24802 5660 24866 5666
rect 23638 5604 23706 5610
rect 23638 5552 23644 5604
rect 23696 5552 23706 5604
rect 23638 5546 23706 5552
rect 24714 5602 24778 5608
rect 24714 5550 24720 5602
rect 24772 5564 24778 5602
rect 24772 5550 24780 5564
rect 23364 5534 23430 5542
rect 23364 5482 23372 5534
rect 23424 5482 23430 5534
rect 23364 5474 23430 5482
rect 23638 5444 23666 5546
rect 24714 5544 24780 5550
rect 15020 5440 22194 5444
rect 22758 5440 24078 5444
rect 24752 5440 24780 5544
rect 25252 5542 25302 5932
rect 25564 5899 25570 5932
rect 25622 5899 25628 5951
rect 25564 5892 25628 5899
rect 25656 5726 25684 6298
rect 25772 6290 25782 6342
rect 25720 6284 25782 6290
rect 25816 6240 25844 6824
rect 25934 6654 25984 7270
rect 26028 7260 26049 7376
rect 26357 7260 26378 7376
rect 27916 7376 28266 7390
rect 26028 7246 26378 7260
rect 27126 7062 27192 7068
rect 27126 7060 27132 7062
rect 26504 7032 27132 7060
rect 25916 6648 25984 6654
rect 25916 6596 25925 6648
rect 25977 6596 25984 6648
rect 25916 6590 25984 6596
rect 26220 6652 26300 6664
rect 26220 6600 26229 6652
rect 26281 6628 26300 6652
rect 26504 6628 26532 7032
rect 27126 7010 27132 7032
rect 27184 7010 27192 7062
rect 27126 7004 27192 7010
rect 26796 6870 26872 6874
rect 26796 6868 26964 6870
rect 26796 6816 26812 6868
rect 26864 6842 26964 6868
rect 26864 6816 26872 6842
rect 26796 6810 26872 6816
rect 26281 6600 26532 6628
rect 26220 6592 26532 6600
rect 25776 6212 25844 6240
rect 25776 6090 25804 6212
rect 25738 6084 25804 6090
rect 25738 6032 25744 6084
rect 25796 6032 25804 6084
rect 25738 6026 25804 6032
rect 26504 5966 26532 6592
rect 26604 6436 26872 6442
rect 26604 6414 26812 6436
rect 26604 6356 26632 6414
rect 26806 6384 26812 6414
rect 26864 6384 26872 6436
rect 26806 6378 26872 6384
rect 26568 6348 26632 6356
rect 26568 6296 26574 6348
rect 26626 6296 26632 6348
rect 26568 6288 26632 6296
rect 25804 5960 26532 5966
rect 25798 5958 26532 5960
rect 25740 5951 26532 5958
rect 25740 5899 25746 5951
rect 25798 5930 26532 5951
rect 25798 5899 25804 5930
rect 25740 5892 25804 5899
rect 25616 5716 25684 5726
rect 26936 5724 26964 6842
rect 27142 6598 27192 7004
rect 27444 6900 27498 6916
rect 27444 6860 27445 6900
rect 27284 6848 27445 6860
rect 27497 6848 27498 6900
rect 27284 6832 27498 6848
rect 27668 6890 27732 6906
rect 27668 6838 27677 6890
rect 27729 6838 27732 6890
rect 27142 6590 27208 6598
rect 27142 6538 27150 6590
rect 27202 6538 27208 6590
rect 27142 6530 27208 6538
rect 27284 6326 27312 6832
rect 27668 6824 27732 6838
rect 27354 6456 27420 6464
rect 27354 6404 27362 6456
rect 27414 6422 27420 6456
rect 27414 6404 27636 6422
rect 27354 6398 27636 6404
rect 27392 6394 27636 6398
rect 27608 6348 27636 6394
rect 27608 6342 27670 6348
rect 27284 6298 27572 6326
rect 27248 6212 27284 6214
rect 27248 6200 27320 6212
rect 27248 6148 27258 6200
rect 27310 6148 27320 6200
rect 27248 6136 27320 6148
rect 27124 6006 27190 6012
rect 27124 5954 27130 6006
rect 27182 5960 27190 6006
rect 27182 5954 27516 5960
rect 27124 5951 27516 5954
rect 27124 5948 27458 5951
rect 27138 5932 27458 5948
rect 25616 5664 25624 5716
rect 25676 5664 25684 5716
rect 25616 5658 25684 5664
rect 26690 5718 26964 5724
rect 26690 5666 26696 5718
rect 26748 5696 26964 5718
rect 26748 5666 26754 5696
rect 26690 5660 26754 5666
rect 25526 5604 25594 5610
rect 25526 5552 25532 5604
rect 25584 5552 25594 5604
rect 25526 5546 25594 5552
rect 26602 5602 26666 5608
rect 26602 5550 26608 5602
rect 26660 5564 26666 5602
rect 26660 5550 26668 5564
rect 25252 5534 25318 5542
rect 25252 5482 25260 5534
rect 25312 5482 25318 5534
rect 25252 5474 25318 5482
rect 25526 5440 25554 5546
rect 26602 5544 26668 5550
rect 26640 5440 26668 5544
rect 27140 5542 27190 5932
rect 27452 5899 27458 5932
rect 27510 5899 27516 5951
rect 27452 5892 27516 5899
rect 27544 5726 27572 6298
rect 27660 6290 27670 6342
rect 27608 6284 27670 6290
rect 27704 6240 27732 6824
rect 27822 6654 27872 7270
rect 27916 7260 27937 7376
rect 28245 7260 28266 7376
rect 29804 7376 30154 7390
rect 27916 7246 28266 7260
rect 29014 7062 29080 7068
rect 29014 7060 29020 7062
rect 28392 7032 29020 7060
rect 27804 6648 27872 6654
rect 27804 6596 27813 6648
rect 27865 6596 27872 6648
rect 27804 6590 27872 6596
rect 28108 6652 28188 6664
rect 28108 6600 28117 6652
rect 28169 6628 28188 6652
rect 28392 6628 28420 7032
rect 29014 7010 29020 7032
rect 29072 7010 29080 7062
rect 29014 7004 29080 7010
rect 28684 6870 28760 6874
rect 28684 6868 28852 6870
rect 28684 6816 28700 6868
rect 28752 6842 28852 6868
rect 28752 6816 28760 6842
rect 28684 6810 28760 6816
rect 28169 6600 28420 6628
rect 28108 6592 28420 6600
rect 27664 6212 27732 6240
rect 27664 6090 27692 6212
rect 27626 6084 27692 6090
rect 27626 6032 27632 6084
rect 27684 6032 27692 6084
rect 27626 6026 27692 6032
rect 28392 5966 28420 6592
rect 28492 6436 28760 6442
rect 28492 6414 28700 6436
rect 28492 6356 28520 6414
rect 28694 6384 28700 6414
rect 28752 6384 28760 6436
rect 28694 6378 28760 6384
rect 28456 6348 28520 6356
rect 28456 6296 28462 6348
rect 28514 6296 28520 6348
rect 28456 6288 28520 6296
rect 27692 5960 28420 5966
rect 27686 5958 28420 5960
rect 27628 5951 28420 5958
rect 27628 5899 27634 5951
rect 27686 5930 28420 5951
rect 27686 5899 27692 5930
rect 27628 5892 27692 5899
rect 27504 5716 27572 5726
rect 28824 5724 28852 6842
rect 29030 6598 29080 7004
rect 29332 6900 29386 6916
rect 29332 6860 29333 6900
rect 29172 6848 29333 6860
rect 29385 6848 29386 6900
rect 29172 6832 29386 6848
rect 29556 6890 29620 6906
rect 29556 6838 29565 6890
rect 29617 6838 29620 6890
rect 29030 6590 29096 6598
rect 29030 6538 29038 6590
rect 29090 6538 29096 6590
rect 29030 6530 29096 6538
rect 29172 6326 29200 6832
rect 29556 6824 29620 6838
rect 29242 6456 29308 6464
rect 29242 6404 29250 6456
rect 29302 6422 29308 6456
rect 29302 6404 29524 6422
rect 29242 6398 29524 6404
rect 29280 6394 29524 6398
rect 29496 6348 29524 6394
rect 29496 6342 29558 6348
rect 29172 6298 29460 6326
rect 29136 6212 29172 6214
rect 29136 6200 29208 6212
rect 29136 6148 29146 6200
rect 29198 6148 29208 6200
rect 29136 6136 29208 6148
rect 29012 6006 29078 6012
rect 29012 5954 29018 6006
rect 29070 5960 29078 6006
rect 29070 5954 29404 5960
rect 29012 5951 29404 5954
rect 29012 5948 29346 5951
rect 29026 5932 29346 5948
rect 27504 5664 27512 5716
rect 27564 5664 27572 5716
rect 27504 5658 27572 5664
rect 28578 5718 28852 5724
rect 28578 5666 28584 5718
rect 28636 5696 28852 5718
rect 28636 5666 28642 5696
rect 28578 5660 28642 5666
rect 27414 5604 27482 5610
rect 27414 5552 27420 5604
rect 27472 5552 27482 5604
rect 27414 5546 27482 5552
rect 28490 5602 28554 5608
rect 28490 5550 28496 5602
rect 28548 5564 28554 5602
rect 28548 5550 28556 5564
rect 27140 5534 27206 5542
rect 27140 5482 27148 5534
rect 27200 5482 27206 5534
rect 27140 5474 27206 5482
rect 27414 5440 27442 5546
rect 28490 5544 28556 5550
rect 28528 5440 28556 5544
rect 29028 5542 29078 5932
rect 29340 5899 29346 5932
rect 29398 5899 29404 5951
rect 29340 5892 29404 5899
rect 29432 5726 29460 6298
rect 29548 6290 29558 6342
rect 29496 6284 29558 6290
rect 29592 6240 29620 6824
rect 29710 6654 29760 7270
rect 29804 7260 29825 7376
rect 30133 7260 30154 7376
rect 31692 7376 32042 7390
rect 29804 7246 30154 7260
rect 30902 7062 30968 7068
rect 30902 7060 30908 7062
rect 30280 7032 30908 7060
rect 29692 6648 29760 6654
rect 29692 6596 29701 6648
rect 29753 6596 29760 6648
rect 29692 6590 29760 6596
rect 29996 6652 30076 6664
rect 29996 6600 30005 6652
rect 30057 6628 30076 6652
rect 30280 6628 30308 7032
rect 30902 7010 30908 7032
rect 30960 7010 30968 7062
rect 30902 7004 30968 7010
rect 30572 6870 30648 6874
rect 30572 6868 30740 6870
rect 30572 6816 30588 6868
rect 30640 6842 30740 6868
rect 30640 6816 30648 6842
rect 30572 6810 30648 6816
rect 30057 6600 30308 6628
rect 29996 6592 30308 6600
rect 29552 6212 29620 6240
rect 29552 6090 29580 6212
rect 29514 6084 29580 6090
rect 29514 6032 29520 6084
rect 29572 6032 29580 6084
rect 29514 6026 29580 6032
rect 30280 5966 30308 6592
rect 30380 6436 30648 6442
rect 30380 6414 30588 6436
rect 30380 6356 30408 6414
rect 30582 6384 30588 6414
rect 30640 6384 30648 6436
rect 30582 6378 30648 6384
rect 30344 6348 30408 6356
rect 30344 6296 30350 6348
rect 30402 6296 30408 6348
rect 30344 6288 30408 6296
rect 29580 5960 30308 5966
rect 29574 5958 30308 5960
rect 29516 5951 30308 5958
rect 29516 5899 29522 5951
rect 29574 5930 30308 5951
rect 29574 5899 29580 5930
rect 29516 5892 29580 5899
rect 29392 5716 29460 5726
rect 30712 5724 30740 6842
rect 30918 6598 30968 7004
rect 31220 6900 31274 6916
rect 31220 6860 31221 6900
rect 31060 6848 31221 6860
rect 31273 6848 31274 6900
rect 31060 6832 31274 6848
rect 31444 6890 31508 6906
rect 31444 6838 31453 6890
rect 31505 6838 31508 6890
rect 30918 6590 30984 6598
rect 30918 6538 30926 6590
rect 30978 6538 30984 6590
rect 30918 6530 30984 6538
rect 31060 6326 31088 6832
rect 31444 6824 31508 6838
rect 31130 6456 31196 6464
rect 31130 6404 31138 6456
rect 31190 6422 31196 6456
rect 31190 6404 31412 6422
rect 31130 6398 31412 6404
rect 31168 6394 31412 6398
rect 31384 6348 31412 6394
rect 31384 6342 31446 6348
rect 31060 6298 31348 6326
rect 31024 6212 31060 6214
rect 31024 6200 31096 6212
rect 31024 6148 31034 6200
rect 31086 6148 31096 6200
rect 31024 6136 31096 6148
rect 30900 6006 30966 6012
rect 30900 5954 30906 6006
rect 30958 5960 30966 6006
rect 30958 5954 31292 5960
rect 30900 5951 31292 5954
rect 30900 5948 31234 5951
rect 30914 5932 31234 5948
rect 29392 5664 29400 5716
rect 29452 5664 29460 5716
rect 29392 5658 29460 5664
rect 30466 5718 30740 5724
rect 30466 5666 30472 5718
rect 30524 5696 30740 5718
rect 30524 5666 30530 5696
rect 30466 5660 30530 5666
rect 29302 5604 29370 5610
rect 29302 5552 29308 5604
rect 29360 5552 29370 5604
rect 29302 5546 29370 5552
rect 30378 5602 30442 5608
rect 30378 5550 30384 5602
rect 30436 5564 30442 5602
rect 30436 5550 30444 5564
rect 29028 5534 29094 5542
rect 29028 5482 29036 5534
rect 29088 5482 29094 5534
rect 29028 5474 29094 5482
rect 29302 5440 29330 5546
rect 30378 5544 30444 5550
rect 30416 5440 30444 5544
rect 30916 5542 30966 5932
rect 31228 5899 31234 5932
rect 31286 5899 31292 5951
rect 31228 5892 31292 5899
rect 31320 5726 31348 6298
rect 31436 6290 31446 6342
rect 31384 6284 31446 6290
rect 31480 6240 31508 6824
rect 31598 6654 31648 7270
rect 31692 7260 31713 7376
rect 32021 7260 32042 7376
rect 33580 7376 33930 7390
rect 31692 7246 32042 7260
rect 32790 7062 32856 7068
rect 32790 7060 32796 7062
rect 32168 7032 32796 7060
rect 31580 6648 31648 6654
rect 31580 6596 31589 6648
rect 31641 6596 31648 6648
rect 31580 6590 31648 6596
rect 31884 6652 31964 6664
rect 31884 6600 31893 6652
rect 31945 6628 31964 6652
rect 32168 6628 32196 7032
rect 32790 7010 32796 7032
rect 32848 7010 32856 7062
rect 32790 7004 32856 7010
rect 32460 6870 32536 6874
rect 32460 6868 32628 6870
rect 32460 6816 32476 6868
rect 32528 6842 32628 6868
rect 32528 6816 32536 6842
rect 32460 6810 32536 6816
rect 31945 6600 32196 6628
rect 31884 6592 32196 6600
rect 31440 6212 31508 6240
rect 31440 6090 31468 6212
rect 31402 6084 31468 6090
rect 31402 6032 31408 6084
rect 31460 6032 31468 6084
rect 31402 6026 31468 6032
rect 32168 5966 32196 6592
rect 32268 6436 32536 6442
rect 32268 6414 32476 6436
rect 32268 6356 32296 6414
rect 32470 6384 32476 6414
rect 32528 6384 32536 6436
rect 32470 6378 32536 6384
rect 32232 6348 32296 6356
rect 32232 6296 32238 6348
rect 32290 6296 32296 6348
rect 32232 6288 32296 6296
rect 31468 5960 32196 5966
rect 31462 5958 32196 5960
rect 31404 5951 32196 5958
rect 31404 5899 31410 5951
rect 31462 5930 32196 5951
rect 31462 5899 31468 5930
rect 31404 5892 31468 5899
rect 31280 5716 31348 5726
rect 32600 5724 32628 6842
rect 32806 6598 32856 7004
rect 33108 6900 33162 6916
rect 33108 6860 33109 6900
rect 32948 6848 33109 6860
rect 33161 6848 33162 6900
rect 32948 6832 33162 6848
rect 33332 6890 33396 6906
rect 33332 6838 33341 6890
rect 33393 6838 33396 6890
rect 32806 6590 32872 6598
rect 32806 6538 32814 6590
rect 32866 6538 32872 6590
rect 32806 6530 32872 6538
rect 32948 6326 32976 6832
rect 33332 6824 33396 6838
rect 33018 6456 33084 6464
rect 33018 6404 33026 6456
rect 33078 6422 33084 6456
rect 33078 6404 33300 6422
rect 33018 6398 33300 6404
rect 33056 6394 33300 6398
rect 33272 6348 33300 6394
rect 33272 6342 33334 6348
rect 32948 6298 33236 6326
rect 32912 6212 32948 6214
rect 32912 6200 32984 6212
rect 32912 6148 32922 6200
rect 32974 6148 32984 6200
rect 32912 6136 32984 6148
rect 32788 6006 32854 6012
rect 32788 5954 32794 6006
rect 32846 5960 32854 6006
rect 32846 5954 33180 5960
rect 32788 5951 33180 5954
rect 32788 5948 33122 5951
rect 32802 5932 33122 5948
rect 31280 5664 31288 5716
rect 31340 5664 31348 5716
rect 31280 5658 31348 5664
rect 32354 5718 32628 5724
rect 32354 5666 32360 5718
rect 32412 5696 32628 5718
rect 32412 5666 32418 5696
rect 32354 5660 32418 5666
rect 31190 5604 31258 5610
rect 31190 5552 31196 5604
rect 31248 5552 31258 5604
rect 31190 5546 31258 5552
rect 32266 5602 32330 5608
rect 32266 5550 32272 5602
rect 32324 5564 32330 5602
rect 32324 5550 32332 5564
rect 30916 5534 30982 5542
rect 30916 5482 30924 5534
rect 30976 5482 30982 5534
rect 30916 5474 30982 5482
rect 31190 5440 31218 5546
rect 32266 5544 32332 5550
rect 32304 5440 32332 5544
rect 32804 5542 32854 5932
rect 33116 5899 33122 5932
rect 33174 5899 33180 5951
rect 33116 5892 33180 5899
rect 33208 5726 33236 6298
rect 33324 6290 33334 6342
rect 33272 6284 33334 6290
rect 33368 6240 33396 6824
rect 33486 6654 33536 7270
rect 33580 7260 33601 7376
rect 33909 7260 33930 7376
rect 35468 7376 35818 7390
rect 33580 7246 33930 7260
rect 34678 7062 34744 7068
rect 34678 7060 34684 7062
rect 34056 7032 34684 7060
rect 33468 6648 33536 6654
rect 33468 6596 33477 6648
rect 33529 6596 33536 6648
rect 33468 6590 33536 6596
rect 33772 6652 33852 6664
rect 33772 6600 33781 6652
rect 33833 6628 33852 6652
rect 34056 6628 34084 7032
rect 34678 7010 34684 7032
rect 34736 7010 34744 7062
rect 34678 7004 34744 7010
rect 34348 6870 34424 6874
rect 34348 6868 34516 6870
rect 34348 6816 34364 6868
rect 34416 6842 34516 6868
rect 34416 6816 34424 6842
rect 34348 6810 34424 6816
rect 33833 6600 34084 6628
rect 33772 6592 34084 6600
rect 33328 6212 33396 6240
rect 33328 6090 33356 6212
rect 33290 6084 33356 6090
rect 33290 6032 33296 6084
rect 33348 6032 33356 6084
rect 33290 6026 33356 6032
rect 34056 5966 34084 6592
rect 34156 6436 34424 6442
rect 34156 6414 34364 6436
rect 34156 6356 34184 6414
rect 34358 6384 34364 6414
rect 34416 6384 34424 6436
rect 34358 6378 34424 6384
rect 34120 6348 34184 6356
rect 34120 6296 34126 6348
rect 34178 6296 34184 6348
rect 34120 6288 34184 6296
rect 33356 5960 34084 5966
rect 33350 5958 34084 5960
rect 33292 5951 34084 5958
rect 33292 5899 33298 5951
rect 33350 5930 34084 5951
rect 33350 5899 33356 5930
rect 33292 5892 33356 5899
rect 33168 5716 33236 5726
rect 34488 5724 34516 6842
rect 34694 6598 34744 7004
rect 34996 6900 35050 6916
rect 34996 6860 34997 6900
rect 34836 6848 34997 6860
rect 35049 6848 35050 6900
rect 34836 6832 35050 6848
rect 35220 6890 35284 6906
rect 35220 6838 35229 6890
rect 35281 6838 35284 6890
rect 34694 6590 34760 6598
rect 34694 6538 34702 6590
rect 34754 6538 34760 6590
rect 34694 6530 34760 6538
rect 34836 6326 34864 6832
rect 35220 6824 35284 6838
rect 34906 6456 34972 6464
rect 34906 6404 34914 6456
rect 34966 6422 34972 6456
rect 34966 6404 35188 6422
rect 34906 6398 35188 6404
rect 34944 6394 35188 6398
rect 35160 6348 35188 6394
rect 35160 6342 35222 6348
rect 34836 6298 35124 6326
rect 34800 6212 34836 6214
rect 34800 6200 34872 6212
rect 34800 6148 34810 6200
rect 34862 6148 34872 6200
rect 34800 6136 34872 6148
rect 34676 6006 34742 6012
rect 34676 5954 34682 6006
rect 34734 5960 34742 6006
rect 34734 5954 35068 5960
rect 34676 5951 35068 5954
rect 34676 5948 35010 5951
rect 34690 5932 35010 5948
rect 33168 5664 33176 5716
rect 33228 5664 33236 5716
rect 33168 5658 33236 5664
rect 34242 5718 34516 5724
rect 34242 5666 34248 5718
rect 34300 5696 34516 5718
rect 34300 5666 34306 5696
rect 34242 5660 34306 5666
rect 33078 5604 33146 5610
rect 33078 5552 33084 5604
rect 33136 5552 33146 5604
rect 33078 5546 33146 5552
rect 34154 5602 34218 5608
rect 34154 5550 34160 5602
rect 34212 5564 34218 5602
rect 34212 5550 34220 5564
rect 32804 5534 32870 5542
rect 32804 5482 32812 5534
rect 32864 5482 32870 5534
rect 32804 5474 32870 5482
rect 33078 5440 33106 5546
rect 34154 5544 34220 5550
rect 34192 5440 34220 5544
rect 34692 5542 34742 5932
rect 35004 5899 35010 5932
rect 35062 5899 35068 5951
rect 35004 5892 35068 5899
rect 35096 5726 35124 6298
rect 35212 6290 35222 6342
rect 35160 6284 35222 6290
rect 35256 6240 35284 6824
rect 35374 6654 35424 7270
rect 35468 7260 35489 7376
rect 35797 7260 35818 7376
rect 37356 7376 37706 7390
rect 35468 7246 35818 7260
rect 36566 7062 36632 7068
rect 36566 7060 36572 7062
rect 35944 7032 36572 7060
rect 35356 6648 35424 6654
rect 35356 6596 35365 6648
rect 35417 6596 35424 6648
rect 35356 6590 35424 6596
rect 35660 6652 35740 6664
rect 35660 6600 35669 6652
rect 35721 6628 35740 6652
rect 35944 6628 35972 7032
rect 36566 7010 36572 7032
rect 36624 7010 36632 7062
rect 36566 7004 36632 7010
rect 36236 6870 36312 6874
rect 36236 6868 36404 6870
rect 36236 6816 36252 6868
rect 36304 6842 36404 6868
rect 36304 6816 36312 6842
rect 36236 6810 36312 6816
rect 35721 6600 35972 6628
rect 35660 6592 35972 6600
rect 35216 6212 35284 6240
rect 35216 6090 35244 6212
rect 35178 6084 35244 6090
rect 35178 6032 35184 6084
rect 35236 6032 35244 6084
rect 35178 6026 35244 6032
rect 35944 5966 35972 6592
rect 36044 6436 36312 6442
rect 36044 6414 36252 6436
rect 36044 6356 36072 6414
rect 36246 6384 36252 6414
rect 36304 6384 36312 6436
rect 36246 6378 36312 6384
rect 36008 6348 36072 6356
rect 36008 6296 36014 6348
rect 36066 6296 36072 6348
rect 36008 6288 36072 6296
rect 35244 5960 35972 5966
rect 35238 5958 35972 5960
rect 35180 5951 35972 5958
rect 35180 5899 35186 5951
rect 35238 5930 35972 5951
rect 35238 5899 35244 5930
rect 35180 5892 35244 5899
rect 35056 5716 35124 5726
rect 36376 5724 36404 6842
rect 36582 6598 36632 7004
rect 36884 6900 36938 6916
rect 36884 6860 36885 6900
rect 36724 6848 36885 6860
rect 36937 6848 36938 6900
rect 36724 6832 36938 6848
rect 37108 6890 37172 6906
rect 37108 6838 37117 6890
rect 37169 6838 37172 6890
rect 36582 6590 36648 6598
rect 36582 6538 36590 6590
rect 36642 6538 36648 6590
rect 36582 6530 36648 6538
rect 36724 6326 36752 6832
rect 37108 6824 37172 6838
rect 36794 6456 36860 6464
rect 36794 6404 36802 6456
rect 36854 6422 36860 6456
rect 36854 6404 37076 6422
rect 36794 6398 37076 6404
rect 36832 6394 37076 6398
rect 37048 6348 37076 6394
rect 37048 6342 37110 6348
rect 36724 6298 37012 6326
rect 36688 6212 36724 6214
rect 36688 6200 36760 6212
rect 36688 6148 36698 6200
rect 36750 6148 36760 6200
rect 36688 6136 36760 6148
rect 36564 6006 36630 6012
rect 36564 5954 36570 6006
rect 36622 5960 36630 6006
rect 36622 5954 36956 5960
rect 36564 5951 36956 5954
rect 36564 5948 36898 5951
rect 36578 5932 36898 5948
rect 35056 5664 35064 5716
rect 35116 5664 35124 5716
rect 35056 5658 35124 5664
rect 36130 5718 36404 5724
rect 36130 5666 36136 5718
rect 36188 5696 36404 5718
rect 36188 5666 36194 5696
rect 36130 5660 36194 5666
rect 34966 5604 35034 5610
rect 34966 5552 34972 5604
rect 35024 5552 35034 5604
rect 34966 5546 35034 5552
rect 36042 5602 36106 5608
rect 36042 5550 36048 5602
rect 36100 5564 36106 5602
rect 36100 5550 36108 5564
rect 34692 5534 34758 5542
rect 34692 5482 34700 5534
rect 34752 5482 34758 5534
rect 34692 5474 34758 5482
rect 34966 5440 34994 5546
rect 36042 5544 36108 5550
rect 36080 5444 36108 5544
rect 36580 5542 36630 5932
rect 36892 5899 36898 5932
rect 36950 5899 36956 5951
rect 36892 5892 36956 5899
rect 36984 5726 37012 6298
rect 37100 6290 37110 6342
rect 37048 6284 37110 6290
rect 37144 6240 37172 6824
rect 37262 6654 37312 7270
rect 37356 7260 37377 7376
rect 37685 7260 37706 7376
rect 39244 7376 39594 7390
rect 37356 7246 37706 7260
rect 38454 7062 38520 7068
rect 38454 7060 38460 7062
rect 37832 7032 38460 7060
rect 37244 6648 37312 6654
rect 37244 6596 37253 6648
rect 37305 6596 37312 6648
rect 37244 6590 37312 6596
rect 37548 6652 37628 6664
rect 37548 6600 37557 6652
rect 37609 6628 37628 6652
rect 37832 6628 37860 7032
rect 38454 7010 38460 7032
rect 38512 7010 38520 7062
rect 38454 7004 38520 7010
rect 38124 6870 38200 6874
rect 38124 6868 38292 6870
rect 38124 6816 38140 6868
rect 38192 6842 38292 6868
rect 38192 6816 38200 6842
rect 38124 6810 38200 6816
rect 37609 6600 37860 6628
rect 37548 6592 37860 6600
rect 37104 6212 37172 6240
rect 37104 6090 37132 6212
rect 37066 6084 37132 6090
rect 37066 6032 37072 6084
rect 37124 6032 37132 6084
rect 37066 6026 37132 6032
rect 37832 5966 37860 6592
rect 37932 6436 38200 6442
rect 37932 6414 38140 6436
rect 37932 6356 37960 6414
rect 38134 6384 38140 6414
rect 38192 6384 38200 6436
rect 38134 6378 38200 6384
rect 37896 6348 37960 6356
rect 37896 6296 37902 6348
rect 37954 6296 37960 6348
rect 37896 6288 37960 6296
rect 37132 5960 37860 5966
rect 37126 5958 37860 5960
rect 37068 5951 37860 5958
rect 37068 5899 37074 5951
rect 37126 5930 37860 5951
rect 37126 5899 37132 5930
rect 37068 5892 37132 5899
rect 36944 5716 37012 5726
rect 38264 5724 38292 6842
rect 38470 6598 38520 7004
rect 38772 6900 38826 6916
rect 38772 6860 38773 6900
rect 38612 6848 38773 6860
rect 38825 6848 38826 6900
rect 38612 6832 38826 6848
rect 38996 6890 39060 6906
rect 38996 6838 39005 6890
rect 39057 6838 39060 6890
rect 38470 6590 38536 6598
rect 38470 6538 38478 6590
rect 38530 6538 38536 6590
rect 38470 6530 38536 6538
rect 38612 6326 38640 6832
rect 38996 6824 39060 6838
rect 38682 6456 38748 6464
rect 38682 6404 38690 6456
rect 38742 6422 38748 6456
rect 38742 6404 38964 6422
rect 38682 6398 38964 6404
rect 38720 6394 38964 6398
rect 38936 6348 38964 6394
rect 38936 6342 38998 6348
rect 38612 6298 38900 6326
rect 38576 6212 38612 6214
rect 38576 6200 38648 6212
rect 38576 6148 38586 6200
rect 38638 6148 38648 6200
rect 38576 6136 38648 6148
rect 38452 6006 38518 6012
rect 38452 5954 38458 6006
rect 38510 5960 38518 6006
rect 38510 5954 38844 5960
rect 38452 5951 38844 5954
rect 38452 5948 38786 5951
rect 38466 5932 38786 5948
rect 36944 5664 36952 5716
rect 37004 5664 37012 5716
rect 36944 5658 37012 5664
rect 38018 5718 38292 5724
rect 38018 5666 38024 5718
rect 38076 5696 38292 5718
rect 38076 5666 38082 5696
rect 38018 5660 38082 5666
rect 36854 5604 36922 5610
rect 36854 5552 36860 5604
rect 36912 5552 36922 5604
rect 36854 5546 36922 5552
rect 37930 5602 37994 5608
rect 37930 5550 37936 5602
rect 37988 5564 37994 5602
rect 37988 5550 37996 5564
rect 36580 5534 36646 5542
rect 36580 5482 36588 5534
rect 36640 5482 36646 5534
rect 36580 5474 36646 5482
rect 36854 5444 36882 5546
rect 37930 5544 37996 5550
rect 37968 5444 37996 5544
rect 38468 5542 38518 5932
rect 38780 5899 38786 5932
rect 38838 5899 38844 5951
rect 38780 5892 38844 5899
rect 38872 5726 38900 6298
rect 38988 6290 38998 6342
rect 38936 6284 38998 6290
rect 39032 6240 39060 6824
rect 39150 6654 39200 7270
rect 39244 7260 39265 7376
rect 39573 7260 39594 7376
rect 41132 7376 41482 7390
rect 39244 7246 39594 7260
rect 40342 7062 40408 7068
rect 40342 7060 40348 7062
rect 39720 7032 40348 7060
rect 39132 6648 39200 6654
rect 39132 6596 39141 6648
rect 39193 6596 39200 6648
rect 39132 6590 39200 6596
rect 39436 6652 39516 6664
rect 39436 6600 39445 6652
rect 39497 6628 39516 6652
rect 39720 6628 39748 7032
rect 40342 7010 40348 7032
rect 40400 7010 40408 7062
rect 40342 7004 40408 7010
rect 40012 6870 40088 6874
rect 40012 6868 40180 6870
rect 40012 6816 40028 6868
rect 40080 6842 40180 6868
rect 40080 6816 40088 6842
rect 40012 6810 40088 6816
rect 39497 6600 39748 6628
rect 39436 6592 39748 6600
rect 38992 6212 39060 6240
rect 38992 6090 39020 6212
rect 38954 6084 39020 6090
rect 38954 6032 38960 6084
rect 39012 6032 39020 6084
rect 38954 6026 39020 6032
rect 39720 5966 39748 6592
rect 39820 6436 40088 6442
rect 39820 6414 40028 6436
rect 39820 6356 39848 6414
rect 40022 6384 40028 6414
rect 40080 6384 40088 6436
rect 40022 6378 40088 6384
rect 39784 6348 39848 6356
rect 39784 6296 39790 6348
rect 39842 6296 39848 6348
rect 39784 6288 39848 6296
rect 39020 5960 39748 5966
rect 39014 5958 39748 5960
rect 38956 5951 39748 5958
rect 38956 5899 38962 5951
rect 39014 5930 39748 5951
rect 39014 5899 39020 5930
rect 38956 5892 39020 5899
rect 38832 5716 38900 5726
rect 40152 5724 40180 6842
rect 40358 6598 40408 7004
rect 40660 6900 40714 6916
rect 40660 6860 40661 6900
rect 40500 6848 40661 6860
rect 40713 6848 40714 6900
rect 40500 6832 40714 6848
rect 40884 6890 40948 6906
rect 40884 6838 40893 6890
rect 40945 6838 40948 6890
rect 40358 6590 40424 6598
rect 40358 6538 40366 6590
rect 40418 6538 40424 6590
rect 40358 6530 40424 6538
rect 40500 6326 40528 6832
rect 40884 6824 40948 6838
rect 40570 6456 40636 6464
rect 40570 6404 40578 6456
rect 40630 6422 40636 6456
rect 40630 6404 40852 6422
rect 40570 6398 40852 6404
rect 40608 6394 40852 6398
rect 40824 6348 40852 6394
rect 40824 6342 40886 6348
rect 40500 6298 40788 6326
rect 40464 6212 40500 6214
rect 40464 6200 40536 6212
rect 40464 6148 40474 6200
rect 40526 6148 40536 6200
rect 40464 6136 40536 6148
rect 40340 6006 40406 6012
rect 40340 5954 40346 6006
rect 40398 5960 40406 6006
rect 40398 5954 40732 5960
rect 40340 5951 40732 5954
rect 40340 5948 40674 5951
rect 40354 5932 40674 5948
rect 38832 5664 38840 5716
rect 38892 5664 38900 5716
rect 38832 5658 38900 5664
rect 39906 5718 40180 5724
rect 39906 5666 39912 5718
rect 39964 5696 40180 5718
rect 39964 5666 39970 5696
rect 39906 5660 39970 5666
rect 38742 5604 38810 5610
rect 38742 5552 38748 5604
rect 38800 5552 38810 5604
rect 38742 5546 38810 5552
rect 39818 5602 39882 5608
rect 39818 5550 39824 5602
rect 39876 5564 39882 5602
rect 39876 5550 39884 5564
rect 38468 5534 38534 5542
rect 38468 5482 38476 5534
rect 38528 5482 38534 5534
rect 38468 5474 38534 5482
rect 38742 5444 38770 5546
rect 39818 5544 39884 5550
rect 35974 5440 37298 5444
rect 37862 5440 39182 5444
rect 39856 5440 39884 5544
rect 40356 5542 40406 5932
rect 40668 5899 40674 5932
rect 40726 5899 40732 5951
rect 40668 5892 40732 5899
rect 40760 5726 40788 6298
rect 40876 6290 40886 6342
rect 40824 6284 40886 6290
rect 40920 6240 40948 6824
rect 41038 6654 41088 7270
rect 41132 7260 41153 7376
rect 41461 7260 41482 7376
rect 43020 7376 43370 7390
rect 41132 7246 41482 7260
rect 42230 7062 42296 7068
rect 42230 7060 42236 7062
rect 41608 7032 42236 7060
rect 41020 6648 41088 6654
rect 41020 6596 41029 6648
rect 41081 6596 41088 6648
rect 41020 6590 41088 6596
rect 41324 6652 41404 6664
rect 41324 6600 41333 6652
rect 41385 6628 41404 6652
rect 41608 6628 41636 7032
rect 42230 7010 42236 7032
rect 42288 7010 42296 7062
rect 42230 7004 42296 7010
rect 41900 6870 41976 6874
rect 41900 6868 42068 6870
rect 41900 6816 41916 6868
rect 41968 6842 42068 6868
rect 41968 6816 41976 6842
rect 41900 6810 41976 6816
rect 41385 6600 41636 6628
rect 41324 6592 41636 6600
rect 40880 6212 40948 6240
rect 40880 6090 40908 6212
rect 40842 6084 40908 6090
rect 40842 6032 40848 6084
rect 40900 6032 40908 6084
rect 40842 6026 40908 6032
rect 41608 5966 41636 6592
rect 41708 6436 41976 6442
rect 41708 6414 41916 6436
rect 41708 6356 41736 6414
rect 41910 6384 41916 6414
rect 41968 6384 41976 6436
rect 41910 6378 41976 6384
rect 41672 6348 41736 6356
rect 41672 6296 41678 6348
rect 41730 6296 41736 6348
rect 41672 6288 41736 6296
rect 40908 5960 41636 5966
rect 40902 5958 41636 5960
rect 40844 5951 41636 5958
rect 40844 5899 40850 5951
rect 40902 5930 41636 5951
rect 40902 5899 40908 5930
rect 40844 5892 40908 5899
rect 40720 5716 40788 5726
rect 42040 5724 42068 6842
rect 42246 6598 42296 7004
rect 42548 6900 42602 6916
rect 42548 6860 42549 6900
rect 42388 6848 42549 6860
rect 42601 6848 42602 6900
rect 42388 6832 42602 6848
rect 42772 6890 42836 6906
rect 42772 6838 42781 6890
rect 42833 6838 42836 6890
rect 42246 6590 42312 6598
rect 42246 6538 42254 6590
rect 42306 6538 42312 6590
rect 42246 6530 42312 6538
rect 42388 6326 42416 6832
rect 42772 6824 42836 6838
rect 42458 6456 42524 6464
rect 42458 6404 42466 6456
rect 42518 6422 42524 6456
rect 42518 6404 42740 6422
rect 42458 6398 42740 6404
rect 42496 6394 42740 6398
rect 42712 6348 42740 6394
rect 42712 6342 42774 6348
rect 42388 6298 42676 6326
rect 42352 6212 42388 6214
rect 42352 6200 42424 6212
rect 42352 6148 42362 6200
rect 42414 6148 42424 6200
rect 42352 6136 42424 6148
rect 42228 6006 42294 6012
rect 42228 5954 42234 6006
rect 42286 5960 42294 6006
rect 42286 5954 42620 5960
rect 42228 5951 42620 5954
rect 42228 5948 42562 5951
rect 42242 5932 42562 5948
rect 40720 5664 40728 5716
rect 40780 5664 40788 5716
rect 40720 5658 40788 5664
rect 41794 5718 42068 5724
rect 41794 5666 41800 5718
rect 41852 5696 42068 5718
rect 41852 5666 41858 5696
rect 41794 5660 41858 5666
rect 40630 5604 40698 5610
rect 40630 5552 40636 5604
rect 40688 5552 40698 5604
rect 40630 5546 40698 5552
rect 41706 5602 41770 5608
rect 41706 5550 41712 5602
rect 41764 5564 41770 5602
rect 41764 5550 41772 5564
rect 40356 5534 40422 5542
rect 40356 5482 40364 5534
rect 40416 5482 40422 5534
rect 40356 5474 40422 5482
rect 40630 5440 40658 5546
rect 41706 5544 41772 5550
rect 41744 5440 41772 5544
rect 42244 5542 42294 5932
rect 42556 5899 42562 5932
rect 42614 5899 42620 5951
rect 42556 5892 42620 5899
rect 42648 5726 42676 6298
rect 42764 6290 42774 6342
rect 42712 6284 42774 6290
rect 42808 6240 42836 6824
rect 42926 6654 42976 7270
rect 43020 7260 43041 7376
rect 43349 7260 43370 7376
rect 44902 7376 45252 7390
rect 43020 7246 43370 7260
rect 44118 7062 44184 7068
rect 44118 7060 44124 7062
rect 43496 7032 44124 7060
rect 42908 6648 42976 6654
rect 42908 6596 42917 6648
rect 42969 6596 42976 6648
rect 42908 6590 42976 6596
rect 43212 6652 43292 6664
rect 43212 6600 43221 6652
rect 43273 6628 43292 6652
rect 43496 6628 43524 7032
rect 44118 7010 44124 7032
rect 44176 7010 44184 7062
rect 44118 7004 44184 7010
rect 43788 6870 43864 6874
rect 43788 6868 43956 6870
rect 43788 6816 43804 6868
rect 43856 6842 43956 6868
rect 43856 6816 43864 6842
rect 43788 6810 43864 6816
rect 43273 6600 43524 6628
rect 43212 6592 43524 6600
rect 42768 6212 42836 6240
rect 42768 6090 42796 6212
rect 42730 6084 42796 6090
rect 42730 6032 42736 6084
rect 42788 6032 42796 6084
rect 42730 6026 42796 6032
rect 43496 5966 43524 6592
rect 43596 6436 43864 6442
rect 43596 6414 43804 6436
rect 43596 6356 43624 6414
rect 43798 6384 43804 6414
rect 43856 6384 43864 6436
rect 43798 6378 43864 6384
rect 43560 6348 43624 6356
rect 43560 6296 43566 6348
rect 43618 6296 43624 6348
rect 43560 6288 43624 6296
rect 42796 5960 43524 5966
rect 42790 5958 43524 5960
rect 42732 5951 43524 5958
rect 42732 5899 42738 5951
rect 42790 5930 43524 5951
rect 42790 5899 42796 5930
rect 42732 5892 42796 5899
rect 42608 5716 42676 5726
rect 43928 5724 43956 6842
rect 44134 6598 44184 7004
rect 44436 6900 44490 6916
rect 44436 6860 44437 6900
rect 44276 6848 44437 6860
rect 44489 6848 44490 6900
rect 44276 6832 44490 6848
rect 44660 6890 44724 6906
rect 44660 6838 44669 6890
rect 44721 6838 44724 6890
rect 44134 6590 44200 6598
rect 44134 6538 44142 6590
rect 44194 6538 44200 6590
rect 44134 6530 44200 6538
rect 44276 6326 44304 6832
rect 44660 6824 44724 6838
rect 44346 6456 44412 6464
rect 44346 6404 44354 6456
rect 44406 6422 44412 6456
rect 44406 6404 44628 6422
rect 44346 6398 44628 6404
rect 44384 6394 44628 6398
rect 44600 6348 44628 6394
rect 44600 6342 44662 6348
rect 44276 6298 44564 6326
rect 44240 6212 44276 6214
rect 44240 6200 44312 6212
rect 44240 6148 44250 6200
rect 44302 6148 44312 6200
rect 44240 6136 44312 6148
rect 44116 6006 44182 6012
rect 44116 5954 44122 6006
rect 44174 5960 44182 6006
rect 44174 5954 44508 5960
rect 44116 5951 44508 5954
rect 44116 5948 44450 5951
rect 44130 5932 44450 5948
rect 42608 5664 42616 5716
rect 42668 5664 42676 5716
rect 42608 5658 42676 5664
rect 43682 5718 43956 5724
rect 43682 5666 43688 5718
rect 43740 5696 43956 5718
rect 43740 5666 43746 5696
rect 43682 5660 43746 5666
rect 42518 5604 42586 5610
rect 42518 5552 42524 5604
rect 42576 5552 42586 5604
rect 42518 5546 42586 5552
rect 43594 5602 43658 5608
rect 43594 5550 43600 5602
rect 43652 5564 43658 5602
rect 43652 5550 43660 5564
rect 42244 5534 42310 5542
rect 42244 5482 42252 5534
rect 42304 5482 42310 5534
rect 42244 5474 42310 5482
rect 42518 5440 42546 5546
rect 43594 5544 43660 5550
rect 43632 5440 43660 5544
rect 44132 5542 44182 5932
rect 44444 5899 44450 5932
rect 44502 5899 44508 5951
rect 44444 5892 44508 5899
rect 44536 5726 44564 6298
rect 44652 6290 44662 6342
rect 44600 6284 44662 6290
rect 44696 6240 44724 6824
rect 44814 6654 44864 7270
rect 44902 7260 44923 7376
rect 45231 7260 45252 7376
rect 46790 7376 47140 7390
rect 44902 7246 45252 7260
rect 46000 7062 46066 7068
rect 46000 7060 46006 7062
rect 45378 7032 46006 7060
rect 44796 6648 44864 6654
rect 44796 6596 44805 6648
rect 44857 6596 44864 6648
rect 44796 6590 44864 6596
rect 45094 6652 45174 6664
rect 45094 6600 45103 6652
rect 45155 6628 45174 6652
rect 45378 6628 45406 7032
rect 46000 7010 46006 7032
rect 46058 7010 46066 7062
rect 46000 7004 46066 7010
rect 45670 6870 45746 6874
rect 45670 6868 45838 6870
rect 45670 6816 45686 6868
rect 45738 6842 45838 6868
rect 45738 6816 45746 6842
rect 45670 6810 45746 6816
rect 45155 6600 45406 6628
rect 45094 6592 45406 6600
rect 44656 6212 44724 6240
rect 44656 6090 44684 6212
rect 44618 6084 44684 6090
rect 44618 6032 44624 6084
rect 44676 6032 44684 6084
rect 44618 6026 44684 6032
rect 45378 5966 45406 6592
rect 45478 6436 45746 6442
rect 45478 6414 45686 6436
rect 45478 6356 45506 6414
rect 45680 6384 45686 6414
rect 45738 6384 45746 6436
rect 45680 6378 45746 6384
rect 45442 6348 45506 6356
rect 45442 6296 45448 6348
rect 45500 6296 45506 6348
rect 45442 6288 45506 6296
rect 44684 5960 45406 5966
rect 44678 5958 45406 5960
rect 44620 5951 45406 5958
rect 44620 5899 44626 5951
rect 44678 5930 45406 5951
rect 44678 5899 44684 5930
rect 44620 5892 44684 5899
rect 44496 5716 44564 5726
rect 45810 5724 45838 6842
rect 46016 6598 46066 7004
rect 46318 6900 46372 6916
rect 46318 6860 46319 6900
rect 46158 6848 46319 6860
rect 46371 6848 46372 6900
rect 46158 6832 46372 6848
rect 46542 6890 46606 6906
rect 46542 6838 46551 6890
rect 46603 6838 46606 6890
rect 46016 6590 46082 6598
rect 46016 6538 46024 6590
rect 46076 6538 46082 6590
rect 46016 6530 46082 6538
rect 46158 6326 46186 6832
rect 46542 6824 46606 6838
rect 46228 6456 46294 6464
rect 46228 6404 46236 6456
rect 46288 6422 46294 6456
rect 46288 6404 46510 6422
rect 46228 6398 46510 6404
rect 46266 6394 46510 6398
rect 46482 6348 46510 6394
rect 46482 6342 46544 6348
rect 46158 6298 46446 6326
rect 46122 6212 46158 6214
rect 46122 6200 46194 6212
rect 46122 6148 46132 6200
rect 46184 6148 46194 6200
rect 46122 6136 46194 6148
rect 45998 6006 46064 6012
rect 45998 5954 46004 6006
rect 46056 5960 46064 6006
rect 46056 5954 46390 5960
rect 45998 5951 46390 5954
rect 45998 5948 46332 5951
rect 46012 5932 46332 5948
rect 44496 5664 44504 5716
rect 44556 5664 44564 5716
rect 44496 5658 44564 5664
rect 45564 5718 45838 5724
rect 45564 5666 45570 5718
rect 45622 5696 45838 5718
rect 45622 5666 45628 5696
rect 45564 5660 45628 5666
rect 44406 5604 44474 5610
rect 44406 5552 44412 5604
rect 44464 5552 44474 5604
rect 44406 5546 44474 5552
rect 45476 5602 45540 5608
rect 45476 5550 45482 5602
rect 45534 5564 45540 5602
rect 45534 5550 45542 5564
rect 44132 5534 44198 5542
rect 44132 5482 44140 5534
rect 44192 5482 44198 5534
rect 44132 5474 44198 5482
rect 44406 5440 44434 5546
rect 45476 5544 45542 5550
rect 45514 5444 45542 5544
rect 46014 5542 46064 5932
rect 46326 5899 46332 5932
rect 46384 5899 46390 5951
rect 46326 5892 46390 5899
rect 46418 5726 46446 6298
rect 46534 6290 46544 6342
rect 46482 6284 46544 6290
rect 46578 6240 46606 6824
rect 46702 6654 46746 7270
rect 46790 7260 46811 7376
rect 47119 7260 47140 7376
rect 48678 7376 49028 7390
rect 46790 7246 47140 7260
rect 47888 7062 47954 7068
rect 47888 7060 47894 7062
rect 47266 7032 47894 7060
rect 46678 6648 46746 6654
rect 46678 6596 46687 6648
rect 46739 6596 46746 6648
rect 46678 6590 46746 6596
rect 46982 6652 47062 6664
rect 46982 6600 46991 6652
rect 47043 6628 47062 6652
rect 47266 6628 47294 7032
rect 47888 7010 47894 7032
rect 47946 7010 47954 7062
rect 47888 7004 47954 7010
rect 47558 6870 47634 6874
rect 47558 6868 47726 6870
rect 47558 6816 47574 6868
rect 47626 6842 47726 6868
rect 47626 6816 47634 6842
rect 47558 6810 47634 6816
rect 47043 6600 47294 6628
rect 46982 6592 47294 6600
rect 46538 6212 46606 6240
rect 46538 6090 46566 6212
rect 46500 6084 46566 6090
rect 46500 6032 46506 6084
rect 46558 6032 46566 6084
rect 46500 6026 46566 6032
rect 47266 5966 47294 6592
rect 47366 6436 47634 6442
rect 47366 6414 47574 6436
rect 47366 6356 47394 6414
rect 47568 6384 47574 6414
rect 47626 6384 47634 6436
rect 47568 6378 47634 6384
rect 47330 6348 47394 6356
rect 47330 6296 47336 6348
rect 47388 6296 47394 6348
rect 47330 6288 47394 6296
rect 46566 5960 47294 5966
rect 46560 5958 47294 5960
rect 46502 5951 47294 5958
rect 46502 5899 46508 5951
rect 46560 5930 47294 5951
rect 46560 5899 46566 5930
rect 46502 5892 46566 5899
rect 46378 5716 46446 5726
rect 47698 5724 47726 6842
rect 47904 6598 47954 7004
rect 48206 6900 48260 6916
rect 48206 6860 48207 6900
rect 48046 6848 48207 6860
rect 48259 6848 48260 6900
rect 48046 6832 48260 6848
rect 48430 6890 48494 6906
rect 48430 6838 48439 6890
rect 48491 6838 48494 6890
rect 47904 6590 47970 6598
rect 47904 6538 47912 6590
rect 47964 6538 47970 6590
rect 47904 6530 47970 6538
rect 48046 6326 48074 6832
rect 48430 6824 48494 6838
rect 48116 6456 48182 6464
rect 48116 6404 48124 6456
rect 48176 6422 48182 6456
rect 48176 6404 48398 6422
rect 48116 6398 48398 6404
rect 48154 6394 48398 6398
rect 48370 6348 48398 6394
rect 48370 6342 48432 6348
rect 48046 6298 48334 6326
rect 48010 6212 48046 6214
rect 48010 6200 48082 6212
rect 48010 6148 48020 6200
rect 48072 6148 48082 6200
rect 48010 6136 48082 6148
rect 47886 6006 47952 6012
rect 47886 5954 47892 6006
rect 47944 5960 47952 6006
rect 47944 5954 48278 5960
rect 47886 5951 48278 5954
rect 47886 5948 48220 5951
rect 47900 5932 48220 5948
rect 46378 5664 46386 5716
rect 46438 5664 46446 5716
rect 46378 5658 46446 5664
rect 47452 5718 47726 5724
rect 47452 5666 47458 5718
rect 47510 5696 47726 5718
rect 47510 5666 47516 5696
rect 47452 5660 47516 5666
rect 46288 5604 46356 5610
rect 46288 5552 46294 5604
rect 46346 5552 46356 5604
rect 46288 5546 46356 5552
rect 47364 5602 47428 5608
rect 47364 5550 47370 5602
rect 47422 5564 47428 5602
rect 47422 5550 47430 5564
rect 46014 5534 46080 5542
rect 46014 5482 46022 5534
rect 46074 5482 46080 5534
rect 46014 5474 46080 5482
rect 46288 5444 46316 5546
rect 47364 5544 47430 5550
rect 47402 5444 47430 5544
rect 47902 5542 47952 5932
rect 48214 5899 48220 5932
rect 48272 5899 48278 5951
rect 48214 5892 48278 5899
rect 48306 5726 48334 6298
rect 48422 6290 48432 6342
rect 48370 6284 48432 6290
rect 48466 6240 48494 6824
rect 48590 6654 48634 7270
rect 48678 7260 48699 7376
rect 49007 7260 49028 7376
rect 50566 7376 50916 7390
rect 48678 7246 49028 7260
rect 49776 7062 49842 7068
rect 49776 7060 49782 7062
rect 49154 7032 49782 7060
rect 48566 6648 48634 6654
rect 48566 6596 48575 6648
rect 48627 6596 48634 6648
rect 48566 6590 48634 6596
rect 48870 6652 48950 6664
rect 48870 6600 48879 6652
rect 48931 6628 48950 6652
rect 49154 6628 49182 7032
rect 49776 7010 49782 7032
rect 49834 7010 49842 7062
rect 49776 7004 49842 7010
rect 49446 6870 49522 6874
rect 49446 6868 49614 6870
rect 49446 6816 49462 6868
rect 49514 6842 49614 6868
rect 49514 6816 49522 6842
rect 49446 6810 49522 6816
rect 48931 6600 49182 6628
rect 48870 6592 49182 6600
rect 48426 6212 48494 6240
rect 48426 6090 48454 6212
rect 48388 6084 48454 6090
rect 48388 6032 48394 6084
rect 48446 6032 48454 6084
rect 48388 6026 48454 6032
rect 49154 5966 49182 6592
rect 49254 6436 49522 6442
rect 49254 6414 49462 6436
rect 49254 6356 49282 6414
rect 49456 6384 49462 6414
rect 49514 6384 49522 6436
rect 49456 6378 49522 6384
rect 49218 6348 49282 6356
rect 49218 6296 49224 6348
rect 49276 6296 49282 6348
rect 49218 6288 49282 6296
rect 48454 5960 49182 5966
rect 48448 5958 49182 5960
rect 48390 5951 49182 5958
rect 48390 5899 48396 5951
rect 48448 5930 49182 5951
rect 48448 5899 48454 5930
rect 48390 5892 48454 5899
rect 48266 5716 48334 5726
rect 49586 5724 49614 6842
rect 49792 6598 49842 7004
rect 50094 6900 50148 6916
rect 50094 6860 50095 6900
rect 49934 6848 50095 6860
rect 50147 6848 50148 6900
rect 49934 6832 50148 6848
rect 50318 6890 50382 6906
rect 50318 6838 50327 6890
rect 50379 6838 50382 6890
rect 49792 6590 49858 6598
rect 49792 6538 49800 6590
rect 49852 6538 49858 6590
rect 49792 6530 49858 6538
rect 49934 6326 49962 6832
rect 50318 6824 50382 6838
rect 50004 6456 50070 6464
rect 50004 6404 50012 6456
rect 50064 6422 50070 6456
rect 50064 6404 50286 6422
rect 50004 6398 50286 6404
rect 50042 6394 50286 6398
rect 50258 6348 50286 6394
rect 50258 6342 50320 6348
rect 49934 6298 50222 6326
rect 49898 6212 49934 6214
rect 49898 6200 49970 6212
rect 49898 6148 49908 6200
rect 49960 6148 49970 6200
rect 49898 6136 49970 6148
rect 49774 6006 49840 6012
rect 49774 5954 49780 6006
rect 49832 5960 49840 6006
rect 49832 5954 50166 5960
rect 49774 5951 50166 5954
rect 49774 5948 50108 5951
rect 49788 5932 50108 5948
rect 48266 5664 48274 5716
rect 48326 5664 48334 5716
rect 48266 5658 48334 5664
rect 49340 5718 49614 5724
rect 49340 5666 49346 5718
rect 49398 5696 49614 5718
rect 49398 5666 49404 5696
rect 49340 5660 49404 5666
rect 48176 5604 48244 5610
rect 48176 5552 48182 5604
rect 48234 5552 48244 5604
rect 48176 5546 48244 5552
rect 49252 5602 49316 5608
rect 49252 5550 49258 5602
rect 49310 5564 49316 5602
rect 49310 5550 49318 5564
rect 47902 5534 47968 5542
rect 47902 5482 47910 5534
rect 47962 5482 47968 5534
rect 47902 5474 47968 5482
rect 48176 5444 48204 5546
rect 49252 5544 49318 5550
rect 49290 5444 49318 5544
rect 49790 5542 49840 5932
rect 50102 5899 50108 5932
rect 50160 5899 50166 5951
rect 50102 5892 50166 5899
rect 50194 5726 50222 6298
rect 50310 6290 50320 6342
rect 50258 6284 50320 6290
rect 50354 6240 50382 6824
rect 50478 6654 50522 7270
rect 50566 7260 50587 7376
rect 50895 7260 50916 7376
rect 52454 7376 52804 7390
rect 50566 7246 50916 7260
rect 51664 7062 51730 7068
rect 51664 7060 51670 7062
rect 51042 7032 51670 7060
rect 50454 6648 50522 6654
rect 50454 6596 50463 6648
rect 50515 6596 50522 6648
rect 50454 6590 50522 6596
rect 50758 6652 50838 6664
rect 50758 6600 50767 6652
rect 50819 6628 50838 6652
rect 51042 6628 51070 7032
rect 51664 7010 51670 7032
rect 51722 7010 51730 7062
rect 51664 7004 51730 7010
rect 51334 6870 51410 6874
rect 51334 6868 51502 6870
rect 51334 6816 51350 6868
rect 51402 6842 51502 6868
rect 51402 6816 51410 6842
rect 51334 6810 51410 6816
rect 50819 6600 51070 6628
rect 50758 6592 51070 6600
rect 50314 6212 50382 6240
rect 50314 6090 50342 6212
rect 50276 6084 50342 6090
rect 50276 6032 50282 6084
rect 50334 6032 50342 6084
rect 50276 6026 50342 6032
rect 51042 5966 51070 6592
rect 51142 6436 51410 6442
rect 51142 6414 51350 6436
rect 51142 6356 51170 6414
rect 51344 6384 51350 6414
rect 51402 6384 51410 6436
rect 51344 6378 51410 6384
rect 51106 6348 51170 6356
rect 51106 6296 51112 6348
rect 51164 6296 51170 6348
rect 51106 6288 51170 6296
rect 50342 5960 51070 5966
rect 50336 5958 51070 5960
rect 50278 5951 51070 5958
rect 50278 5899 50284 5951
rect 50336 5930 51070 5951
rect 50336 5899 50342 5930
rect 50278 5892 50342 5899
rect 50154 5716 50222 5726
rect 51474 5724 51502 6842
rect 51680 6598 51730 7004
rect 51982 6900 52036 6916
rect 51982 6860 51983 6900
rect 51822 6848 51983 6860
rect 52035 6848 52036 6900
rect 51822 6832 52036 6848
rect 52206 6890 52270 6906
rect 52206 6838 52215 6890
rect 52267 6838 52270 6890
rect 51680 6590 51746 6598
rect 51680 6538 51688 6590
rect 51740 6538 51746 6590
rect 51680 6530 51746 6538
rect 51822 6326 51850 6832
rect 52206 6824 52270 6838
rect 51892 6456 51958 6464
rect 51892 6404 51900 6456
rect 51952 6422 51958 6456
rect 51952 6404 52174 6422
rect 51892 6398 52174 6404
rect 51930 6394 52174 6398
rect 52146 6348 52174 6394
rect 52146 6342 52208 6348
rect 51822 6298 52110 6326
rect 51786 6212 51822 6214
rect 51786 6200 51858 6212
rect 51786 6148 51796 6200
rect 51848 6148 51858 6200
rect 51786 6136 51858 6148
rect 51662 6006 51728 6012
rect 51662 5954 51668 6006
rect 51720 5960 51728 6006
rect 51720 5954 52054 5960
rect 51662 5951 52054 5954
rect 51662 5948 51996 5951
rect 51676 5932 51996 5948
rect 50154 5664 50162 5716
rect 50214 5664 50222 5716
rect 50154 5658 50222 5664
rect 51228 5718 51502 5724
rect 51228 5666 51234 5718
rect 51286 5696 51502 5718
rect 51286 5666 51292 5696
rect 51228 5660 51292 5666
rect 50064 5604 50132 5610
rect 50064 5552 50070 5604
rect 50122 5552 50132 5604
rect 50064 5546 50132 5552
rect 51140 5602 51204 5608
rect 51140 5550 51146 5602
rect 51198 5564 51204 5602
rect 51198 5550 51206 5564
rect 49790 5534 49856 5542
rect 49790 5482 49798 5534
rect 49850 5482 49856 5534
rect 49790 5474 49856 5482
rect 50064 5444 50092 5546
rect 51140 5544 51206 5550
rect 51178 5444 51206 5544
rect 51678 5542 51728 5932
rect 51990 5899 51996 5932
rect 52048 5899 52054 5951
rect 51990 5892 52054 5899
rect 52082 5726 52110 6298
rect 52198 6290 52208 6342
rect 52146 6284 52208 6290
rect 52242 6240 52270 6824
rect 52366 6654 52410 7270
rect 52454 7260 52475 7376
rect 52783 7260 52804 7376
rect 54342 7376 54692 7390
rect 52454 7246 52804 7260
rect 53552 7062 53618 7068
rect 53552 7060 53558 7062
rect 52930 7032 53558 7060
rect 52342 6648 52410 6654
rect 52342 6596 52351 6648
rect 52403 6596 52410 6648
rect 52342 6590 52410 6596
rect 52646 6652 52726 6664
rect 52646 6600 52655 6652
rect 52707 6628 52726 6652
rect 52930 6628 52958 7032
rect 53552 7010 53558 7032
rect 53610 7010 53618 7062
rect 53552 7004 53618 7010
rect 53222 6870 53298 6874
rect 53222 6868 53390 6870
rect 53222 6816 53238 6868
rect 53290 6842 53390 6868
rect 53290 6816 53298 6842
rect 53222 6810 53298 6816
rect 52707 6600 52958 6628
rect 52646 6592 52958 6600
rect 52202 6212 52270 6240
rect 52202 6090 52230 6212
rect 52164 6084 52230 6090
rect 52164 6032 52170 6084
rect 52222 6032 52230 6084
rect 52164 6026 52230 6032
rect 52930 5966 52958 6592
rect 53030 6436 53298 6442
rect 53030 6414 53238 6436
rect 53030 6356 53058 6414
rect 53232 6384 53238 6414
rect 53290 6384 53298 6436
rect 53232 6378 53298 6384
rect 52994 6348 53058 6356
rect 52994 6296 53000 6348
rect 53052 6296 53058 6348
rect 52994 6288 53058 6296
rect 52230 5960 52958 5966
rect 52224 5958 52958 5960
rect 52166 5951 52958 5958
rect 52166 5899 52172 5951
rect 52224 5930 52958 5951
rect 52224 5899 52230 5930
rect 52166 5892 52230 5899
rect 52042 5716 52110 5726
rect 53362 5724 53390 6842
rect 53568 6598 53618 7004
rect 53870 6900 53924 6916
rect 53870 6860 53871 6900
rect 53710 6848 53871 6860
rect 53923 6848 53924 6900
rect 53710 6832 53924 6848
rect 54094 6890 54158 6906
rect 54094 6838 54103 6890
rect 54155 6838 54158 6890
rect 53568 6590 53634 6598
rect 53568 6538 53576 6590
rect 53628 6538 53634 6590
rect 53568 6530 53634 6538
rect 53710 6326 53738 6832
rect 54094 6824 54158 6838
rect 53780 6456 53846 6464
rect 53780 6404 53788 6456
rect 53840 6422 53846 6456
rect 53840 6404 54062 6422
rect 53780 6398 54062 6404
rect 53818 6394 54062 6398
rect 54034 6348 54062 6394
rect 54034 6342 54096 6348
rect 53710 6298 53998 6326
rect 53674 6212 53710 6214
rect 53674 6200 53746 6212
rect 53674 6148 53684 6200
rect 53736 6148 53746 6200
rect 53674 6136 53746 6148
rect 53550 6006 53616 6012
rect 53550 5954 53556 6006
rect 53608 5960 53616 6006
rect 53608 5954 53942 5960
rect 53550 5951 53942 5954
rect 53550 5948 53884 5951
rect 53564 5932 53884 5948
rect 52042 5664 52050 5716
rect 52102 5664 52110 5716
rect 52042 5658 52110 5664
rect 53116 5718 53390 5724
rect 53116 5666 53122 5718
rect 53174 5696 53390 5718
rect 53174 5666 53180 5696
rect 53116 5660 53180 5666
rect 51952 5604 52020 5610
rect 51952 5552 51958 5604
rect 52010 5552 52020 5604
rect 51952 5546 52020 5552
rect 53028 5602 53092 5608
rect 53028 5550 53034 5602
rect 53086 5564 53092 5602
rect 53086 5550 53094 5564
rect 51678 5534 51744 5542
rect 51678 5482 51686 5534
rect 51738 5482 51744 5534
rect 51678 5474 51744 5482
rect 51952 5444 51980 5546
rect 53028 5544 53094 5550
rect 53066 5444 53094 5544
rect 53566 5542 53616 5932
rect 53878 5899 53884 5932
rect 53936 5899 53942 5951
rect 53878 5892 53942 5899
rect 53970 5726 53998 6298
rect 54086 6290 54096 6342
rect 54034 6284 54096 6290
rect 54130 6240 54158 6824
rect 54254 6654 54298 7270
rect 54342 7260 54363 7376
rect 54671 7260 54692 7376
rect 56230 7376 56580 7390
rect 54342 7246 54692 7260
rect 55440 7062 55506 7068
rect 55440 7060 55446 7062
rect 54818 7032 55446 7060
rect 54230 6648 54298 6654
rect 54230 6596 54239 6648
rect 54291 6596 54298 6648
rect 54230 6590 54298 6596
rect 54534 6652 54614 6664
rect 54534 6600 54543 6652
rect 54595 6628 54614 6652
rect 54818 6628 54846 7032
rect 55440 7010 55446 7032
rect 55498 7010 55506 7062
rect 55440 7004 55506 7010
rect 55110 6870 55186 6874
rect 55110 6868 55278 6870
rect 55110 6816 55126 6868
rect 55178 6842 55278 6868
rect 55178 6816 55186 6842
rect 55110 6810 55186 6816
rect 54595 6600 54846 6628
rect 54534 6592 54846 6600
rect 54090 6212 54158 6240
rect 54090 6090 54118 6212
rect 54052 6084 54118 6090
rect 54052 6032 54058 6084
rect 54110 6032 54118 6084
rect 54052 6026 54118 6032
rect 54818 5966 54846 6592
rect 54918 6436 55186 6442
rect 54918 6414 55126 6436
rect 54918 6356 54946 6414
rect 55120 6384 55126 6414
rect 55178 6384 55186 6436
rect 55120 6378 55186 6384
rect 54882 6348 54946 6356
rect 54882 6296 54888 6348
rect 54940 6296 54946 6348
rect 54882 6288 54946 6296
rect 54118 5960 54846 5966
rect 54112 5958 54846 5960
rect 54054 5951 54846 5958
rect 54054 5899 54060 5951
rect 54112 5930 54846 5951
rect 54112 5899 54118 5930
rect 54054 5892 54118 5899
rect 53930 5716 53998 5726
rect 55250 5724 55278 6842
rect 55456 6598 55506 7004
rect 55758 6900 55812 6916
rect 55758 6860 55759 6900
rect 55598 6848 55759 6860
rect 55811 6848 55812 6900
rect 55598 6832 55812 6848
rect 55982 6890 56046 6906
rect 55982 6838 55991 6890
rect 56043 6838 56046 6890
rect 55456 6590 55522 6598
rect 55456 6538 55464 6590
rect 55516 6538 55522 6590
rect 55456 6530 55522 6538
rect 55598 6326 55626 6832
rect 55982 6824 56046 6838
rect 55668 6456 55734 6464
rect 55668 6404 55676 6456
rect 55728 6422 55734 6456
rect 55728 6404 55950 6422
rect 55668 6398 55950 6404
rect 55706 6394 55950 6398
rect 55922 6348 55950 6394
rect 55922 6342 55984 6348
rect 55598 6298 55886 6326
rect 55562 6212 55598 6214
rect 55562 6200 55634 6212
rect 55562 6148 55572 6200
rect 55624 6148 55634 6200
rect 55562 6136 55634 6148
rect 55438 6006 55504 6012
rect 55438 5954 55444 6006
rect 55496 5960 55504 6006
rect 55496 5954 55830 5960
rect 55438 5951 55830 5954
rect 55438 5948 55772 5951
rect 55452 5932 55772 5948
rect 53930 5664 53938 5716
rect 53990 5664 53998 5716
rect 53930 5658 53998 5664
rect 55004 5718 55278 5724
rect 55004 5666 55010 5718
rect 55062 5696 55278 5718
rect 55062 5666 55068 5696
rect 55004 5660 55068 5666
rect 53840 5604 53908 5610
rect 53840 5552 53846 5604
rect 53898 5552 53908 5604
rect 53840 5546 53908 5552
rect 54916 5602 54980 5608
rect 54916 5550 54922 5602
rect 54974 5564 54980 5602
rect 54974 5550 54982 5564
rect 53566 5534 53632 5542
rect 53566 5482 53574 5534
rect 53626 5482 53632 5534
rect 53566 5474 53632 5482
rect 53840 5444 53868 5546
rect 54916 5544 54982 5550
rect 45222 5440 52396 5444
rect 52960 5440 54280 5444
rect 54954 5440 54982 5544
rect 55454 5542 55504 5932
rect 55766 5899 55772 5932
rect 55824 5899 55830 5951
rect 55766 5892 55830 5899
rect 55858 5726 55886 6298
rect 55974 6290 55984 6342
rect 55922 6284 55984 6290
rect 56018 6240 56046 6824
rect 56142 6654 56186 7270
rect 56230 7260 56251 7376
rect 56559 7260 56580 7376
rect 58118 7376 58468 7390
rect 56230 7246 56580 7260
rect 57328 7062 57394 7068
rect 57328 7060 57334 7062
rect 56706 7032 57334 7060
rect 56118 6648 56186 6654
rect 56118 6596 56127 6648
rect 56179 6596 56186 6648
rect 56118 6590 56186 6596
rect 56422 6652 56502 6664
rect 56422 6600 56431 6652
rect 56483 6628 56502 6652
rect 56706 6628 56734 7032
rect 57328 7010 57334 7032
rect 57386 7010 57394 7062
rect 57328 7004 57394 7010
rect 56998 6870 57074 6874
rect 56998 6868 57166 6870
rect 56998 6816 57014 6868
rect 57066 6842 57166 6868
rect 57066 6816 57074 6842
rect 56998 6810 57074 6816
rect 56483 6600 56734 6628
rect 56422 6592 56734 6600
rect 55978 6212 56046 6240
rect 55978 6090 56006 6212
rect 55940 6084 56006 6090
rect 55940 6032 55946 6084
rect 55998 6032 56006 6084
rect 55940 6026 56006 6032
rect 56706 5966 56734 6592
rect 56806 6436 57074 6442
rect 56806 6414 57014 6436
rect 56806 6356 56834 6414
rect 57008 6384 57014 6414
rect 57066 6384 57074 6436
rect 57008 6378 57074 6384
rect 56770 6348 56834 6356
rect 56770 6296 56776 6348
rect 56828 6296 56834 6348
rect 56770 6288 56834 6296
rect 56006 5960 56734 5966
rect 56000 5958 56734 5960
rect 55942 5951 56734 5958
rect 55942 5899 55948 5951
rect 56000 5930 56734 5951
rect 56000 5899 56006 5930
rect 55942 5892 56006 5899
rect 55818 5716 55886 5726
rect 57138 5724 57166 6842
rect 57344 6598 57394 7004
rect 57646 6900 57700 6916
rect 57646 6860 57647 6900
rect 57486 6848 57647 6860
rect 57699 6848 57700 6900
rect 57486 6832 57700 6848
rect 57870 6890 57934 6906
rect 57870 6838 57879 6890
rect 57931 6838 57934 6890
rect 57344 6590 57410 6598
rect 57344 6538 57352 6590
rect 57404 6538 57410 6590
rect 57344 6530 57410 6538
rect 57486 6326 57514 6832
rect 57870 6824 57934 6838
rect 57556 6456 57622 6464
rect 57556 6404 57564 6456
rect 57616 6422 57622 6456
rect 57616 6404 57838 6422
rect 57556 6398 57838 6404
rect 57594 6394 57838 6398
rect 57810 6348 57838 6394
rect 57810 6342 57872 6348
rect 57486 6298 57774 6326
rect 57450 6212 57486 6214
rect 57450 6200 57522 6212
rect 57450 6148 57460 6200
rect 57512 6148 57522 6200
rect 57450 6136 57522 6148
rect 57326 6006 57392 6012
rect 57326 5954 57332 6006
rect 57384 5960 57392 6006
rect 57384 5954 57718 5960
rect 57326 5951 57718 5954
rect 57326 5948 57660 5951
rect 57340 5932 57660 5948
rect 55818 5664 55826 5716
rect 55878 5664 55886 5716
rect 55818 5658 55886 5664
rect 56892 5718 57166 5724
rect 56892 5666 56898 5718
rect 56950 5696 57166 5718
rect 56950 5666 56956 5696
rect 56892 5660 56956 5666
rect 55728 5604 55796 5610
rect 55728 5552 55734 5604
rect 55786 5552 55796 5604
rect 55728 5546 55796 5552
rect 56804 5602 56868 5608
rect 56804 5550 56810 5602
rect 56862 5564 56868 5602
rect 56862 5550 56870 5564
rect 55454 5534 55520 5542
rect 55454 5482 55462 5534
rect 55514 5482 55520 5534
rect 55454 5474 55520 5482
rect 55728 5440 55756 5546
rect 56804 5544 56870 5550
rect 56842 5440 56870 5544
rect 57342 5542 57392 5932
rect 57654 5899 57660 5932
rect 57712 5899 57718 5951
rect 57654 5892 57718 5899
rect 57746 5726 57774 6298
rect 57862 6290 57872 6342
rect 57810 6284 57872 6290
rect 57906 6240 57934 6824
rect 58030 6654 58074 7270
rect 58118 7260 58139 7376
rect 58447 7260 58468 7376
rect 58118 7246 58468 7260
rect 59216 7062 59282 7068
rect 59216 7060 59222 7062
rect 58594 7032 59222 7060
rect 58006 6648 58074 6654
rect 58006 6596 58015 6648
rect 58067 6596 58074 6648
rect 58006 6590 58074 6596
rect 58310 6652 58390 6664
rect 58310 6600 58319 6652
rect 58371 6628 58390 6652
rect 58594 6628 58622 7032
rect 59216 7010 59222 7032
rect 59274 7010 59282 7062
rect 59216 7004 59282 7010
rect 58886 6870 58962 6874
rect 58886 6868 59054 6870
rect 58886 6816 58902 6868
rect 58954 6842 59054 6868
rect 58954 6816 58962 6842
rect 58886 6810 58962 6816
rect 58371 6600 58622 6628
rect 58310 6592 58622 6600
rect 57866 6212 57934 6240
rect 57866 6090 57894 6212
rect 57828 6084 57894 6090
rect 57828 6032 57834 6084
rect 57886 6032 57894 6084
rect 57828 6026 57894 6032
rect 58594 5966 58622 6592
rect 58694 6436 58962 6442
rect 58694 6414 58902 6436
rect 58694 6356 58722 6414
rect 58896 6384 58902 6414
rect 58954 6384 58962 6436
rect 58896 6378 58962 6384
rect 58658 6348 58722 6356
rect 58658 6296 58664 6348
rect 58716 6296 58722 6348
rect 58658 6288 58722 6296
rect 57894 5960 58622 5966
rect 57888 5958 58622 5960
rect 57830 5951 58622 5958
rect 57830 5899 57836 5951
rect 57888 5930 58622 5951
rect 57888 5899 57894 5930
rect 57830 5892 57894 5899
rect 57706 5716 57774 5726
rect 59026 5724 59054 6842
rect 59232 6598 59282 7004
rect 59534 6900 59588 6916
rect 59534 6860 59535 6900
rect 59374 6848 59535 6860
rect 59587 6848 59588 6900
rect 59374 6832 59588 6848
rect 59758 6890 59822 6906
rect 59758 6838 59767 6890
rect 59819 6838 59822 6890
rect 59232 6590 59298 6598
rect 59232 6538 59240 6590
rect 59292 6538 59298 6590
rect 59232 6530 59298 6538
rect 59374 6326 59402 6832
rect 59758 6824 59822 6838
rect 59444 6456 59510 6464
rect 59444 6404 59452 6456
rect 59504 6422 59510 6456
rect 59504 6404 59726 6422
rect 59444 6398 59726 6404
rect 59482 6394 59726 6398
rect 59698 6348 59726 6394
rect 59698 6342 59760 6348
rect 59374 6298 59662 6326
rect 59338 6212 59374 6214
rect 59338 6200 59410 6212
rect 59338 6148 59348 6200
rect 59400 6148 59410 6200
rect 59338 6136 59410 6148
rect 59214 6006 59280 6012
rect 59214 5954 59220 6006
rect 59272 5960 59280 6006
rect 59272 5954 59606 5960
rect 59214 5951 59606 5954
rect 59214 5948 59548 5951
rect 59228 5932 59548 5948
rect 57706 5664 57714 5716
rect 57766 5664 57774 5716
rect 57706 5658 57774 5664
rect 58780 5718 59054 5724
rect 58780 5666 58786 5718
rect 58838 5696 59054 5718
rect 58838 5666 58844 5696
rect 58780 5660 58844 5666
rect 57616 5604 57684 5610
rect 57616 5552 57622 5604
rect 57674 5552 57684 5604
rect 57616 5546 57684 5552
rect 58692 5602 58756 5608
rect 58692 5550 58698 5602
rect 58750 5564 58756 5602
rect 58750 5550 58758 5564
rect 57342 5534 57408 5542
rect 57342 5482 57350 5534
rect 57402 5482 57408 5534
rect 57342 5474 57408 5482
rect 57616 5440 57644 5546
rect 58692 5544 58758 5550
rect 58730 5440 58758 5544
rect 59230 5542 59280 5932
rect 59542 5899 59548 5932
rect 59600 5899 59606 5951
rect 59542 5892 59606 5899
rect 59634 5726 59662 6298
rect 59750 6290 59760 6342
rect 59698 6284 59760 6290
rect 59794 6240 59822 6824
rect 59918 6654 59962 7270
rect 59894 6648 59962 6654
rect 59894 6596 59903 6648
rect 59955 6596 59962 6648
rect 59894 6590 59962 6596
rect 59754 6212 59822 6240
rect 59754 6090 59782 6212
rect 59716 6084 59782 6090
rect 59716 6032 59722 6084
rect 59774 6032 59782 6084
rect 59716 6026 59782 6032
rect 60491 5966 60605 6013
rect 59782 5960 60605 5966
rect 59776 5958 60605 5960
rect 59718 5951 60605 5958
rect 59718 5899 59724 5951
rect 59776 5930 60605 5951
rect 59776 5899 59782 5930
rect 59718 5892 59782 5899
rect 59594 5716 59662 5726
rect 59594 5664 59602 5716
rect 59654 5664 59662 5716
rect 59594 5658 59662 5664
rect 59504 5604 59572 5610
rect 59504 5552 59510 5604
rect 59562 5552 59572 5604
rect 59504 5546 59572 5552
rect 59230 5534 59296 5542
rect 59230 5482 59238 5534
rect 59290 5482 59296 5534
rect 59230 5474 59296 5482
rect 59504 5440 59532 5546
rect -78 5412 14674 5440
rect -78 5378 14666 5412
rect -79 5331 14666 5378
rect 15020 5378 29772 5440
rect 30124 5412 44876 5440
rect 30124 5378 44868 5412
rect 15020 5335 22194 5378
rect -398 5252 -48 5266
rect -398 5136 -377 5252
rect -69 5136 -48 5252
rect -398 5122 -48 5136
rect 211 5074 1237 5331
rect 1490 5252 1840 5266
rect 1490 5136 1511 5252
rect 1819 5136 1840 5252
rect 1490 5122 1840 5136
rect 2087 5074 3113 5331
rect 3378 5252 3728 5266
rect 3378 5136 3399 5252
rect 3707 5136 3728 5252
rect 3378 5122 3728 5136
rect 3991 5074 5017 5331
rect 5266 5252 5616 5266
rect 5266 5136 5287 5252
rect 5595 5136 5616 5252
rect 5266 5122 5616 5136
rect 5772 5082 7096 5331
rect 7154 5252 7504 5266
rect 7154 5136 7175 5252
rect 7483 5136 7504 5252
rect 7154 5122 7504 5136
rect 7660 5082 8980 5331
rect 9042 5252 9392 5266
rect 9042 5136 9063 5252
rect 9371 5136 9392 5252
rect 9042 5122 9392 5136
rect 5772 5074 8980 5082
rect 9658 5074 10684 5331
rect 10930 5252 11280 5266
rect 10930 5136 10951 5252
rect 11259 5136 11280 5252
rect 10930 5122 11280 5136
rect 11559 5074 12585 5331
rect 12818 5252 13168 5266
rect 12818 5136 12839 5252
rect 13147 5136 13168 5252
rect 12818 5122 13168 5136
rect 13446 5074 14472 5331
rect 14700 5252 15050 5266
rect 14700 5136 14721 5252
rect 15029 5136 15050 5252
rect 14700 5122 15050 5136
rect 15323 5074 16349 5335
rect 16588 5252 16938 5266
rect 16588 5136 16609 5252
rect 16917 5136 16938 5252
rect 16588 5122 16938 5136
rect 17192 5074 18218 5335
rect 18476 5252 18826 5266
rect 18476 5136 18497 5252
rect 18805 5136 18826 5252
rect 18476 5122 18826 5136
rect 19087 5074 20113 5335
rect 20364 5252 20714 5266
rect 20364 5136 20385 5252
rect 20693 5136 20714 5252
rect 20364 5122 20714 5136
rect 20870 5082 22194 5335
rect 22758 5331 29772 5378
rect 30123 5331 44868 5378
rect 45222 5378 59974 5440
rect 45222 5335 52396 5378
rect 22252 5252 22602 5266
rect 22252 5136 22273 5252
rect 22581 5136 22602 5252
rect 22252 5122 22602 5136
rect 22758 5082 24078 5331
rect 24140 5252 24490 5266
rect 24140 5136 24161 5252
rect 24469 5136 24490 5252
rect 24140 5122 24490 5136
rect 20870 5074 24078 5082
rect 24756 5074 25782 5331
rect 26028 5252 26378 5266
rect 26028 5136 26049 5252
rect 26357 5136 26378 5252
rect 26028 5122 26378 5136
rect 26641 5074 27667 5331
rect 27916 5252 28266 5266
rect 27916 5136 27937 5252
rect 28245 5136 28266 5252
rect 27916 5122 28266 5136
rect 28528 5074 29554 5331
rect 29804 5252 30154 5266
rect 29804 5136 29825 5252
rect 30133 5136 30154 5252
rect 29804 5122 30154 5136
rect 30413 5074 31439 5331
rect 31692 5252 32042 5266
rect 31692 5136 31713 5252
rect 32021 5136 32042 5252
rect 31692 5122 32042 5136
rect 32289 5074 33315 5331
rect 33580 5252 33930 5266
rect 33580 5136 33601 5252
rect 33909 5136 33930 5252
rect 33580 5122 33930 5136
rect 34193 5074 35219 5331
rect 35468 5252 35818 5266
rect 35468 5136 35489 5252
rect 35797 5136 35818 5252
rect 35468 5122 35818 5136
rect 35974 5082 37298 5331
rect 37356 5252 37706 5266
rect 37356 5136 37377 5252
rect 37685 5136 37706 5252
rect 37356 5122 37706 5136
rect 37862 5082 39182 5331
rect 39244 5252 39594 5266
rect 39244 5136 39265 5252
rect 39573 5136 39594 5252
rect 39244 5122 39594 5136
rect 35974 5074 39182 5082
rect 39860 5074 40886 5331
rect 41132 5252 41482 5266
rect 41132 5136 41153 5252
rect 41461 5136 41482 5252
rect 41132 5122 41482 5136
rect 41761 5074 42787 5331
rect 43020 5252 43370 5266
rect 43020 5136 43041 5252
rect 43349 5136 43370 5252
rect 43020 5122 43370 5136
rect 43648 5074 44674 5331
rect 44902 5252 45252 5266
rect 44902 5136 44923 5252
rect 45231 5136 45252 5252
rect 44902 5122 45252 5136
rect 45525 5074 46551 5335
rect 46790 5252 47140 5266
rect 46790 5136 46811 5252
rect 47119 5136 47140 5252
rect 46790 5122 47140 5136
rect 47394 5074 48420 5335
rect 48678 5252 49028 5266
rect 48678 5136 48699 5252
rect 49007 5136 49028 5252
rect 48678 5122 49028 5136
rect 49289 5074 50315 5335
rect 50566 5252 50916 5266
rect 50566 5136 50587 5252
rect 50895 5136 50916 5252
rect 50566 5122 50916 5136
rect 51072 5082 52396 5335
rect 52960 5331 59974 5378
rect 52454 5252 52804 5266
rect 52454 5136 52475 5252
rect 52783 5136 52804 5252
rect 52454 5122 52804 5136
rect 52960 5082 54280 5331
rect 54342 5252 54692 5266
rect 54342 5136 54363 5252
rect 54671 5136 54692 5252
rect 54342 5122 54692 5136
rect 51072 5074 54280 5082
rect 54958 5074 55984 5331
rect 56230 5252 56580 5266
rect 56230 5136 56251 5252
rect 56559 5136 56580 5252
rect 56230 5122 56580 5136
rect 56843 5074 57869 5331
rect 58118 5252 58468 5266
rect 58118 5136 58139 5252
rect 58447 5136 58468 5252
rect 58118 5122 58468 5136
rect 58730 5074 59756 5331
rect -80 5019 14666 5074
rect -80 4967 5864 5019
rect 5916 4967 5979 5019
rect 6031 4967 6106 5019
rect 6158 4967 6223 5019
rect 6275 4967 6337 5019
rect 6389 5018 14666 5019
rect 6389 4967 6456 5018
rect -80 4966 6456 4967
rect 6508 4966 6554 5018
rect 6606 4966 6650 5018
rect 6702 4966 6758 5018
rect 6810 4966 6857 5018
rect 6909 4966 6951 5018
rect 7003 5017 14666 5018
rect 7003 4966 7665 5017
rect -80 4965 7665 4966
rect 7717 4965 7761 5017
rect 7813 5016 14666 5017
rect 7813 4965 7850 5016
rect -80 4964 7850 4965
rect 7902 4964 7950 5016
rect 8002 4964 8047 5016
rect 8099 4964 8184 5016
rect 8236 4964 8338 5016
rect 8390 5014 14666 5016
rect 8390 4964 8464 5014
rect -80 4962 8464 4964
rect 8516 4962 8566 5014
rect 8618 4962 8673 5014
rect 8725 5012 14666 5014
rect 15020 5021 29772 5074
rect 15020 5020 21676 5021
rect 8725 4962 8785 5012
rect -80 4960 8785 4962
rect 8837 4960 14665 5012
rect -80 4948 14665 4960
rect 15020 4968 20891 5020
rect 20943 4968 20988 5020
rect 21040 4968 21085 5020
rect 21137 4968 21191 5020
rect 21243 4968 21296 5020
rect 21348 4968 21413 5020
rect 21465 5019 21676 5020
rect 21465 4968 21547 5019
rect 21599 5018 21676 5019
rect 15020 4967 21547 4968
rect 21606 4969 21676 5018
rect 21728 4969 21792 5021
rect 21844 4969 21898 5021
rect 21950 4969 22005 5021
rect 22057 5018 29772 5021
rect 22057 5017 23565 5018
rect 22057 4969 22780 5017
rect 15020 4966 21554 4967
rect 21606 4966 22780 4969
rect 15020 4965 22780 4966
rect 22832 4965 22877 5017
rect 22929 4965 22974 5017
rect 23026 4965 23080 5017
rect 23132 4965 23185 5017
rect 23237 4965 23302 5017
rect 23354 5016 23565 5017
rect 23354 4965 23436 5016
rect 15020 4964 23436 4965
rect 23488 4966 23565 5016
rect 23617 4966 23681 5018
rect 23733 4966 23787 5018
rect 23839 4966 23894 5018
rect 23946 4966 29772 5018
rect 23488 4964 29772 4966
rect 15020 4948 29772 4964
rect 30122 5019 44868 5074
rect 30122 4967 36066 5019
rect 36118 4967 36181 5019
rect 36233 4967 36308 5019
rect 36360 4967 36425 5019
rect 36477 4967 36539 5019
rect 36591 5018 44868 5019
rect 36591 4967 36658 5018
rect 30122 4966 36658 4967
rect 36710 4966 36756 5018
rect 36808 4966 36852 5018
rect 36904 4966 36960 5018
rect 37012 4966 37059 5018
rect 37111 4966 37153 5018
rect 37205 5017 44868 5018
rect 37205 4966 37867 5017
rect 30122 4965 37867 4966
rect 37919 4965 37963 5017
rect 38015 5016 44868 5017
rect 38015 4965 38052 5016
rect 30122 4964 38052 4965
rect 38104 4964 38152 5016
rect 38204 4964 38249 5016
rect 38301 4964 38386 5016
rect 38438 4964 38540 5016
rect 38592 5014 44868 5016
rect 38592 4964 38666 5014
rect 30122 4962 38666 4964
rect 38718 4962 38768 5014
rect 38820 4962 38875 5014
rect 38927 5012 44868 5014
rect 45222 5021 59974 5074
rect 45222 5020 51878 5021
rect 38927 4962 38987 5012
rect 30122 4960 38987 4962
rect 39039 4960 44867 5012
rect 30122 4948 44867 4960
rect 45222 4968 51093 5020
rect 51145 4968 51190 5020
rect 51242 4968 51287 5020
rect 51339 4968 51393 5020
rect 51445 4968 51498 5020
rect 51550 4968 51615 5020
rect 51667 5019 51878 5020
rect 51667 4968 51749 5019
rect 51801 5018 51878 5019
rect 45222 4967 51749 4968
rect 51808 4969 51878 5018
rect 51930 4969 51994 5021
rect 52046 4969 52100 5021
rect 52152 4969 52207 5021
rect 52259 5018 59974 5021
rect 52259 5017 53767 5018
rect 52259 4969 52982 5017
rect 45222 4966 51756 4967
rect 51808 4966 52982 4969
rect 45222 4965 52982 4966
rect 53034 4965 53079 5017
rect 53131 4965 53176 5017
rect 53228 4965 53282 5017
rect 53334 4965 53387 5017
rect 53439 4965 53504 5017
rect 53556 5016 53767 5017
rect 53556 4965 53638 5016
rect 45222 4964 53638 4965
rect 53690 4966 53767 5016
rect 53819 4966 53883 5018
rect 53935 4966 53989 5018
rect 54041 4966 54096 5018
rect 54148 4966 59974 5018
rect 53690 4964 59974 4966
rect 45222 4948 59974 4964
rect -80 4886 14666 4948
rect 15020 4886 29774 4948
rect 30122 4886 44868 4948
rect 45222 4886 59976 4948
rect 2087 4885 3113 4886
rect 3991 4882 5017 4886
rect 9658 4885 10684 4886
rect 11559 4884 12585 4886
rect 24756 4884 25782 4886
rect 26641 4885 27667 4886
rect 32289 4885 33315 4886
rect 34193 4882 35219 4886
rect 39860 4885 40886 4886
rect 41761 4884 42787 4886
rect 54958 4884 55984 4886
rect 56843 4885 57869 4886
rect 7240 4813 7429 4843
rect 7240 4761 7264 4813
rect 7316 4812 7429 4813
rect 7316 4761 7345 4812
rect 7240 4760 7345 4761
rect 7397 4760 7429 4812
rect 6208 4670 6692 4719
rect 6208 4669 6581 4670
rect 6208 4667 6379 4669
rect 6208 4615 6272 4667
rect 6324 4617 6379 4667
rect 6431 4617 6481 4669
rect 6533 4618 6581 4669
rect 6633 4618 6692 4670
rect 6533 4617 6692 4618
rect 6324 4615 6692 4617
rect 6208 3372 6692 4615
rect 6208 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6692 3372
rect 6208 3257 6692 3316
rect 6208 3201 6275 3257
rect 6331 3201 6389 3257
rect 6445 3201 6503 3257
rect 6559 3201 6692 3257
rect 6208 3142 6692 3201
rect 6208 3086 6275 3142
rect 6331 3086 6389 3142
rect 6445 3086 6503 3142
rect 6559 3086 6692 3142
rect 6208 2817 6692 3086
rect 6208 2765 6266 2817
rect 6318 2765 6364 2817
rect 6416 2765 6459 2817
rect 6511 2765 6564 2817
rect 6616 2765 6692 2817
rect 6208 2729 6692 2765
rect 7240 3558 7429 4760
rect 14423 4747 14683 4818
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14683 4747
rect 22351 4810 22540 4833
rect 22351 4758 22380 4810
rect 22432 4758 22475 4810
rect 22527 4758 22540 4810
rect 14423 3770 14683 4695
rect 14423 3718 14467 3770
rect 14519 3718 14590 3770
rect 14642 3718 14683 3770
rect 14423 3674 14683 3718
rect 21264 4673 21731 4697
rect 21264 4621 21302 4673
rect 21354 4621 21405 4673
rect 21457 4621 21488 4673
rect 21540 4621 21589 4673
rect 21641 4621 21676 4673
rect 21728 4621 21731 4673
rect 7240 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3506 7429 3558
rect 7240 2675 7429 3506
rect 14848 3413 15054 3458
rect 14848 3409 14986 3413
rect 14848 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3361 15054 3413
rect 14933 3357 15054 3361
rect 7240 2623 7265 2675
rect 7317 2673 7429 2675
rect 7317 2623 7345 2673
rect 7240 2621 7345 2623
rect 7397 2621 7429 2673
rect 13629 3222 13982 3268
rect 13629 3221 13857 3222
rect 13629 3169 13680 3221
rect 13732 3169 13764 3221
rect 13816 3170 13857 3221
rect 13909 3170 13982 3222
rect 13816 3169 13982 3170
rect 13629 2811 13982 3169
rect 14848 2992 15054 3357
rect 14848 2940 14885 2992
rect 14937 2987 15054 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 15054 2987
rect 14848 2914 15054 2935
rect 14848 2912 14979 2914
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 15054 2914
rect 14937 2860 15054 2862
rect 14848 2831 15054 2860
rect 21264 3282 21731 4621
rect 21264 3226 21314 3282
rect 21370 3226 21418 3282
rect 21474 3226 21522 3282
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21264 3166 21731 3226
rect 21264 3110 21314 3166
rect 21370 3110 21418 3166
rect 21474 3110 21522 3166
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3050 21731 3110
rect 21264 2994 21314 3050
rect 21370 2994 21418 3050
rect 21474 2994 21522 3050
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 13629 2755 13669 2811
rect 13725 2755 13777 2811
rect 13833 2755 13885 2811
rect 13941 2755 13982 2811
rect 13629 2717 13982 2755
rect 21264 2822 21731 2994
rect 21264 2770 21316 2822
rect 21368 2770 21416 2822
rect 21468 2770 21515 2822
rect 21567 2770 21618 2822
rect 21670 2770 21731 2822
rect 21264 2746 21731 2770
rect 22351 3556 22540 4758
rect 30356 4770 30691 4813
rect 30356 4718 30402 4770
rect 30454 4718 30515 4770
rect 30567 4718 30616 4770
rect 30668 4718 30691 4770
rect 30356 4150 30691 4718
rect 37442 4812 37629 4831
rect 37442 4760 37457 4812
rect 37509 4760 37559 4812
rect 37611 4760 37629 4812
rect 30356 4147 30517 4150
rect 30356 4095 30414 4147
rect 30466 4098 30517 4147
rect 30569 4098 30618 4150
rect 30670 4098 30691 4150
rect 30466 4095 30691 4098
rect 30356 4063 30691 4095
rect 36380 4674 36680 4695
rect 36380 4669 36607 4674
rect 36380 4617 36434 4669
rect 36486 4617 36522 4669
rect 36574 4622 36607 4669
rect 36659 4622 36680 4674
rect 36574 4617 36680 4622
rect 31127 3741 31666 3764
rect 31127 3689 31195 3741
rect 31247 3689 31355 3741
rect 31407 3689 31488 3741
rect 31540 3689 31601 3741
rect 31653 3689 31666 3741
rect 22351 3549 22475 3556
rect 22351 3497 22376 3549
rect 22428 3504 22475 3549
rect 22527 3504 22540 3556
rect 22428 3497 22540 3504
rect 13629 2661 13669 2717
rect 13725 2661 13777 2717
rect 13833 2661 13885 2717
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 22351 2690 22540 3497
rect 30318 3600 30743 3618
rect 30318 3597 30577 3600
rect 30318 3595 30466 3597
rect 30318 3543 30370 3595
rect 30422 3545 30466 3595
rect 30518 3548 30577 3597
rect 30629 3597 30743 3600
rect 30629 3548 30669 3597
rect 30518 3545 30669 3548
rect 30721 3545 30743 3597
rect 30422 3543 30743 3545
rect 30318 2931 30743 3543
rect 31127 3173 31666 3689
rect 31127 3121 31184 3173
rect 31236 3121 31328 3173
rect 31380 3121 31472 3173
rect 31524 3121 31666 3173
rect 31127 3089 31666 3121
rect 31127 3037 31183 3089
rect 31235 3037 31327 3089
rect 31379 3037 31471 3089
rect 31523 3037 31666 3089
rect 31127 2963 31666 3037
rect 36380 3631 36680 4617
rect 36380 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36680 3631
rect 36380 3543 36680 3575
rect 36380 3487 36401 3543
rect 36457 3487 36495 3543
rect 36551 3487 36589 3543
rect 36645 3487 36680 3543
rect 36380 3455 36680 3487
rect 36380 3399 36401 3455
rect 36457 3399 36495 3455
rect 36551 3399 36589 3455
rect 36645 3399 36680 3455
rect 30318 2875 30364 2931
rect 30420 2875 30489 2931
rect 30545 2875 30614 2931
rect 30670 2875 30743 2931
rect 30318 2835 30743 2875
rect 30318 2779 30364 2835
rect 30420 2779 30489 2835
rect 30545 2779 30614 2835
rect 30670 2779 30743 2835
rect 30318 2747 30743 2779
rect 36380 2816 36680 3399
rect 36380 2764 36424 2816
rect 36476 2764 36512 2816
rect 36564 2812 36680 2816
rect 36564 2764 36610 2812
rect 36380 2760 36610 2764
rect 36662 2760 36680 2812
rect 36380 2743 36680 2760
rect 37442 3714 37629 4760
rect 44571 4747 44790 4800
rect 44571 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 44571 3923 44790 4695
rect 44571 3922 44690 3923
rect 44571 3870 44600 3922
rect 44652 3871 44690 3922
rect 44742 3871 44790 3923
rect 44652 3870 44790 3871
rect 44571 3835 44790 3870
rect 52546 4785 52735 4808
rect 52546 4733 52575 4785
rect 52627 4733 52670 4785
rect 52722 4733 52735 4785
rect 37442 3713 37563 3714
rect 37442 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3662 37629 3714
rect 37512 3661 37629 3662
rect 22351 2638 22381 2690
rect 22433 2638 22464 2690
rect 22516 2638 22540 2690
rect 22351 2625 22540 2638
rect 37442 2680 37629 3661
rect 52546 3714 52735 4733
rect 52546 3709 52664 3714
rect 52546 3657 52573 3709
rect 52625 3662 52664 3709
rect 52716 3662 52735 3714
rect 52625 3657 52735 3662
rect 44990 3573 45196 3618
rect 44990 3569 45128 3573
rect 44990 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3521 45196 3573
rect 45075 3517 45196 3521
rect 44990 3175 45196 3517
rect 44990 3172 45120 3175
rect 44990 3120 45031 3172
rect 45083 3123 45120 3172
rect 45172 3123 45196 3175
rect 45083 3120 45196 3123
rect 44990 3096 45196 3120
rect 44990 3044 45031 3096
rect 45083 3044 45124 3096
rect 45176 3044 45196 3096
rect 44990 3001 45196 3044
rect 45998 3383 46412 3405
rect 45998 3382 46127 3383
rect 45998 3330 46035 3382
rect 46087 3331 46127 3382
rect 46179 3382 46412 3383
rect 46179 3331 46217 3382
rect 46087 3330 46217 3331
rect 46269 3381 46412 3382
rect 46269 3330 46305 3381
rect 45998 3329 46305 3330
rect 46357 3329 46412 3381
rect 37442 2628 37459 2680
rect 37511 2628 37550 2680
rect 37602 2628 37629 2680
rect 7240 2603 7429 2621
rect 37442 2620 37629 2628
rect 45998 2784 46412 3329
rect 45998 2728 46035 2784
rect 46091 2728 46128 2784
rect 46184 2728 46221 2784
rect 46277 2728 46314 2784
rect 46370 2728 46412 2784
rect 45998 2702 46412 2728
rect 45998 2646 46035 2702
rect 46091 2646 46128 2702
rect 46184 2646 46221 2702
rect 46277 2646 46314 2702
rect 46370 2646 46412 2702
rect 45998 2609 46412 2646
rect 52546 2665 52735 3657
rect 53311 4666 53732 4695
rect 53311 4614 53350 4666
rect 53402 4614 53444 4666
rect 53496 4614 53521 4666
rect 53573 4665 53675 4666
rect 53573 4614 53601 4665
rect 53311 4613 53601 4614
rect 53653 4614 53675 4665
rect 53727 4614 53732 4666
rect 53653 4613 53732 4614
rect 53311 3176 53732 4613
rect 53311 3120 53348 3176
rect 53404 3120 53452 3176
rect 53508 3120 53556 3176
rect 53612 3120 53660 3176
rect 53716 3120 53732 3176
rect 53311 3086 53732 3120
rect 53311 3030 53348 3086
rect 53404 3030 53452 3086
rect 53508 3030 53556 3086
rect 53612 3030 53660 3086
rect 53716 3030 53732 3086
rect 53311 2813 53732 3030
rect 53311 2761 53346 2813
rect 53398 2761 53434 2813
rect 53486 2761 53517 2813
rect 53569 2761 53604 2813
rect 53656 2761 53732 2813
rect 53311 2745 53732 2761
rect 52546 2613 52576 2665
rect 52628 2613 52659 2665
rect 52711 2613 52735 2665
rect 52546 2600 52735 2613
rect 2113 2554 3139 2555
rect 3998 2554 5024 2556
rect 17195 2554 18221 2556
rect 19096 2554 20122 2555
rect 24763 2554 25789 2558
rect 26667 2554 27693 2555
rect 32315 2554 33341 2555
rect 34200 2554 35226 2556
rect 47397 2554 48423 2556
rect 49298 2554 50324 2555
rect 54965 2554 55991 2558
rect 56869 2554 57895 2555
rect 6 2492 14760 2554
rect 15114 2492 29860 2554
rect 30208 2492 44962 2554
rect 45316 2492 60062 2554
rect 8 2476 14760 2492
rect 8 2474 6292 2476
rect 8 2422 5834 2474
rect 5886 2422 5941 2474
rect 5993 2422 6047 2474
rect 6099 2422 6163 2474
rect 6215 2424 6292 2474
rect 6344 2475 14760 2476
rect 6344 2424 6426 2475
rect 6215 2423 6426 2424
rect 6478 2423 6543 2475
rect 6595 2423 6648 2475
rect 6700 2423 6754 2475
rect 6806 2423 6851 2475
rect 6903 2423 6948 2475
rect 7000 2474 14760 2475
rect 7000 2471 8174 2474
rect 8226 2473 14760 2474
rect 7000 2423 7723 2471
rect 6215 2422 7723 2423
rect 8 2419 7723 2422
rect 7775 2419 7830 2471
rect 7882 2419 7936 2471
rect 7988 2419 8052 2471
rect 8104 2422 8174 2471
rect 8233 2472 14760 2473
rect 8104 2421 8181 2422
rect 8233 2421 8315 2472
rect 8104 2420 8315 2421
rect 8367 2420 8432 2472
rect 8484 2420 8537 2472
rect 8589 2420 8643 2472
rect 8695 2420 8740 2472
rect 8792 2420 8837 2472
rect 8889 2420 14760 2472
rect 15115 2480 29860 2492
rect 15115 2428 20943 2480
rect 20995 2478 29860 2480
rect 20995 2428 21055 2478
rect 8104 2419 14760 2420
rect 8 2366 14760 2419
rect 15114 2426 21055 2428
rect 21107 2426 21162 2478
rect 21214 2426 21264 2478
rect 21316 2476 29860 2478
rect 21316 2426 21390 2476
rect 15114 2424 21390 2426
rect 21442 2424 21544 2476
rect 21596 2424 21681 2476
rect 21733 2424 21778 2476
rect 21830 2424 21878 2476
rect 21930 2475 29860 2476
rect 21930 2424 21967 2475
rect 15114 2423 21967 2424
rect 22019 2423 22063 2475
rect 22115 2474 29860 2475
rect 22115 2423 22777 2474
rect 15114 2422 22777 2423
rect 22829 2422 22871 2474
rect 22923 2422 22970 2474
rect 23022 2422 23078 2474
rect 23130 2422 23174 2474
rect 23226 2422 23272 2474
rect 23324 2473 29860 2474
rect 23324 2422 23391 2473
rect 15114 2421 23391 2422
rect 23443 2421 23505 2473
rect 23557 2421 23622 2473
rect 23674 2421 23749 2473
rect 23801 2421 23864 2473
rect 23916 2421 29860 2473
rect 15114 2366 29860 2421
rect 30210 2476 44962 2492
rect 30210 2474 36494 2476
rect 30210 2422 36036 2474
rect 36088 2422 36143 2474
rect 36195 2422 36249 2474
rect 36301 2422 36365 2474
rect 36417 2424 36494 2474
rect 36546 2475 44962 2476
rect 36546 2424 36628 2475
rect 36417 2423 36628 2424
rect 36680 2423 36745 2475
rect 36797 2423 36850 2475
rect 36902 2423 36956 2475
rect 37008 2423 37053 2475
rect 37105 2423 37150 2475
rect 37202 2474 44962 2475
rect 37202 2471 38376 2474
rect 38428 2473 44962 2474
rect 37202 2423 37925 2471
rect 36417 2422 37925 2423
rect 30210 2419 37925 2422
rect 37977 2419 38032 2471
rect 38084 2419 38138 2471
rect 38190 2419 38254 2471
rect 38306 2422 38376 2471
rect 38435 2472 44962 2473
rect 38306 2421 38383 2422
rect 38435 2421 38517 2472
rect 38306 2420 38517 2421
rect 38569 2420 38634 2472
rect 38686 2420 38739 2472
rect 38791 2420 38845 2472
rect 38897 2420 38942 2472
rect 38994 2420 39039 2472
rect 39091 2420 44962 2472
rect 45317 2480 60062 2492
rect 45317 2428 51145 2480
rect 51197 2478 60062 2480
rect 51197 2428 51257 2478
rect 38306 2419 44962 2420
rect 30210 2366 44962 2419
rect 45316 2426 51257 2428
rect 51309 2426 51364 2478
rect 51416 2426 51466 2478
rect 51518 2476 60062 2478
rect 51518 2426 51592 2476
rect 45316 2424 51592 2426
rect 51644 2424 51746 2476
rect 51798 2424 51883 2476
rect 51935 2424 51980 2476
rect 52032 2424 52080 2476
rect 52132 2475 60062 2476
rect 52132 2424 52169 2475
rect 45316 2423 52169 2424
rect 52221 2423 52265 2475
rect 52317 2474 60062 2475
rect 52317 2423 52979 2474
rect 45316 2422 52979 2423
rect 53031 2422 53073 2474
rect 53125 2422 53172 2474
rect 53224 2422 53280 2474
rect 53332 2422 53376 2474
rect 53428 2422 53474 2474
rect 53526 2473 60062 2474
rect 53526 2422 53593 2473
rect 45316 2421 53593 2422
rect 53645 2421 53707 2473
rect 53759 2421 53824 2473
rect 53876 2421 53951 2473
rect 54003 2421 54066 2473
rect 54118 2421 60062 2473
rect 45316 2366 60062 2421
rect 226 2109 1252 2366
rect 1514 2304 1864 2318
rect 1514 2188 1535 2304
rect 1843 2188 1864 2304
rect 1514 2174 1864 2188
rect 2113 2109 3139 2366
rect 3402 2304 3752 2318
rect 3402 2188 3423 2304
rect 3731 2188 3752 2304
rect 3402 2174 3752 2188
rect 3998 2109 5024 2366
rect 5702 2358 8910 2366
rect 5290 2304 5640 2318
rect 5290 2188 5311 2304
rect 5619 2188 5640 2304
rect 5290 2174 5640 2188
rect 5702 2109 7022 2358
rect 7178 2304 7528 2318
rect 7178 2188 7199 2304
rect 7507 2188 7528 2304
rect 7178 2174 7528 2188
rect 8 2062 7022 2109
rect 7586 2105 8910 2358
rect 9066 2304 9416 2318
rect 9066 2188 9087 2304
rect 9395 2188 9416 2304
rect 9066 2174 9416 2188
rect 9667 2105 10693 2366
rect 10954 2304 11304 2318
rect 10954 2188 10975 2304
rect 11283 2188 11304 2304
rect 10954 2174 11304 2188
rect 11562 2105 12588 2366
rect 12842 2304 13192 2318
rect 12842 2188 12863 2304
rect 13171 2188 13192 2304
rect 12842 2174 13192 2188
rect 13431 2105 14457 2366
rect 14730 2304 15080 2318
rect 14730 2188 14751 2304
rect 15059 2188 15080 2304
rect 14730 2174 15080 2188
rect 15308 2109 16334 2366
rect 16612 2304 16962 2318
rect 16612 2188 16633 2304
rect 16941 2188 16962 2304
rect 16612 2174 16962 2188
rect 17195 2109 18221 2366
rect 18500 2304 18850 2318
rect 18500 2188 18521 2304
rect 18829 2188 18850 2304
rect 18500 2174 18850 2188
rect 19096 2109 20122 2366
rect 20800 2358 24008 2366
rect 20388 2304 20738 2318
rect 20388 2188 20409 2304
rect 20717 2188 20738 2304
rect 20388 2174 20738 2188
rect 20800 2109 22120 2358
rect 22276 2304 22626 2318
rect 22276 2188 22297 2304
rect 22605 2188 22626 2304
rect 22276 2174 22626 2188
rect 22684 2109 24008 2358
rect 24164 2304 24514 2318
rect 24164 2188 24185 2304
rect 24493 2188 24514 2304
rect 24164 2174 24514 2188
rect 24763 2109 25789 2366
rect 26052 2304 26402 2318
rect 26052 2188 26073 2304
rect 26381 2188 26402 2304
rect 26052 2174 26402 2188
rect 26667 2109 27693 2366
rect 27940 2304 28290 2318
rect 27940 2188 27961 2304
rect 28269 2188 28290 2304
rect 27940 2174 28290 2188
rect 28543 2109 29569 2366
rect 29828 2304 30178 2318
rect 29828 2188 29849 2304
rect 30157 2188 30178 2304
rect 29828 2174 30178 2188
rect 30428 2109 31454 2366
rect 31716 2304 32066 2318
rect 31716 2188 31737 2304
rect 32045 2188 32066 2304
rect 31716 2174 32066 2188
rect 32315 2109 33341 2366
rect 33604 2304 33954 2318
rect 33604 2188 33625 2304
rect 33933 2188 33954 2304
rect 33604 2174 33954 2188
rect 34200 2109 35226 2366
rect 35904 2358 39112 2366
rect 35492 2304 35842 2318
rect 35492 2188 35513 2304
rect 35821 2188 35842 2304
rect 35492 2174 35842 2188
rect 35904 2109 37224 2358
rect 37380 2304 37730 2318
rect 37380 2188 37401 2304
rect 37709 2188 37730 2304
rect 37380 2174 37730 2188
rect 7586 2062 14760 2105
rect 8 2000 14760 2062
rect 15114 2062 29859 2109
rect 30210 2062 37224 2109
rect 37788 2105 39112 2358
rect 39268 2304 39618 2318
rect 39268 2188 39289 2304
rect 39597 2188 39618 2304
rect 39268 2174 39618 2188
rect 39869 2105 40895 2366
rect 41156 2304 41506 2318
rect 41156 2188 41177 2304
rect 41485 2188 41506 2304
rect 41156 2174 41506 2188
rect 41764 2105 42790 2366
rect 43044 2304 43394 2318
rect 43044 2188 43065 2304
rect 43373 2188 43394 2304
rect 43044 2174 43394 2188
rect 43633 2105 44659 2366
rect 44932 2304 45282 2318
rect 44932 2188 44953 2304
rect 45261 2188 45282 2304
rect 44932 2174 45282 2188
rect 45510 2109 46536 2366
rect 46814 2304 47164 2318
rect 46814 2188 46835 2304
rect 47143 2188 47164 2304
rect 46814 2174 47164 2188
rect 47397 2109 48423 2366
rect 48702 2304 49052 2318
rect 48702 2188 48723 2304
rect 49031 2188 49052 2304
rect 48702 2174 49052 2188
rect 49298 2109 50324 2366
rect 51002 2358 54210 2366
rect 50590 2304 50940 2318
rect 50590 2188 50611 2304
rect 50919 2188 50940 2304
rect 50590 2174 50940 2188
rect 51002 2109 52322 2358
rect 52478 2304 52828 2318
rect 52478 2188 52499 2304
rect 52807 2188 52828 2304
rect 52478 2174 52828 2188
rect 52886 2109 54210 2358
rect 54366 2304 54716 2318
rect 54366 2188 54387 2304
rect 54695 2188 54716 2304
rect 54366 2174 54716 2188
rect 54965 2109 55991 2366
rect 56254 2304 56604 2318
rect 56254 2188 56275 2304
rect 56583 2188 56604 2304
rect 56254 2174 56604 2188
rect 56869 2109 57895 2366
rect 58142 2304 58492 2318
rect 58142 2188 58163 2304
rect 58471 2188 58492 2304
rect 58142 2174 58492 2188
rect 58745 2109 59771 2366
rect 60030 2304 60380 2318
rect 60030 2188 60051 2304
rect 60359 2188 60380 2304
rect 60030 2174 60380 2188
rect 37788 2062 44962 2105
rect 15114 2028 29858 2062
rect 15106 2000 29858 2028
rect 30210 2000 44962 2062
rect 45316 2062 60061 2109
rect 45316 2028 60060 2062
rect 45308 2000 60060 2028
rect 450 1894 478 2000
rect 686 1958 752 1966
rect 686 1906 692 1958
rect 744 1906 752 1958
rect 686 1898 752 1906
rect 410 1888 478 1894
rect 410 1836 420 1888
rect 472 1836 478 1888
rect 410 1830 478 1836
rect 320 1776 388 1782
rect 320 1724 328 1776
rect 380 1724 388 1776
rect 320 1714 388 1724
rect 200 1541 264 1548
rect 200 1510 206 1541
rect -634 1489 206 1510
rect 258 1489 264 1541
rect -634 1482 264 1489
rect -634 1480 206 1482
rect -634 1474 200 1480
rect -629 1391 -539 1474
rect 200 1408 266 1414
rect 200 1356 208 1408
rect 260 1356 266 1408
rect 200 1350 266 1356
rect 200 1228 228 1350
rect 160 1200 228 1228
rect 20 844 88 850
rect 20 792 27 844
rect 79 792 88 844
rect 20 786 88 792
rect 20 170 64 786
rect 160 616 188 1200
rect 222 1150 284 1156
rect 222 1098 232 1150
rect 320 1142 348 1714
rect 376 1541 440 1548
rect 376 1489 382 1541
rect 434 1508 440 1541
rect 702 1508 752 1898
rect 1224 1896 1252 2000
rect 1224 1890 1290 1896
rect 2338 1894 2366 2000
rect 2574 1958 2640 1966
rect 2574 1906 2580 1958
rect 2632 1906 2640 1958
rect 2574 1898 2640 1906
rect 1224 1876 1232 1890
rect 1226 1838 1232 1876
rect 1284 1838 1290 1890
rect 1226 1832 1290 1838
rect 2298 1888 2366 1894
rect 2298 1836 2308 1888
rect 2360 1836 2366 1888
rect 2298 1830 2366 1836
rect 1138 1774 1202 1780
rect 1138 1744 1144 1774
rect 928 1722 1144 1744
rect 1196 1722 1202 1774
rect 928 1716 1202 1722
rect 2208 1776 2276 1782
rect 2208 1724 2216 1776
rect 2268 1724 2276 1776
rect 434 1492 754 1508
rect 434 1489 768 1492
rect 376 1486 768 1489
rect 376 1480 710 1486
rect 702 1434 710 1480
rect 762 1434 768 1486
rect 702 1428 768 1434
rect 572 1292 644 1304
rect 572 1240 582 1292
rect 634 1240 644 1292
rect 572 1228 644 1240
rect 608 1226 644 1228
rect 320 1114 608 1142
rect 222 1092 284 1098
rect 256 1046 284 1092
rect 256 1042 500 1046
rect 256 1036 538 1042
rect 256 1018 478 1036
rect 472 984 478 1018
rect 530 984 538 1036
rect 472 976 538 984
rect 160 602 224 616
rect 580 608 608 1114
rect 684 902 750 910
rect 684 850 690 902
rect 742 850 750 902
rect 684 842 750 850
rect 160 550 163 602
rect 215 550 224 602
rect 160 534 224 550
rect 394 592 608 608
rect 394 540 395 592
rect 447 580 608 592
rect 447 540 448 580
rect 394 524 448 540
rect 700 436 750 842
rect 928 598 956 1716
rect 2208 1714 2276 1724
rect 2088 1541 2152 1548
rect 2088 1510 2094 1541
rect 1360 1489 2094 1510
rect 2146 1489 2152 1541
rect 1360 1482 2152 1489
rect 1360 1480 2094 1482
rect 1360 1474 2088 1480
rect 1260 1144 1324 1152
rect 1260 1092 1266 1144
rect 1318 1092 1324 1144
rect 1260 1084 1324 1092
rect 1020 1056 1086 1062
rect 1020 1004 1028 1056
rect 1080 1026 1086 1056
rect 1260 1026 1288 1084
rect 1080 1004 1288 1026
rect 1020 998 1288 1004
rect 1360 848 1388 1474
rect 2088 1408 2154 1414
rect 2088 1356 2096 1408
rect 2148 1356 2154 1408
rect 2088 1350 2154 1356
rect 2088 1228 2116 1350
rect 2048 1200 2116 1228
rect 1360 840 1672 848
rect 1360 812 1611 840
rect 1020 624 1096 630
rect 1020 598 1028 624
rect 928 572 1028 598
rect 1080 572 1096 624
rect 928 570 1096 572
rect 1020 566 1096 570
rect 700 430 766 436
rect 700 378 708 430
rect 760 408 766 430
rect 1360 408 1388 812
rect 1592 788 1611 812
rect 1663 788 1672 840
rect 1592 776 1672 788
rect 1908 844 1976 850
rect 1908 792 1915 844
rect 1967 792 1976 844
rect 1908 786 1976 792
rect 760 380 1388 408
rect 760 378 766 380
rect 700 372 766 378
rect 1514 180 1864 194
rect 1514 64 1535 180
rect 1843 64 1864 180
rect 1908 170 1952 786
rect 2048 616 2076 1200
rect 2110 1150 2172 1156
rect 2110 1098 2120 1150
rect 2208 1142 2236 1714
rect 2264 1541 2328 1548
rect 2264 1489 2270 1541
rect 2322 1508 2328 1541
rect 2590 1508 2640 1898
rect 3112 1896 3140 2000
rect 3112 1890 3178 1896
rect 4226 1894 4254 2000
rect 4462 1958 4528 1966
rect 4462 1906 4468 1958
rect 4520 1906 4528 1958
rect 4462 1898 4528 1906
rect 3112 1876 3120 1890
rect 3114 1838 3120 1876
rect 3172 1838 3178 1890
rect 3114 1832 3178 1838
rect 4186 1888 4254 1894
rect 4186 1836 4196 1888
rect 4248 1836 4254 1888
rect 4186 1830 4254 1836
rect 3026 1774 3090 1780
rect 3026 1744 3032 1774
rect 2816 1722 3032 1744
rect 3084 1722 3090 1774
rect 2816 1716 3090 1722
rect 4096 1776 4164 1782
rect 4096 1724 4104 1776
rect 4156 1724 4164 1776
rect 2322 1492 2642 1508
rect 2322 1489 2656 1492
rect 2264 1486 2656 1489
rect 2264 1480 2598 1486
rect 2590 1434 2598 1480
rect 2650 1434 2656 1486
rect 2590 1428 2656 1434
rect 2460 1292 2532 1304
rect 2460 1240 2470 1292
rect 2522 1240 2532 1292
rect 2460 1228 2532 1240
rect 2496 1226 2532 1228
rect 2208 1114 2496 1142
rect 2110 1092 2172 1098
rect 2144 1046 2172 1092
rect 2144 1042 2388 1046
rect 2144 1036 2426 1042
rect 2144 1018 2366 1036
rect 2360 984 2366 1018
rect 2418 984 2426 1036
rect 2360 976 2426 984
rect 2048 602 2112 616
rect 2468 608 2496 1114
rect 2572 902 2638 910
rect 2572 850 2578 902
rect 2630 850 2638 902
rect 2572 842 2638 850
rect 2048 550 2051 602
rect 2103 550 2112 602
rect 2048 534 2112 550
rect 2282 592 2496 608
rect 2282 540 2283 592
rect 2335 580 2496 592
rect 2335 540 2336 580
rect 2282 524 2336 540
rect 2588 436 2638 842
rect 2816 598 2844 1716
rect 4096 1714 4164 1724
rect 3976 1541 4040 1548
rect 3976 1510 3982 1541
rect 3248 1489 3982 1510
rect 4034 1489 4040 1541
rect 3248 1482 4040 1489
rect 3248 1480 3982 1482
rect 3248 1474 3976 1480
rect 3148 1144 3212 1152
rect 3148 1092 3154 1144
rect 3206 1092 3212 1144
rect 3148 1084 3212 1092
rect 2908 1056 2974 1062
rect 2908 1004 2916 1056
rect 2968 1026 2974 1056
rect 3148 1026 3176 1084
rect 2968 1004 3176 1026
rect 2908 998 3176 1004
rect 3248 848 3276 1474
rect 3976 1408 4042 1414
rect 3976 1356 3984 1408
rect 4036 1356 4042 1408
rect 3976 1350 4042 1356
rect 3976 1228 4004 1350
rect 3936 1200 4004 1228
rect 3248 840 3560 848
rect 3248 812 3499 840
rect 2908 624 2984 630
rect 2908 598 2916 624
rect 2816 572 2916 598
rect 2968 572 2984 624
rect 2816 570 2984 572
rect 2908 566 2984 570
rect 2588 430 2654 436
rect 2588 378 2596 430
rect 2648 408 2654 430
rect 3248 408 3276 812
rect 3480 788 3499 812
rect 3551 788 3560 840
rect 3480 776 3560 788
rect 3796 844 3864 850
rect 3796 792 3803 844
rect 3855 792 3864 844
rect 3796 786 3864 792
rect 2648 380 3276 408
rect 2648 378 2654 380
rect 2588 372 2654 378
rect 3402 180 3752 194
rect 1514 50 1864 64
rect 3402 64 3423 180
rect 3731 64 3752 180
rect 3796 170 3840 786
rect 3936 616 3964 1200
rect 3998 1150 4060 1156
rect 3998 1098 4008 1150
rect 4096 1142 4124 1714
rect 4152 1541 4216 1548
rect 4152 1489 4158 1541
rect 4210 1508 4216 1541
rect 4478 1508 4528 1898
rect 5000 1896 5028 2000
rect 5702 1996 7022 2000
rect 7586 1996 14760 2000
rect 5000 1890 5066 1896
rect 6114 1894 6142 1996
rect 6350 1958 6416 1966
rect 6350 1906 6356 1958
rect 6408 1906 6416 1958
rect 6350 1898 6416 1906
rect 5000 1876 5008 1890
rect 5002 1838 5008 1876
rect 5060 1838 5066 1890
rect 5002 1832 5066 1838
rect 6074 1888 6142 1894
rect 6074 1836 6084 1888
rect 6136 1836 6142 1888
rect 6074 1830 6142 1836
rect 4914 1774 4978 1780
rect 4914 1744 4920 1774
rect 4704 1722 4920 1744
rect 4972 1722 4978 1774
rect 4704 1716 4978 1722
rect 5984 1776 6052 1782
rect 5984 1724 5992 1776
rect 6044 1724 6052 1776
rect 4210 1492 4530 1508
rect 4210 1489 4544 1492
rect 4152 1486 4544 1489
rect 4152 1480 4486 1486
rect 4478 1434 4486 1480
rect 4538 1434 4544 1486
rect 4478 1428 4544 1434
rect 4348 1292 4420 1304
rect 4348 1240 4358 1292
rect 4410 1240 4420 1292
rect 4348 1228 4420 1240
rect 4384 1226 4420 1228
rect 4096 1114 4384 1142
rect 3998 1092 4060 1098
rect 4032 1046 4060 1092
rect 4032 1042 4276 1046
rect 4032 1036 4314 1042
rect 4032 1018 4254 1036
rect 4248 984 4254 1018
rect 4306 984 4314 1036
rect 4248 976 4314 984
rect 3936 602 4000 616
rect 4356 608 4384 1114
rect 4460 902 4526 910
rect 4460 850 4466 902
rect 4518 850 4526 902
rect 4460 842 4526 850
rect 3936 550 3939 602
rect 3991 550 4000 602
rect 3936 534 4000 550
rect 4170 592 4384 608
rect 4170 540 4171 592
rect 4223 580 4384 592
rect 4223 540 4224 580
rect 4170 524 4224 540
rect 4476 436 4526 842
rect 4704 598 4732 1716
rect 5984 1714 6052 1724
rect 5864 1541 5928 1548
rect 5864 1510 5870 1541
rect 5136 1489 5870 1510
rect 5922 1489 5928 1541
rect 5136 1482 5928 1489
rect 5136 1480 5870 1482
rect 5136 1474 5864 1480
rect 5036 1144 5100 1152
rect 5036 1092 5042 1144
rect 5094 1092 5100 1144
rect 5036 1084 5100 1092
rect 4796 1056 4862 1062
rect 4796 1004 4804 1056
rect 4856 1026 4862 1056
rect 5036 1026 5064 1084
rect 4856 1004 5064 1026
rect 4796 998 5064 1004
rect 5136 848 5164 1474
rect 5864 1408 5930 1414
rect 5864 1356 5872 1408
rect 5924 1356 5930 1408
rect 5864 1350 5930 1356
rect 5864 1228 5892 1350
rect 5824 1200 5892 1228
rect 5136 840 5448 848
rect 5136 812 5387 840
rect 4796 624 4872 630
rect 4796 598 4804 624
rect 4704 572 4804 598
rect 4856 572 4872 624
rect 4704 570 4872 572
rect 4796 566 4872 570
rect 4476 430 4542 436
rect 4476 378 4484 430
rect 4536 408 4542 430
rect 5136 408 5164 812
rect 5368 788 5387 812
rect 5439 788 5448 840
rect 5368 776 5448 788
rect 5684 844 5752 850
rect 5684 792 5691 844
rect 5743 792 5752 844
rect 5684 786 5752 792
rect 4536 380 5164 408
rect 4536 378 4542 380
rect 4476 372 4542 378
rect 5290 180 5640 194
rect 3402 50 3752 64
rect 5290 64 5311 180
rect 5619 64 5640 180
rect 5684 170 5728 786
rect 5824 616 5852 1200
rect 5886 1150 5948 1156
rect 5886 1098 5896 1150
rect 5984 1142 6012 1714
rect 6040 1541 6104 1548
rect 6040 1489 6046 1541
rect 6098 1508 6104 1541
rect 6366 1508 6416 1898
rect 6888 1896 6916 1996
rect 6888 1890 6954 1896
rect 8002 1894 8030 1996
rect 8238 1958 8304 1966
rect 8238 1906 8244 1958
rect 8296 1906 8304 1958
rect 8238 1898 8304 1906
rect 6888 1876 6896 1890
rect 6890 1838 6896 1876
rect 6948 1838 6954 1890
rect 6890 1832 6954 1838
rect 7962 1888 8030 1894
rect 7962 1836 7972 1888
rect 8024 1836 8030 1888
rect 7962 1830 8030 1836
rect 6802 1774 6866 1780
rect 6802 1744 6808 1774
rect 6592 1722 6808 1744
rect 6860 1722 6866 1774
rect 6592 1716 6866 1722
rect 7872 1776 7940 1782
rect 7872 1724 7880 1776
rect 7932 1724 7940 1776
rect 6098 1492 6418 1508
rect 6098 1489 6432 1492
rect 6040 1486 6432 1489
rect 6040 1480 6374 1486
rect 6366 1434 6374 1480
rect 6426 1434 6432 1486
rect 6366 1428 6432 1434
rect 6236 1292 6308 1304
rect 6236 1240 6246 1292
rect 6298 1240 6308 1292
rect 6236 1228 6308 1240
rect 6272 1226 6308 1228
rect 5984 1114 6272 1142
rect 5886 1092 5948 1098
rect 5920 1046 5948 1092
rect 5920 1042 6164 1046
rect 5920 1036 6202 1042
rect 5920 1018 6142 1036
rect 6136 984 6142 1018
rect 6194 984 6202 1036
rect 6136 976 6202 984
rect 5824 602 5888 616
rect 6244 608 6272 1114
rect 6348 902 6414 910
rect 6348 850 6354 902
rect 6406 850 6414 902
rect 6348 842 6414 850
rect 5824 550 5827 602
rect 5879 550 5888 602
rect 5824 534 5888 550
rect 6058 592 6272 608
rect 6058 540 6059 592
rect 6111 580 6272 592
rect 6111 540 6112 580
rect 6058 524 6112 540
rect 6364 436 6414 842
rect 6592 598 6620 1716
rect 7872 1714 7940 1724
rect 7752 1541 7816 1548
rect 7752 1510 7758 1541
rect 7024 1489 7758 1510
rect 7810 1489 7816 1541
rect 7024 1482 7816 1489
rect 7024 1480 7758 1482
rect 7024 1474 7752 1480
rect 6924 1144 6988 1152
rect 6924 1092 6930 1144
rect 6982 1092 6988 1144
rect 6924 1084 6988 1092
rect 6684 1056 6750 1062
rect 6684 1004 6692 1056
rect 6744 1026 6750 1056
rect 6924 1026 6952 1084
rect 6744 1004 6952 1026
rect 6684 998 6952 1004
rect 7024 848 7052 1474
rect 7752 1408 7818 1414
rect 7752 1356 7760 1408
rect 7812 1356 7818 1408
rect 7752 1350 7818 1356
rect 7752 1228 7780 1350
rect 7712 1200 7780 1228
rect 7024 840 7336 848
rect 7024 812 7275 840
rect 6684 624 6760 630
rect 6684 598 6692 624
rect 6592 572 6692 598
rect 6744 572 6760 624
rect 6592 570 6760 572
rect 6684 566 6760 570
rect 6364 430 6430 436
rect 6364 378 6372 430
rect 6424 408 6430 430
rect 7024 408 7052 812
rect 7256 788 7275 812
rect 7327 788 7336 840
rect 7256 776 7336 788
rect 7572 844 7640 850
rect 7572 792 7579 844
rect 7631 792 7640 844
rect 7572 786 7640 792
rect 6424 380 7052 408
rect 6424 378 6430 380
rect 6364 372 6430 378
rect 7178 180 7528 194
rect 5290 50 5640 64
rect 7178 64 7199 180
rect 7507 64 7528 180
rect 7572 170 7616 786
rect 7712 616 7740 1200
rect 7774 1150 7836 1156
rect 7774 1098 7784 1150
rect 7872 1142 7900 1714
rect 7928 1541 7992 1548
rect 7928 1489 7934 1541
rect 7986 1508 7992 1541
rect 8254 1508 8304 1898
rect 8776 1896 8804 1996
rect 8776 1890 8842 1896
rect 9890 1894 9918 1996
rect 10126 1958 10192 1966
rect 10126 1906 10132 1958
rect 10184 1906 10192 1958
rect 10126 1898 10192 1906
rect 8776 1876 8784 1890
rect 8778 1838 8784 1876
rect 8836 1838 8842 1890
rect 8778 1832 8842 1838
rect 9850 1888 9918 1894
rect 9850 1836 9860 1888
rect 9912 1836 9918 1888
rect 9850 1830 9918 1836
rect 8690 1774 8754 1780
rect 8690 1744 8696 1774
rect 8480 1722 8696 1744
rect 8748 1722 8754 1774
rect 8480 1716 8754 1722
rect 9760 1776 9828 1782
rect 9760 1724 9768 1776
rect 9820 1724 9828 1776
rect 7986 1492 8306 1508
rect 7986 1489 8320 1492
rect 7928 1486 8320 1489
rect 7928 1480 8262 1486
rect 8254 1434 8262 1480
rect 8314 1434 8320 1486
rect 8254 1428 8320 1434
rect 8124 1292 8196 1304
rect 8124 1240 8134 1292
rect 8186 1240 8196 1292
rect 8124 1228 8196 1240
rect 8160 1226 8196 1228
rect 7872 1114 8160 1142
rect 7774 1092 7836 1098
rect 7808 1046 7836 1092
rect 7808 1042 8052 1046
rect 7808 1036 8090 1042
rect 7808 1018 8030 1036
rect 8024 984 8030 1018
rect 8082 984 8090 1036
rect 8024 976 8090 984
rect 7712 602 7776 616
rect 8132 608 8160 1114
rect 8236 902 8302 910
rect 8236 850 8242 902
rect 8294 850 8302 902
rect 8236 842 8302 850
rect 7712 550 7715 602
rect 7767 550 7776 602
rect 7712 534 7776 550
rect 7946 592 8160 608
rect 7946 540 7947 592
rect 7999 580 8160 592
rect 7999 540 8000 580
rect 7946 524 8000 540
rect 8252 436 8302 842
rect 8480 598 8508 1716
rect 9760 1714 9828 1724
rect 9640 1541 9704 1548
rect 9640 1510 9646 1541
rect 8912 1489 9646 1510
rect 9698 1489 9704 1541
rect 8912 1482 9704 1489
rect 8912 1480 9646 1482
rect 8912 1474 9640 1480
rect 8812 1144 8876 1152
rect 8812 1092 8818 1144
rect 8870 1092 8876 1144
rect 8812 1084 8876 1092
rect 8572 1056 8638 1062
rect 8572 1004 8580 1056
rect 8632 1026 8638 1056
rect 8812 1026 8840 1084
rect 8632 1004 8840 1026
rect 8572 998 8840 1004
rect 8912 848 8940 1474
rect 9640 1408 9706 1414
rect 9640 1356 9648 1408
rect 9700 1356 9706 1408
rect 9640 1350 9706 1356
rect 9640 1228 9668 1350
rect 9600 1200 9668 1228
rect 8912 840 9224 848
rect 8912 812 9163 840
rect 8572 624 8648 630
rect 8572 598 8580 624
rect 8480 572 8580 598
rect 8632 572 8648 624
rect 8480 570 8648 572
rect 8572 566 8648 570
rect 8252 430 8318 436
rect 8252 378 8260 430
rect 8312 408 8318 430
rect 8912 408 8940 812
rect 9144 788 9163 812
rect 9215 788 9224 840
rect 9144 776 9224 788
rect 9460 844 9528 850
rect 9460 792 9467 844
rect 9519 792 9528 844
rect 9460 786 9528 792
rect 8312 380 8940 408
rect 8312 378 8318 380
rect 8252 372 8318 378
rect 9066 180 9416 194
rect 7178 50 7528 64
rect 9066 64 9087 180
rect 9395 64 9416 180
rect 9460 170 9504 786
rect 9600 616 9628 1200
rect 9662 1150 9724 1156
rect 9662 1098 9672 1150
rect 9760 1142 9788 1714
rect 9816 1541 9880 1548
rect 9816 1489 9822 1541
rect 9874 1508 9880 1541
rect 10142 1508 10192 1898
rect 10664 1896 10692 1996
rect 10664 1890 10730 1896
rect 11778 1894 11806 1996
rect 12014 1958 12080 1966
rect 12014 1906 12020 1958
rect 12072 1906 12080 1958
rect 12014 1898 12080 1906
rect 10664 1876 10672 1890
rect 10666 1838 10672 1876
rect 10724 1838 10730 1890
rect 10666 1832 10730 1838
rect 11738 1888 11806 1894
rect 11738 1836 11748 1888
rect 11800 1836 11806 1888
rect 11738 1830 11806 1836
rect 10578 1774 10642 1780
rect 10578 1744 10584 1774
rect 10368 1722 10584 1744
rect 10636 1722 10642 1774
rect 10368 1716 10642 1722
rect 11648 1776 11716 1782
rect 11648 1724 11656 1776
rect 11708 1724 11716 1776
rect 9874 1492 10194 1508
rect 9874 1489 10208 1492
rect 9816 1486 10208 1489
rect 9816 1480 10150 1486
rect 10142 1434 10150 1480
rect 10202 1434 10208 1486
rect 10142 1428 10208 1434
rect 10012 1292 10084 1304
rect 10012 1240 10022 1292
rect 10074 1240 10084 1292
rect 10012 1228 10084 1240
rect 10048 1226 10084 1228
rect 9760 1114 10048 1142
rect 9662 1092 9724 1098
rect 9696 1046 9724 1092
rect 9696 1042 9940 1046
rect 9696 1036 9978 1042
rect 9696 1018 9918 1036
rect 9912 984 9918 1018
rect 9970 984 9978 1036
rect 9912 976 9978 984
rect 9600 602 9664 616
rect 10020 608 10048 1114
rect 10124 902 10190 910
rect 10124 850 10130 902
rect 10182 850 10190 902
rect 10124 842 10190 850
rect 9600 550 9603 602
rect 9655 550 9664 602
rect 9600 534 9664 550
rect 9834 592 10048 608
rect 9834 540 9835 592
rect 9887 580 10048 592
rect 9887 540 9888 580
rect 9834 524 9888 540
rect 10140 436 10190 842
rect 10368 598 10396 1716
rect 11648 1714 11716 1724
rect 11528 1541 11592 1548
rect 11528 1510 11534 1541
rect 10800 1489 11534 1510
rect 11586 1489 11592 1541
rect 10800 1482 11592 1489
rect 10800 1480 11534 1482
rect 10800 1474 11528 1480
rect 10700 1144 10764 1152
rect 10700 1092 10706 1144
rect 10758 1092 10764 1144
rect 10700 1084 10764 1092
rect 10460 1056 10526 1062
rect 10460 1004 10468 1056
rect 10520 1026 10526 1056
rect 10700 1026 10728 1084
rect 10520 1004 10728 1026
rect 10460 998 10728 1004
rect 10800 848 10828 1474
rect 11528 1408 11594 1414
rect 11528 1356 11536 1408
rect 11588 1356 11594 1408
rect 11528 1350 11594 1356
rect 11528 1228 11556 1350
rect 11488 1200 11556 1228
rect 10800 840 11112 848
rect 10800 812 11051 840
rect 10460 624 10536 630
rect 10460 598 10468 624
rect 10368 572 10468 598
rect 10520 572 10536 624
rect 10368 570 10536 572
rect 10460 566 10536 570
rect 10140 430 10206 436
rect 10140 378 10148 430
rect 10200 408 10206 430
rect 10800 408 10828 812
rect 11032 788 11051 812
rect 11103 788 11112 840
rect 11032 776 11112 788
rect 11348 844 11416 850
rect 11348 792 11355 844
rect 11407 792 11416 844
rect 11348 786 11416 792
rect 10200 380 10828 408
rect 10200 378 10206 380
rect 10140 372 10206 378
rect 10954 180 11304 194
rect 9066 50 9416 64
rect 10954 64 10975 180
rect 11283 64 11304 180
rect 11348 170 11392 786
rect 11488 616 11516 1200
rect 11550 1150 11612 1156
rect 11550 1098 11560 1150
rect 11648 1142 11676 1714
rect 11704 1541 11768 1548
rect 11704 1489 11710 1541
rect 11762 1508 11768 1541
rect 12030 1508 12080 1898
rect 12552 1896 12580 1996
rect 12552 1890 12618 1896
rect 13666 1894 13694 1996
rect 13902 1958 13968 1966
rect 13902 1906 13908 1958
rect 13960 1906 13968 1958
rect 13902 1898 13968 1906
rect 12552 1876 12560 1890
rect 12554 1838 12560 1876
rect 12612 1838 12618 1890
rect 12554 1832 12618 1838
rect 13626 1888 13694 1894
rect 13626 1836 13636 1888
rect 13688 1836 13694 1888
rect 13626 1830 13694 1836
rect 12466 1774 12530 1780
rect 12466 1744 12472 1774
rect 12256 1722 12472 1744
rect 12524 1722 12530 1774
rect 12256 1716 12530 1722
rect 13536 1776 13604 1782
rect 13536 1724 13544 1776
rect 13596 1724 13604 1776
rect 11762 1492 12082 1508
rect 11762 1489 12096 1492
rect 11704 1486 12096 1489
rect 11704 1480 12038 1486
rect 12030 1434 12038 1480
rect 12090 1434 12096 1486
rect 12030 1428 12096 1434
rect 11900 1292 11972 1304
rect 11900 1240 11910 1292
rect 11962 1240 11972 1292
rect 11900 1228 11972 1240
rect 11936 1226 11972 1228
rect 11648 1114 11936 1142
rect 11550 1092 11612 1098
rect 11584 1046 11612 1092
rect 11584 1042 11828 1046
rect 11584 1036 11866 1042
rect 11584 1018 11806 1036
rect 11800 984 11806 1018
rect 11858 984 11866 1036
rect 11800 976 11866 984
rect 11488 602 11552 616
rect 11908 608 11936 1114
rect 12012 902 12078 910
rect 12012 850 12018 902
rect 12070 850 12078 902
rect 12012 842 12078 850
rect 11488 550 11491 602
rect 11543 550 11552 602
rect 11488 534 11552 550
rect 11722 592 11936 608
rect 11722 540 11723 592
rect 11775 580 11936 592
rect 11775 540 11776 580
rect 11722 524 11776 540
rect 12028 436 12078 842
rect 12256 598 12284 1716
rect 13536 1714 13604 1724
rect 13416 1541 13480 1548
rect 13416 1510 13422 1541
rect 12688 1489 13422 1510
rect 13474 1489 13480 1541
rect 12688 1482 13480 1489
rect 12688 1480 13422 1482
rect 12688 1474 13416 1480
rect 12588 1144 12652 1152
rect 12588 1092 12594 1144
rect 12646 1092 12652 1144
rect 12588 1084 12652 1092
rect 12348 1056 12414 1062
rect 12348 1004 12356 1056
rect 12408 1026 12414 1056
rect 12588 1026 12616 1084
rect 12408 1004 12616 1026
rect 12348 998 12616 1004
rect 12688 848 12716 1474
rect 13416 1408 13482 1414
rect 13416 1356 13424 1408
rect 13476 1356 13482 1408
rect 13416 1350 13482 1356
rect 13416 1228 13444 1350
rect 13376 1200 13444 1228
rect 12688 840 13000 848
rect 12688 812 12939 840
rect 12348 624 12424 630
rect 12348 598 12356 624
rect 12256 572 12356 598
rect 12408 572 12424 624
rect 12256 570 12424 572
rect 12348 566 12424 570
rect 12028 430 12094 436
rect 12028 378 12036 430
rect 12088 408 12094 430
rect 12688 408 12716 812
rect 12920 788 12939 812
rect 12991 788 13000 840
rect 12920 776 13000 788
rect 13236 844 13304 850
rect 13236 792 13243 844
rect 13295 792 13304 844
rect 13236 786 13304 792
rect 12088 380 12716 408
rect 12088 378 12094 380
rect 12028 372 12094 378
rect 12842 180 13192 194
rect 10954 50 11304 64
rect 12842 64 12863 180
rect 13171 64 13192 180
rect 13236 170 13280 786
rect 13376 616 13404 1200
rect 13438 1150 13500 1156
rect 13438 1098 13448 1150
rect 13536 1142 13564 1714
rect 13592 1541 13656 1548
rect 13592 1489 13598 1541
rect 13650 1508 13656 1541
rect 13918 1508 13968 1898
rect 14440 1896 14468 1996
rect 14440 1890 14506 1896
rect 15548 1894 15576 2000
rect 15784 1958 15850 1966
rect 15784 1906 15790 1958
rect 15842 1906 15850 1958
rect 15784 1898 15850 1906
rect 14440 1876 14448 1890
rect 14442 1838 14448 1876
rect 14500 1838 14506 1890
rect 14442 1832 14506 1838
rect 15508 1888 15576 1894
rect 15508 1836 15518 1888
rect 15570 1836 15576 1888
rect 15508 1830 15576 1836
rect 14354 1774 14418 1780
rect 14354 1744 14360 1774
rect 14144 1722 14360 1744
rect 14412 1722 14418 1774
rect 14144 1716 14418 1722
rect 15418 1776 15486 1782
rect 15418 1724 15426 1776
rect 15478 1724 15486 1776
rect 13650 1492 13970 1508
rect 13650 1489 13984 1492
rect 13592 1486 13984 1489
rect 13592 1480 13926 1486
rect 13918 1434 13926 1480
rect 13978 1434 13984 1486
rect 13918 1428 13984 1434
rect 13788 1292 13860 1304
rect 13788 1240 13798 1292
rect 13850 1240 13860 1292
rect 13788 1228 13860 1240
rect 13824 1226 13860 1228
rect 13536 1114 13824 1142
rect 13438 1092 13500 1098
rect 13472 1046 13500 1092
rect 13472 1042 13716 1046
rect 13472 1036 13754 1042
rect 13472 1018 13694 1036
rect 13688 984 13694 1018
rect 13746 984 13754 1036
rect 13688 976 13754 984
rect 13376 602 13440 616
rect 13796 608 13824 1114
rect 13900 902 13966 910
rect 13900 850 13906 902
rect 13958 850 13966 902
rect 13900 842 13966 850
rect 13376 550 13379 602
rect 13431 550 13440 602
rect 13376 534 13440 550
rect 13610 592 13824 608
rect 13610 540 13611 592
rect 13663 580 13824 592
rect 13663 540 13664 580
rect 13610 524 13664 540
rect 13916 436 13966 842
rect 14144 598 14172 1716
rect 15418 1714 15486 1724
rect 15298 1541 15362 1548
rect 15298 1510 15304 1541
rect 14576 1489 15304 1510
rect 15356 1489 15362 1541
rect 14576 1482 15362 1489
rect 14576 1480 15304 1482
rect 14576 1474 15298 1480
rect 14476 1144 14540 1152
rect 14476 1092 14482 1144
rect 14534 1092 14540 1144
rect 14476 1084 14540 1092
rect 14236 1056 14302 1062
rect 14236 1004 14244 1056
rect 14296 1026 14302 1056
rect 14476 1026 14504 1084
rect 14296 1004 14504 1026
rect 14236 998 14504 1004
rect 14576 848 14604 1474
rect 15298 1408 15364 1414
rect 15298 1356 15306 1408
rect 15358 1356 15364 1408
rect 15298 1350 15364 1356
rect 15298 1228 15326 1350
rect 15258 1200 15326 1228
rect 14576 840 14888 848
rect 14576 812 14827 840
rect 14236 624 14312 630
rect 14236 598 14244 624
rect 14144 572 14244 598
rect 14296 572 14312 624
rect 14144 570 14312 572
rect 14236 566 14312 570
rect 13916 430 13982 436
rect 13916 378 13924 430
rect 13976 408 13982 430
rect 14576 408 14604 812
rect 14808 788 14827 812
rect 14879 788 14888 840
rect 14808 776 14888 788
rect 15118 844 15186 850
rect 15118 792 15125 844
rect 15177 792 15186 844
rect 15118 786 15186 792
rect 13976 380 14604 408
rect 13976 378 13982 380
rect 13916 372 13982 378
rect 14730 180 15080 194
rect 12842 50 13192 64
rect 14730 64 14751 180
rect 15059 64 15080 180
rect 15118 170 15168 786
rect 15258 616 15286 1200
rect 15320 1150 15382 1156
rect 15320 1098 15330 1150
rect 15418 1142 15446 1714
rect 15474 1541 15538 1548
rect 15474 1489 15480 1541
rect 15532 1508 15538 1541
rect 15800 1508 15850 1898
rect 16322 1896 16350 2000
rect 16322 1890 16388 1896
rect 17436 1894 17464 2000
rect 17672 1958 17738 1966
rect 17672 1906 17678 1958
rect 17730 1906 17738 1958
rect 17672 1898 17738 1906
rect 16322 1876 16330 1890
rect 16324 1838 16330 1876
rect 16382 1838 16388 1890
rect 16324 1832 16388 1838
rect 17396 1888 17464 1894
rect 17396 1836 17406 1888
rect 17458 1836 17464 1888
rect 17396 1830 17464 1836
rect 16236 1774 16300 1780
rect 16236 1744 16242 1774
rect 16026 1722 16242 1744
rect 16294 1722 16300 1774
rect 16026 1716 16300 1722
rect 17306 1776 17374 1782
rect 17306 1724 17314 1776
rect 17366 1724 17374 1776
rect 15532 1492 15852 1508
rect 15532 1489 15866 1492
rect 15474 1486 15866 1489
rect 15474 1480 15808 1486
rect 15800 1434 15808 1480
rect 15860 1434 15866 1486
rect 15800 1428 15866 1434
rect 15670 1292 15742 1304
rect 15670 1240 15680 1292
rect 15732 1240 15742 1292
rect 15670 1228 15742 1240
rect 15706 1226 15742 1228
rect 15418 1114 15706 1142
rect 15320 1092 15382 1098
rect 15354 1046 15382 1092
rect 15354 1042 15598 1046
rect 15354 1036 15636 1042
rect 15354 1018 15576 1036
rect 15570 984 15576 1018
rect 15628 984 15636 1036
rect 15570 976 15636 984
rect 15258 602 15322 616
rect 15678 608 15706 1114
rect 15782 902 15848 910
rect 15782 850 15788 902
rect 15840 850 15848 902
rect 15782 842 15848 850
rect 15258 550 15261 602
rect 15313 550 15322 602
rect 15258 534 15322 550
rect 15492 592 15706 608
rect 15492 540 15493 592
rect 15545 580 15706 592
rect 15545 540 15546 580
rect 15492 524 15546 540
rect 15798 436 15848 842
rect 16026 598 16054 1716
rect 17306 1714 17374 1724
rect 17186 1541 17250 1548
rect 17186 1510 17192 1541
rect 16458 1489 17192 1510
rect 17244 1489 17250 1541
rect 16458 1482 17250 1489
rect 16458 1480 17192 1482
rect 16458 1474 17186 1480
rect 16358 1144 16422 1152
rect 16358 1092 16364 1144
rect 16416 1092 16422 1144
rect 16358 1084 16422 1092
rect 16118 1056 16184 1062
rect 16118 1004 16126 1056
rect 16178 1026 16184 1056
rect 16358 1026 16386 1084
rect 16178 1004 16386 1026
rect 16118 998 16386 1004
rect 16458 848 16486 1474
rect 17186 1408 17252 1414
rect 17186 1356 17194 1408
rect 17246 1356 17252 1408
rect 17186 1350 17252 1356
rect 17186 1228 17214 1350
rect 17146 1200 17214 1228
rect 16458 840 16770 848
rect 16458 812 16709 840
rect 16118 624 16194 630
rect 16118 598 16126 624
rect 16026 572 16126 598
rect 16178 572 16194 624
rect 16026 570 16194 572
rect 16118 566 16194 570
rect 15798 430 15864 436
rect 15798 378 15806 430
rect 15858 408 15864 430
rect 16458 408 16486 812
rect 16690 788 16709 812
rect 16761 788 16770 840
rect 16690 776 16770 788
rect 17006 844 17074 850
rect 17006 792 17013 844
rect 17065 792 17074 844
rect 17006 786 17074 792
rect 15858 380 16486 408
rect 15858 378 15864 380
rect 15798 372 15864 378
rect 16612 180 16962 194
rect 14730 50 15080 64
rect 16612 64 16633 180
rect 16941 64 16962 180
rect 17006 170 17056 786
rect 17146 616 17174 1200
rect 17208 1150 17270 1156
rect 17208 1098 17218 1150
rect 17306 1142 17334 1714
rect 17362 1541 17426 1548
rect 17362 1489 17368 1541
rect 17420 1508 17426 1541
rect 17688 1508 17738 1898
rect 18210 1896 18238 2000
rect 18210 1890 18276 1896
rect 19324 1894 19352 2000
rect 19560 1958 19626 1966
rect 19560 1906 19566 1958
rect 19618 1906 19626 1958
rect 19560 1898 19626 1906
rect 18210 1876 18218 1890
rect 18212 1838 18218 1876
rect 18270 1838 18276 1890
rect 18212 1832 18276 1838
rect 19284 1888 19352 1894
rect 19284 1836 19294 1888
rect 19346 1836 19352 1888
rect 19284 1830 19352 1836
rect 18124 1774 18188 1780
rect 18124 1744 18130 1774
rect 17914 1722 18130 1744
rect 18182 1722 18188 1774
rect 17914 1716 18188 1722
rect 19194 1776 19262 1782
rect 19194 1724 19202 1776
rect 19254 1724 19262 1776
rect 17420 1492 17740 1508
rect 17420 1489 17754 1492
rect 17362 1486 17754 1489
rect 17362 1480 17696 1486
rect 17688 1434 17696 1480
rect 17748 1434 17754 1486
rect 17688 1428 17754 1434
rect 17558 1292 17630 1304
rect 17558 1240 17568 1292
rect 17620 1240 17630 1292
rect 17558 1228 17630 1240
rect 17594 1226 17630 1228
rect 17306 1114 17594 1142
rect 17208 1092 17270 1098
rect 17242 1046 17270 1092
rect 17242 1042 17486 1046
rect 17242 1036 17524 1042
rect 17242 1018 17464 1036
rect 17458 984 17464 1018
rect 17516 984 17524 1036
rect 17458 976 17524 984
rect 17146 602 17210 616
rect 17566 608 17594 1114
rect 17670 902 17736 910
rect 17670 850 17676 902
rect 17728 850 17736 902
rect 17670 842 17736 850
rect 17146 550 17149 602
rect 17201 550 17210 602
rect 17146 534 17210 550
rect 17380 592 17594 608
rect 17380 540 17381 592
rect 17433 580 17594 592
rect 17433 540 17434 580
rect 17380 524 17434 540
rect 17686 436 17736 842
rect 17914 598 17942 1716
rect 19194 1714 19262 1724
rect 19074 1541 19138 1548
rect 19074 1510 19080 1541
rect 18346 1489 19080 1510
rect 19132 1489 19138 1541
rect 18346 1482 19138 1489
rect 18346 1480 19080 1482
rect 18346 1474 19074 1480
rect 18246 1144 18310 1152
rect 18246 1092 18252 1144
rect 18304 1092 18310 1144
rect 18246 1084 18310 1092
rect 18006 1056 18072 1062
rect 18006 1004 18014 1056
rect 18066 1026 18072 1056
rect 18246 1026 18274 1084
rect 18066 1004 18274 1026
rect 18006 998 18274 1004
rect 18346 848 18374 1474
rect 19074 1408 19140 1414
rect 19074 1356 19082 1408
rect 19134 1356 19140 1408
rect 19074 1350 19140 1356
rect 19074 1228 19102 1350
rect 19034 1200 19102 1228
rect 18346 840 18658 848
rect 18346 812 18597 840
rect 18006 624 18082 630
rect 18006 598 18014 624
rect 17914 572 18014 598
rect 18066 572 18082 624
rect 17914 570 18082 572
rect 18006 566 18082 570
rect 17686 430 17752 436
rect 17686 378 17694 430
rect 17746 408 17752 430
rect 18346 408 18374 812
rect 18578 788 18597 812
rect 18649 788 18658 840
rect 18578 776 18658 788
rect 18894 844 18962 850
rect 18894 792 18901 844
rect 18953 792 18962 844
rect 18894 786 18962 792
rect 17746 380 18374 408
rect 17746 378 17752 380
rect 17686 372 17752 378
rect 18500 180 18850 194
rect 16612 50 16962 64
rect 18500 64 18521 180
rect 18829 64 18850 180
rect 18894 170 18944 786
rect 19034 616 19062 1200
rect 19096 1150 19158 1156
rect 19096 1098 19106 1150
rect 19194 1142 19222 1714
rect 19250 1541 19314 1548
rect 19250 1489 19256 1541
rect 19308 1508 19314 1541
rect 19576 1508 19626 1898
rect 20098 1896 20126 2000
rect 20800 1996 22120 2000
rect 22684 1996 24008 2000
rect 20098 1890 20164 1896
rect 21212 1894 21240 1996
rect 21448 1958 21514 1966
rect 21448 1906 21454 1958
rect 21506 1906 21514 1958
rect 21448 1898 21514 1906
rect 20098 1876 20106 1890
rect 20100 1838 20106 1876
rect 20158 1838 20164 1890
rect 20100 1832 20164 1838
rect 21172 1888 21240 1894
rect 21172 1836 21182 1888
rect 21234 1836 21240 1888
rect 21172 1830 21240 1836
rect 20012 1774 20076 1780
rect 20012 1744 20018 1774
rect 19802 1722 20018 1744
rect 20070 1722 20076 1774
rect 19802 1716 20076 1722
rect 21082 1776 21150 1782
rect 21082 1724 21090 1776
rect 21142 1724 21150 1776
rect 19308 1492 19628 1508
rect 19308 1489 19642 1492
rect 19250 1486 19642 1489
rect 19250 1480 19584 1486
rect 19576 1434 19584 1480
rect 19636 1434 19642 1486
rect 19576 1428 19642 1434
rect 19446 1292 19518 1304
rect 19446 1240 19456 1292
rect 19508 1240 19518 1292
rect 19446 1228 19518 1240
rect 19482 1226 19518 1228
rect 19194 1114 19482 1142
rect 19096 1092 19158 1098
rect 19130 1046 19158 1092
rect 19130 1042 19374 1046
rect 19130 1036 19412 1042
rect 19130 1018 19352 1036
rect 19346 984 19352 1018
rect 19404 984 19412 1036
rect 19346 976 19412 984
rect 19034 602 19098 616
rect 19454 608 19482 1114
rect 19558 902 19624 910
rect 19558 850 19564 902
rect 19616 850 19624 902
rect 19558 842 19624 850
rect 19034 550 19037 602
rect 19089 550 19098 602
rect 19034 534 19098 550
rect 19268 592 19482 608
rect 19268 540 19269 592
rect 19321 580 19482 592
rect 19321 540 19322 580
rect 19268 524 19322 540
rect 19574 436 19624 842
rect 19802 598 19830 1716
rect 21082 1714 21150 1724
rect 20962 1541 21026 1548
rect 20962 1510 20968 1541
rect 20234 1489 20968 1510
rect 21020 1489 21026 1541
rect 20234 1482 21026 1489
rect 20234 1480 20968 1482
rect 20234 1474 20962 1480
rect 20134 1144 20198 1152
rect 20134 1092 20140 1144
rect 20192 1092 20198 1144
rect 20134 1084 20198 1092
rect 19894 1056 19960 1062
rect 19894 1004 19902 1056
rect 19954 1026 19960 1056
rect 20134 1026 20162 1084
rect 19954 1004 20162 1026
rect 19894 998 20162 1004
rect 20234 848 20262 1474
rect 20962 1408 21028 1414
rect 20962 1356 20970 1408
rect 21022 1356 21028 1408
rect 20962 1350 21028 1356
rect 20962 1228 20990 1350
rect 20922 1200 20990 1228
rect 20234 840 20546 848
rect 20234 812 20485 840
rect 19894 624 19970 630
rect 19894 598 19902 624
rect 19802 572 19902 598
rect 19954 572 19970 624
rect 19802 570 19970 572
rect 19894 566 19970 570
rect 19574 430 19640 436
rect 19574 378 19582 430
rect 19634 408 19640 430
rect 20234 408 20262 812
rect 20466 788 20485 812
rect 20537 788 20546 840
rect 20466 776 20546 788
rect 20782 844 20850 850
rect 20782 792 20789 844
rect 20841 792 20850 844
rect 20782 786 20850 792
rect 19634 380 20262 408
rect 19634 378 19640 380
rect 19574 372 19640 378
rect 20388 180 20738 194
rect 18500 50 18850 64
rect 20388 64 20409 180
rect 20717 64 20738 180
rect 20782 170 20832 786
rect 20922 616 20950 1200
rect 20984 1150 21046 1156
rect 20984 1098 20994 1150
rect 21082 1142 21110 1714
rect 21138 1541 21202 1548
rect 21138 1489 21144 1541
rect 21196 1508 21202 1541
rect 21464 1508 21514 1898
rect 21986 1896 22014 1996
rect 21986 1890 22052 1896
rect 23100 1894 23128 1996
rect 23336 1958 23402 1966
rect 23336 1906 23342 1958
rect 23394 1906 23402 1958
rect 23336 1898 23402 1906
rect 21986 1876 21994 1890
rect 21988 1838 21994 1876
rect 22046 1838 22052 1890
rect 21988 1832 22052 1838
rect 23060 1888 23128 1894
rect 23060 1836 23070 1888
rect 23122 1836 23128 1888
rect 23060 1830 23128 1836
rect 21900 1774 21964 1780
rect 21900 1744 21906 1774
rect 21690 1722 21906 1744
rect 21958 1722 21964 1774
rect 21690 1716 21964 1722
rect 22970 1776 23038 1782
rect 22970 1724 22978 1776
rect 23030 1724 23038 1776
rect 21196 1492 21516 1508
rect 21196 1489 21530 1492
rect 21138 1486 21530 1489
rect 21138 1480 21472 1486
rect 21464 1434 21472 1480
rect 21524 1434 21530 1486
rect 21464 1428 21530 1434
rect 21334 1292 21406 1304
rect 21334 1240 21344 1292
rect 21396 1240 21406 1292
rect 21334 1228 21406 1240
rect 21370 1226 21406 1228
rect 21082 1114 21370 1142
rect 20984 1092 21046 1098
rect 21018 1046 21046 1092
rect 21018 1042 21262 1046
rect 21018 1036 21300 1042
rect 21018 1018 21240 1036
rect 21234 984 21240 1018
rect 21292 984 21300 1036
rect 21234 976 21300 984
rect 20922 602 20986 616
rect 21342 608 21370 1114
rect 21446 902 21512 910
rect 21446 850 21452 902
rect 21504 850 21512 902
rect 21446 842 21512 850
rect 20922 550 20925 602
rect 20977 550 20986 602
rect 20922 534 20986 550
rect 21156 592 21370 608
rect 21156 540 21157 592
rect 21209 580 21370 592
rect 21209 540 21210 580
rect 21156 524 21210 540
rect 21462 436 21512 842
rect 21690 598 21718 1716
rect 22970 1714 23038 1724
rect 22850 1541 22914 1548
rect 22850 1510 22856 1541
rect 22122 1489 22856 1510
rect 22908 1489 22914 1541
rect 22122 1482 22914 1489
rect 22122 1480 22856 1482
rect 22122 1474 22850 1480
rect 22022 1144 22086 1152
rect 22022 1092 22028 1144
rect 22080 1092 22086 1144
rect 22022 1084 22086 1092
rect 21782 1056 21848 1062
rect 21782 1004 21790 1056
rect 21842 1026 21848 1056
rect 22022 1026 22050 1084
rect 21842 1004 22050 1026
rect 21782 998 22050 1004
rect 22122 848 22150 1474
rect 22850 1408 22916 1414
rect 22850 1356 22858 1408
rect 22910 1356 22916 1408
rect 22850 1350 22916 1356
rect 22850 1228 22878 1350
rect 22810 1200 22878 1228
rect 22122 840 22434 848
rect 22122 812 22373 840
rect 21782 624 21858 630
rect 21782 598 21790 624
rect 21690 572 21790 598
rect 21842 572 21858 624
rect 21690 570 21858 572
rect 21782 566 21858 570
rect 21462 430 21528 436
rect 21462 378 21470 430
rect 21522 408 21528 430
rect 22122 408 22150 812
rect 22354 788 22373 812
rect 22425 788 22434 840
rect 22354 776 22434 788
rect 22670 844 22738 850
rect 22670 792 22677 844
rect 22729 792 22738 844
rect 22670 786 22738 792
rect 21522 380 22150 408
rect 21522 378 21528 380
rect 21462 372 21528 378
rect 22276 180 22626 194
rect 20388 50 20738 64
rect 22276 64 22297 180
rect 22605 64 22626 180
rect 22670 170 22720 786
rect 22810 616 22838 1200
rect 22872 1150 22934 1156
rect 22872 1098 22882 1150
rect 22970 1142 22998 1714
rect 23026 1541 23090 1548
rect 23026 1489 23032 1541
rect 23084 1508 23090 1541
rect 23352 1508 23402 1898
rect 23874 1896 23902 1996
rect 23874 1890 23940 1896
rect 24988 1894 25016 2000
rect 25224 1958 25290 1966
rect 25224 1906 25230 1958
rect 25282 1906 25290 1958
rect 25224 1898 25290 1906
rect 23874 1876 23882 1890
rect 23876 1838 23882 1876
rect 23934 1838 23940 1890
rect 23876 1832 23940 1838
rect 24948 1888 25016 1894
rect 24948 1836 24958 1888
rect 25010 1836 25016 1888
rect 24948 1830 25016 1836
rect 23788 1774 23852 1780
rect 23788 1744 23794 1774
rect 23578 1722 23794 1744
rect 23846 1722 23852 1774
rect 23578 1716 23852 1722
rect 24858 1776 24926 1782
rect 24858 1724 24866 1776
rect 24918 1724 24926 1776
rect 23084 1492 23404 1508
rect 23084 1489 23418 1492
rect 23026 1486 23418 1489
rect 23026 1480 23360 1486
rect 23352 1434 23360 1480
rect 23412 1434 23418 1486
rect 23352 1428 23418 1434
rect 23222 1292 23294 1304
rect 23222 1240 23232 1292
rect 23284 1240 23294 1292
rect 23222 1228 23294 1240
rect 23258 1226 23294 1228
rect 22970 1114 23258 1142
rect 22872 1092 22934 1098
rect 22906 1046 22934 1092
rect 22906 1042 23150 1046
rect 22906 1036 23188 1042
rect 22906 1018 23128 1036
rect 23122 984 23128 1018
rect 23180 984 23188 1036
rect 23122 976 23188 984
rect 22810 602 22874 616
rect 23230 608 23258 1114
rect 23334 902 23400 910
rect 23334 850 23340 902
rect 23392 850 23400 902
rect 23334 842 23400 850
rect 22810 550 22813 602
rect 22865 550 22874 602
rect 22810 534 22874 550
rect 23044 592 23258 608
rect 23044 540 23045 592
rect 23097 580 23258 592
rect 23097 540 23098 580
rect 23044 524 23098 540
rect 23350 436 23400 842
rect 23578 598 23606 1716
rect 24858 1714 24926 1724
rect 24738 1541 24802 1548
rect 24738 1510 24744 1541
rect 24010 1489 24744 1510
rect 24796 1489 24802 1541
rect 24010 1482 24802 1489
rect 24010 1480 24744 1482
rect 24010 1474 24738 1480
rect 23910 1144 23974 1152
rect 23910 1092 23916 1144
rect 23968 1092 23974 1144
rect 23910 1084 23974 1092
rect 23670 1056 23736 1062
rect 23670 1004 23678 1056
rect 23730 1026 23736 1056
rect 23910 1026 23938 1084
rect 23730 1004 23938 1026
rect 23670 998 23938 1004
rect 24010 848 24038 1474
rect 24738 1408 24804 1414
rect 24738 1356 24746 1408
rect 24798 1356 24804 1408
rect 24738 1350 24804 1356
rect 24738 1228 24766 1350
rect 24698 1200 24766 1228
rect 24010 840 24322 848
rect 24010 812 24261 840
rect 23670 624 23746 630
rect 23670 598 23678 624
rect 23578 572 23678 598
rect 23730 572 23746 624
rect 23578 570 23746 572
rect 23670 566 23746 570
rect 23350 430 23416 436
rect 23350 378 23358 430
rect 23410 408 23416 430
rect 24010 408 24038 812
rect 24242 788 24261 812
rect 24313 788 24322 840
rect 24242 776 24322 788
rect 24558 844 24626 850
rect 24558 792 24565 844
rect 24617 792 24626 844
rect 24558 786 24626 792
rect 23410 380 24038 408
rect 23410 378 23416 380
rect 23350 372 23416 378
rect 24164 180 24514 194
rect 22276 50 22626 64
rect 24164 64 24185 180
rect 24493 64 24514 180
rect 24558 170 24608 786
rect 24698 616 24726 1200
rect 24760 1150 24822 1156
rect 24760 1098 24770 1150
rect 24858 1142 24886 1714
rect 24914 1541 24978 1548
rect 24914 1489 24920 1541
rect 24972 1508 24978 1541
rect 25240 1508 25290 1898
rect 25762 1896 25790 2000
rect 25762 1890 25828 1896
rect 26876 1894 26904 2000
rect 27112 1958 27178 1966
rect 27112 1906 27118 1958
rect 27170 1906 27178 1958
rect 27112 1898 27178 1906
rect 25762 1876 25770 1890
rect 25764 1838 25770 1876
rect 25822 1838 25828 1890
rect 25764 1832 25828 1838
rect 26836 1888 26904 1894
rect 26836 1836 26846 1888
rect 26898 1836 26904 1888
rect 26836 1830 26904 1836
rect 25676 1774 25740 1780
rect 25676 1744 25682 1774
rect 25466 1722 25682 1744
rect 25734 1722 25740 1774
rect 25466 1716 25740 1722
rect 26746 1776 26814 1782
rect 26746 1724 26754 1776
rect 26806 1724 26814 1776
rect 24972 1492 25292 1508
rect 24972 1489 25306 1492
rect 24914 1486 25306 1489
rect 24914 1480 25248 1486
rect 25240 1434 25248 1480
rect 25300 1434 25306 1486
rect 25240 1428 25306 1434
rect 25110 1292 25182 1304
rect 25110 1240 25120 1292
rect 25172 1240 25182 1292
rect 25110 1228 25182 1240
rect 25146 1226 25182 1228
rect 24858 1114 25146 1142
rect 24760 1092 24822 1098
rect 24794 1046 24822 1092
rect 24794 1042 25038 1046
rect 24794 1036 25076 1042
rect 24794 1018 25016 1036
rect 25010 984 25016 1018
rect 25068 984 25076 1036
rect 25010 976 25076 984
rect 24698 602 24762 616
rect 25118 608 25146 1114
rect 25222 902 25288 910
rect 25222 850 25228 902
rect 25280 850 25288 902
rect 25222 842 25288 850
rect 24698 550 24701 602
rect 24753 550 24762 602
rect 24698 534 24762 550
rect 24932 592 25146 608
rect 24932 540 24933 592
rect 24985 580 25146 592
rect 24985 540 24986 580
rect 24932 524 24986 540
rect 25238 436 25288 842
rect 25466 598 25494 1716
rect 26746 1714 26814 1724
rect 26626 1541 26690 1548
rect 26626 1510 26632 1541
rect 25898 1489 26632 1510
rect 26684 1489 26690 1541
rect 25898 1482 26690 1489
rect 25898 1480 26632 1482
rect 25898 1474 26626 1480
rect 25798 1144 25862 1152
rect 25798 1092 25804 1144
rect 25856 1092 25862 1144
rect 25798 1084 25862 1092
rect 25558 1056 25624 1062
rect 25558 1004 25566 1056
rect 25618 1026 25624 1056
rect 25798 1026 25826 1084
rect 25618 1004 25826 1026
rect 25558 998 25826 1004
rect 25898 848 25926 1474
rect 26626 1408 26692 1414
rect 26626 1356 26634 1408
rect 26686 1356 26692 1408
rect 26626 1350 26692 1356
rect 26626 1228 26654 1350
rect 26586 1200 26654 1228
rect 25898 840 26210 848
rect 25898 812 26149 840
rect 25558 624 25634 630
rect 25558 598 25566 624
rect 25466 572 25566 598
rect 25618 572 25634 624
rect 25466 570 25634 572
rect 25558 566 25634 570
rect 25238 430 25304 436
rect 25238 378 25246 430
rect 25298 408 25304 430
rect 25898 408 25926 812
rect 26130 788 26149 812
rect 26201 788 26210 840
rect 26130 776 26210 788
rect 26446 844 26514 850
rect 26446 792 26453 844
rect 26505 792 26514 844
rect 26446 786 26514 792
rect 25298 380 25926 408
rect 25298 378 25304 380
rect 25238 372 25304 378
rect 26052 180 26402 194
rect 24164 50 24514 64
rect 26052 64 26073 180
rect 26381 64 26402 180
rect 26446 170 26496 786
rect 26586 616 26614 1200
rect 26648 1150 26710 1156
rect 26648 1098 26658 1150
rect 26746 1142 26774 1714
rect 26802 1541 26866 1548
rect 26802 1489 26808 1541
rect 26860 1508 26866 1541
rect 27128 1508 27178 1898
rect 27650 1896 27678 2000
rect 27650 1890 27716 1896
rect 28764 1894 28792 2000
rect 29000 1958 29066 1966
rect 29000 1906 29006 1958
rect 29058 1906 29066 1958
rect 29000 1898 29066 1906
rect 27650 1876 27658 1890
rect 27652 1838 27658 1876
rect 27710 1838 27716 1890
rect 27652 1832 27716 1838
rect 28724 1888 28792 1894
rect 28724 1836 28734 1888
rect 28786 1836 28792 1888
rect 28724 1830 28792 1836
rect 27564 1774 27628 1780
rect 27564 1744 27570 1774
rect 27354 1722 27570 1744
rect 27622 1722 27628 1774
rect 27354 1716 27628 1722
rect 28634 1776 28702 1782
rect 28634 1724 28642 1776
rect 28694 1724 28702 1776
rect 26860 1492 27180 1508
rect 26860 1489 27194 1492
rect 26802 1486 27194 1489
rect 26802 1480 27136 1486
rect 27128 1434 27136 1480
rect 27188 1434 27194 1486
rect 27128 1428 27194 1434
rect 26998 1292 27070 1304
rect 26998 1240 27008 1292
rect 27060 1240 27070 1292
rect 26998 1228 27070 1240
rect 27034 1226 27070 1228
rect 26746 1114 27034 1142
rect 26648 1092 26710 1098
rect 26682 1046 26710 1092
rect 26682 1042 26926 1046
rect 26682 1036 26964 1042
rect 26682 1018 26904 1036
rect 26898 984 26904 1018
rect 26956 984 26964 1036
rect 26898 976 26964 984
rect 26586 602 26650 616
rect 27006 608 27034 1114
rect 27110 902 27176 910
rect 27110 850 27116 902
rect 27168 850 27176 902
rect 27110 842 27176 850
rect 26586 550 26589 602
rect 26641 550 26650 602
rect 26586 534 26650 550
rect 26820 592 27034 608
rect 26820 540 26821 592
rect 26873 580 27034 592
rect 26873 540 26874 580
rect 26820 524 26874 540
rect 27126 436 27176 842
rect 27354 598 27382 1716
rect 28634 1714 28702 1724
rect 28514 1541 28578 1548
rect 28514 1510 28520 1541
rect 27786 1489 28520 1510
rect 28572 1489 28578 1541
rect 27786 1482 28578 1489
rect 27786 1480 28520 1482
rect 27786 1474 28514 1480
rect 27686 1144 27750 1152
rect 27686 1092 27692 1144
rect 27744 1092 27750 1144
rect 27686 1084 27750 1092
rect 27446 1056 27512 1062
rect 27446 1004 27454 1056
rect 27506 1026 27512 1056
rect 27686 1026 27714 1084
rect 27506 1004 27714 1026
rect 27446 998 27714 1004
rect 27786 848 27814 1474
rect 28514 1408 28580 1414
rect 28514 1356 28522 1408
rect 28574 1356 28580 1408
rect 28514 1350 28580 1356
rect 28514 1228 28542 1350
rect 28474 1200 28542 1228
rect 27786 840 28098 848
rect 27786 812 28037 840
rect 27446 624 27522 630
rect 27446 598 27454 624
rect 27354 572 27454 598
rect 27506 572 27522 624
rect 27354 570 27522 572
rect 27446 566 27522 570
rect 27126 430 27192 436
rect 27126 378 27134 430
rect 27186 408 27192 430
rect 27786 408 27814 812
rect 28018 788 28037 812
rect 28089 788 28098 840
rect 28018 776 28098 788
rect 28334 844 28402 850
rect 28334 792 28341 844
rect 28393 792 28402 844
rect 28334 786 28402 792
rect 27186 380 27814 408
rect 27186 378 27192 380
rect 27126 372 27192 378
rect 27940 180 28290 194
rect 26052 50 26402 64
rect 27940 64 27961 180
rect 28269 64 28290 180
rect 28334 170 28384 786
rect 28474 616 28502 1200
rect 28536 1150 28598 1156
rect 28536 1098 28546 1150
rect 28634 1142 28662 1714
rect 28690 1541 28754 1548
rect 28690 1489 28696 1541
rect 28748 1508 28754 1541
rect 29016 1508 29066 1898
rect 29538 1896 29566 2000
rect 29538 1890 29604 1896
rect 30652 1894 30680 2000
rect 30888 1958 30954 1966
rect 30888 1906 30894 1958
rect 30946 1906 30954 1958
rect 30888 1898 30954 1906
rect 29538 1876 29546 1890
rect 29540 1838 29546 1876
rect 29598 1838 29604 1890
rect 29540 1832 29604 1838
rect 30612 1888 30680 1894
rect 30612 1836 30622 1888
rect 30674 1836 30680 1888
rect 30612 1830 30680 1836
rect 29452 1774 29516 1780
rect 29452 1744 29458 1774
rect 29242 1722 29458 1744
rect 29510 1722 29516 1774
rect 29242 1716 29516 1722
rect 30522 1776 30590 1782
rect 30522 1724 30530 1776
rect 30582 1724 30590 1776
rect 28748 1492 29068 1508
rect 28748 1489 29082 1492
rect 28690 1486 29082 1489
rect 28690 1480 29024 1486
rect 29016 1434 29024 1480
rect 29076 1434 29082 1486
rect 29016 1428 29082 1434
rect 28886 1292 28958 1304
rect 28886 1240 28896 1292
rect 28948 1240 28958 1292
rect 28886 1228 28958 1240
rect 28922 1226 28958 1228
rect 28634 1114 28922 1142
rect 28536 1092 28598 1098
rect 28570 1046 28598 1092
rect 28570 1042 28814 1046
rect 28570 1036 28852 1042
rect 28570 1018 28792 1036
rect 28786 984 28792 1018
rect 28844 984 28852 1036
rect 28786 976 28852 984
rect 28474 602 28538 616
rect 28894 608 28922 1114
rect 28998 902 29064 910
rect 28998 850 29004 902
rect 29056 850 29064 902
rect 28998 842 29064 850
rect 28474 550 28477 602
rect 28529 550 28538 602
rect 28474 534 28538 550
rect 28708 592 28922 608
rect 28708 540 28709 592
rect 28761 580 28922 592
rect 28761 540 28762 580
rect 28708 524 28762 540
rect 29014 436 29064 842
rect 29242 598 29270 1716
rect 30522 1714 30590 1724
rect 30402 1541 30466 1548
rect 30402 1510 30408 1541
rect 29674 1489 30408 1510
rect 30460 1489 30466 1541
rect 29674 1482 30466 1489
rect 29674 1480 30408 1482
rect 29674 1474 30402 1480
rect 29574 1144 29638 1152
rect 29574 1092 29580 1144
rect 29632 1092 29638 1144
rect 29574 1084 29638 1092
rect 29334 1056 29400 1062
rect 29334 1004 29342 1056
rect 29394 1026 29400 1056
rect 29574 1026 29602 1084
rect 29394 1004 29602 1026
rect 29334 998 29602 1004
rect 29674 848 29702 1474
rect 30402 1408 30468 1414
rect 30402 1356 30410 1408
rect 30462 1356 30468 1408
rect 30402 1350 30468 1356
rect 30402 1228 30430 1350
rect 30362 1200 30430 1228
rect 29674 840 29986 848
rect 29674 812 29925 840
rect 29334 624 29410 630
rect 29334 598 29342 624
rect 29242 572 29342 598
rect 29394 572 29410 624
rect 29242 570 29410 572
rect 29334 566 29410 570
rect 29014 430 29080 436
rect 29014 378 29022 430
rect 29074 408 29080 430
rect 29674 408 29702 812
rect 29906 788 29925 812
rect 29977 788 29986 840
rect 29906 776 29986 788
rect 30222 844 30290 850
rect 30222 792 30229 844
rect 30281 792 30290 844
rect 30222 786 30290 792
rect 29074 380 29702 408
rect 29074 378 29080 380
rect 29014 372 29080 378
rect 29828 180 30178 194
rect 27940 50 28290 64
rect 29828 64 29849 180
rect 30157 64 30178 180
rect 30222 170 30272 786
rect 30362 616 30390 1200
rect 30424 1150 30486 1156
rect 30424 1098 30434 1150
rect 30522 1142 30550 1714
rect 30578 1541 30642 1548
rect 30578 1489 30584 1541
rect 30636 1508 30642 1541
rect 30904 1508 30954 1898
rect 31426 1896 31454 2000
rect 31426 1890 31492 1896
rect 32540 1894 32568 2000
rect 32776 1958 32842 1966
rect 32776 1906 32782 1958
rect 32834 1906 32842 1958
rect 32776 1898 32842 1906
rect 31426 1876 31434 1890
rect 31428 1838 31434 1876
rect 31486 1838 31492 1890
rect 31428 1832 31492 1838
rect 32500 1888 32568 1894
rect 32500 1836 32510 1888
rect 32562 1836 32568 1888
rect 32500 1830 32568 1836
rect 31340 1774 31404 1780
rect 31340 1744 31346 1774
rect 31130 1722 31346 1744
rect 31398 1722 31404 1774
rect 31130 1716 31404 1722
rect 32410 1776 32478 1782
rect 32410 1724 32418 1776
rect 32470 1724 32478 1776
rect 30636 1492 30956 1508
rect 30636 1489 30970 1492
rect 30578 1486 30970 1489
rect 30578 1480 30912 1486
rect 30904 1434 30912 1480
rect 30964 1434 30970 1486
rect 30904 1428 30970 1434
rect 30774 1292 30846 1304
rect 30774 1240 30784 1292
rect 30836 1240 30846 1292
rect 30774 1228 30846 1240
rect 30810 1226 30846 1228
rect 30522 1114 30810 1142
rect 30424 1092 30486 1098
rect 30458 1046 30486 1092
rect 30458 1042 30702 1046
rect 30458 1036 30740 1042
rect 30458 1018 30680 1036
rect 30674 984 30680 1018
rect 30732 984 30740 1036
rect 30674 976 30740 984
rect 30362 602 30426 616
rect 30782 608 30810 1114
rect 30886 902 30952 910
rect 30886 850 30892 902
rect 30944 850 30952 902
rect 30886 842 30952 850
rect 30362 550 30365 602
rect 30417 550 30426 602
rect 30362 534 30426 550
rect 30596 592 30810 608
rect 30596 540 30597 592
rect 30649 580 30810 592
rect 30649 540 30650 580
rect 30596 524 30650 540
rect 30902 436 30952 842
rect 31130 598 31158 1716
rect 32410 1714 32478 1724
rect 32290 1541 32354 1548
rect 32290 1510 32296 1541
rect 31562 1489 32296 1510
rect 32348 1489 32354 1541
rect 31562 1482 32354 1489
rect 31562 1480 32296 1482
rect 31562 1474 32290 1480
rect 31462 1144 31526 1152
rect 31462 1092 31468 1144
rect 31520 1092 31526 1144
rect 31462 1084 31526 1092
rect 31222 1056 31288 1062
rect 31222 1004 31230 1056
rect 31282 1026 31288 1056
rect 31462 1026 31490 1084
rect 31282 1004 31490 1026
rect 31222 998 31490 1004
rect 31562 848 31590 1474
rect 32290 1408 32356 1414
rect 32290 1356 32298 1408
rect 32350 1356 32356 1408
rect 32290 1350 32356 1356
rect 32290 1228 32318 1350
rect 32250 1200 32318 1228
rect 31562 840 31874 848
rect 31562 812 31813 840
rect 31222 624 31298 630
rect 31222 598 31230 624
rect 31130 572 31230 598
rect 31282 572 31298 624
rect 31130 570 31298 572
rect 31222 566 31298 570
rect 30902 430 30968 436
rect 30902 378 30910 430
rect 30962 408 30968 430
rect 31562 408 31590 812
rect 31794 788 31813 812
rect 31865 788 31874 840
rect 31794 776 31874 788
rect 32110 844 32178 850
rect 32110 792 32117 844
rect 32169 792 32178 844
rect 32110 786 32178 792
rect 30962 380 31590 408
rect 30962 378 30968 380
rect 30902 372 30968 378
rect 31716 180 32066 194
rect 29828 50 30178 64
rect 31716 64 31737 180
rect 32045 64 32066 180
rect 32110 170 32160 786
rect 32250 616 32278 1200
rect 32312 1150 32374 1156
rect 32312 1098 32322 1150
rect 32410 1142 32438 1714
rect 32466 1541 32530 1548
rect 32466 1489 32472 1541
rect 32524 1508 32530 1541
rect 32792 1508 32842 1898
rect 33314 1896 33342 2000
rect 33314 1890 33380 1896
rect 34428 1894 34456 2000
rect 34664 1958 34730 1966
rect 34664 1906 34670 1958
rect 34722 1906 34730 1958
rect 34664 1898 34730 1906
rect 33314 1876 33322 1890
rect 33316 1838 33322 1876
rect 33374 1838 33380 1890
rect 33316 1832 33380 1838
rect 34388 1888 34456 1894
rect 34388 1836 34398 1888
rect 34450 1836 34456 1888
rect 34388 1830 34456 1836
rect 33228 1774 33292 1780
rect 33228 1744 33234 1774
rect 33018 1722 33234 1744
rect 33286 1722 33292 1774
rect 33018 1716 33292 1722
rect 34298 1776 34366 1782
rect 34298 1724 34306 1776
rect 34358 1724 34366 1776
rect 32524 1492 32844 1508
rect 32524 1489 32858 1492
rect 32466 1486 32858 1489
rect 32466 1480 32800 1486
rect 32792 1434 32800 1480
rect 32852 1434 32858 1486
rect 32792 1428 32858 1434
rect 32662 1292 32734 1304
rect 32662 1240 32672 1292
rect 32724 1240 32734 1292
rect 32662 1228 32734 1240
rect 32698 1226 32734 1228
rect 32410 1114 32698 1142
rect 32312 1092 32374 1098
rect 32346 1046 32374 1092
rect 32346 1042 32590 1046
rect 32346 1036 32628 1042
rect 32346 1018 32568 1036
rect 32562 984 32568 1018
rect 32620 984 32628 1036
rect 32562 976 32628 984
rect 32250 602 32314 616
rect 32670 608 32698 1114
rect 32774 902 32840 910
rect 32774 850 32780 902
rect 32832 850 32840 902
rect 32774 842 32840 850
rect 32250 550 32253 602
rect 32305 550 32314 602
rect 32250 534 32314 550
rect 32484 592 32698 608
rect 32484 540 32485 592
rect 32537 580 32698 592
rect 32537 540 32538 580
rect 32484 524 32538 540
rect 32790 436 32840 842
rect 33018 598 33046 1716
rect 34298 1714 34366 1724
rect 34178 1541 34242 1548
rect 34178 1510 34184 1541
rect 33450 1489 34184 1510
rect 34236 1489 34242 1541
rect 33450 1482 34242 1489
rect 33450 1480 34184 1482
rect 33450 1474 34178 1480
rect 33350 1144 33414 1152
rect 33350 1092 33356 1144
rect 33408 1092 33414 1144
rect 33350 1084 33414 1092
rect 33110 1056 33176 1062
rect 33110 1004 33118 1056
rect 33170 1026 33176 1056
rect 33350 1026 33378 1084
rect 33170 1004 33378 1026
rect 33110 998 33378 1004
rect 33450 848 33478 1474
rect 34178 1408 34244 1414
rect 34178 1356 34186 1408
rect 34238 1356 34244 1408
rect 34178 1350 34244 1356
rect 34178 1228 34206 1350
rect 34138 1200 34206 1228
rect 33450 840 33762 848
rect 33450 812 33701 840
rect 33110 624 33186 630
rect 33110 598 33118 624
rect 33018 572 33118 598
rect 33170 572 33186 624
rect 33018 570 33186 572
rect 33110 566 33186 570
rect 32790 430 32856 436
rect 32790 378 32798 430
rect 32850 408 32856 430
rect 33450 408 33478 812
rect 33682 788 33701 812
rect 33753 788 33762 840
rect 33682 776 33762 788
rect 33998 844 34066 850
rect 33998 792 34005 844
rect 34057 792 34066 844
rect 33998 786 34066 792
rect 32850 380 33478 408
rect 32850 378 32856 380
rect 32790 372 32856 378
rect 33604 180 33954 194
rect 31716 50 32066 64
rect 33604 64 33625 180
rect 33933 64 33954 180
rect 33998 170 34048 786
rect 34138 616 34166 1200
rect 34200 1150 34262 1156
rect 34200 1098 34210 1150
rect 34298 1142 34326 1714
rect 34354 1541 34418 1548
rect 34354 1489 34360 1541
rect 34412 1508 34418 1541
rect 34680 1508 34730 1898
rect 35202 1896 35230 2000
rect 35904 1996 37224 2000
rect 37788 1996 44962 2000
rect 35202 1890 35268 1896
rect 36316 1894 36344 1996
rect 36552 1958 36618 1966
rect 36552 1906 36558 1958
rect 36610 1906 36618 1958
rect 36552 1898 36618 1906
rect 35202 1876 35210 1890
rect 35204 1838 35210 1876
rect 35262 1838 35268 1890
rect 35204 1832 35268 1838
rect 36276 1888 36344 1894
rect 36276 1836 36286 1888
rect 36338 1836 36344 1888
rect 36276 1830 36344 1836
rect 35116 1774 35180 1780
rect 35116 1744 35122 1774
rect 34906 1722 35122 1744
rect 35174 1722 35180 1774
rect 34906 1716 35180 1722
rect 36186 1776 36254 1782
rect 36186 1724 36194 1776
rect 36246 1724 36254 1776
rect 34412 1492 34732 1508
rect 34412 1489 34746 1492
rect 34354 1486 34746 1489
rect 34354 1480 34688 1486
rect 34680 1434 34688 1480
rect 34740 1434 34746 1486
rect 34680 1428 34746 1434
rect 34550 1292 34622 1304
rect 34550 1240 34560 1292
rect 34612 1240 34622 1292
rect 34550 1228 34622 1240
rect 34586 1226 34622 1228
rect 34298 1114 34586 1142
rect 34200 1092 34262 1098
rect 34234 1046 34262 1092
rect 34234 1042 34478 1046
rect 34234 1036 34516 1042
rect 34234 1018 34456 1036
rect 34450 984 34456 1018
rect 34508 984 34516 1036
rect 34450 976 34516 984
rect 34138 602 34202 616
rect 34558 608 34586 1114
rect 34662 902 34728 910
rect 34662 850 34668 902
rect 34720 850 34728 902
rect 34662 842 34728 850
rect 34138 550 34141 602
rect 34193 550 34202 602
rect 34138 534 34202 550
rect 34372 592 34586 608
rect 34372 540 34373 592
rect 34425 580 34586 592
rect 34425 540 34426 580
rect 34372 524 34426 540
rect 34678 436 34728 842
rect 34906 598 34934 1716
rect 36186 1714 36254 1724
rect 36066 1541 36130 1548
rect 36066 1510 36072 1541
rect 35338 1489 36072 1510
rect 36124 1489 36130 1541
rect 35338 1482 36130 1489
rect 35338 1480 36072 1482
rect 35338 1474 36066 1480
rect 35238 1144 35302 1152
rect 35238 1092 35244 1144
rect 35296 1092 35302 1144
rect 35238 1084 35302 1092
rect 34998 1056 35064 1062
rect 34998 1004 35006 1056
rect 35058 1026 35064 1056
rect 35238 1026 35266 1084
rect 35058 1004 35266 1026
rect 34998 998 35266 1004
rect 35338 848 35366 1474
rect 36066 1408 36132 1414
rect 36066 1356 36074 1408
rect 36126 1356 36132 1408
rect 36066 1350 36132 1356
rect 36066 1228 36094 1350
rect 36026 1200 36094 1228
rect 35338 840 35650 848
rect 35338 812 35589 840
rect 34998 624 35074 630
rect 34998 598 35006 624
rect 34906 572 35006 598
rect 35058 572 35074 624
rect 34906 570 35074 572
rect 34998 566 35074 570
rect 34678 430 34744 436
rect 34678 378 34686 430
rect 34738 408 34744 430
rect 35338 408 35366 812
rect 35570 788 35589 812
rect 35641 788 35650 840
rect 35570 776 35650 788
rect 35886 844 35954 850
rect 35886 792 35893 844
rect 35945 792 35954 844
rect 35886 786 35954 792
rect 34738 380 35366 408
rect 34738 378 34744 380
rect 34678 372 34744 378
rect 35492 180 35842 194
rect 33604 50 33954 64
rect 35492 64 35513 180
rect 35821 64 35842 180
rect 35886 170 35936 786
rect 36026 616 36054 1200
rect 36088 1150 36150 1156
rect 36088 1098 36098 1150
rect 36186 1142 36214 1714
rect 36242 1541 36306 1548
rect 36242 1489 36248 1541
rect 36300 1508 36306 1541
rect 36568 1508 36618 1898
rect 37090 1896 37118 1996
rect 37090 1890 37156 1896
rect 38204 1894 38232 1996
rect 38440 1958 38506 1966
rect 38440 1906 38446 1958
rect 38498 1906 38506 1958
rect 38440 1898 38506 1906
rect 37090 1876 37098 1890
rect 37092 1838 37098 1876
rect 37150 1838 37156 1890
rect 37092 1832 37156 1838
rect 38164 1888 38232 1894
rect 38164 1836 38174 1888
rect 38226 1836 38232 1888
rect 38164 1830 38232 1836
rect 37004 1774 37068 1780
rect 37004 1744 37010 1774
rect 36794 1722 37010 1744
rect 37062 1722 37068 1774
rect 36794 1716 37068 1722
rect 38074 1776 38142 1782
rect 38074 1724 38082 1776
rect 38134 1724 38142 1776
rect 36300 1492 36620 1508
rect 36300 1489 36634 1492
rect 36242 1486 36634 1489
rect 36242 1480 36576 1486
rect 36568 1434 36576 1480
rect 36628 1434 36634 1486
rect 36568 1428 36634 1434
rect 36438 1292 36510 1304
rect 36438 1240 36448 1292
rect 36500 1240 36510 1292
rect 36438 1228 36510 1240
rect 36474 1226 36510 1228
rect 36186 1114 36474 1142
rect 36088 1092 36150 1098
rect 36122 1046 36150 1092
rect 36122 1042 36366 1046
rect 36122 1036 36404 1042
rect 36122 1018 36344 1036
rect 36338 984 36344 1018
rect 36396 984 36404 1036
rect 36338 976 36404 984
rect 36026 602 36090 616
rect 36446 608 36474 1114
rect 36550 902 36616 910
rect 36550 850 36556 902
rect 36608 850 36616 902
rect 36550 842 36616 850
rect 36026 550 36029 602
rect 36081 550 36090 602
rect 36026 534 36090 550
rect 36260 592 36474 608
rect 36260 540 36261 592
rect 36313 580 36474 592
rect 36313 540 36314 580
rect 36260 524 36314 540
rect 36566 436 36616 842
rect 36794 598 36822 1716
rect 38074 1714 38142 1724
rect 37954 1541 38018 1548
rect 37954 1510 37960 1541
rect 37226 1489 37960 1510
rect 38012 1489 38018 1541
rect 37226 1482 38018 1489
rect 37226 1480 37960 1482
rect 37226 1474 37954 1480
rect 37126 1144 37190 1152
rect 37126 1092 37132 1144
rect 37184 1092 37190 1144
rect 37126 1084 37190 1092
rect 36886 1056 36952 1062
rect 36886 1004 36894 1056
rect 36946 1026 36952 1056
rect 37126 1026 37154 1084
rect 36946 1004 37154 1026
rect 36886 998 37154 1004
rect 37226 848 37254 1474
rect 37954 1408 38020 1414
rect 37954 1356 37962 1408
rect 38014 1356 38020 1408
rect 37954 1350 38020 1356
rect 37954 1228 37982 1350
rect 37914 1200 37982 1228
rect 37226 840 37538 848
rect 37226 812 37477 840
rect 36886 624 36962 630
rect 36886 598 36894 624
rect 36794 572 36894 598
rect 36946 572 36962 624
rect 36794 570 36962 572
rect 36886 566 36962 570
rect 36566 430 36632 436
rect 36566 378 36574 430
rect 36626 408 36632 430
rect 37226 408 37254 812
rect 37458 788 37477 812
rect 37529 788 37538 840
rect 37458 776 37538 788
rect 37774 844 37842 850
rect 37774 792 37781 844
rect 37833 792 37842 844
rect 37774 786 37842 792
rect 36626 380 37254 408
rect 36626 378 36632 380
rect 36566 372 36632 378
rect 37380 180 37730 194
rect 35492 50 35842 64
rect 37380 64 37401 180
rect 37709 64 37730 180
rect 37774 170 37824 786
rect 37914 616 37942 1200
rect 37976 1150 38038 1156
rect 37976 1098 37986 1150
rect 38074 1142 38102 1714
rect 38130 1541 38194 1548
rect 38130 1489 38136 1541
rect 38188 1508 38194 1541
rect 38456 1508 38506 1898
rect 38978 1896 39006 1996
rect 38978 1890 39044 1896
rect 40092 1894 40120 1996
rect 40328 1958 40394 1966
rect 40328 1906 40334 1958
rect 40386 1906 40394 1958
rect 40328 1898 40394 1906
rect 38978 1876 38986 1890
rect 38980 1838 38986 1876
rect 39038 1838 39044 1890
rect 38980 1832 39044 1838
rect 40052 1888 40120 1894
rect 40052 1836 40062 1888
rect 40114 1836 40120 1888
rect 40052 1830 40120 1836
rect 38892 1774 38956 1780
rect 38892 1744 38898 1774
rect 38682 1722 38898 1744
rect 38950 1722 38956 1774
rect 38682 1716 38956 1722
rect 39962 1776 40030 1782
rect 39962 1724 39970 1776
rect 40022 1724 40030 1776
rect 38188 1492 38508 1508
rect 38188 1489 38522 1492
rect 38130 1486 38522 1489
rect 38130 1480 38464 1486
rect 38456 1434 38464 1480
rect 38516 1434 38522 1486
rect 38456 1428 38522 1434
rect 38326 1292 38398 1304
rect 38326 1240 38336 1292
rect 38388 1240 38398 1292
rect 38326 1228 38398 1240
rect 38362 1226 38398 1228
rect 38074 1114 38362 1142
rect 37976 1092 38038 1098
rect 38010 1046 38038 1092
rect 38010 1042 38254 1046
rect 38010 1036 38292 1042
rect 38010 1018 38232 1036
rect 38226 984 38232 1018
rect 38284 984 38292 1036
rect 38226 976 38292 984
rect 37914 602 37978 616
rect 38334 608 38362 1114
rect 38438 902 38504 910
rect 38438 850 38444 902
rect 38496 850 38504 902
rect 38438 842 38504 850
rect 37914 550 37917 602
rect 37969 550 37978 602
rect 37914 534 37978 550
rect 38148 592 38362 608
rect 38148 540 38149 592
rect 38201 580 38362 592
rect 38201 540 38202 580
rect 38148 524 38202 540
rect 38454 436 38504 842
rect 38682 598 38710 1716
rect 39962 1714 40030 1724
rect 39842 1541 39906 1548
rect 39842 1510 39848 1541
rect 39114 1489 39848 1510
rect 39900 1489 39906 1541
rect 39114 1482 39906 1489
rect 39114 1480 39848 1482
rect 39114 1474 39842 1480
rect 39014 1144 39078 1152
rect 39014 1092 39020 1144
rect 39072 1092 39078 1144
rect 39014 1084 39078 1092
rect 38774 1056 38840 1062
rect 38774 1004 38782 1056
rect 38834 1026 38840 1056
rect 39014 1026 39042 1084
rect 38834 1004 39042 1026
rect 38774 998 39042 1004
rect 39114 848 39142 1474
rect 39842 1408 39908 1414
rect 39842 1356 39850 1408
rect 39902 1356 39908 1408
rect 39842 1350 39908 1356
rect 39842 1228 39870 1350
rect 39802 1200 39870 1228
rect 39114 840 39426 848
rect 39114 812 39365 840
rect 38774 624 38850 630
rect 38774 598 38782 624
rect 38682 572 38782 598
rect 38834 572 38850 624
rect 38682 570 38850 572
rect 38774 566 38850 570
rect 38454 430 38520 436
rect 38454 378 38462 430
rect 38514 408 38520 430
rect 39114 408 39142 812
rect 39346 788 39365 812
rect 39417 788 39426 840
rect 39346 776 39426 788
rect 39662 844 39730 850
rect 39662 792 39669 844
rect 39721 792 39730 844
rect 39662 786 39730 792
rect 38514 380 39142 408
rect 38514 378 38520 380
rect 38454 372 38520 378
rect 39268 180 39618 194
rect 37380 50 37730 64
rect 39268 64 39289 180
rect 39597 64 39618 180
rect 39662 170 39712 786
rect 39802 616 39830 1200
rect 39864 1150 39926 1156
rect 39864 1098 39874 1150
rect 39962 1142 39990 1714
rect 40018 1541 40082 1548
rect 40018 1489 40024 1541
rect 40076 1508 40082 1541
rect 40344 1508 40394 1898
rect 40866 1896 40894 1996
rect 40866 1890 40932 1896
rect 41980 1894 42008 1996
rect 42216 1958 42282 1966
rect 42216 1906 42222 1958
rect 42274 1906 42282 1958
rect 42216 1898 42282 1906
rect 40866 1876 40874 1890
rect 40868 1838 40874 1876
rect 40926 1838 40932 1890
rect 40868 1832 40932 1838
rect 41940 1888 42008 1894
rect 41940 1836 41950 1888
rect 42002 1836 42008 1888
rect 41940 1830 42008 1836
rect 40780 1774 40844 1780
rect 40780 1744 40786 1774
rect 40570 1722 40786 1744
rect 40838 1722 40844 1774
rect 40570 1716 40844 1722
rect 41850 1776 41918 1782
rect 41850 1724 41858 1776
rect 41910 1724 41918 1776
rect 40076 1492 40396 1508
rect 40076 1489 40410 1492
rect 40018 1486 40410 1489
rect 40018 1480 40352 1486
rect 40344 1434 40352 1480
rect 40404 1434 40410 1486
rect 40344 1428 40410 1434
rect 40214 1292 40286 1304
rect 40214 1240 40224 1292
rect 40276 1240 40286 1292
rect 40214 1228 40286 1240
rect 40250 1226 40286 1228
rect 39962 1114 40250 1142
rect 39864 1092 39926 1098
rect 39898 1046 39926 1092
rect 39898 1042 40142 1046
rect 39898 1036 40180 1042
rect 39898 1018 40120 1036
rect 40114 984 40120 1018
rect 40172 984 40180 1036
rect 40114 976 40180 984
rect 39802 602 39866 616
rect 40222 608 40250 1114
rect 40326 902 40392 910
rect 40326 850 40332 902
rect 40384 850 40392 902
rect 40326 842 40392 850
rect 39802 550 39805 602
rect 39857 550 39866 602
rect 39802 534 39866 550
rect 40036 592 40250 608
rect 40036 540 40037 592
rect 40089 580 40250 592
rect 40089 540 40090 580
rect 40036 524 40090 540
rect 40342 436 40392 842
rect 40570 598 40598 1716
rect 41850 1714 41918 1724
rect 41730 1541 41794 1548
rect 41730 1510 41736 1541
rect 41002 1489 41736 1510
rect 41788 1489 41794 1541
rect 41002 1482 41794 1489
rect 41002 1480 41736 1482
rect 41002 1474 41730 1480
rect 40902 1144 40966 1152
rect 40902 1092 40908 1144
rect 40960 1092 40966 1144
rect 40902 1084 40966 1092
rect 40662 1056 40728 1062
rect 40662 1004 40670 1056
rect 40722 1026 40728 1056
rect 40902 1026 40930 1084
rect 40722 1004 40930 1026
rect 40662 998 40930 1004
rect 41002 848 41030 1474
rect 41730 1408 41796 1414
rect 41730 1356 41738 1408
rect 41790 1356 41796 1408
rect 41730 1350 41796 1356
rect 41730 1228 41758 1350
rect 41690 1200 41758 1228
rect 41002 840 41314 848
rect 41002 812 41253 840
rect 40662 624 40738 630
rect 40662 598 40670 624
rect 40570 572 40670 598
rect 40722 572 40738 624
rect 40570 570 40738 572
rect 40662 566 40738 570
rect 40342 430 40408 436
rect 40342 378 40350 430
rect 40402 408 40408 430
rect 41002 408 41030 812
rect 41234 788 41253 812
rect 41305 788 41314 840
rect 41234 776 41314 788
rect 41550 844 41618 850
rect 41550 792 41557 844
rect 41609 792 41618 844
rect 41550 786 41618 792
rect 40402 380 41030 408
rect 40402 378 40408 380
rect 40342 372 40408 378
rect 41156 180 41506 194
rect 39268 50 39618 64
rect 41156 64 41177 180
rect 41485 64 41506 180
rect 41550 170 41600 786
rect 41690 616 41718 1200
rect 41752 1150 41814 1156
rect 41752 1098 41762 1150
rect 41850 1142 41878 1714
rect 41906 1541 41970 1548
rect 41906 1489 41912 1541
rect 41964 1508 41970 1541
rect 42232 1508 42282 1898
rect 42754 1896 42782 1996
rect 42754 1890 42820 1896
rect 43868 1894 43896 1996
rect 44104 1958 44170 1966
rect 44104 1906 44110 1958
rect 44162 1906 44170 1958
rect 44104 1898 44170 1906
rect 42754 1876 42762 1890
rect 42756 1838 42762 1876
rect 42814 1838 42820 1890
rect 42756 1832 42820 1838
rect 43828 1888 43896 1894
rect 43828 1836 43838 1888
rect 43890 1836 43896 1888
rect 43828 1830 43896 1836
rect 42668 1774 42732 1780
rect 42668 1744 42674 1774
rect 42458 1722 42674 1744
rect 42726 1722 42732 1774
rect 42458 1716 42732 1722
rect 43738 1776 43806 1782
rect 43738 1724 43746 1776
rect 43798 1724 43806 1776
rect 41964 1492 42284 1508
rect 41964 1489 42298 1492
rect 41906 1486 42298 1489
rect 41906 1480 42240 1486
rect 42232 1434 42240 1480
rect 42292 1434 42298 1486
rect 42232 1428 42298 1434
rect 42102 1292 42174 1304
rect 42102 1240 42112 1292
rect 42164 1240 42174 1292
rect 42102 1228 42174 1240
rect 42138 1226 42174 1228
rect 41850 1114 42138 1142
rect 41752 1092 41814 1098
rect 41786 1046 41814 1092
rect 41786 1042 42030 1046
rect 41786 1036 42068 1042
rect 41786 1018 42008 1036
rect 42002 984 42008 1018
rect 42060 984 42068 1036
rect 42002 976 42068 984
rect 41690 602 41754 616
rect 42110 608 42138 1114
rect 42214 902 42280 910
rect 42214 850 42220 902
rect 42272 850 42280 902
rect 42214 842 42280 850
rect 41690 550 41693 602
rect 41745 550 41754 602
rect 41690 534 41754 550
rect 41924 592 42138 608
rect 41924 540 41925 592
rect 41977 580 42138 592
rect 41977 540 41978 580
rect 41924 524 41978 540
rect 42230 436 42280 842
rect 42458 598 42486 1716
rect 43738 1714 43806 1724
rect 43618 1541 43682 1548
rect 43618 1510 43624 1541
rect 42890 1489 43624 1510
rect 43676 1489 43682 1541
rect 42890 1482 43682 1489
rect 42890 1480 43624 1482
rect 42890 1474 43618 1480
rect 42790 1144 42854 1152
rect 42790 1092 42796 1144
rect 42848 1092 42854 1144
rect 42790 1084 42854 1092
rect 42550 1056 42616 1062
rect 42550 1004 42558 1056
rect 42610 1026 42616 1056
rect 42790 1026 42818 1084
rect 42610 1004 42818 1026
rect 42550 998 42818 1004
rect 42890 848 42918 1474
rect 43618 1408 43684 1414
rect 43618 1356 43626 1408
rect 43678 1356 43684 1408
rect 43618 1350 43684 1356
rect 43618 1228 43646 1350
rect 43578 1200 43646 1228
rect 42890 840 43202 848
rect 42890 812 43141 840
rect 42550 624 42626 630
rect 42550 598 42558 624
rect 42458 572 42558 598
rect 42610 572 42626 624
rect 42458 570 42626 572
rect 42550 566 42626 570
rect 42230 430 42296 436
rect 42230 378 42238 430
rect 42290 408 42296 430
rect 42890 408 42918 812
rect 43122 788 43141 812
rect 43193 788 43202 840
rect 43122 776 43202 788
rect 43438 844 43506 850
rect 43438 792 43445 844
rect 43497 792 43506 844
rect 43438 786 43506 792
rect 42290 380 42918 408
rect 42290 378 42296 380
rect 42230 372 42296 378
rect 43044 180 43394 194
rect 41156 50 41506 64
rect 43044 64 43065 180
rect 43373 64 43394 180
rect 43438 170 43488 786
rect 43578 616 43606 1200
rect 43640 1150 43702 1156
rect 43640 1098 43650 1150
rect 43738 1142 43766 1714
rect 43794 1541 43858 1548
rect 43794 1489 43800 1541
rect 43852 1508 43858 1541
rect 44120 1508 44170 1898
rect 44642 1896 44670 1996
rect 44642 1890 44708 1896
rect 45750 1894 45778 2000
rect 45986 1958 46052 1966
rect 45986 1906 45992 1958
rect 46044 1906 46052 1958
rect 45986 1898 46052 1906
rect 44642 1876 44650 1890
rect 44644 1838 44650 1876
rect 44702 1838 44708 1890
rect 44644 1832 44708 1838
rect 45710 1888 45778 1894
rect 45710 1836 45720 1888
rect 45772 1836 45778 1888
rect 45710 1830 45778 1836
rect 44556 1774 44620 1780
rect 44556 1744 44562 1774
rect 44346 1722 44562 1744
rect 44614 1722 44620 1774
rect 44346 1716 44620 1722
rect 45620 1776 45688 1782
rect 45620 1724 45628 1776
rect 45680 1724 45688 1776
rect 43852 1492 44172 1508
rect 43852 1489 44186 1492
rect 43794 1486 44186 1489
rect 43794 1480 44128 1486
rect 44120 1434 44128 1480
rect 44180 1434 44186 1486
rect 44120 1428 44186 1434
rect 43990 1292 44062 1304
rect 43990 1240 44000 1292
rect 44052 1240 44062 1292
rect 43990 1228 44062 1240
rect 44026 1226 44062 1228
rect 43738 1114 44026 1142
rect 43640 1092 43702 1098
rect 43674 1046 43702 1092
rect 43674 1042 43918 1046
rect 43674 1036 43956 1042
rect 43674 1018 43896 1036
rect 43890 984 43896 1018
rect 43948 984 43956 1036
rect 43890 976 43956 984
rect 43578 602 43642 616
rect 43998 608 44026 1114
rect 44102 902 44168 910
rect 44102 850 44108 902
rect 44160 850 44168 902
rect 44102 842 44168 850
rect 43578 550 43581 602
rect 43633 550 43642 602
rect 43578 534 43642 550
rect 43812 592 44026 608
rect 43812 540 43813 592
rect 43865 580 44026 592
rect 43865 540 43866 580
rect 43812 524 43866 540
rect 44118 436 44168 842
rect 44346 598 44374 1716
rect 45620 1714 45688 1724
rect 45500 1541 45564 1548
rect 45500 1510 45506 1541
rect 44778 1489 45506 1510
rect 45558 1489 45564 1541
rect 44778 1482 45564 1489
rect 44778 1480 45506 1482
rect 44778 1474 45500 1480
rect 44678 1144 44742 1152
rect 44678 1092 44684 1144
rect 44736 1092 44742 1144
rect 44678 1084 44742 1092
rect 44438 1056 44504 1062
rect 44438 1004 44446 1056
rect 44498 1026 44504 1056
rect 44678 1026 44706 1084
rect 44498 1004 44706 1026
rect 44438 998 44706 1004
rect 44778 848 44806 1474
rect 45500 1408 45566 1414
rect 45500 1356 45508 1408
rect 45560 1356 45566 1408
rect 45500 1350 45566 1356
rect 45500 1228 45528 1350
rect 45460 1200 45528 1228
rect 44778 840 45090 848
rect 44778 812 45029 840
rect 44438 624 44514 630
rect 44438 598 44446 624
rect 44346 572 44446 598
rect 44498 572 44514 624
rect 44346 570 44514 572
rect 44438 566 44514 570
rect 44118 430 44184 436
rect 44118 378 44126 430
rect 44178 408 44184 430
rect 44778 408 44806 812
rect 45010 788 45029 812
rect 45081 788 45090 840
rect 45010 776 45090 788
rect 45320 844 45388 850
rect 45320 792 45327 844
rect 45379 792 45388 844
rect 45320 786 45388 792
rect 44178 380 44806 408
rect 44178 378 44184 380
rect 44118 372 44184 378
rect 44932 180 45282 194
rect 43044 50 43394 64
rect 44932 64 44953 180
rect 45261 64 45282 180
rect 45320 170 45376 786
rect 45460 616 45488 1200
rect 45522 1150 45584 1156
rect 45522 1098 45532 1150
rect 45620 1142 45648 1714
rect 45676 1541 45740 1548
rect 45676 1489 45682 1541
rect 45734 1508 45740 1541
rect 46002 1508 46052 1898
rect 46524 1896 46552 2000
rect 46524 1890 46590 1896
rect 47638 1894 47666 2000
rect 47874 1958 47940 1966
rect 47874 1906 47880 1958
rect 47932 1906 47940 1958
rect 47874 1898 47940 1906
rect 46524 1876 46532 1890
rect 46526 1838 46532 1876
rect 46584 1838 46590 1890
rect 46526 1832 46590 1838
rect 47598 1888 47666 1894
rect 47598 1836 47608 1888
rect 47660 1836 47666 1888
rect 47598 1830 47666 1836
rect 46438 1774 46502 1780
rect 46438 1744 46444 1774
rect 46228 1722 46444 1744
rect 46496 1722 46502 1774
rect 46228 1716 46502 1722
rect 47508 1776 47576 1782
rect 47508 1724 47516 1776
rect 47568 1724 47576 1776
rect 45734 1492 46054 1508
rect 45734 1489 46068 1492
rect 45676 1486 46068 1489
rect 45676 1480 46010 1486
rect 46002 1434 46010 1480
rect 46062 1434 46068 1486
rect 46002 1428 46068 1434
rect 45872 1292 45944 1304
rect 45872 1240 45882 1292
rect 45934 1240 45944 1292
rect 45872 1228 45944 1240
rect 45908 1226 45944 1228
rect 45620 1114 45908 1142
rect 45522 1092 45584 1098
rect 45556 1046 45584 1092
rect 45556 1042 45800 1046
rect 45556 1036 45838 1042
rect 45556 1018 45778 1036
rect 45772 984 45778 1018
rect 45830 984 45838 1036
rect 45772 976 45838 984
rect 45460 602 45524 616
rect 45880 608 45908 1114
rect 45984 902 46050 910
rect 45984 850 45990 902
rect 46042 850 46050 902
rect 45984 842 46050 850
rect 45460 550 45463 602
rect 45515 550 45524 602
rect 45460 534 45524 550
rect 45694 592 45908 608
rect 45694 540 45695 592
rect 45747 580 45908 592
rect 45747 540 45748 580
rect 45694 524 45748 540
rect 46000 436 46050 842
rect 46228 598 46256 1716
rect 47508 1714 47576 1724
rect 47388 1541 47452 1548
rect 47388 1510 47394 1541
rect 46660 1489 47394 1510
rect 47446 1489 47452 1541
rect 46660 1482 47452 1489
rect 46660 1480 47394 1482
rect 46660 1474 47388 1480
rect 46560 1144 46624 1152
rect 46560 1092 46566 1144
rect 46618 1092 46624 1144
rect 46560 1084 46624 1092
rect 46320 1056 46386 1062
rect 46320 1004 46328 1056
rect 46380 1026 46386 1056
rect 46560 1026 46588 1084
rect 46380 1004 46588 1026
rect 46320 998 46588 1004
rect 46660 848 46688 1474
rect 47388 1408 47454 1414
rect 47388 1356 47396 1408
rect 47448 1356 47454 1408
rect 47388 1350 47454 1356
rect 47388 1228 47416 1350
rect 47348 1200 47416 1228
rect 46660 840 46972 848
rect 46660 812 46911 840
rect 46320 624 46396 630
rect 46320 598 46328 624
rect 46228 572 46328 598
rect 46380 572 46396 624
rect 46228 570 46396 572
rect 46320 566 46396 570
rect 46000 430 46066 436
rect 46000 378 46008 430
rect 46060 408 46066 430
rect 46660 408 46688 812
rect 46892 788 46911 812
rect 46963 788 46972 840
rect 46892 776 46972 788
rect 47208 844 47276 850
rect 47208 792 47215 844
rect 47267 792 47276 844
rect 47208 786 47276 792
rect 46060 380 46688 408
rect 46060 378 46066 380
rect 46000 372 46066 378
rect 46814 180 47164 194
rect 44932 50 45282 64
rect 46814 64 46835 180
rect 47143 64 47164 180
rect 47208 170 47264 786
rect 47348 616 47376 1200
rect 47410 1150 47472 1156
rect 47410 1098 47420 1150
rect 47508 1142 47536 1714
rect 47564 1541 47628 1548
rect 47564 1489 47570 1541
rect 47622 1508 47628 1541
rect 47890 1508 47940 1898
rect 48412 1896 48440 2000
rect 48412 1890 48478 1896
rect 49526 1894 49554 2000
rect 49762 1958 49828 1966
rect 49762 1906 49768 1958
rect 49820 1906 49828 1958
rect 49762 1898 49828 1906
rect 48412 1876 48420 1890
rect 48414 1838 48420 1876
rect 48472 1838 48478 1890
rect 48414 1832 48478 1838
rect 49486 1888 49554 1894
rect 49486 1836 49496 1888
rect 49548 1836 49554 1888
rect 49486 1830 49554 1836
rect 48326 1774 48390 1780
rect 48326 1744 48332 1774
rect 48116 1722 48332 1744
rect 48384 1722 48390 1774
rect 48116 1716 48390 1722
rect 49396 1776 49464 1782
rect 49396 1724 49404 1776
rect 49456 1724 49464 1776
rect 47622 1492 47942 1508
rect 47622 1489 47956 1492
rect 47564 1486 47956 1489
rect 47564 1480 47898 1486
rect 47890 1434 47898 1480
rect 47950 1434 47956 1486
rect 47890 1428 47956 1434
rect 47760 1292 47832 1304
rect 47760 1240 47770 1292
rect 47822 1240 47832 1292
rect 47760 1228 47832 1240
rect 47796 1226 47832 1228
rect 47508 1114 47796 1142
rect 47410 1092 47472 1098
rect 47444 1046 47472 1092
rect 47444 1042 47688 1046
rect 47444 1036 47726 1042
rect 47444 1018 47666 1036
rect 47660 984 47666 1018
rect 47718 984 47726 1036
rect 47660 976 47726 984
rect 47348 602 47412 616
rect 47768 608 47796 1114
rect 47872 902 47938 910
rect 47872 850 47878 902
rect 47930 850 47938 902
rect 47872 842 47938 850
rect 47348 550 47351 602
rect 47403 550 47412 602
rect 47348 534 47412 550
rect 47582 592 47796 608
rect 47582 540 47583 592
rect 47635 580 47796 592
rect 47635 540 47636 580
rect 47582 524 47636 540
rect 47888 436 47938 842
rect 48116 598 48144 1716
rect 49396 1714 49464 1724
rect 49276 1541 49340 1548
rect 49276 1510 49282 1541
rect 48548 1489 49282 1510
rect 49334 1489 49340 1541
rect 48548 1482 49340 1489
rect 48548 1480 49282 1482
rect 48548 1474 49276 1480
rect 48448 1144 48512 1152
rect 48448 1092 48454 1144
rect 48506 1092 48512 1144
rect 48448 1084 48512 1092
rect 48208 1056 48274 1062
rect 48208 1004 48216 1056
rect 48268 1026 48274 1056
rect 48448 1026 48476 1084
rect 48268 1004 48476 1026
rect 48208 998 48476 1004
rect 48548 848 48576 1474
rect 49276 1408 49342 1414
rect 49276 1356 49284 1408
rect 49336 1356 49342 1408
rect 49276 1350 49342 1356
rect 49276 1228 49304 1350
rect 49236 1200 49304 1228
rect 48548 840 48860 848
rect 48548 812 48799 840
rect 48208 624 48284 630
rect 48208 598 48216 624
rect 48116 572 48216 598
rect 48268 572 48284 624
rect 48116 570 48284 572
rect 48208 566 48284 570
rect 47888 430 47954 436
rect 47888 378 47896 430
rect 47948 408 47954 430
rect 48548 408 48576 812
rect 48780 788 48799 812
rect 48851 788 48860 840
rect 48780 776 48860 788
rect 49096 844 49164 850
rect 49096 792 49103 844
rect 49155 792 49164 844
rect 49096 786 49164 792
rect 47948 380 48576 408
rect 47948 378 47954 380
rect 47888 372 47954 378
rect 48702 180 49052 194
rect 46814 50 47164 64
rect 48702 64 48723 180
rect 49031 64 49052 180
rect 49096 170 49152 786
rect 49236 616 49264 1200
rect 49298 1150 49360 1156
rect 49298 1098 49308 1150
rect 49396 1142 49424 1714
rect 49452 1541 49516 1548
rect 49452 1489 49458 1541
rect 49510 1508 49516 1541
rect 49778 1508 49828 1898
rect 50300 1896 50328 2000
rect 51002 1996 52322 2000
rect 52886 1996 54210 2000
rect 50300 1890 50366 1896
rect 51414 1894 51442 1996
rect 51650 1958 51716 1966
rect 51650 1906 51656 1958
rect 51708 1906 51716 1958
rect 51650 1898 51716 1906
rect 50300 1876 50308 1890
rect 50302 1838 50308 1876
rect 50360 1838 50366 1890
rect 50302 1832 50366 1838
rect 51374 1888 51442 1894
rect 51374 1836 51384 1888
rect 51436 1836 51442 1888
rect 51374 1830 51442 1836
rect 50214 1774 50278 1780
rect 50214 1744 50220 1774
rect 50004 1722 50220 1744
rect 50272 1722 50278 1774
rect 50004 1716 50278 1722
rect 51284 1776 51352 1782
rect 51284 1724 51292 1776
rect 51344 1724 51352 1776
rect 49510 1492 49830 1508
rect 49510 1489 49844 1492
rect 49452 1486 49844 1489
rect 49452 1480 49786 1486
rect 49778 1434 49786 1480
rect 49838 1434 49844 1486
rect 49778 1428 49844 1434
rect 49648 1292 49720 1304
rect 49648 1240 49658 1292
rect 49710 1240 49720 1292
rect 49648 1228 49720 1240
rect 49684 1226 49720 1228
rect 49396 1114 49684 1142
rect 49298 1092 49360 1098
rect 49332 1046 49360 1092
rect 49332 1042 49576 1046
rect 49332 1036 49614 1042
rect 49332 1018 49554 1036
rect 49548 984 49554 1018
rect 49606 984 49614 1036
rect 49548 976 49614 984
rect 49236 602 49300 616
rect 49656 608 49684 1114
rect 49760 902 49826 910
rect 49760 850 49766 902
rect 49818 850 49826 902
rect 49760 842 49826 850
rect 49236 550 49239 602
rect 49291 550 49300 602
rect 49236 534 49300 550
rect 49470 592 49684 608
rect 49470 540 49471 592
rect 49523 580 49684 592
rect 49523 540 49524 580
rect 49470 524 49524 540
rect 49776 436 49826 842
rect 50004 598 50032 1716
rect 51284 1714 51352 1724
rect 51164 1541 51228 1548
rect 51164 1510 51170 1541
rect 50436 1489 51170 1510
rect 51222 1489 51228 1541
rect 50436 1482 51228 1489
rect 50436 1480 51170 1482
rect 50436 1474 51164 1480
rect 50336 1144 50400 1152
rect 50336 1092 50342 1144
rect 50394 1092 50400 1144
rect 50336 1084 50400 1092
rect 50096 1056 50162 1062
rect 50096 1004 50104 1056
rect 50156 1026 50162 1056
rect 50336 1026 50364 1084
rect 50156 1004 50364 1026
rect 50096 998 50364 1004
rect 50436 848 50464 1474
rect 51164 1408 51230 1414
rect 51164 1356 51172 1408
rect 51224 1356 51230 1408
rect 51164 1350 51230 1356
rect 51164 1228 51192 1350
rect 51124 1200 51192 1228
rect 50436 840 50748 848
rect 50436 812 50687 840
rect 50096 624 50172 630
rect 50096 598 50104 624
rect 50004 572 50104 598
rect 50156 572 50172 624
rect 50004 570 50172 572
rect 50096 566 50172 570
rect 49776 430 49842 436
rect 49776 378 49784 430
rect 49836 408 49842 430
rect 50436 408 50464 812
rect 50668 788 50687 812
rect 50739 788 50748 840
rect 50668 776 50748 788
rect 50984 844 51052 850
rect 50984 792 50991 844
rect 51043 792 51052 844
rect 50984 786 51052 792
rect 49836 380 50464 408
rect 49836 378 49842 380
rect 49776 372 49842 378
rect 50590 180 50940 194
rect 48702 50 49052 64
rect 50590 64 50611 180
rect 50919 64 50940 180
rect 50984 170 51040 786
rect 51124 616 51152 1200
rect 51186 1150 51248 1156
rect 51186 1098 51196 1150
rect 51284 1142 51312 1714
rect 51340 1541 51404 1548
rect 51340 1489 51346 1541
rect 51398 1508 51404 1541
rect 51666 1508 51716 1898
rect 52188 1896 52216 1996
rect 52188 1890 52254 1896
rect 53302 1894 53330 1996
rect 53538 1958 53604 1966
rect 53538 1906 53544 1958
rect 53596 1906 53604 1958
rect 53538 1898 53604 1906
rect 52188 1876 52196 1890
rect 52190 1838 52196 1876
rect 52248 1838 52254 1890
rect 52190 1832 52254 1838
rect 53262 1888 53330 1894
rect 53262 1836 53272 1888
rect 53324 1836 53330 1888
rect 53262 1830 53330 1836
rect 52102 1774 52166 1780
rect 52102 1744 52108 1774
rect 51892 1722 52108 1744
rect 52160 1722 52166 1774
rect 51892 1716 52166 1722
rect 53172 1776 53240 1782
rect 53172 1724 53180 1776
rect 53232 1724 53240 1776
rect 51398 1492 51718 1508
rect 51398 1489 51732 1492
rect 51340 1486 51732 1489
rect 51340 1480 51674 1486
rect 51666 1434 51674 1480
rect 51726 1434 51732 1486
rect 51666 1428 51732 1434
rect 51536 1292 51608 1304
rect 51536 1240 51546 1292
rect 51598 1240 51608 1292
rect 51536 1228 51608 1240
rect 51572 1226 51608 1228
rect 51284 1114 51572 1142
rect 51186 1092 51248 1098
rect 51220 1046 51248 1092
rect 51220 1042 51464 1046
rect 51220 1036 51502 1042
rect 51220 1018 51442 1036
rect 51436 984 51442 1018
rect 51494 984 51502 1036
rect 51436 976 51502 984
rect 51124 602 51188 616
rect 51544 608 51572 1114
rect 51648 902 51714 910
rect 51648 850 51654 902
rect 51706 850 51714 902
rect 51648 842 51714 850
rect 51124 550 51127 602
rect 51179 550 51188 602
rect 51124 534 51188 550
rect 51358 592 51572 608
rect 51358 540 51359 592
rect 51411 580 51572 592
rect 51411 540 51412 580
rect 51358 524 51412 540
rect 51664 436 51714 842
rect 51892 598 51920 1716
rect 53172 1714 53240 1724
rect 53052 1541 53116 1548
rect 53052 1510 53058 1541
rect 52324 1489 53058 1510
rect 53110 1489 53116 1541
rect 52324 1482 53116 1489
rect 52324 1480 53058 1482
rect 52324 1474 53052 1480
rect 52224 1144 52288 1152
rect 52224 1092 52230 1144
rect 52282 1092 52288 1144
rect 52224 1084 52288 1092
rect 51984 1056 52050 1062
rect 51984 1004 51992 1056
rect 52044 1026 52050 1056
rect 52224 1026 52252 1084
rect 52044 1004 52252 1026
rect 51984 998 52252 1004
rect 52324 848 52352 1474
rect 53052 1408 53118 1414
rect 53052 1356 53060 1408
rect 53112 1356 53118 1408
rect 53052 1350 53118 1356
rect 53052 1228 53080 1350
rect 53012 1200 53080 1228
rect 52324 840 52636 848
rect 52324 812 52575 840
rect 51984 624 52060 630
rect 51984 598 51992 624
rect 51892 572 51992 598
rect 52044 572 52060 624
rect 51892 570 52060 572
rect 51984 566 52060 570
rect 51664 430 51730 436
rect 51664 378 51672 430
rect 51724 408 51730 430
rect 52324 408 52352 812
rect 52556 788 52575 812
rect 52627 788 52636 840
rect 52556 776 52636 788
rect 52872 844 52940 850
rect 52872 792 52879 844
rect 52931 792 52940 844
rect 52872 786 52940 792
rect 51724 380 52352 408
rect 51724 378 51730 380
rect 51664 372 51730 378
rect 52478 180 52828 194
rect 50590 50 50940 64
rect 52478 64 52499 180
rect 52807 64 52828 180
rect 52872 170 52928 786
rect 53012 616 53040 1200
rect 53074 1150 53136 1156
rect 53074 1098 53084 1150
rect 53172 1142 53200 1714
rect 53228 1541 53292 1548
rect 53228 1489 53234 1541
rect 53286 1508 53292 1541
rect 53554 1508 53604 1898
rect 54076 1896 54104 1996
rect 54076 1890 54142 1896
rect 55190 1894 55218 2000
rect 55426 1958 55492 1966
rect 55426 1906 55432 1958
rect 55484 1906 55492 1958
rect 55426 1898 55492 1906
rect 54076 1876 54084 1890
rect 54078 1838 54084 1876
rect 54136 1838 54142 1890
rect 54078 1832 54142 1838
rect 55150 1888 55218 1894
rect 55150 1836 55160 1888
rect 55212 1836 55218 1888
rect 55150 1830 55218 1836
rect 53990 1774 54054 1780
rect 53990 1744 53996 1774
rect 53780 1722 53996 1744
rect 54048 1722 54054 1774
rect 53780 1716 54054 1722
rect 55060 1776 55128 1782
rect 55060 1724 55068 1776
rect 55120 1724 55128 1776
rect 53286 1492 53606 1508
rect 53286 1489 53620 1492
rect 53228 1486 53620 1489
rect 53228 1480 53562 1486
rect 53554 1434 53562 1480
rect 53614 1434 53620 1486
rect 53554 1428 53620 1434
rect 53424 1292 53496 1304
rect 53424 1240 53434 1292
rect 53486 1240 53496 1292
rect 53424 1228 53496 1240
rect 53460 1226 53496 1228
rect 53172 1114 53460 1142
rect 53074 1092 53136 1098
rect 53108 1046 53136 1092
rect 53108 1042 53352 1046
rect 53108 1036 53390 1042
rect 53108 1018 53330 1036
rect 53324 984 53330 1018
rect 53382 984 53390 1036
rect 53324 976 53390 984
rect 53012 602 53076 616
rect 53432 608 53460 1114
rect 53536 902 53602 910
rect 53536 850 53542 902
rect 53594 850 53602 902
rect 53536 842 53602 850
rect 53012 550 53015 602
rect 53067 550 53076 602
rect 53012 534 53076 550
rect 53246 592 53460 608
rect 53246 540 53247 592
rect 53299 580 53460 592
rect 53299 540 53300 580
rect 53246 524 53300 540
rect 53552 436 53602 842
rect 53780 598 53808 1716
rect 55060 1714 55128 1724
rect 54940 1541 55004 1548
rect 54940 1510 54946 1541
rect 54212 1489 54946 1510
rect 54998 1489 55004 1541
rect 54212 1482 55004 1489
rect 54212 1480 54946 1482
rect 54212 1474 54940 1480
rect 54112 1144 54176 1152
rect 54112 1092 54118 1144
rect 54170 1092 54176 1144
rect 54112 1084 54176 1092
rect 53872 1056 53938 1062
rect 53872 1004 53880 1056
rect 53932 1026 53938 1056
rect 54112 1026 54140 1084
rect 53932 1004 54140 1026
rect 53872 998 54140 1004
rect 54212 848 54240 1474
rect 54940 1408 55006 1414
rect 54940 1356 54948 1408
rect 55000 1356 55006 1408
rect 54940 1350 55006 1356
rect 54940 1228 54968 1350
rect 54900 1200 54968 1228
rect 54212 840 54524 848
rect 54212 812 54463 840
rect 53872 624 53948 630
rect 53872 598 53880 624
rect 53780 572 53880 598
rect 53932 572 53948 624
rect 53780 570 53948 572
rect 53872 566 53948 570
rect 53552 430 53618 436
rect 53552 378 53560 430
rect 53612 408 53618 430
rect 54212 408 54240 812
rect 54444 788 54463 812
rect 54515 788 54524 840
rect 54444 776 54524 788
rect 54760 844 54828 850
rect 54760 792 54767 844
rect 54819 792 54828 844
rect 54760 786 54828 792
rect 53612 380 54240 408
rect 53612 378 53618 380
rect 53552 372 53618 378
rect 54366 180 54716 194
rect 52478 50 52828 64
rect 54366 64 54387 180
rect 54695 64 54716 180
rect 54760 170 54816 786
rect 54900 616 54928 1200
rect 54962 1150 55024 1156
rect 54962 1098 54972 1150
rect 55060 1142 55088 1714
rect 55116 1541 55180 1548
rect 55116 1489 55122 1541
rect 55174 1508 55180 1541
rect 55442 1508 55492 1898
rect 55964 1896 55992 2000
rect 55964 1890 56030 1896
rect 57078 1894 57106 2000
rect 57314 1958 57380 1966
rect 57314 1906 57320 1958
rect 57372 1906 57380 1958
rect 57314 1898 57380 1906
rect 55964 1876 55972 1890
rect 55966 1838 55972 1876
rect 56024 1838 56030 1890
rect 55966 1832 56030 1838
rect 57038 1888 57106 1894
rect 57038 1836 57048 1888
rect 57100 1836 57106 1888
rect 57038 1830 57106 1836
rect 55878 1774 55942 1780
rect 55878 1744 55884 1774
rect 55668 1722 55884 1744
rect 55936 1722 55942 1774
rect 55668 1716 55942 1722
rect 56948 1776 57016 1782
rect 56948 1724 56956 1776
rect 57008 1724 57016 1776
rect 55174 1492 55494 1508
rect 55174 1489 55508 1492
rect 55116 1486 55508 1489
rect 55116 1480 55450 1486
rect 55442 1434 55450 1480
rect 55502 1434 55508 1486
rect 55442 1428 55508 1434
rect 55312 1292 55384 1304
rect 55312 1240 55322 1292
rect 55374 1240 55384 1292
rect 55312 1228 55384 1240
rect 55348 1226 55384 1228
rect 55060 1114 55348 1142
rect 54962 1092 55024 1098
rect 54996 1046 55024 1092
rect 54996 1042 55240 1046
rect 54996 1036 55278 1042
rect 54996 1018 55218 1036
rect 55212 984 55218 1018
rect 55270 984 55278 1036
rect 55212 976 55278 984
rect 54900 602 54964 616
rect 55320 608 55348 1114
rect 55424 902 55490 910
rect 55424 850 55430 902
rect 55482 850 55490 902
rect 55424 842 55490 850
rect 54900 550 54903 602
rect 54955 550 54964 602
rect 54900 534 54964 550
rect 55134 592 55348 608
rect 55134 540 55135 592
rect 55187 580 55348 592
rect 55187 540 55188 580
rect 55134 524 55188 540
rect 55440 436 55490 842
rect 55668 598 55696 1716
rect 56948 1714 57016 1724
rect 56828 1541 56892 1548
rect 56828 1510 56834 1541
rect 56100 1489 56834 1510
rect 56886 1489 56892 1541
rect 56100 1482 56892 1489
rect 56100 1480 56834 1482
rect 56100 1474 56828 1480
rect 56000 1144 56064 1152
rect 56000 1092 56006 1144
rect 56058 1092 56064 1144
rect 56000 1084 56064 1092
rect 55760 1056 55826 1062
rect 55760 1004 55768 1056
rect 55820 1026 55826 1056
rect 56000 1026 56028 1084
rect 55820 1004 56028 1026
rect 55760 998 56028 1004
rect 56100 848 56128 1474
rect 56828 1408 56894 1414
rect 56828 1356 56836 1408
rect 56888 1356 56894 1408
rect 56828 1350 56894 1356
rect 56828 1228 56856 1350
rect 56788 1200 56856 1228
rect 56100 840 56412 848
rect 56100 812 56351 840
rect 55760 624 55836 630
rect 55760 598 55768 624
rect 55668 572 55768 598
rect 55820 572 55836 624
rect 55668 570 55836 572
rect 55760 566 55836 570
rect 55440 430 55506 436
rect 55440 378 55448 430
rect 55500 408 55506 430
rect 56100 408 56128 812
rect 56332 788 56351 812
rect 56403 788 56412 840
rect 56332 776 56412 788
rect 56648 844 56716 850
rect 56648 792 56655 844
rect 56707 792 56716 844
rect 56648 786 56716 792
rect 55500 380 56128 408
rect 55500 378 55506 380
rect 55440 372 55506 378
rect 56254 180 56604 194
rect 54366 50 54716 64
rect 56254 64 56275 180
rect 56583 64 56604 180
rect 56648 170 56704 786
rect 56788 616 56816 1200
rect 56850 1150 56912 1156
rect 56850 1098 56860 1150
rect 56948 1142 56976 1714
rect 57004 1541 57068 1548
rect 57004 1489 57010 1541
rect 57062 1508 57068 1541
rect 57330 1508 57380 1898
rect 57852 1896 57880 2000
rect 57852 1890 57918 1896
rect 58966 1894 58994 2000
rect 59202 1958 59268 1966
rect 59202 1906 59208 1958
rect 59260 1906 59268 1958
rect 59202 1898 59268 1906
rect 57852 1876 57860 1890
rect 57854 1838 57860 1876
rect 57912 1838 57918 1890
rect 57854 1832 57918 1838
rect 58926 1888 58994 1894
rect 58926 1836 58936 1888
rect 58988 1836 58994 1888
rect 58926 1830 58994 1836
rect 57766 1774 57830 1780
rect 57766 1744 57772 1774
rect 57556 1722 57772 1744
rect 57824 1722 57830 1774
rect 57556 1716 57830 1722
rect 58836 1776 58904 1782
rect 58836 1724 58844 1776
rect 58896 1724 58904 1776
rect 57062 1492 57382 1508
rect 57062 1489 57396 1492
rect 57004 1486 57396 1489
rect 57004 1480 57338 1486
rect 57330 1434 57338 1480
rect 57390 1434 57396 1486
rect 57330 1428 57396 1434
rect 57200 1292 57272 1304
rect 57200 1240 57210 1292
rect 57262 1240 57272 1292
rect 57200 1228 57272 1240
rect 57236 1226 57272 1228
rect 56948 1114 57236 1142
rect 56850 1092 56912 1098
rect 56884 1046 56912 1092
rect 56884 1042 57128 1046
rect 56884 1036 57166 1042
rect 56884 1018 57106 1036
rect 57100 984 57106 1018
rect 57158 984 57166 1036
rect 57100 976 57166 984
rect 56788 602 56852 616
rect 57208 608 57236 1114
rect 57312 902 57378 910
rect 57312 850 57318 902
rect 57370 850 57378 902
rect 57312 842 57378 850
rect 56788 550 56791 602
rect 56843 550 56852 602
rect 56788 534 56852 550
rect 57022 592 57236 608
rect 57022 540 57023 592
rect 57075 580 57236 592
rect 57075 540 57076 580
rect 57022 524 57076 540
rect 57328 436 57378 842
rect 57556 598 57584 1716
rect 58836 1714 58904 1724
rect 58716 1541 58780 1548
rect 58716 1510 58722 1541
rect 57988 1489 58722 1510
rect 58774 1489 58780 1541
rect 57988 1482 58780 1489
rect 57988 1480 58722 1482
rect 57988 1474 58716 1480
rect 57888 1144 57952 1152
rect 57888 1092 57894 1144
rect 57946 1092 57952 1144
rect 57888 1084 57952 1092
rect 57648 1056 57714 1062
rect 57648 1004 57656 1056
rect 57708 1026 57714 1056
rect 57888 1026 57916 1084
rect 57708 1004 57916 1026
rect 57648 998 57916 1004
rect 57988 848 58016 1474
rect 58716 1408 58782 1414
rect 58716 1356 58724 1408
rect 58776 1356 58782 1408
rect 58716 1350 58782 1356
rect 58716 1228 58744 1350
rect 58676 1200 58744 1228
rect 57988 840 58300 848
rect 57988 812 58239 840
rect 57648 624 57724 630
rect 57648 598 57656 624
rect 57556 572 57656 598
rect 57708 572 57724 624
rect 57556 570 57724 572
rect 57648 566 57724 570
rect 57328 430 57394 436
rect 57328 378 57336 430
rect 57388 408 57394 430
rect 57988 408 58016 812
rect 58220 788 58239 812
rect 58291 788 58300 840
rect 58220 776 58300 788
rect 58536 844 58604 850
rect 58536 792 58543 844
rect 58595 792 58604 844
rect 58536 786 58604 792
rect 57388 380 58016 408
rect 57388 378 57394 380
rect 57328 372 57394 378
rect 58142 180 58492 194
rect 56254 50 56604 64
rect 58142 64 58163 180
rect 58471 64 58492 180
rect 58536 170 58592 786
rect 58676 616 58704 1200
rect 58738 1150 58800 1156
rect 58738 1098 58748 1150
rect 58836 1142 58864 1714
rect 58892 1541 58956 1548
rect 58892 1489 58898 1541
rect 58950 1508 58956 1541
rect 59218 1508 59268 1898
rect 59740 1896 59768 2000
rect 59740 1890 59806 1896
rect 59740 1876 59748 1890
rect 59742 1838 59748 1876
rect 59800 1838 59806 1890
rect 59742 1832 59806 1838
rect 59654 1774 59718 1780
rect 59654 1744 59660 1774
rect 59444 1722 59660 1744
rect 59712 1722 59718 1774
rect 59444 1716 59718 1722
rect 58950 1492 59270 1508
rect 58950 1489 59284 1492
rect 58892 1486 59284 1489
rect 58892 1480 59226 1486
rect 59218 1434 59226 1480
rect 59278 1434 59284 1486
rect 59218 1428 59284 1434
rect 59088 1292 59160 1304
rect 59088 1240 59098 1292
rect 59150 1240 59160 1292
rect 59088 1228 59160 1240
rect 59124 1226 59160 1228
rect 58836 1114 59124 1142
rect 58738 1092 58800 1098
rect 58772 1046 58800 1092
rect 58772 1042 59016 1046
rect 58772 1036 59054 1042
rect 58772 1018 58994 1036
rect 58988 984 58994 1018
rect 59046 984 59054 1036
rect 58988 976 59054 984
rect 58676 602 58740 616
rect 59096 608 59124 1114
rect 59200 902 59266 910
rect 59200 850 59206 902
rect 59258 850 59266 902
rect 59200 842 59266 850
rect 58676 550 58679 602
rect 58731 550 58740 602
rect 58676 534 58740 550
rect 58910 592 59124 608
rect 58910 540 58911 592
rect 58963 580 59124 592
rect 58963 540 58964 580
rect 58910 524 58964 540
rect 59216 436 59266 842
rect 59444 598 59472 1716
rect 60491 1588 60605 5930
rect 60448 1510 60642 1588
rect 59876 1474 60642 1510
rect 59776 1144 59840 1152
rect 59776 1092 59782 1144
rect 59834 1092 59840 1144
rect 59776 1084 59840 1092
rect 59536 1056 59602 1062
rect 59536 1004 59544 1056
rect 59596 1026 59602 1056
rect 59776 1026 59804 1084
rect 59596 1004 59804 1026
rect 59536 998 59804 1004
rect 59876 848 59904 1474
rect 59876 840 60188 848
rect 59876 812 60127 840
rect 59536 624 59612 630
rect 59536 598 59544 624
rect 59444 572 59544 598
rect 59596 572 59612 624
rect 59444 570 59612 572
rect 59536 566 59612 570
rect 59216 430 59282 436
rect 59216 378 59224 430
rect 59276 408 59282 430
rect 59876 408 59904 812
rect 60108 788 60127 812
rect 60179 788 60188 840
rect 60108 776 60188 788
rect 59276 380 59904 408
rect 59276 378 59282 380
rect 59216 372 59282 378
rect 60030 180 60380 194
rect 58142 50 58492 64
rect 60030 64 60051 180
rect 60359 64 60380 180
rect 60030 50 60380 64
<< via2 >>
rect -371 7290 -315 7346
rect -291 7290 -235 7346
rect -211 7290 -155 7346
rect -131 7290 -75 7346
rect 1517 7290 1573 7346
rect 1597 7290 1653 7346
rect 1677 7290 1733 7346
rect 1757 7290 1813 7346
rect 3405 7290 3461 7346
rect 3485 7290 3541 7346
rect 3565 7290 3621 7346
rect 3645 7290 3701 7346
rect 5293 7290 5349 7346
rect 5373 7290 5429 7346
rect 5453 7290 5509 7346
rect 5533 7290 5589 7346
rect 7181 7290 7237 7346
rect 7261 7290 7317 7346
rect 7341 7290 7397 7346
rect 7421 7290 7477 7346
rect 9069 7290 9125 7346
rect 9149 7290 9205 7346
rect 9229 7290 9285 7346
rect 9309 7290 9365 7346
rect 10957 7290 11013 7346
rect 11037 7290 11093 7346
rect 11117 7290 11173 7346
rect 11197 7290 11253 7346
rect 12845 7290 12901 7346
rect 12925 7290 12981 7346
rect 13005 7290 13061 7346
rect 13085 7290 13141 7346
rect 14727 7290 14783 7346
rect 14807 7290 14863 7346
rect 14887 7290 14943 7346
rect 14967 7290 15023 7346
rect 16615 7290 16671 7346
rect 16695 7290 16751 7346
rect 16775 7290 16831 7346
rect 16855 7290 16911 7346
rect 18503 7290 18559 7346
rect 18583 7290 18639 7346
rect 18663 7290 18719 7346
rect 18743 7290 18799 7346
rect 20391 7290 20447 7346
rect 20471 7290 20527 7346
rect 20551 7290 20607 7346
rect 20631 7290 20687 7346
rect 22279 7290 22335 7346
rect 22359 7290 22415 7346
rect 22439 7290 22495 7346
rect 22519 7290 22575 7346
rect 24167 7290 24223 7346
rect 24247 7290 24303 7346
rect 24327 7290 24383 7346
rect 24407 7290 24463 7346
rect 26055 7290 26111 7346
rect 26135 7290 26191 7346
rect 26215 7290 26271 7346
rect 26295 7290 26351 7346
rect 27943 7290 27999 7346
rect 28023 7290 28079 7346
rect 28103 7290 28159 7346
rect 28183 7290 28239 7346
rect 29831 7290 29887 7346
rect 29911 7290 29967 7346
rect 29991 7290 30047 7346
rect 30071 7290 30127 7346
rect 31719 7290 31775 7346
rect 31799 7290 31855 7346
rect 31879 7290 31935 7346
rect 31959 7290 32015 7346
rect 33607 7290 33663 7346
rect 33687 7290 33743 7346
rect 33767 7290 33823 7346
rect 33847 7290 33903 7346
rect 35495 7290 35551 7346
rect 35575 7290 35631 7346
rect 35655 7290 35711 7346
rect 35735 7290 35791 7346
rect 37383 7290 37439 7346
rect 37463 7290 37519 7346
rect 37543 7290 37599 7346
rect 37623 7290 37679 7346
rect 39271 7290 39327 7346
rect 39351 7290 39407 7346
rect 39431 7290 39487 7346
rect 39511 7290 39567 7346
rect 41159 7290 41215 7346
rect 41239 7290 41295 7346
rect 41319 7290 41375 7346
rect 41399 7290 41455 7346
rect 43047 7290 43103 7346
rect 43127 7290 43183 7346
rect 43207 7290 43263 7346
rect 43287 7290 43343 7346
rect 44929 7290 44985 7346
rect 45009 7290 45065 7346
rect 45089 7290 45145 7346
rect 45169 7290 45225 7346
rect 46817 7290 46873 7346
rect 46897 7290 46953 7346
rect 46977 7290 47033 7346
rect 47057 7290 47113 7346
rect 48705 7290 48761 7346
rect 48785 7290 48841 7346
rect 48865 7290 48921 7346
rect 48945 7290 49001 7346
rect 50593 7290 50649 7346
rect 50673 7290 50729 7346
rect 50753 7290 50809 7346
rect 50833 7290 50889 7346
rect 52481 7290 52537 7346
rect 52561 7290 52617 7346
rect 52641 7290 52697 7346
rect 52721 7290 52777 7346
rect 54369 7290 54425 7346
rect 54449 7290 54505 7346
rect 54529 7290 54585 7346
rect 54609 7290 54665 7346
rect 56257 7290 56313 7346
rect 56337 7290 56393 7346
rect 56417 7290 56473 7346
rect 56497 7290 56553 7346
rect 58145 7290 58201 7346
rect 58225 7290 58281 7346
rect 58305 7290 58361 7346
rect 58385 7290 58441 7346
rect -371 5166 -315 5222
rect -291 5166 -235 5222
rect -211 5166 -155 5222
rect -131 5166 -75 5222
rect 1517 5166 1573 5222
rect 1597 5166 1653 5222
rect 1677 5166 1733 5222
rect 1757 5166 1813 5222
rect 3405 5166 3461 5222
rect 3485 5166 3541 5222
rect 3565 5166 3621 5222
rect 3645 5166 3701 5222
rect 5293 5166 5349 5222
rect 5373 5166 5429 5222
rect 5453 5166 5509 5222
rect 5533 5166 5589 5222
rect 7181 5166 7237 5222
rect 7261 5166 7317 5222
rect 7341 5166 7397 5222
rect 7421 5166 7477 5222
rect 9069 5166 9125 5222
rect 9149 5166 9205 5222
rect 9229 5166 9285 5222
rect 9309 5166 9365 5222
rect 10957 5166 11013 5222
rect 11037 5166 11093 5222
rect 11117 5166 11173 5222
rect 11197 5166 11253 5222
rect 12845 5166 12901 5222
rect 12925 5166 12981 5222
rect 13005 5166 13061 5222
rect 13085 5166 13141 5222
rect 14727 5166 14783 5222
rect 14807 5166 14863 5222
rect 14887 5166 14943 5222
rect 14967 5166 15023 5222
rect 16615 5166 16671 5222
rect 16695 5166 16751 5222
rect 16775 5166 16831 5222
rect 16855 5166 16911 5222
rect 18503 5166 18559 5222
rect 18583 5166 18639 5222
rect 18663 5166 18719 5222
rect 18743 5166 18799 5222
rect 20391 5166 20447 5222
rect 20471 5166 20527 5222
rect 20551 5166 20607 5222
rect 20631 5166 20687 5222
rect 22279 5166 22335 5222
rect 22359 5166 22415 5222
rect 22439 5166 22495 5222
rect 22519 5166 22575 5222
rect 24167 5166 24223 5222
rect 24247 5166 24303 5222
rect 24327 5166 24383 5222
rect 24407 5166 24463 5222
rect 26055 5166 26111 5222
rect 26135 5166 26191 5222
rect 26215 5166 26271 5222
rect 26295 5166 26351 5222
rect 27943 5166 27999 5222
rect 28023 5166 28079 5222
rect 28103 5166 28159 5222
rect 28183 5166 28239 5222
rect 29831 5166 29887 5222
rect 29911 5166 29967 5222
rect 29991 5166 30047 5222
rect 30071 5166 30127 5222
rect 31719 5166 31775 5222
rect 31799 5166 31855 5222
rect 31879 5166 31935 5222
rect 31959 5166 32015 5222
rect 33607 5166 33663 5222
rect 33687 5166 33743 5222
rect 33767 5166 33823 5222
rect 33847 5166 33903 5222
rect 35495 5166 35551 5222
rect 35575 5166 35631 5222
rect 35655 5166 35711 5222
rect 35735 5166 35791 5222
rect 37383 5166 37439 5222
rect 37463 5166 37519 5222
rect 37543 5166 37599 5222
rect 37623 5166 37679 5222
rect 39271 5166 39327 5222
rect 39351 5166 39407 5222
rect 39431 5166 39487 5222
rect 39511 5166 39567 5222
rect 41159 5166 41215 5222
rect 41239 5166 41295 5222
rect 41319 5166 41375 5222
rect 41399 5166 41455 5222
rect 43047 5166 43103 5222
rect 43127 5166 43183 5222
rect 43207 5166 43263 5222
rect 43287 5166 43343 5222
rect 44929 5166 44985 5222
rect 45009 5166 45065 5222
rect 45089 5166 45145 5222
rect 45169 5166 45225 5222
rect 46817 5166 46873 5222
rect 46897 5166 46953 5222
rect 46977 5166 47033 5222
rect 47057 5166 47113 5222
rect 48705 5166 48761 5222
rect 48785 5166 48841 5222
rect 48865 5166 48921 5222
rect 48945 5166 49001 5222
rect 50593 5166 50649 5222
rect 50673 5166 50729 5222
rect 50753 5166 50809 5222
rect 50833 5166 50889 5222
rect 52481 5166 52537 5222
rect 52561 5166 52617 5222
rect 52641 5166 52697 5222
rect 52721 5166 52777 5222
rect 54369 5166 54425 5222
rect 54449 5166 54505 5222
rect 54529 5166 54585 5222
rect 54609 5166 54665 5222
rect 56257 5166 56313 5222
rect 56337 5166 56393 5222
rect 56417 5166 56473 5222
rect 56497 5166 56553 5222
rect 58145 5166 58201 5222
rect 58225 5166 58281 5222
rect 58305 5166 58361 5222
rect 58385 5166 58441 5222
rect 6275 3316 6331 3372
rect 6389 3316 6445 3372
rect 6503 3316 6559 3372
rect 6275 3201 6331 3257
rect 6389 3201 6445 3257
rect 6503 3201 6559 3257
rect 6275 3086 6331 3142
rect 6389 3086 6445 3142
rect 6503 3086 6559 3142
rect 21314 3226 21370 3282
rect 21418 3226 21474 3282
rect 21522 3226 21578 3282
rect 21626 3226 21682 3282
rect 21314 3110 21370 3166
rect 21418 3110 21474 3166
rect 21522 3110 21578 3166
rect 21626 3110 21682 3166
rect 21314 2994 21370 3050
rect 21418 2994 21474 3050
rect 21522 2994 21578 3050
rect 21626 2994 21682 3050
rect 13669 2755 13725 2811
rect 13777 2755 13833 2811
rect 13885 2755 13941 2811
rect 13669 2661 13725 2717
rect 13777 2661 13833 2717
rect 13885 2661 13941 2717
rect 36401 3575 36457 3631
rect 36495 3575 36551 3631
rect 36589 3575 36645 3631
rect 36401 3487 36457 3543
rect 36495 3487 36551 3543
rect 36589 3487 36645 3543
rect 36401 3399 36457 3455
rect 36495 3399 36551 3455
rect 36589 3399 36645 3455
rect 30364 2875 30420 2931
rect 30489 2875 30545 2931
rect 30614 2875 30670 2931
rect 30364 2779 30420 2835
rect 30489 2779 30545 2835
rect 30614 2779 30670 2835
rect 46035 2728 46091 2784
rect 46128 2728 46184 2784
rect 46221 2728 46277 2784
rect 46314 2728 46370 2784
rect 46035 2646 46091 2702
rect 46128 2646 46184 2702
rect 46221 2646 46277 2702
rect 46314 2646 46370 2702
rect 53348 3120 53404 3176
rect 53452 3120 53508 3176
rect 53556 3120 53612 3176
rect 53660 3120 53716 3176
rect 53348 3030 53404 3086
rect 53452 3030 53508 3086
rect 53556 3030 53612 3086
rect 53660 3030 53716 3086
rect 1541 2218 1597 2274
rect 1621 2218 1677 2274
rect 1701 2218 1757 2274
rect 1781 2218 1837 2274
rect 3429 2218 3485 2274
rect 3509 2218 3565 2274
rect 3589 2218 3645 2274
rect 3669 2218 3725 2274
rect 5317 2218 5373 2274
rect 5397 2218 5453 2274
rect 5477 2218 5533 2274
rect 5557 2218 5613 2274
rect 7205 2218 7261 2274
rect 7285 2218 7341 2274
rect 7365 2218 7421 2274
rect 7445 2218 7501 2274
rect 9093 2218 9149 2274
rect 9173 2218 9229 2274
rect 9253 2218 9309 2274
rect 9333 2218 9389 2274
rect 10981 2218 11037 2274
rect 11061 2218 11117 2274
rect 11141 2218 11197 2274
rect 11221 2218 11277 2274
rect 12869 2218 12925 2274
rect 12949 2218 13005 2274
rect 13029 2218 13085 2274
rect 13109 2218 13165 2274
rect 14757 2218 14813 2274
rect 14837 2218 14893 2274
rect 14917 2218 14973 2274
rect 14997 2218 15053 2274
rect 16639 2218 16695 2274
rect 16719 2218 16775 2274
rect 16799 2218 16855 2274
rect 16879 2218 16935 2274
rect 18527 2218 18583 2274
rect 18607 2218 18663 2274
rect 18687 2218 18743 2274
rect 18767 2218 18823 2274
rect 20415 2218 20471 2274
rect 20495 2218 20551 2274
rect 20575 2218 20631 2274
rect 20655 2218 20711 2274
rect 22303 2218 22359 2274
rect 22383 2218 22439 2274
rect 22463 2218 22519 2274
rect 22543 2218 22599 2274
rect 24191 2218 24247 2274
rect 24271 2218 24327 2274
rect 24351 2218 24407 2274
rect 24431 2218 24487 2274
rect 26079 2218 26135 2274
rect 26159 2218 26215 2274
rect 26239 2218 26295 2274
rect 26319 2218 26375 2274
rect 27967 2218 28023 2274
rect 28047 2218 28103 2274
rect 28127 2218 28183 2274
rect 28207 2218 28263 2274
rect 29855 2218 29911 2274
rect 29935 2218 29991 2274
rect 30015 2218 30071 2274
rect 30095 2218 30151 2274
rect 31743 2218 31799 2274
rect 31823 2218 31879 2274
rect 31903 2218 31959 2274
rect 31983 2218 32039 2274
rect 33631 2218 33687 2274
rect 33711 2218 33767 2274
rect 33791 2218 33847 2274
rect 33871 2218 33927 2274
rect 35519 2218 35575 2274
rect 35599 2218 35655 2274
rect 35679 2218 35735 2274
rect 35759 2218 35815 2274
rect 37407 2218 37463 2274
rect 37487 2218 37543 2274
rect 37567 2218 37623 2274
rect 37647 2218 37703 2274
rect 39295 2218 39351 2274
rect 39375 2218 39431 2274
rect 39455 2218 39511 2274
rect 39535 2218 39591 2274
rect 41183 2218 41239 2274
rect 41263 2218 41319 2274
rect 41343 2218 41399 2274
rect 41423 2218 41479 2274
rect 43071 2218 43127 2274
rect 43151 2218 43207 2274
rect 43231 2218 43287 2274
rect 43311 2218 43367 2274
rect 44959 2218 45015 2274
rect 45039 2218 45095 2274
rect 45119 2218 45175 2274
rect 45199 2218 45255 2274
rect 46841 2218 46897 2274
rect 46921 2218 46977 2274
rect 47001 2218 47057 2274
rect 47081 2218 47137 2274
rect 48729 2218 48785 2274
rect 48809 2218 48865 2274
rect 48889 2218 48945 2274
rect 48969 2218 49025 2274
rect 50617 2218 50673 2274
rect 50697 2218 50753 2274
rect 50777 2218 50833 2274
rect 50857 2218 50913 2274
rect 52505 2218 52561 2274
rect 52585 2218 52641 2274
rect 52665 2218 52721 2274
rect 52745 2218 52801 2274
rect 54393 2218 54449 2274
rect 54473 2218 54529 2274
rect 54553 2218 54609 2274
rect 54633 2218 54689 2274
rect 56281 2218 56337 2274
rect 56361 2218 56417 2274
rect 56441 2218 56497 2274
rect 56521 2218 56577 2274
rect 58169 2218 58225 2274
rect 58249 2218 58305 2274
rect 58329 2218 58385 2274
rect 58409 2218 58465 2274
rect 60057 2218 60113 2274
rect 60137 2218 60193 2274
rect 60217 2218 60273 2274
rect 60297 2218 60353 2274
rect 1541 94 1597 150
rect 1621 94 1677 150
rect 1701 94 1757 150
rect 1781 94 1837 150
rect 3429 94 3485 150
rect 3509 94 3565 150
rect 3589 94 3645 150
rect 3669 94 3725 150
rect 5317 94 5373 150
rect 5397 94 5453 150
rect 5477 94 5533 150
rect 5557 94 5613 150
rect 7205 94 7261 150
rect 7285 94 7341 150
rect 7365 94 7421 150
rect 7445 94 7501 150
rect 9093 94 9149 150
rect 9173 94 9229 150
rect 9253 94 9309 150
rect 9333 94 9389 150
rect 10981 94 11037 150
rect 11061 94 11117 150
rect 11141 94 11197 150
rect 11221 94 11277 150
rect 12869 94 12925 150
rect 12949 94 13005 150
rect 13029 94 13085 150
rect 13109 94 13165 150
rect 14757 94 14813 150
rect 14837 94 14893 150
rect 14917 94 14973 150
rect 14997 94 15053 150
rect 16639 94 16695 150
rect 16719 94 16775 150
rect 16799 94 16855 150
rect 16879 94 16935 150
rect 18527 94 18583 150
rect 18607 94 18663 150
rect 18687 94 18743 150
rect 18767 94 18823 150
rect 20415 94 20471 150
rect 20495 94 20551 150
rect 20575 94 20631 150
rect 20655 94 20711 150
rect 22303 94 22359 150
rect 22383 94 22439 150
rect 22463 94 22519 150
rect 22543 94 22599 150
rect 24191 94 24247 150
rect 24271 94 24327 150
rect 24351 94 24407 150
rect 24431 94 24487 150
rect 26079 94 26135 150
rect 26159 94 26215 150
rect 26239 94 26295 150
rect 26319 94 26375 150
rect 27967 94 28023 150
rect 28047 94 28103 150
rect 28127 94 28183 150
rect 28207 94 28263 150
rect 29855 94 29911 150
rect 29935 94 29991 150
rect 30015 94 30071 150
rect 30095 94 30151 150
rect 31743 94 31799 150
rect 31823 94 31879 150
rect 31903 94 31959 150
rect 31983 94 32039 150
rect 33631 94 33687 150
rect 33711 94 33767 150
rect 33791 94 33847 150
rect 33871 94 33927 150
rect 35519 94 35575 150
rect 35599 94 35655 150
rect 35679 94 35735 150
rect 35759 94 35815 150
rect 37407 94 37463 150
rect 37487 94 37543 150
rect 37567 94 37623 150
rect 37647 94 37703 150
rect 39295 94 39351 150
rect 39375 94 39431 150
rect 39455 94 39511 150
rect 39535 94 39591 150
rect 41183 94 41239 150
rect 41263 94 41319 150
rect 41343 94 41399 150
rect 41423 94 41479 150
rect 43071 94 43127 150
rect 43151 94 43207 150
rect 43231 94 43287 150
rect 43311 94 43367 150
rect 44959 94 45015 150
rect 45039 94 45095 150
rect 45119 94 45175 150
rect 45199 94 45255 150
rect 46841 94 46897 150
rect 46921 94 46977 150
rect 47001 94 47057 150
rect 47081 94 47137 150
rect 48729 94 48785 150
rect 48809 94 48865 150
rect 48889 94 48945 150
rect 48969 94 49025 150
rect 50617 94 50673 150
rect 50697 94 50753 150
rect 50777 94 50833 150
rect 50857 94 50913 150
rect 52505 94 52561 150
rect 52585 94 52641 150
rect 52665 94 52721 150
rect 52745 94 52801 150
rect 54393 94 54449 150
rect 54473 94 54529 150
rect 54553 94 54609 150
rect 54633 94 54689 150
rect 56281 94 56337 150
rect 56361 94 56417 150
rect 56441 94 56497 150
rect 56521 94 56577 150
rect 58169 94 58225 150
rect 58249 94 58305 150
rect 58329 94 58385 150
rect 58409 94 58465 150
rect 60057 94 60113 150
rect 60137 94 60193 150
rect 60217 94 60273 150
rect 60297 94 60353 150
<< metal3 >>
rect 1458 7440 14674 7441
rect 16556 7440 29772 7441
rect 31660 7440 44876 7441
rect 46758 7440 59974 7441
rect -430 7390 59974 7440
rect -430 7389 3073 7390
rect -430 7346 2518 7389
rect -430 7290 -371 7346
rect -315 7290 -291 7346
rect -235 7290 -211 7346
rect -155 7290 -131 7346
rect -75 7290 1517 7346
rect 1573 7290 1597 7346
rect 1653 7290 1677 7346
rect 1733 7290 1757 7346
rect 1813 7290 2518 7346
rect -430 7211 2518 7290
rect 2624 7388 3073 7389
rect 2624 7211 2727 7388
rect -430 7210 2727 7211
rect 2833 7210 2893 7388
rect 2999 7212 3073 7388
rect 3179 7346 59974 7390
rect 3179 7290 3405 7346
rect 3461 7290 3485 7346
rect 3541 7290 3565 7346
rect 3621 7290 3645 7346
rect 3701 7290 5293 7346
rect 5349 7290 5373 7346
rect 5429 7290 5453 7346
rect 5509 7290 5533 7346
rect 5589 7290 7181 7346
rect 7237 7290 7261 7346
rect 7317 7290 7341 7346
rect 7397 7290 7421 7346
rect 7477 7290 9069 7346
rect 9125 7290 9149 7346
rect 9205 7290 9229 7346
rect 9285 7290 9309 7346
rect 9365 7290 10957 7346
rect 11013 7290 11037 7346
rect 11093 7290 11117 7346
rect 11173 7290 11197 7346
rect 11253 7290 12845 7346
rect 12901 7290 12925 7346
rect 12981 7290 13005 7346
rect 13061 7290 13085 7346
rect 13141 7290 14727 7346
rect 14783 7290 14807 7346
rect 14863 7290 14887 7346
rect 14943 7290 14967 7346
rect 15023 7290 16615 7346
rect 16671 7290 16695 7346
rect 16751 7290 16775 7346
rect 16831 7290 16855 7346
rect 16911 7290 18503 7346
rect 18559 7290 18583 7346
rect 18639 7290 18663 7346
rect 18719 7290 18743 7346
rect 18799 7290 20391 7346
rect 20447 7290 20471 7346
rect 20527 7290 20551 7346
rect 20607 7290 20631 7346
rect 20687 7290 22279 7346
rect 22335 7290 22359 7346
rect 22415 7290 22439 7346
rect 22495 7290 22519 7346
rect 22575 7290 24167 7346
rect 24223 7290 24247 7346
rect 24303 7290 24327 7346
rect 24383 7290 24407 7346
rect 24463 7290 26055 7346
rect 26111 7290 26135 7346
rect 26191 7290 26215 7346
rect 26271 7290 26295 7346
rect 26351 7290 27943 7346
rect 27999 7290 28023 7346
rect 28079 7290 28103 7346
rect 28159 7290 28183 7346
rect 28239 7290 29831 7346
rect 29887 7290 29911 7346
rect 29967 7290 29991 7346
rect 30047 7290 30071 7346
rect 30127 7290 31719 7346
rect 31775 7290 31799 7346
rect 31855 7290 31879 7346
rect 31935 7290 31959 7346
rect 32015 7290 33607 7346
rect 33663 7290 33687 7346
rect 33743 7290 33767 7346
rect 33823 7290 33847 7346
rect 33903 7290 35495 7346
rect 35551 7290 35575 7346
rect 35631 7290 35655 7346
rect 35711 7290 35735 7346
rect 35791 7290 37383 7346
rect 37439 7290 37463 7346
rect 37519 7290 37543 7346
rect 37599 7290 37623 7346
rect 37679 7290 39271 7346
rect 39327 7290 39351 7346
rect 39407 7290 39431 7346
rect 39487 7290 39511 7346
rect 39567 7290 41159 7346
rect 41215 7290 41239 7346
rect 41295 7290 41319 7346
rect 41375 7290 41399 7346
rect 41455 7290 43047 7346
rect 43103 7290 43127 7346
rect 43183 7290 43207 7346
rect 43263 7290 43287 7346
rect 43343 7290 44929 7346
rect 44985 7290 45009 7346
rect 45065 7290 45089 7346
rect 45145 7290 45169 7346
rect 45225 7290 46817 7346
rect 46873 7290 46897 7346
rect 46953 7290 46977 7346
rect 47033 7290 47057 7346
rect 47113 7290 48705 7346
rect 48761 7290 48785 7346
rect 48841 7290 48865 7346
rect 48921 7290 48945 7346
rect 49001 7290 50593 7346
rect 50649 7290 50673 7346
rect 50729 7290 50753 7346
rect 50809 7290 50833 7346
rect 50889 7290 52481 7346
rect 52537 7290 52561 7346
rect 52617 7290 52641 7346
rect 52697 7290 52721 7346
rect 52777 7290 54369 7346
rect 54425 7290 54449 7346
rect 54505 7290 54529 7346
rect 54585 7290 54609 7346
rect 54665 7290 56257 7346
rect 56313 7290 56337 7346
rect 56393 7290 56417 7346
rect 56473 7290 56497 7346
rect 56553 7290 58145 7346
rect 58201 7290 58225 7346
rect 58281 7290 58305 7346
rect 58361 7290 58385 7346
rect 58441 7290 59974 7346
rect 3179 7212 59974 7290
rect 2999 7210 59974 7212
rect -430 7186 59974 7210
rect -430 5272 59982 5318
rect -430 5271 1456 5272
rect -430 5222 1284 5271
rect -430 5166 -371 5222
rect -315 5166 -291 5222
rect -235 5166 -211 5222
rect -155 5166 -131 5222
rect -75 5166 1284 5222
rect -430 5093 1284 5166
rect 1390 5094 1456 5271
rect 1562 5271 59982 5272
rect 1562 5222 1630 5271
rect 1736 5222 59982 5271
rect 1573 5166 1597 5222
rect 1736 5166 1757 5222
rect 1813 5166 3405 5222
rect 3461 5166 3485 5222
rect 3541 5166 3565 5222
rect 3621 5166 3645 5222
rect 3701 5166 5293 5222
rect 5349 5166 5373 5222
rect 5429 5166 5453 5222
rect 5509 5166 5533 5222
rect 5589 5166 7181 5222
rect 7237 5166 7261 5222
rect 7317 5166 7341 5222
rect 7397 5166 7421 5222
rect 7477 5166 9069 5222
rect 9125 5166 9149 5222
rect 9205 5166 9229 5222
rect 9285 5166 9309 5222
rect 9365 5166 10957 5222
rect 11013 5166 11037 5222
rect 11093 5166 11117 5222
rect 11173 5166 11197 5222
rect 11253 5166 12845 5222
rect 12901 5166 12925 5222
rect 12981 5166 13005 5222
rect 13061 5166 13085 5222
rect 13141 5166 14727 5222
rect 14783 5166 14807 5222
rect 14863 5166 14887 5222
rect 14943 5166 14967 5222
rect 15023 5166 16615 5222
rect 16671 5166 16695 5222
rect 16751 5166 16775 5222
rect 16831 5166 16855 5222
rect 16911 5166 18503 5222
rect 18559 5166 18583 5222
rect 18639 5166 18663 5222
rect 18719 5166 18743 5222
rect 18799 5166 20391 5222
rect 20447 5166 20471 5222
rect 20527 5166 20551 5222
rect 20607 5166 20631 5222
rect 20687 5166 22279 5222
rect 22335 5166 22359 5222
rect 22415 5166 22439 5222
rect 22495 5166 22519 5222
rect 22575 5166 24167 5222
rect 24223 5166 24247 5222
rect 24303 5166 24327 5222
rect 24383 5166 24407 5222
rect 24463 5166 26055 5222
rect 26111 5166 26135 5222
rect 26191 5166 26215 5222
rect 26271 5166 26295 5222
rect 26351 5166 27943 5222
rect 27999 5166 28023 5222
rect 28079 5166 28103 5222
rect 28159 5166 28183 5222
rect 28239 5166 29831 5222
rect 29887 5166 29911 5222
rect 29967 5166 29991 5222
rect 30047 5166 30071 5222
rect 30127 5166 31719 5222
rect 31775 5166 31799 5222
rect 31855 5166 31879 5222
rect 31935 5166 31959 5222
rect 32015 5166 33607 5222
rect 33663 5166 33687 5222
rect 33743 5166 33767 5222
rect 33823 5166 33847 5222
rect 33903 5166 35495 5222
rect 35551 5166 35575 5222
rect 35631 5166 35655 5222
rect 35711 5166 35735 5222
rect 35791 5166 37383 5222
rect 37439 5166 37463 5222
rect 37519 5166 37543 5222
rect 37599 5166 37623 5222
rect 37679 5166 39271 5222
rect 39327 5166 39351 5222
rect 39407 5166 39431 5222
rect 39487 5166 39511 5222
rect 39567 5166 41159 5222
rect 41215 5166 41239 5222
rect 41295 5166 41319 5222
rect 41375 5166 41399 5222
rect 41455 5166 43047 5222
rect 43103 5166 43127 5222
rect 43183 5166 43207 5222
rect 43263 5166 43287 5222
rect 43343 5166 44929 5222
rect 44985 5166 45009 5222
rect 45065 5166 45089 5222
rect 45145 5166 45169 5222
rect 45225 5166 46817 5222
rect 46873 5166 46897 5222
rect 46953 5166 46977 5222
rect 47033 5166 47057 5222
rect 47113 5166 48705 5222
rect 48761 5166 48785 5222
rect 48841 5166 48865 5222
rect 48921 5166 48945 5222
rect 49001 5166 50593 5222
rect 50649 5166 50673 5222
rect 50729 5166 50753 5222
rect 50809 5166 50833 5222
rect 50889 5166 52481 5222
rect 52537 5166 52561 5222
rect 52617 5166 52641 5222
rect 52697 5166 52721 5222
rect 52777 5166 54369 5222
rect 54425 5166 54449 5222
rect 54505 5166 54529 5222
rect 54585 5166 54609 5222
rect 54665 5166 56257 5222
rect 56313 5166 56337 5222
rect 56393 5166 56417 5222
rect 56473 5166 56497 5222
rect 56553 5166 58145 5222
rect 58201 5166 58225 5222
rect 58281 5166 58305 5222
rect 58361 5166 58385 5222
rect 58441 5166 59982 5222
rect 1562 5094 1630 5166
rect 1390 5093 1630 5094
rect 1736 5093 59982 5166
rect -430 5064 59982 5093
rect 36378 3631 36682 3645
rect 36378 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36682 3631
rect 36378 3543 36682 3575
rect 36378 3487 36401 3543
rect 36457 3532 36495 3543
rect 36551 3533 36589 3543
rect 36645 3533 36682 3543
rect 36551 3487 36568 3533
rect 36378 3455 36414 3487
rect 36501 3455 36568 3487
rect 6274 3398 6616 3431
rect 36378 3399 36401 3455
rect 36551 3421 36568 3455
rect 36655 3421 36682 3533
rect 36457 3399 36495 3420
rect 36551 3399 36589 3421
rect 36645 3399 36682 3421
rect 6206 3372 6695 3398
rect 36378 3379 36682 3399
rect 6206 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6695 3372
rect 6206 3257 6695 3316
rect 6206 3229 6275 3257
rect 6331 3229 6389 3257
rect 6445 3235 6503 3257
rect 6559 3235 6695 3257
rect 6206 3138 6272 3229
rect 6358 3201 6389 3229
rect 6559 3201 6568 3235
rect 6358 3144 6423 3201
rect 6509 3144 6568 3201
rect 6654 3144 6695 3235
rect 6358 3142 6695 3144
rect 6358 3138 6389 3142
rect 6206 3086 6275 3138
rect 6331 3086 6389 3138
rect 6445 3086 6503 3142
rect 6559 3086 6695 3142
rect 6206 3031 6695 3086
rect 21264 3282 21731 3336
rect 21264 3239 21314 3282
rect 21370 3239 21418 3282
rect 21264 3155 21312 3239
rect 21405 3226 21418 3239
rect 21474 3239 21522 3282
rect 21474 3226 21479 3239
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21405 3166 21479 3226
rect 21572 3166 21731 3226
rect 21405 3155 21418 3166
rect 21264 3110 21314 3155
rect 21370 3110 21418 3155
rect 21474 3155 21479 3166
rect 21474 3110 21522 3155
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3078 21731 3110
rect 21264 2994 21312 3078
rect 21405 3050 21479 3078
rect 21572 3050 21731 3078
rect 21405 2994 21418 3050
rect 21474 2994 21479 3050
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 53311 3183 53733 3204
rect 53311 3176 53355 3183
rect 53439 3176 53476 3183
rect 53560 3176 53614 3183
rect 53698 3176 53733 3183
rect 53311 3120 53348 3176
rect 53439 3120 53452 3176
rect 53612 3120 53614 3176
rect 53716 3120 53733 3176
rect 53311 3086 53355 3120
rect 53439 3086 53476 3120
rect 53560 3086 53614 3120
rect 53698 3086 53733 3120
rect 53311 3030 53348 3086
rect 53439 3030 53452 3086
rect 53612 3030 53614 3086
rect 53716 3030 53733 3086
rect 53311 3025 53355 3030
rect 53439 3025 53476 3030
rect 53560 3025 53614 3030
rect 53698 3025 53733 3030
rect 53311 2996 53733 3025
rect 21264 2950 21731 2994
rect 30316 2931 30741 2969
rect 30316 2892 30364 2931
rect 30420 2892 30489 2931
rect 30545 2892 30614 2931
rect 30670 2892 30741 2931
rect 13629 2811 13982 2834
rect 13629 2763 13669 2811
rect 13725 2763 13777 2811
rect 13833 2763 13885 2811
rect 13629 2694 13653 2763
rect 13730 2694 13756 2763
rect 13833 2694 13859 2763
rect 13941 2755 13982 2811
rect 13936 2717 13982 2755
rect 30316 2780 30362 2892
rect 30449 2780 30481 2892
rect 30568 2780 30600 2892
rect 30687 2780 30741 2892
rect 30316 2779 30364 2780
rect 30420 2779 30489 2780
rect 30545 2779 30614 2780
rect 30670 2779 30741 2780
rect 30316 2742 30741 2779
rect 45998 2808 46413 2851
rect 45998 2807 46176 2808
rect 45998 2784 46036 2807
rect 46120 2784 46176 2807
rect 46260 2784 46304 2808
rect 13629 2661 13669 2694
rect 13725 2661 13777 2694
rect 13833 2661 13885 2694
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 45998 2728 46035 2784
rect 46120 2728 46128 2784
rect 46277 2728 46304 2784
rect 45998 2702 46036 2728
rect 46120 2702 46176 2728
rect 46260 2702 46304 2728
rect 45998 2646 46035 2702
rect 46120 2649 46128 2702
rect 46277 2650 46304 2702
rect 46388 2650 46413 2808
rect 46091 2646 46128 2649
rect 46184 2646 46221 2650
rect 46277 2646 46314 2650
rect 46370 2646 46413 2650
rect 45998 2610 46413 2646
rect 0 2325 60412 2376
rect 0 2323 1491 2325
rect 0 2145 1286 2323
rect 1392 2147 1491 2323
rect 1597 2274 1690 2325
rect 1796 2274 60412 2325
rect 1597 2218 1621 2274
rect 1677 2218 1690 2274
rect 1837 2218 3429 2274
rect 3485 2218 3509 2274
rect 3565 2218 3589 2274
rect 3645 2218 3669 2274
rect 3725 2218 5317 2274
rect 5373 2218 5397 2274
rect 5453 2218 5477 2274
rect 5533 2218 5557 2274
rect 5613 2218 7205 2274
rect 7261 2218 7285 2274
rect 7341 2218 7365 2274
rect 7421 2218 7445 2274
rect 7501 2218 9093 2274
rect 9149 2218 9173 2274
rect 9229 2218 9253 2274
rect 9309 2218 9333 2274
rect 9389 2218 10981 2274
rect 11037 2218 11061 2274
rect 11117 2218 11141 2274
rect 11197 2218 11221 2274
rect 11277 2218 12869 2274
rect 12925 2218 12949 2274
rect 13005 2218 13029 2274
rect 13085 2218 13109 2274
rect 13165 2218 14757 2274
rect 14813 2218 14837 2274
rect 14893 2218 14917 2274
rect 14973 2218 14997 2274
rect 15053 2218 16639 2274
rect 16695 2218 16719 2274
rect 16775 2218 16799 2274
rect 16855 2218 16879 2274
rect 16935 2218 18527 2274
rect 18583 2218 18607 2274
rect 18663 2218 18687 2274
rect 18743 2218 18767 2274
rect 18823 2218 20415 2274
rect 20471 2218 20495 2274
rect 20551 2218 20575 2274
rect 20631 2218 20655 2274
rect 20711 2218 22303 2274
rect 22359 2218 22383 2274
rect 22439 2218 22463 2274
rect 22519 2218 22543 2274
rect 22599 2218 24191 2274
rect 24247 2218 24271 2274
rect 24327 2218 24351 2274
rect 24407 2218 24431 2274
rect 24487 2218 26079 2274
rect 26135 2218 26159 2274
rect 26215 2218 26239 2274
rect 26295 2218 26319 2274
rect 26375 2218 27967 2274
rect 28023 2218 28047 2274
rect 28103 2218 28127 2274
rect 28183 2218 28207 2274
rect 28263 2218 29855 2274
rect 29911 2218 29935 2274
rect 29991 2218 30015 2274
rect 30071 2218 30095 2274
rect 30151 2218 31743 2274
rect 31799 2218 31823 2274
rect 31879 2218 31903 2274
rect 31959 2218 31983 2274
rect 32039 2218 33631 2274
rect 33687 2218 33711 2274
rect 33767 2218 33791 2274
rect 33847 2218 33871 2274
rect 33927 2218 35519 2274
rect 35575 2218 35599 2274
rect 35655 2218 35679 2274
rect 35735 2218 35759 2274
rect 35815 2218 37407 2274
rect 37463 2218 37487 2274
rect 37543 2218 37567 2274
rect 37623 2218 37647 2274
rect 37703 2218 39295 2274
rect 39351 2218 39375 2274
rect 39431 2218 39455 2274
rect 39511 2218 39535 2274
rect 39591 2218 41183 2274
rect 41239 2218 41263 2274
rect 41319 2218 41343 2274
rect 41399 2218 41423 2274
rect 41479 2218 43071 2274
rect 43127 2218 43151 2274
rect 43207 2218 43231 2274
rect 43287 2218 43311 2274
rect 43367 2218 44959 2274
rect 45015 2218 45039 2274
rect 45095 2218 45119 2274
rect 45175 2218 45199 2274
rect 45255 2218 46841 2274
rect 46897 2218 46921 2274
rect 46977 2218 47001 2274
rect 47057 2218 47081 2274
rect 47137 2218 48729 2274
rect 48785 2218 48809 2274
rect 48865 2218 48889 2274
rect 48945 2218 48969 2274
rect 49025 2218 50617 2274
rect 50673 2218 50697 2274
rect 50753 2218 50777 2274
rect 50833 2218 50857 2274
rect 50913 2218 52505 2274
rect 52561 2218 52585 2274
rect 52641 2218 52665 2274
rect 52721 2218 52745 2274
rect 52801 2218 54393 2274
rect 54449 2218 54473 2274
rect 54529 2218 54553 2274
rect 54609 2218 54633 2274
rect 54689 2218 56281 2274
rect 56337 2218 56361 2274
rect 56417 2218 56441 2274
rect 56497 2218 56521 2274
rect 56577 2218 58169 2274
rect 58225 2218 58249 2274
rect 58305 2218 58329 2274
rect 58385 2218 58409 2274
rect 58465 2218 60057 2274
rect 60113 2218 60137 2274
rect 60193 2218 60217 2274
rect 60273 2218 60297 2274
rect 60353 2218 60412 2274
rect 1597 2147 1690 2218
rect 1796 2147 60412 2218
rect 1392 2145 60412 2147
rect 0 2122 60412 2145
rect 8 212 60412 254
rect 8 150 2532 212
rect 8 94 1541 150
rect 1597 94 1621 150
rect 1677 94 1701 150
rect 1757 94 1781 150
rect 1837 94 2532 150
rect 8 34 2532 94
rect 2638 34 2753 212
rect 2859 34 2962 212
rect 3068 34 3136 212
rect 3242 209 60412 212
rect 3242 157 13779 209
rect 3242 150 6260 157
rect 3242 94 3429 150
rect 3485 94 3509 150
rect 3565 94 3589 150
rect 3645 94 3669 150
rect 3725 94 5317 150
rect 5373 94 5397 150
rect 5453 94 5477 150
rect 5533 94 5557 150
rect 5613 94 6260 150
rect 3242 66 6260 94
rect 6346 66 6408 157
rect 6494 66 6556 157
rect 6642 150 13779 157
rect 6642 94 7205 150
rect 7261 94 7285 150
rect 7341 94 7365 150
rect 7421 94 7445 150
rect 7501 94 9093 150
rect 9149 94 9173 150
rect 9229 94 9253 150
rect 9309 94 9333 150
rect 9389 94 10981 150
rect 11037 94 11061 150
rect 11117 94 11141 150
rect 11197 94 11221 150
rect 11277 94 12869 150
rect 12925 94 12949 150
rect 13005 94 13029 150
rect 13085 94 13109 150
rect 13165 140 13779 150
rect 13856 200 60412 209
rect 13856 190 53361 200
rect 13856 169 46038 190
rect 13856 150 21317 169
rect 13856 140 14757 150
rect 13165 94 14757 140
rect 14813 94 14837 150
rect 14893 94 14917 150
rect 14973 94 14997 150
rect 15053 94 16639 150
rect 16695 94 16719 150
rect 16775 94 16799 150
rect 16855 94 16879 150
rect 16935 94 18527 150
rect 18583 94 18607 150
rect 18663 94 18687 150
rect 18743 94 18767 150
rect 18823 94 20415 150
rect 20471 94 20495 150
rect 20551 94 20575 150
rect 20631 94 20655 150
rect 20711 94 21317 150
rect 6642 90 21317 94
rect 6642 66 13802 90
rect 3242 34 13802 66
rect 8 21 13802 34
rect 13879 61 21317 90
rect 21413 61 21450 169
rect 21546 61 21583 169
rect 21679 160 46038 169
rect 21679 150 30383 160
rect 21679 94 22303 150
rect 22359 94 22383 150
rect 22439 94 22463 150
rect 22519 94 22543 150
rect 22599 94 24191 150
rect 24247 94 24271 150
rect 24327 94 24351 150
rect 24407 94 24431 150
rect 24487 94 26079 150
rect 26135 94 26159 150
rect 26215 94 26239 150
rect 26295 94 26319 150
rect 26375 94 27967 150
rect 28023 94 28047 150
rect 28103 94 28127 150
rect 28183 94 28207 150
rect 28263 94 29855 150
rect 29911 94 29935 150
rect 29991 94 30015 150
rect 30071 94 30095 150
rect 30151 94 30383 150
rect 21679 61 30383 94
rect 13879 48 30383 61
rect 30470 48 30506 160
rect 30593 48 30638 160
rect 30725 157 46038 160
rect 30725 150 36412 157
rect 30725 94 31743 150
rect 31799 94 31823 150
rect 31879 94 31903 150
rect 31959 94 31983 150
rect 32039 94 33631 150
rect 33687 94 33711 150
rect 33767 94 33791 150
rect 33847 94 33871 150
rect 33927 94 35519 150
rect 35575 94 35599 150
rect 35655 94 35679 150
rect 35735 94 35759 150
rect 35815 94 36412 150
rect 30725 48 36412 94
rect 13879 45 36412 48
rect 36499 45 36581 157
rect 36668 150 46038 157
rect 36668 94 37407 150
rect 37463 94 37487 150
rect 37543 94 37567 150
rect 37623 94 37647 150
rect 37703 94 39295 150
rect 39351 94 39375 150
rect 39431 94 39455 150
rect 39511 94 39535 150
rect 39591 94 41183 150
rect 41239 94 41263 150
rect 41319 94 41343 150
rect 41399 94 41423 150
rect 41479 94 43071 150
rect 43127 94 43151 150
rect 43207 94 43231 150
rect 43287 94 43311 150
rect 43367 94 44959 150
rect 45015 94 45039 150
rect 45095 94 45119 150
rect 45175 94 45199 150
rect 45255 94 46038 150
rect 36668 45 46038 94
rect 13879 32 46038 45
rect 46122 32 46151 190
rect 46235 32 46266 190
rect 46350 150 53361 190
rect 46350 94 46841 150
rect 46897 94 46921 150
rect 46977 94 47001 150
rect 47057 94 47081 150
rect 47137 94 48729 150
rect 48785 94 48809 150
rect 48865 94 48889 150
rect 48945 94 48969 150
rect 49025 94 50617 150
rect 50673 94 50697 150
rect 50753 94 50777 150
rect 50833 94 50857 150
rect 50913 94 52505 150
rect 52561 94 52585 150
rect 52641 94 52665 150
rect 52721 94 52745 150
rect 52801 94 53361 150
rect 46350 42 53361 94
rect 53445 42 53480 200
rect 53564 42 53609 200
rect 53693 150 60412 200
rect 53693 94 54393 150
rect 54449 94 54473 150
rect 54529 94 54553 150
rect 54609 94 54633 150
rect 54689 94 56281 150
rect 56337 94 56361 150
rect 56417 94 56441 150
rect 56497 94 56521 150
rect 56577 94 58169 150
rect 58225 94 58249 150
rect 58305 94 58329 150
rect 58385 94 58409 150
rect 58465 94 60057 150
rect 60113 94 60137 150
rect 60193 94 60217 150
rect 60273 94 60297 150
rect 60353 94 60412 150
rect 53693 42 60412 94
rect 46350 32 60412 42
rect 13879 21 60412 32
rect 8 0 60412 21
rect 8 -1 13224 0
rect 15106 -1 28322 0
rect 30210 -1 43426 0
rect 45308 -1 58524 0
<< via3 >>
rect 2518 7211 2624 7389
rect 2727 7210 2833 7388
rect 2893 7210 2999 7388
rect 3073 7212 3179 7390
rect 1284 5093 1390 5271
rect 1456 5222 1562 5272
rect 1630 5222 1736 5271
rect 1456 5166 1517 5222
rect 1517 5166 1562 5222
rect 1630 5166 1653 5222
rect 1653 5166 1677 5222
rect 1677 5166 1733 5222
rect 1733 5166 1736 5222
rect 1456 5094 1562 5166
rect 1630 5093 1736 5166
rect 36414 3487 36457 3532
rect 36457 3487 36495 3532
rect 36495 3487 36501 3532
rect 36568 3487 36589 3533
rect 36589 3487 36645 3533
rect 36645 3487 36655 3533
rect 36414 3455 36501 3487
rect 36568 3455 36655 3487
rect 36414 3420 36457 3455
rect 36457 3420 36495 3455
rect 36495 3420 36501 3455
rect 36568 3421 36589 3455
rect 36589 3421 36645 3455
rect 36645 3421 36655 3455
rect 6272 3201 6275 3229
rect 6275 3201 6331 3229
rect 6331 3201 6358 3229
rect 6423 3201 6445 3235
rect 6445 3201 6503 3235
rect 6503 3201 6509 3235
rect 6272 3142 6358 3201
rect 6423 3144 6509 3201
rect 6568 3144 6654 3235
rect 6272 3138 6275 3142
rect 6275 3138 6331 3142
rect 6331 3138 6358 3142
rect 21312 3226 21314 3239
rect 21314 3226 21370 3239
rect 21370 3226 21405 3239
rect 21479 3226 21522 3239
rect 21522 3226 21572 3239
rect 21312 3166 21405 3226
rect 21479 3166 21572 3226
rect 21312 3155 21314 3166
rect 21314 3155 21370 3166
rect 21370 3155 21405 3166
rect 21479 3155 21522 3166
rect 21522 3155 21572 3166
rect 21312 3050 21405 3078
rect 21479 3050 21572 3078
rect 21312 2994 21314 3050
rect 21314 2994 21370 3050
rect 21370 2994 21405 3050
rect 21479 2994 21522 3050
rect 21522 2994 21572 3050
rect 53355 3176 53439 3183
rect 53476 3176 53560 3183
rect 53614 3176 53698 3183
rect 53355 3120 53404 3176
rect 53404 3120 53439 3176
rect 53476 3120 53508 3176
rect 53508 3120 53556 3176
rect 53556 3120 53560 3176
rect 53614 3120 53660 3176
rect 53660 3120 53698 3176
rect 53355 3086 53439 3120
rect 53476 3086 53560 3120
rect 53614 3086 53698 3120
rect 53355 3030 53404 3086
rect 53404 3030 53439 3086
rect 53476 3030 53508 3086
rect 53508 3030 53556 3086
rect 53556 3030 53560 3086
rect 53614 3030 53660 3086
rect 53660 3030 53698 3086
rect 53355 3025 53439 3030
rect 53476 3025 53560 3030
rect 53614 3025 53698 3030
rect 13653 2755 13669 2763
rect 13669 2755 13725 2763
rect 13725 2755 13730 2763
rect 13653 2717 13730 2755
rect 13653 2694 13669 2717
rect 13669 2694 13725 2717
rect 13725 2694 13730 2717
rect 13756 2755 13777 2763
rect 13777 2755 13833 2763
rect 13756 2717 13833 2755
rect 13756 2694 13777 2717
rect 13777 2694 13833 2717
rect 13859 2755 13885 2763
rect 13885 2755 13936 2763
rect 13859 2717 13936 2755
rect 30362 2875 30364 2892
rect 30364 2875 30420 2892
rect 30420 2875 30449 2892
rect 30362 2835 30449 2875
rect 30362 2780 30364 2835
rect 30364 2780 30420 2835
rect 30420 2780 30449 2835
rect 30481 2875 30489 2892
rect 30489 2875 30545 2892
rect 30545 2875 30568 2892
rect 30481 2835 30568 2875
rect 30481 2780 30489 2835
rect 30489 2780 30545 2835
rect 30545 2780 30568 2835
rect 30600 2875 30614 2892
rect 30614 2875 30670 2892
rect 30670 2875 30687 2892
rect 30600 2835 30687 2875
rect 30600 2780 30614 2835
rect 30614 2780 30670 2835
rect 30670 2780 30687 2835
rect 46036 2784 46120 2807
rect 46176 2784 46260 2808
rect 46304 2784 46388 2808
rect 13859 2694 13885 2717
rect 13885 2694 13936 2717
rect 46036 2728 46091 2784
rect 46091 2728 46120 2784
rect 46176 2728 46184 2784
rect 46184 2728 46221 2784
rect 46221 2728 46260 2784
rect 46304 2728 46314 2784
rect 46314 2728 46370 2784
rect 46370 2728 46388 2784
rect 46036 2702 46120 2728
rect 46176 2702 46260 2728
rect 46304 2702 46388 2728
rect 46036 2649 46091 2702
rect 46091 2649 46120 2702
rect 46176 2650 46184 2702
rect 46184 2650 46221 2702
rect 46221 2650 46260 2702
rect 46304 2650 46314 2702
rect 46314 2650 46370 2702
rect 46370 2650 46388 2702
rect 1286 2145 1392 2323
rect 1491 2274 1597 2325
rect 1690 2274 1796 2325
rect 1491 2218 1541 2274
rect 1541 2218 1597 2274
rect 1690 2218 1701 2274
rect 1701 2218 1757 2274
rect 1757 2218 1781 2274
rect 1781 2218 1796 2274
rect 1491 2147 1597 2218
rect 1690 2147 1796 2218
rect 2532 34 2638 212
rect 2753 34 2859 212
rect 2962 34 3068 212
rect 3136 34 3242 212
rect 6260 66 6346 157
rect 6408 66 6494 157
rect 6556 66 6642 157
rect 13779 140 13856 209
rect 13802 21 13879 90
rect 21317 61 21413 169
rect 21450 61 21546 169
rect 21583 61 21679 169
rect 30383 48 30470 160
rect 30506 48 30593 160
rect 30638 48 30725 160
rect 36412 45 36499 157
rect 36581 45 36668 157
rect 46038 32 46122 190
rect 46151 32 46235 190
rect 46266 32 46350 190
rect 53361 42 53445 200
rect 53480 42 53564 200
rect 53609 42 53693 200
<< metal4 >>
rect 2467 7390 3251 7443
rect 2467 7389 3073 7390
rect 2467 7211 2518 7389
rect 2624 7388 3073 7389
rect 2624 7211 2727 7388
rect 2467 7210 2727 7211
rect 2833 7210 2893 7388
rect 2999 7212 3073 7388
rect 3179 7212 3251 7390
rect 2999 7210 3251 7212
rect 1234 5272 1852 5401
rect 1234 5271 1456 5272
rect 1234 5093 1284 5271
rect 1390 5094 1456 5271
rect 1562 5271 1852 5272
rect 1562 5094 1630 5271
rect 1390 5093 1630 5094
rect 1736 5093 1852 5271
rect 1234 2325 1852 5093
rect 1234 2323 1491 2325
rect 1234 2145 1286 2323
rect 1392 2147 1491 2323
rect 1597 2147 1690 2325
rect 1796 2147 1852 2325
rect 1392 2145 1852 2147
rect 1234 2095 1852 2145
rect 2467 212 3251 7210
rect 36378 3533 36683 3690
rect 36378 3532 36568 3533
rect 36378 3420 36414 3532
rect 36501 3421 36568 3532
rect 36655 3421 36683 3533
rect 36501 3420 36683 3421
rect 2467 34 2532 212
rect 2638 34 2753 212
rect 2859 34 2962 212
rect 3068 34 3136 212
rect 3242 34 3251 212
rect 2467 -55 3251 34
rect 6214 3235 6683 3350
rect 6214 3229 6423 3235
rect 6214 3138 6272 3229
rect 6358 3144 6423 3229
rect 6509 3144 6568 3235
rect 6654 3144 6683 3235
rect 6358 3138 6683 3144
rect 6214 157 6683 3138
rect 21264 3239 21731 3364
rect 21264 3155 21312 3239
rect 21405 3155 21479 3239
rect 21572 3155 21731 3239
rect 21264 3078 21731 3155
rect 21264 2994 21312 3078
rect 21405 2994 21479 3078
rect 21572 2994 21731 3078
rect 13629 2763 13983 2835
rect 13629 2694 13653 2763
rect 13730 2694 13756 2763
rect 13833 2694 13859 2763
rect 13936 2694 13983 2763
rect 13629 2634 13983 2694
rect 6214 66 6260 157
rect 6346 66 6408 157
rect 6494 66 6556 157
rect 6642 66 6683 157
rect 6214 -33 6683 66
rect 13705 209 13906 2634
rect 13705 140 13779 209
rect 13856 140 13906 209
rect 13705 90 13906 140
rect 13705 21 13802 90
rect 13879 21 13906 90
rect 13705 -58 13906 21
rect 21264 169 21731 2994
rect 21264 61 21317 169
rect 21413 61 21450 169
rect 21546 61 21583 169
rect 21679 61 21731 169
rect 21264 -8 21731 61
rect 30316 2892 30741 2971
rect 30316 2780 30362 2892
rect 30449 2780 30481 2892
rect 30568 2780 30600 2892
rect 30687 2780 30741 2892
rect 30316 160 30741 2780
rect 30316 48 30383 160
rect 30470 48 30506 160
rect 30593 48 30638 160
rect 30725 48 30741 160
rect 30316 6 30741 48
rect 36378 157 36683 3420
rect 53311 3183 53736 3206
rect 53311 3025 53355 3183
rect 53439 3025 53476 3183
rect 53560 3025 53614 3183
rect 53698 3025 53736 3183
rect 36378 45 36412 157
rect 36499 45 36581 157
rect 36668 45 36683 157
rect 36378 -3 36683 45
rect 45998 2808 46412 2897
rect 45998 2807 46176 2808
rect 45998 2649 46036 2807
rect 46120 2650 46176 2807
rect 46260 2650 46304 2808
rect 46388 2650 46412 2808
rect 46120 2649 46412 2650
rect 45998 190 46412 2649
rect 45998 32 46038 190
rect 46122 32 46151 190
rect 46235 32 46266 190
rect 46350 32 46412 190
rect 45998 -56 46412 32
rect 53311 200 53736 3025
rect 53311 42 53361 200
rect 53445 42 53480 200
rect 53564 42 53609 200
rect 53693 42 53736 200
rect 53311 -44 53736 42
<< labels >>
flabel metal4 1234 2325 1852 5093 1 FreeSans 1600 0 0 0 VDD
port 1 n
flabel metal4 2467 212 3251 7210 1 FreeSans 1600 0 0 0 VSS
port 2 n
flabel locali 29711 3786 30067 3836 1 FreeSans 1600 0 0 0 RESET
port 68 n
flabel metal1 60382 780 60604 858 1 FreeSans 1600 0 0 0 OUT
port 3 n
flabel metal2 59918 6648 59962 7270 1 FreeSans 800 0 0 0 C[0]
port 67 n
flabel metal2 58030 6648 58074 7270 1 FreeSans 800 0 0 0 C[1]
port 66 n
flabel metal2 56142 6648 56186 7270 1 FreeSans 800 0 0 0 C[2]
port 65 n
flabel metal2 54254 6648 54298 7270 1 FreeSans 800 0 0 0 C[3]
port 64 n
flabel metal2 52366 6648 52410 7270 1 FreeSans 800 0 0 0 C[4]
port 63 n
flabel metal2 50478 6648 50522 7270 1 FreeSans 800 0 0 0 C[5]
port 62 n
flabel metal2 48590 6648 48634 7270 1 FreeSans 800 0 0 0 C[6]
port 61 n
flabel metal2 46702 6648 46746 7270 1 FreeSans 800 0 0 0 C[7]
port 60 n
flabel metal2 44814 6648 44858 7270 1 FreeSans 800 0 0 0 C[8]
port 59 n
flabel metal2 42926 6648 42970 7270 1 FreeSans 800 0 0 0 C[9]
port 58 n
flabel metal2 41038 6648 41082 7270 1 FreeSans 800 0 0 0 C[10]
port 57 n
flabel metal2 39150 6648 39194 7270 1 FreeSans 800 0 0 0 C[11]
port 56 n
flabel metal2 37262 6648 37306 7270 1 FreeSans 800 0 0 0 C[12]
port 55 n
flabel metal2 35374 6648 35418 7270 1 FreeSans 800 0 0 0 C[13]
port 54 n
flabel metal2 33486 6648 33530 7270 1 FreeSans 800 0 0 0 C[14]
port 53 n
flabel metal2 31598 6648 31642 7270 1 FreeSans 800 0 0 0 C[15]
port 52 n
flabel metal2 29710 6648 29754 7270 1 FreeSans 800 0 0 0 C[16]
port 51 n
flabel metal2 27822 6648 27866 7270 1 FreeSans 800 0 0 0 C[17]
port 50 n
flabel metal2 25934 6648 25978 7270 1 FreeSans 800 0 0 0 C[18]
port 49 n
flabel metal2 24046 6648 24090 7270 1 FreeSans 800 0 0 0 C[19]
port 48 n
flabel metal2 22158 6648 22202 7270 1 FreeSans 800 0 0 0 C[20]
port 47 n
flabel metal2 20270 6648 20314 7270 1 FreeSans 800 0 0 0 C[21]
port 46 n
flabel metal2 18382 6648 18426 7270 1 FreeSans 800 0 0 0 C[22]
port 45 n
flabel metal2 16494 6648 16538 7270 1 FreeSans 800 0 0 0 C[23]
port 44 n
flabel metal2 14606 6648 14650 7270 1 FreeSans 800 0 0 0 C[24]
port 43 n
flabel metal2 12718 6648 12762 7270 1 FreeSans 800 0 0 0 C[25]
port 42 n
flabel metal2 10830 6648 10874 7270 1 FreeSans 800 0 0 0 C[26]
port 41 n
flabel metal2 8942 6648 8986 7270 1 FreeSans 800 0 0 0 C[27]
port 40 n
flabel metal2 7054 6648 7098 7270 1 FreeSans 800 0 0 0 C[28]
port 39 n
flabel metal2 5166 6648 5210 7270 1 FreeSans 800 0 0 0 C[29]
port 38 n
flabel metal2 3278 6648 3322 7270 1 FreeSans 800 0 0 0 C[30]
port 37 n
flabel metal2 1390 6648 1434 7270 1 FreeSans 800 0 0 0 C[31]
port 36 n
flabel metal2 20 170 64 792 1 FreeSans 800 0 0 0 C[32]
port 35 n
flabel metal2 1908 170 1952 792 1 FreeSans 800 0 0 0 C[33]
port 34 n
flabel metal2 3796 170 3840 792 1 FreeSans 800 0 0 0 C[34]
port 33 n
flabel metal2 5684 170 5728 792 1 FreeSans 800 0 0 0 C[35]
port 32 n
flabel metal2 7572 170 7616 792 1 FreeSans 800 0 0 0 C[36]
port 31 n
flabel metal2 9460 170 9504 792 1 FreeSans 800 0 0 0 C[37]
port 30 n
flabel metal2 11348 170 11392 792 1 FreeSans 800 0 0 0 C[38]
port 29 n
flabel metal2 13236 170 13280 792 1 FreeSans 800 0 0 0 C[39]
port 28 n
flabel metal2 15124 170 15168 792 1 FreeSans 800 0 0 0 C[40]
port 27 n
flabel metal2 17012 170 17056 792 1 FreeSans 800 0 0 0 C[41]
port 26 n
flabel metal2 18900 170 18944 792 1 FreeSans 800 0 0 0 C[42]
port 25 n
flabel metal2 20788 170 20832 792 1 FreeSans 800 0 0 0 C[43]
port 24 n
flabel metal2 22676 170 22720 792 1 FreeSans 800 0 0 0 C[44]
port 23 n
flabel metal2 24564 170 24608 792 1 FreeSans 800 0 0 0 C[45]
port 22 n
flabel metal2 26452 170 26496 792 1 FreeSans 800 0 0 0 C[46]
port 21 n
flabel metal2 28340 170 28384 792 1 FreeSans 800 0 0 0 C[47]
port 20 n
flabel metal2 30228 170 30272 792 1 FreeSans 800 0 0 0 C[48]
port 19 n
flabel metal2 32116 170 32160 792 1 FreeSans 800 0 0 0 C[49]
port 18 n
flabel metal2 34004 170 34048 792 1 FreeSans 800 0 0 0 C[50]
port 17 n
flabel metal2 35892 170 35936 792 1 FreeSans 800 0 0 0 C[51]
port 16 n
flabel metal2 37780 170 37824 792 1 FreeSans 800 0 0 0 C[52]
port 15 n
flabel metal2 39668 170 39712 792 1 FreeSans 800 0 0 0 C[53]
port 14 n
flabel metal2 41556 170 41600 792 1 FreeSans 800 0 0 0 C[54]
port 13 n
flabel metal2 43444 170 43488 792 1 FreeSans 800 0 0 0 C[55]
port 12 n
flabel metal2 45332 170 45376 792 1 FreeSans 800 0 0 0 C[56]
port 11 n
flabel metal2 47220 170 47264 792 1 FreeSans 800 0 0 0 C[57]
port 10 n
flabel metal2 49108 170 49152 792 1 FreeSans 800 0 0 0 C[58]
port 9 n
flabel metal2 50996 170 51040 792 1 FreeSans 800 0 0 0 C[59]
port 8 n
flabel metal2 52884 170 52928 792 1 FreeSans 800 0 0 0 C[60]
port 7 n
flabel metal2 54772 170 54816 792 1 FreeSans 800 0 0 0 C[61]
port 6 n
flabel metal2 56660 170 56704 792 1 FreeSans 800 0 0 0 C[62]
port 5 n
flabel metal2 58548 170 58592 792 1 FreeSans 800 0 0 0 C[63]
port 4 n
flabel locali 30424 3724 30458 3758 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 30424 3792 30458 3826 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 30424 3860 30458 3894 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/Y
flabel locali 30056 3792 30090 3826 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali 30148 3792 30182 3826 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali 30240 3792 30274 3826 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel locali 30332 3792 30366 3826 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0/A
flabel nwell 30056 4098 30090 4132 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VPB
flabel pwell 30056 3554 30090 3588 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VNB
flabel metal1 30056 4098 30090 4132 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VPWR
flabel metal1 30056 3554 30090 3588 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0/VGND
rlabel comment 30027 3571 30027 3571 4 sky130_fd_sc_hd__inv_4_0/inv_4
<< end >>
