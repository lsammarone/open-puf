magic
tech sky130B
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_0
timestamp 1648127584
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_1
timestamp 1648127584
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_2
timestamp 1648127584
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_3
timestamp 1648127584
transform 1 0 648 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_4
timestamp 1648127584
transform 1 0 824 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_5
timestamp 1648127584
transform 1 0 1000 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_6
timestamp 1648127584
transform 1 0 1176 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_7
timestamp 1648127584
transform 1 0 1352 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_8
timestamp 1648127584
transform 1 0 1528 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_9
timestamp 1648127584
transform 1 0 1704 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_10
timestamp 1648127584
transform 1 0 1880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_11
timestamp 1648127584
transform 1 0 2056 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_12
timestamp 1648127584
transform 1 0 2232 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_13
timestamp 1648127584
transform 1 0 2408 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_14
timestamp 1648127584
transform 1 0 2584 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_15
timestamp 1648127584
transform 1 0 2760 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808370  sky130_fd_pr__hvdfl1sd__example_55959141808370_0
timestamp 1648127584
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 2788 63 2788 63 0 FreeSans 300 0 0 0 S
flabel comment s 2612 63 2612 63 0 FreeSans 300 0 0 0 D
flabel comment s 2436 63 2436 63 0 FreeSans 300 0 0 0 S
flabel comment s 2260 63 2260 63 0 FreeSans 300 0 0 0 D
flabel comment s 2084 63 2084 63 0 FreeSans 300 0 0 0 S
flabel comment s 1908 63 1908 63 0 FreeSans 300 0 0 0 D
flabel comment s 1732 63 1732 63 0 FreeSans 300 0 0 0 S
flabel comment s 1556 63 1556 63 0 FreeSans 300 0 0 0 D
flabel comment s 1380 63 1380 63 0 FreeSans 300 0 0 0 S
flabel comment s 1204 63 1204 63 0 FreeSans 300 0 0 0 D
flabel comment s 1028 63 1028 63 0 FreeSans 300 0 0 0 S
flabel comment s 852 63 852 63 0 FreeSans 300 0 0 0 D
flabel comment s 676 63 676 63 0 FreeSans 300 0 0 0 S
flabel comment s 500 63 500 63 0 FreeSans 300 0 0 0 D
flabel comment s 324 63 324 63 0 FreeSans 300 0 0 0 S
flabel comment s 148 63 148 63 0 FreeSans 300 0 0 0 D
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 35724170
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35714384
<< end >>
