magic
tech sky130A
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__dfl1sd2__example_55959141808515  sky130_fd_pr__dfl1sd2__example_55959141808515_0
timestamp 1648127584
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808515  sky130_fd_pr__dfl1sd2__example_55959141808515_1
timestamp 1648127584
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808515  sky130_fd_pr__dfl1sd2__example_55959141808515_2
timestamp 1648127584
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808340  sky130_fd_pr__dfl1sd__example_55959141808340_0
timestamp 1648127584
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808340  sky130_fd_pr__dfl1sd__example_55959141808340_1
timestamp 1648127584
transform 1 0 568 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 596 981 596 981 0 FreeSans 300 0 0 0 S
flabel comment s 440 981 440 981 0 FreeSans 300 0 0 0 D
flabel comment s 284 981 284 981 0 FreeSans 300 0 0 0 S
flabel comment s 128 981 128 981 0 FreeSans 300 0 0 0 D
flabel comment s -28 981 -28 981 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 47734064
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47731466
<< end >>
