magic
tech sky130A
magscale 1 2
timestamp 1654402208
<< nwell >>
rect 8774 6644 9298 6822
<< pwell >>
rect 3212 6750 3442 6868
rect 18250 6754 18478 6880
<< psubdiff >>
rect 3238 6826 3416 6842
rect 3238 6792 3276 6826
rect 3310 6792 3344 6826
rect 3378 6792 3416 6826
rect 3238 6776 3416 6792
rect 18276 6834 18452 6854
rect 18276 6800 18313 6834
rect 18347 6800 18381 6834
rect 18415 6800 18452 6834
rect 18276 6780 18452 6800
<< nsubdiff >>
rect 8866 6739 9074 6756
rect 8866 6705 8919 6739
rect 8953 6705 8987 6739
rect 9021 6705 9074 6739
rect 8866 6688 9074 6705
<< psubdiffcont >>
rect 3276 6792 3310 6826
rect 3344 6792 3378 6826
rect 18313 6800 18347 6834
rect 18381 6800 18415 6834
<< nsubdiffcont >>
rect 8919 6705 8953 6739
rect 8987 6705 9021 6739
<< locali >>
rect 3110 6826 3408 6842
rect 3110 6792 3276 6826
rect 3310 6792 3344 6826
rect 3378 6792 3408 6826
rect 3110 6776 3408 6792
rect 18284 6834 18444 6854
rect 18284 6800 18313 6834
rect 18347 6800 18381 6834
rect 18415 6800 18444 6834
rect 18284 6780 18444 6800
rect 8874 6739 9066 6756
rect 8874 6705 8919 6739
rect 8953 6705 8987 6739
rect 9021 6705 9066 6739
rect 8874 6660 9066 6705
rect 8944 6444 8982 6448
rect 8944 6410 8946 6444
rect 8980 6410 8982 6444
rect 8944 6406 8982 6410
rect 10300 6357 10346 6360
rect 10300 6323 10306 6357
rect 10340 6323 10346 6357
rect 10300 6320 10346 6323
rect 12826 6350 12864 6354
rect 12826 6316 12828 6350
rect 12862 6316 12864 6350
rect 12826 6312 12864 6316
<< viali >>
rect 8946 6410 8980 6444
rect 10306 6323 10340 6357
rect 12828 6316 12862 6350
<< metal1 >>
rect 16594 6954 16654 6956
rect 3458 6952 3543 6954
rect 3458 6906 5188 6952
rect 3016 6506 3762 6744
rect 3016 6390 3170 6506
rect 3478 6390 3762 6506
rect 3016 5974 3762 6390
rect 5128 6392 5188 6906
rect 16594 6908 18335 6954
rect 8852 6672 9096 6690
rect 8852 6620 8884 6672
rect 8936 6620 8948 6672
rect 9000 6620 9012 6672
rect 9064 6620 9096 6672
rect 8852 6602 9096 6620
rect 12618 6684 12862 6692
rect 12618 6674 12886 6684
rect 12618 6622 12650 6674
rect 12702 6622 12714 6674
rect 12766 6622 12778 6674
rect 12830 6622 12886 6674
rect 12618 6612 12886 6622
rect 12618 6604 12862 6612
rect 12898 6598 13098 6694
rect 8938 6444 8994 6460
rect 8938 6410 8946 6444
rect 8980 6410 8994 6444
rect 8938 6392 8994 6410
rect 5128 6332 8994 6392
rect 10284 6366 10358 6376
rect 16594 6366 16654 6908
rect 5128 5812 5188 6332
rect 10284 6314 10296 6366
rect 10348 6314 10358 6366
rect 10284 6308 10358 6314
rect 12816 6350 16654 6366
rect 12816 6316 12828 6350
rect 12862 6316 16654 6350
rect 12816 6306 16654 6316
rect 12820 6300 12870 6306
rect 10716 6130 11000 6148
rect 10716 6078 10736 6130
rect 10788 6078 10800 6130
rect 10852 6078 10864 6130
rect 10916 6078 10928 6130
rect 10980 6078 11000 6130
rect 10716 6060 11000 6078
rect 12904 6054 13104 6150
rect 3217 5766 5188 5812
rect 16594 5814 16654 6306
rect 18108 6548 18848 6744
rect 18108 6432 18258 6548
rect 18566 6432 18848 6548
rect 18108 5980 18848 6432
rect 16594 5768 18445 5814
rect 26100 4032 26132 4062
<< via1 >>
rect 3170 6390 3478 6506
rect 8884 6620 8936 6672
rect 8948 6620 9000 6672
rect 9012 6620 9064 6672
rect 12650 6622 12702 6674
rect 12714 6622 12766 6674
rect 12778 6622 12830 6674
rect 10296 6357 10348 6366
rect 10296 6323 10306 6357
rect 10306 6323 10340 6357
rect 10340 6323 10348 6357
rect 10296 6314 10348 6323
rect 10736 6078 10788 6130
rect 10800 6078 10852 6130
rect 10864 6078 10916 6130
rect 10928 6078 10980 6130
rect 18258 6432 18566 6548
<< metal2 >>
rect -2574 9408 -2540 9468
rect -682 9384 -648 9444
rect 1204 9406 1238 9466
rect 3094 9396 3128 9456
rect 4980 9402 5014 9462
rect 6866 9392 6900 9452
rect 8758 9406 8792 9466
rect 10646 9402 10680 9462
rect 12526 9398 12560 9458
rect 14412 9392 14446 9452
rect 16300 9398 16334 9458
rect 18188 9392 18222 9452
rect 20082 9386 20116 9446
rect 21964 9386 21998 9446
rect 23854 9392 23888 9452
rect -6146 7978 -4356 8014
rect 23862 7978 26352 8014
rect -6146 4742 -6110 7978
rect 8862 6674 9086 6700
rect 8862 6618 8866 6674
rect 8922 6672 8946 6674
rect 9002 6672 9026 6674
rect 8936 6620 8946 6672
rect 9002 6620 9012 6672
rect 8922 6618 8946 6620
rect 9002 6618 9026 6620
rect 9082 6618 9086 6674
rect 8862 6592 9086 6618
rect 12628 6676 12852 6702
rect 12628 6620 12632 6676
rect 12688 6674 12712 6676
rect 12768 6674 12792 6676
rect 12702 6622 12712 6674
rect 12768 6622 12778 6674
rect 12688 6620 12712 6622
rect 12768 6620 12792 6622
rect 12848 6620 12852 6676
rect 12628 6594 12852 6620
rect 18258 6548 18566 6558
rect 3170 6506 3478 6516
rect 18258 6422 18566 6432
rect 3170 6380 3478 6390
rect 10290 6366 10354 6376
rect 10290 6334 10296 6366
rect -6072 6314 10296 6334
rect 10348 6314 10354 6366
rect -6072 6302 10354 6314
rect 10726 6132 10990 6158
rect 10726 6130 10750 6132
rect 10806 6130 10830 6132
rect 10886 6130 10910 6132
rect 10966 6130 10990 6132
rect 10726 6078 10736 6130
rect 10980 6078 10990 6130
rect 10726 6076 10750 6078
rect 10806 6076 10830 6078
rect 10886 6076 10910 6078
rect 10966 6076 10990 6078
rect 10726 6050 10990 6076
rect -5702 5786 -4676 5787
rect -3812 5786 -2786 5787
rect -5922 5598 -1960 5786
rect -5702 5341 -4676 5598
rect -3812 5341 -2786 5598
rect -5922 5232 -2039 5341
rect 26316 4742 26352 7978
rect -6146 4706 -5878 4742
rect 26102 4706 26354 4742
rect -5896 3240 -5862 3300
rect -4008 3240 -3974 3300
rect -2122 3240 -2088 3300
rect -232 3248 -198 3308
rect 1654 3246 1688 3306
rect 3546 3242 3580 3302
rect 5432 3246 5466 3306
rect 7322 3246 7356 3306
rect 9206 3246 9240 3306
rect 11088 3250 11122 3310
rect 12978 3250 13012 3310
rect 14866 3246 14900 3306
rect 16756 3246 16790 3306
rect 18640 3246 18674 3306
rect 20532 3254 20566 3314
rect 22418 3246 22452 3306
rect 24306 3244 24340 3304
<< via2 >>
rect 8866 6672 8922 6674
rect 8946 6672 9002 6674
rect 9026 6672 9082 6674
rect 8866 6620 8884 6672
rect 8884 6620 8922 6672
rect 8946 6620 8948 6672
rect 8948 6620 9000 6672
rect 9000 6620 9002 6672
rect 9026 6620 9064 6672
rect 9064 6620 9082 6672
rect 8866 6618 8922 6620
rect 8946 6618 9002 6620
rect 9026 6618 9082 6620
rect 12632 6674 12688 6676
rect 12712 6674 12768 6676
rect 12792 6674 12848 6676
rect 12632 6622 12650 6674
rect 12650 6622 12688 6674
rect 12712 6622 12714 6674
rect 12714 6622 12766 6674
rect 12766 6622 12768 6674
rect 12792 6622 12830 6674
rect 12830 6622 12848 6674
rect 12632 6620 12688 6622
rect 12712 6620 12768 6622
rect 12792 6620 12848 6622
rect 3176 6420 3232 6476
rect 3256 6420 3312 6476
rect 3336 6420 3392 6476
rect 3416 6420 3472 6476
rect 18264 6462 18320 6518
rect 18344 6462 18400 6518
rect 18424 6462 18480 6518
rect 18504 6462 18560 6518
rect 10750 6130 10806 6132
rect 10830 6130 10886 6132
rect 10910 6130 10966 6132
rect 10750 6078 10788 6130
rect 10788 6078 10800 6130
rect 10800 6078 10806 6130
rect 10830 6078 10852 6130
rect 10852 6078 10864 6130
rect 10864 6078 10886 6130
rect 10910 6078 10916 6130
rect 10916 6078 10928 6130
rect 10928 6078 10966 6130
rect 10750 6076 10806 6078
rect 10830 6076 10886 6078
rect 10910 6076 10966 6078
<< metal3 >>
rect -4367 9398 -4039 9424
rect -4367 9334 -4355 9398
rect -4291 9334 -4275 9398
rect -4211 9334 -4195 9398
rect -4131 9334 -4115 9398
rect -4051 9334 -4039 9398
rect -4367 9308 -4039 9334
rect -591 9398 -263 9424
rect -591 9334 -579 9398
rect -515 9334 -499 9398
rect -435 9334 -419 9398
rect -355 9334 -339 9398
rect -275 9334 -263 9398
rect -591 9308 -263 9334
rect 3185 9398 3513 9424
rect 3185 9334 3197 9398
rect 3261 9334 3277 9398
rect 3341 9334 3357 9398
rect 3421 9334 3437 9398
rect 3501 9334 3513 9398
rect 3185 9308 3513 9334
rect 6961 9398 7289 9424
rect 6961 9334 6973 9398
rect 7037 9334 7053 9398
rect 7117 9334 7133 9398
rect 7197 9334 7213 9398
rect 7277 9334 7289 9398
rect 6961 9308 7289 9334
rect 10731 9398 11059 9424
rect 10731 9334 10743 9398
rect 10807 9334 10823 9398
rect 10887 9334 10903 9398
rect 10967 9334 10983 9398
rect 11047 9334 11059 9398
rect 10731 9308 11059 9334
rect 14507 9398 14835 9424
rect 14507 9334 14519 9398
rect 14583 9334 14599 9398
rect 14663 9334 14679 9398
rect 14743 9334 14759 9398
rect 14823 9334 14835 9398
rect 14507 9308 14835 9334
rect 18283 9398 18611 9424
rect 18283 9334 18295 9398
rect 18359 9334 18375 9398
rect 18439 9334 18455 9398
rect 18519 9334 18535 9398
rect 18599 9334 18611 9398
rect 18283 9308 18611 9334
rect 22059 9398 22387 9424
rect 22059 9334 22071 9398
rect 22135 9334 22151 9398
rect 22215 9334 22231 9398
rect 22295 9334 22311 9398
rect 22375 9334 22387 9398
rect 22059 9308 22387 9334
rect -2479 7274 -2151 7300
rect -2479 7210 -2467 7274
rect -2403 7210 -2387 7274
rect -2323 7210 -2307 7274
rect -2243 7210 -2227 7274
rect -2163 7210 -2151 7274
rect -2479 7184 -2151 7210
rect 1297 7274 1625 7300
rect 1297 7210 1309 7274
rect 1373 7210 1389 7274
rect 1453 7210 1469 7274
rect 1533 7210 1549 7274
rect 1613 7210 1625 7274
rect 1297 7184 1625 7210
rect 5073 7274 5401 7300
rect 5073 7210 5085 7274
rect 5149 7210 5165 7274
rect 5229 7210 5245 7274
rect 5309 7210 5325 7274
rect 5389 7210 5401 7274
rect 5073 7184 5401 7210
rect 8849 7274 9177 7300
rect 8849 7210 8861 7274
rect 8925 7210 8941 7274
rect 9005 7210 9021 7274
rect 9085 7210 9101 7274
rect 9165 7210 9177 7274
rect 8849 7184 9177 7210
rect 12619 7274 12947 7300
rect 12619 7210 12631 7274
rect 12695 7210 12711 7274
rect 12775 7210 12791 7274
rect 12855 7210 12871 7274
rect 12935 7210 12947 7274
rect 12619 7184 12947 7210
rect 16395 7274 16723 7300
rect 16395 7210 16407 7274
rect 16471 7210 16487 7274
rect 16551 7210 16567 7274
rect 16631 7210 16647 7274
rect 16711 7210 16723 7274
rect 16395 7184 16723 7210
rect 20171 7274 20499 7300
rect 20171 7210 20183 7274
rect 20247 7210 20263 7274
rect 20327 7210 20343 7274
rect 20407 7210 20423 7274
rect 20487 7210 20499 7274
rect 20171 7184 20499 7210
rect 8852 6678 9096 6695
rect 8852 6614 8862 6678
rect 8926 6614 8942 6678
rect 9006 6614 9022 6678
rect 9086 6614 9096 6678
rect 8852 6597 9096 6614
rect 12618 6680 12862 6697
rect 12618 6616 12628 6680
rect 12692 6616 12708 6680
rect 12772 6616 12788 6680
rect 12852 6616 12862 6680
rect 12618 6599 12862 6616
rect 18248 6522 18576 6553
rect 3160 6480 3488 6511
rect 3160 6416 3172 6480
rect 3236 6416 3252 6480
rect 3316 6416 3332 6480
rect 3396 6416 3412 6480
rect 3476 6416 3488 6480
rect 18248 6458 18260 6522
rect 18324 6458 18340 6522
rect 18404 6458 18420 6522
rect 18484 6458 18500 6522
rect 18564 6458 18576 6522
rect 18248 6427 18576 6458
rect 3160 6385 3488 6416
rect 10716 6136 11000 6153
rect 10716 6072 10746 6136
rect 10810 6072 10826 6136
rect 10890 6072 10906 6136
rect 10970 6072 11000 6136
rect 10716 6055 11000 6072
rect -2509 5510 -2181 5536
rect -2509 5446 -2497 5510
rect -2433 5446 -2417 5510
rect -2353 5446 -2337 5510
rect -2273 5446 -2257 5510
rect -2193 5446 -2181 5510
rect -2509 5420 -2181 5446
rect 1267 5510 1595 5536
rect 1267 5446 1279 5510
rect 1343 5446 1359 5510
rect 1423 5446 1439 5510
rect 1503 5446 1519 5510
rect 1583 5446 1595 5510
rect 1267 5420 1595 5446
rect 5043 5510 5371 5536
rect 5043 5446 5055 5510
rect 5119 5446 5135 5510
rect 5199 5446 5215 5510
rect 5279 5446 5295 5510
rect 5359 5446 5371 5510
rect 5043 5420 5371 5446
rect 8819 5510 9147 5536
rect 8819 5446 8831 5510
rect 8895 5446 8911 5510
rect 8975 5446 8991 5510
rect 9055 5446 9071 5510
rect 9135 5446 9147 5510
rect 8819 5420 9147 5446
rect 12589 5510 12917 5536
rect 12589 5446 12601 5510
rect 12665 5446 12681 5510
rect 12745 5446 12761 5510
rect 12825 5446 12841 5510
rect 12905 5446 12917 5510
rect 12589 5420 12917 5446
rect 16365 5510 16693 5536
rect 16365 5446 16377 5510
rect 16441 5446 16457 5510
rect 16521 5446 16537 5510
rect 16601 5446 16617 5510
rect 16681 5446 16693 5510
rect 16365 5420 16693 5446
rect 20141 5510 20469 5536
rect 20141 5446 20153 5510
rect 20217 5446 20233 5510
rect 20297 5446 20313 5510
rect 20377 5446 20393 5510
rect 20457 5446 20469 5510
rect 20141 5420 20469 5446
rect -4397 3386 -4069 3412
rect -4397 3322 -4385 3386
rect -4321 3322 -4305 3386
rect -4241 3322 -4225 3386
rect -4161 3322 -4145 3386
rect -4081 3322 -4069 3386
rect -4397 3296 -4069 3322
rect -621 3386 -293 3412
rect -621 3322 -609 3386
rect -545 3322 -529 3386
rect -465 3322 -449 3386
rect -385 3322 -369 3386
rect -305 3322 -293 3386
rect -621 3296 -293 3322
rect 3155 3386 3483 3412
rect 3155 3322 3167 3386
rect 3231 3322 3247 3386
rect 3311 3322 3327 3386
rect 3391 3322 3407 3386
rect 3471 3322 3483 3386
rect 3155 3296 3483 3322
rect 6931 3386 7259 3412
rect 6931 3322 6943 3386
rect 7007 3322 7023 3386
rect 7087 3322 7103 3386
rect 7167 3322 7183 3386
rect 7247 3322 7259 3386
rect 6931 3296 7259 3322
rect 10707 3386 11035 3412
rect 10707 3322 10719 3386
rect 10783 3322 10799 3386
rect 10863 3322 10879 3386
rect 10943 3322 10959 3386
rect 11023 3322 11035 3386
rect 10707 3296 11035 3322
rect 14477 3386 14805 3412
rect 14477 3322 14489 3386
rect 14553 3322 14569 3386
rect 14633 3322 14649 3386
rect 14713 3322 14729 3386
rect 14793 3322 14805 3386
rect 14477 3296 14805 3322
rect 18253 3386 18581 3412
rect 18253 3322 18265 3386
rect 18329 3322 18345 3386
rect 18409 3322 18425 3386
rect 18489 3322 18505 3386
rect 18569 3322 18581 3386
rect 18253 3296 18581 3322
rect 22029 3386 22357 3412
rect 22029 3322 22041 3386
rect 22105 3322 22121 3386
rect 22185 3322 22201 3386
rect 22265 3322 22281 3386
rect 22345 3322 22357 3386
rect 22029 3296 22357 3322
<< via3 >>
rect -4355 9334 -4291 9398
rect -4275 9334 -4211 9398
rect -4195 9334 -4131 9398
rect -4115 9334 -4051 9398
rect -579 9334 -515 9398
rect -499 9334 -435 9398
rect -419 9334 -355 9398
rect -339 9334 -275 9398
rect 3197 9334 3261 9398
rect 3277 9334 3341 9398
rect 3357 9334 3421 9398
rect 3437 9334 3501 9398
rect 6973 9334 7037 9398
rect 7053 9334 7117 9398
rect 7133 9334 7197 9398
rect 7213 9334 7277 9398
rect 10743 9334 10807 9398
rect 10823 9334 10887 9398
rect 10903 9334 10967 9398
rect 10983 9334 11047 9398
rect 14519 9334 14583 9398
rect 14599 9334 14663 9398
rect 14679 9334 14743 9398
rect 14759 9334 14823 9398
rect 18295 9334 18359 9398
rect 18375 9334 18439 9398
rect 18455 9334 18519 9398
rect 18535 9334 18599 9398
rect 22071 9334 22135 9398
rect 22151 9334 22215 9398
rect 22231 9334 22295 9398
rect 22311 9334 22375 9398
rect -2467 7210 -2403 7274
rect -2387 7210 -2323 7274
rect -2307 7210 -2243 7274
rect -2227 7210 -2163 7274
rect 1309 7210 1373 7274
rect 1389 7210 1453 7274
rect 1469 7210 1533 7274
rect 1549 7210 1613 7274
rect 5085 7210 5149 7274
rect 5165 7210 5229 7274
rect 5245 7210 5309 7274
rect 5325 7210 5389 7274
rect 8861 7210 8925 7274
rect 8941 7210 9005 7274
rect 9021 7210 9085 7274
rect 9101 7210 9165 7274
rect 12631 7210 12695 7274
rect 12711 7210 12775 7274
rect 12791 7210 12855 7274
rect 12871 7210 12935 7274
rect 16407 7210 16471 7274
rect 16487 7210 16551 7274
rect 16567 7210 16631 7274
rect 16647 7210 16711 7274
rect 20183 7210 20247 7274
rect 20263 7210 20327 7274
rect 20343 7210 20407 7274
rect 20423 7210 20487 7274
rect 8862 6674 8926 6678
rect 8862 6618 8866 6674
rect 8866 6618 8922 6674
rect 8922 6618 8926 6674
rect 8862 6614 8926 6618
rect 8942 6674 9006 6678
rect 8942 6618 8946 6674
rect 8946 6618 9002 6674
rect 9002 6618 9006 6674
rect 8942 6614 9006 6618
rect 9022 6674 9086 6678
rect 9022 6618 9026 6674
rect 9026 6618 9082 6674
rect 9082 6618 9086 6674
rect 9022 6614 9086 6618
rect 12628 6676 12692 6680
rect 12628 6620 12632 6676
rect 12632 6620 12688 6676
rect 12688 6620 12692 6676
rect 12628 6616 12692 6620
rect 12708 6676 12772 6680
rect 12708 6620 12712 6676
rect 12712 6620 12768 6676
rect 12768 6620 12772 6676
rect 12708 6616 12772 6620
rect 12788 6676 12852 6680
rect 12788 6620 12792 6676
rect 12792 6620 12848 6676
rect 12848 6620 12852 6676
rect 12788 6616 12852 6620
rect 3172 6476 3236 6480
rect 3172 6420 3176 6476
rect 3176 6420 3232 6476
rect 3232 6420 3236 6476
rect 3172 6416 3236 6420
rect 3252 6476 3316 6480
rect 3252 6420 3256 6476
rect 3256 6420 3312 6476
rect 3312 6420 3316 6476
rect 3252 6416 3316 6420
rect 3332 6476 3396 6480
rect 3332 6420 3336 6476
rect 3336 6420 3392 6476
rect 3392 6420 3396 6476
rect 3332 6416 3396 6420
rect 3412 6476 3476 6480
rect 3412 6420 3416 6476
rect 3416 6420 3472 6476
rect 3472 6420 3476 6476
rect 3412 6416 3476 6420
rect 18260 6518 18324 6522
rect 18260 6462 18264 6518
rect 18264 6462 18320 6518
rect 18320 6462 18324 6518
rect 18260 6458 18324 6462
rect 18340 6518 18404 6522
rect 18340 6462 18344 6518
rect 18344 6462 18400 6518
rect 18400 6462 18404 6518
rect 18340 6458 18404 6462
rect 18420 6518 18484 6522
rect 18420 6462 18424 6518
rect 18424 6462 18480 6518
rect 18480 6462 18484 6518
rect 18420 6458 18484 6462
rect 18500 6518 18564 6522
rect 18500 6462 18504 6518
rect 18504 6462 18560 6518
rect 18560 6462 18564 6518
rect 18500 6458 18564 6462
rect 10746 6132 10810 6136
rect 10746 6076 10750 6132
rect 10750 6076 10806 6132
rect 10806 6076 10810 6132
rect 10746 6072 10810 6076
rect 10826 6132 10890 6136
rect 10826 6076 10830 6132
rect 10830 6076 10886 6132
rect 10886 6076 10890 6132
rect 10826 6072 10890 6076
rect 10906 6132 10970 6136
rect 10906 6076 10910 6132
rect 10910 6076 10966 6132
rect 10966 6076 10970 6132
rect 10906 6072 10970 6076
rect -2497 5446 -2433 5510
rect -2417 5446 -2353 5510
rect -2337 5446 -2273 5510
rect -2257 5446 -2193 5510
rect 1279 5446 1343 5510
rect 1359 5446 1423 5510
rect 1439 5446 1503 5510
rect 1519 5446 1583 5510
rect 5055 5446 5119 5510
rect 5135 5446 5199 5510
rect 5215 5446 5279 5510
rect 5295 5446 5359 5510
rect 8831 5446 8895 5510
rect 8911 5446 8975 5510
rect 8991 5446 9055 5510
rect 9071 5446 9135 5510
rect 12601 5446 12665 5510
rect 12681 5446 12745 5510
rect 12761 5446 12825 5510
rect 12841 5446 12905 5510
rect 16377 5446 16441 5510
rect 16457 5446 16521 5510
rect 16537 5446 16601 5510
rect 16617 5446 16681 5510
rect 20153 5446 20217 5510
rect 20233 5446 20297 5510
rect 20313 5446 20377 5510
rect 20393 5446 20457 5510
rect -4385 3322 -4321 3386
rect -4305 3322 -4241 3386
rect -4225 3322 -4161 3386
rect -4145 3322 -4081 3386
rect -609 3322 -545 3386
rect -529 3322 -465 3386
rect -449 3322 -385 3386
rect -369 3322 -305 3386
rect 3167 3322 3231 3386
rect 3247 3322 3311 3386
rect 3327 3322 3391 3386
rect 3407 3322 3471 3386
rect 6943 3322 7007 3386
rect 7023 3322 7087 3386
rect 7103 3322 7167 3386
rect 7183 3322 7247 3386
rect 10719 3322 10783 3386
rect 10799 3322 10863 3386
rect 10879 3322 10943 3386
rect 10959 3322 11023 3386
rect 14489 3322 14553 3386
rect 14569 3322 14633 3386
rect 14649 3322 14713 3386
rect 14729 3322 14793 3386
rect 18265 3322 18329 3386
rect 18345 3322 18409 3386
rect 18425 3322 18489 3386
rect 18505 3322 18569 3386
rect 22041 3322 22105 3386
rect 22121 3322 22185 3386
rect 22201 3322 22265 3386
rect 22281 3322 22345 3386
<< metal4 >>
rect -4400 9425 -4062 9488
rect -4400 9398 -4048 9425
rect -4400 9334 -4355 9398
rect -4291 9334 -4275 9398
rect -4211 9334 -4195 9398
rect -4131 9334 -4115 9398
rect -4051 9334 -4048 9398
rect -4400 9307 -4048 9334
rect -4400 3386 -4062 9307
rect -4400 3322 -4385 3386
rect -4321 3322 -4305 3386
rect -4241 3322 -4225 3386
rect -4161 3322 -4145 3386
rect -4081 3322 -4062 3386
rect -4400 3232 -4062 3322
rect -2502 7301 -2164 9488
rect -616 9425 -278 9488
rect -616 9398 -272 9425
rect -616 9334 -579 9398
rect -515 9334 -499 9398
rect -435 9334 -419 9398
rect -355 9334 -339 9398
rect -275 9334 -272 9398
rect -616 9307 -272 9334
rect -2502 7274 -2160 7301
rect -2502 7210 -2467 7274
rect -2403 7210 -2387 7274
rect -2323 7210 -2307 7274
rect -2243 7210 -2227 7274
rect -2163 7210 -2160 7274
rect -2502 7183 -2160 7210
rect -2502 5510 -2164 7183
rect -2502 5446 -2497 5510
rect -2433 5446 -2417 5510
rect -2353 5446 -2337 5510
rect -2273 5446 -2257 5510
rect -2193 5446 -2164 5510
rect -2502 3232 -2164 5446
rect -616 3386 -278 9307
rect -616 3322 -609 3386
rect -545 3322 -529 3386
rect -465 3322 -449 3386
rect -385 3322 -369 3386
rect -305 3322 -278 3386
rect -616 3232 -278 3322
rect 1274 7301 1612 9488
rect 3158 9425 3492 9488
rect 3158 9398 3504 9425
rect 3158 9334 3197 9398
rect 3261 9334 3277 9398
rect 3341 9334 3357 9398
rect 3421 9334 3437 9398
rect 3501 9334 3504 9398
rect 3158 9307 3504 9334
rect 1274 7274 1616 7301
rect 1274 7210 1309 7274
rect 1373 7210 1389 7274
rect 1453 7210 1469 7274
rect 1533 7210 1549 7274
rect 1613 7210 1616 7274
rect 1274 7183 1616 7210
rect 1274 5510 1612 7183
rect 1274 5446 1279 5510
rect 1343 5446 1359 5510
rect 1423 5446 1439 5510
rect 1503 5446 1519 5510
rect 1583 5446 1612 5510
rect 1274 3232 1612 5446
rect 3158 6480 3492 9307
rect 3158 6416 3172 6480
rect 3236 6416 3252 6480
rect 3316 6416 3332 6480
rect 3396 6416 3412 6480
rect 3476 6416 3492 6480
rect 3158 3386 3492 6416
rect 3158 3322 3167 3386
rect 3231 3322 3247 3386
rect 3311 3322 3327 3386
rect 3391 3322 3407 3386
rect 3471 3322 3492 3386
rect 3158 3232 3492 3322
rect 5044 7301 5382 9488
rect 6936 9425 7274 9488
rect 6936 9398 7280 9425
rect 6936 9334 6973 9398
rect 7037 9334 7053 9398
rect 7117 9334 7133 9398
rect 7197 9334 7213 9398
rect 7277 9334 7280 9398
rect 6936 9307 7280 9334
rect 5044 7274 5392 7301
rect 5044 7210 5085 7274
rect 5149 7210 5165 7274
rect 5229 7210 5245 7274
rect 5309 7210 5325 7274
rect 5389 7210 5392 7274
rect 5044 7183 5392 7210
rect 5044 5510 5382 7183
rect 5044 5446 5055 5510
rect 5119 5446 5135 5510
rect 5199 5446 5215 5510
rect 5279 5446 5295 5510
rect 5359 5446 5382 5510
rect 5044 3232 5382 5446
rect 6936 3386 7274 9307
rect 6936 3322 6943 3386
rect 7007 3322 7023 3386
rect 7087 3322 7103 3386
rect 7167 3322 7183 3386
rect 7247 3322 7274 3386
rect 6936 3232 7274 3322
rect 8812 7301 9150 9488
rect 10704 9425 11042 9488
rect 10704 9398 11050 9425
rect 10704 9334 10743 9398
rect 10807 9334 10823 9398
rect 10887 9334 10903 9398
rect 10967 9334 10983 9398
rect 11047 9334 11050 9398
rect 10704 9307 11050 9334
rect 8812 7274 9168 7301
rect 8812 7210 8861 7274
rect 8925 7210 8941 7274
rect 9005 7210 9021 7274
rect 9085 7210 9101 7274
rect 9165 7210 9168 7274
rect 8812 7183 9168 7210
rect 8812 6678 9150 7183
rect 8812 6614 8862 6678
rect 8926 6614 8942 6678
rect 9006 6614 9022 6678
rect 9086 6614 9150 6678
rect 8812 5510 9150 6614
rect 8812 5446 8831 5510
rect 8895 5446 8911 5510
rect 8975 5446 8991 5510
rect 9055 5446 9071 5510
rect 9135 5446 9150 5510
rect 8812 3232 9150 5446
rect 10704 6136 11042 9307
rect 10704 6072 10746 6136
rect 10810 6072 10826 6136
rect 10890 6072 10906 6136
rect 10970 6072 11042 6136
rect 10704 3386 11042 6072
rect 10704 3322 10719 3386
rect 10783 3322 10799 3386
rect 10863 3322 10879 3386
rect 10943 3322 10959 3386
rect 11023 3322 11042 3386
rect 10704 3232 11042 3322
rect 12584 7301 12922 9488
rect 14476 9425 14814 9488
rect 14476 9398 14826 9425
rect 14476 9334 14519 9398
rect 14583 9334 14599 9398
rect 14663 9334 14679 9398
rect 14743 9334 14759 9398
rect 14823 9334 14826 9398
rect 14476 9307 14826 9334
rect 12584 7274 12938 7301
rect 12584 7210 12631 7274
rect 12695 7210 12711 7274
rect 12775 7210 12791 7274
rect 12855 7210 12871 7274
rect 12935 7210 12938 7274
rect 12584 7183 12938 7210
rect 12584 6680 12922 7183
rect 12584 6616 12628 6680
rect 12692 6616 12708 6680
rect 12772 6616 12788 6680
rect 12852 6616 12922 6680
rect 12584 5510 12922 6616
rect 12584 5446 12601 5510
rect 12665 5446 12681 5510
rect 12745 5446 12761 5510
rect 12825 5446 12841 5510
rect 12905 5446 12922 5510
rect 12584 3232 12922 5446
rect 14476 3386 14814 9307
rect 14476 3322 14489 3386
rect 14553 3322 14569 3386
rect 14633 3322 14649 3386
rect 14713 3322 14729 3386
rect 14793 3322 14814 3386
rect 14476 3232 14814 3322
rect 16352 7301 16690 9488
rect 18246 9425 18584 9488
rect 18246 9398 18602 9425
rect 18246 9334 18295 9398
rect 18359 9334 18375 9398
rect 18439 9334 18455 9398
rect 18519 9334 18535 9398
rect 18599 9334 18602 9398
rect 18246 9307 18602 9334
rect 16352 7274 16714 7301
rect 16352 7210 16407 7274
rect 16471 7210 16487 7274
rect 16551 7210 16567 7274
rect 16631 7210 16647 7274
rect 16711 7210 16714 7274
rect 16352 7183 16714 7210
rect 16352 5510 16690 7183
rect 16352 5446 16377 5510
rect 16441 5446 16457 5510
rect 16521 5446 16537 5510
rect 16601 5446 16617 5510
rect 16681 5446 16690 5510
rect 16352 3232 16690 5446
rect 18246 6522 18584 9307
rect 18246 6458 18260 6522
rect 18324 6458 18340 6522
rect 18404 6458 18420 6522
rect 18484 6458 18500 6522
rect 18564 6458 18584 6522
rect 18246 3386 18584 6458
rect 18246 3322 18265 3386
rect 18329 3322 18345 3386
rect 18409 3322 18425 3386
rect 18489 3322 18505 3386
rect 18569 3322 18584 3386
rect 18246 3232 18584 3322
rect 20148 7301 20486 9488
rect 22034 9425 22372 9488
rect 22034 9398 22378 9425
rect 22034 9334 22071 9398
rect 22135 9334 22151 9398
rect 22215 9334 22231 9398
rect 22295 9334 22311 9398
rect 22375 9334 22378 9398
rect 22034 9307 22378 9334
rect 20148 7274 20490 7301
rect 20148 7210 20183 7274
rect 20247 7210 20263 7274
rect 20327 7210 20343 7274
rect 20407 7210 20423 7274
rect 20487 7210 20490 7274
rect 20148 7183 20490 7210
rect 20148 5510 20486 7183
rect 20148 5446 20153 5510
rect 20217 5446 20233 5510
rect 20297 5446 20313 5510
rect 20377 5446 20393 5510
rect 20457 5446 20486 5510
rect 20148 3232 20486 5446
rect 22034 3386 22372 9307
rect 22034 3322 22041 3386
rect 22105 3322 22121 3386
rect 22185 3322 22201 3386
rect 22265 3322 22281 3386
rect 22345 3322 22372 3386
rect 22034 3232 22372 3322
use brbufhalf_32  brbufhalf_32_0
timestamp 1654402208
transform 1 0 -482 0 1 704
box -1666 2527 26746 5370
use brbufhalf_32  brbufhalf_32_1
timestamp 1654402208
transform -1 0 22247 0 -1 12016
box -1666 2527 26746 5370
use invcell  invcell_0
timestamp 1654402208
transform 1 0 -218 0 1 -832
box 8992 6886 13248 7528
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1654402208
transform 1 0 13048 0 1 6102
box -38 -48 130 592
use unitcell2buf_32  unitcell2buf_32_0
timestamp 1654402208
transform 1 0 -5348 0 1 4416
box -574 -1185 1322 1192
use unitcell2buf_32  unitcell2buf_32_1
timestamp 1654402208
transform 1 0 -3460 0 1 4416
box -574 -1185 1322 1192
<< labels >>
flabel metal4 s -2424 9032 -2268 9232 1 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 26100 4032 26132 4062 1 FreeSans 500 0 0 0 OUT
port 2 nsew
flabel metal2 s 6866 9392 6900 9452 1 FreeSans 500 0 0 0 C9
port 3 nsew
flabel metal2 s 4980 9402 5014 9462 1 FreeSans 500 0 0 0 C10
port 4 nsew
flabel metal2 s 3094 9396 3128 9456 1 FreeSans 500 0 0 0 C11
port 5 nsew
flabel metal2 s 1204 9406 1238 9466 1 FreeSans 500 0 0 0 C12
port 6 nsew
flabel metal2 s -682 9384 -648 9444 1 FreeSans 500 0 0 0 C13
port 7 nsew
flabel metal2 s -2574 9408 -2540 9468 1 FreeSans 500 0 0 0 C14
port 8 nsew
flabel metal2 s -5896 3240 -5862 3300 1 FreeSans 500 0 0 0 C15
port 9 nsew
flabel metal2 s -4008 3240 -3974 3300 1 FreeSans 500 0 0 0 C16
port 10 nsew
flabel metal2 s -2122 3240 -2088 3300 1 FreeSans 500 0 0 0 C17
port 11 nsew
flabel metal2 s -232 3248 -198 3308 1 FreeSans 500 0 0 0 C18
port 12 nsew
flabel metal2 s 1654 3246 1688 3306 1 FreeSans 500 0 0 0 C19
port 13 nsew
flabel metal2 s 3546 3242 3580 3302 1 FreeSans 500 0 0 0 C20
port 14 nsew
flabel metal2 s 5432 3246 5466 3306 1 FreeSans 500 0 0 0 C21
port 15 nsew
flabel metal2 s 7322 3246 7356 3306 1 FreeSans 500 0 0 0 C22
port 16 nsew
flabel metal2 s 9206 3246 9240 3306 1 FreeSans 500 0 0 0 C23
port 17 nsew
flabel metal2 s 11088 3250 11122 3310 1 FreeSans 500 0 0 0 C24
port 18 nsew
flabel metal2 s 12978 3250 13012 3310 1 FreeSans 500 0 0 0 C25
port 19 nsew
flabel metal2 s 14866 3246 14900 3306 1 FreeSans 500 0 0 0 C26
port 20 nsew
flabel metal2 s 16756 3246 16790 3306 1 FreeSans 500 0 0 0 C27
port 21 nsew
flabel metal2 s 18640 3246 18674 3306 1 FreeSans 500 0 0 0 C28
port 22 nsew
flabel metal2 s 20532 3254 20566 3314 1 FreeSans 500 0 0 0 C29
port 23 nsew
flabel metal2 s 22418 3246 22452 3306 1 FreeSans 500 0 0 0 C30
port 24 nsew
flabel metal2 s 24306 3244 24340 3304 1 FreeSans 500 0 0 0 C31
port 25 nsew
flabel metal2 s 21964 9386 21998 9446 1 FreeSans 500 0 0 0 C1
port 26 nsew
flabel metal2 s 20082 9386 20116 9446 1 FreeSans 500 0 0 0 C2
port 27 nsew
flabel metal2 s 18188 9392 18222 9452 1 FreeSans 500 0 0 0 C3
port 28 nsew
flabel metal2 s 16300 9398 16334 9458 1 FreeSans 500 0 0 0 C4
port 29 nsew
flabel metal2 s 14412 9392 14446 9452 1 FreeSans 500 0 0 0 C5
port 30 nsew
flabel metal2 s 12526 9398 12560 9458 1 FreeSans 500 0 0 0 C6
port 31 nsew
flabel metal2 s 10646 9402 10680 9462 1 FreeSans 500 0 0 0 C7
port 32 nsew
flabel metal2 s 8758 9406 8792 9466 1 FreeSans 500 0 0 0 C8
port 33 nsew
flabel metal2 s -6046 6308 -5968 6326 1 FreeSans 500 0 0 0 RESET
port 34 nsew
flabel metal4 s -4316 9038 -4160 9238 1 FreeSans 500 0 0 0 VSS
port 35 nsew
flabel metal2 s 23854 9392 23888 9452 1 FreeSans 500 0 0 0 C0
port 36 nsew
<< end >>
