magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 551 157
rect 29 -17 63 21
<< locali >>
rect 94 240 179 391
rect 213 331 261 493
rect 213 240 322 331
rect 263 51 322 240
rect 356 153 434 323
rect 468 153 523 287
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 417 71 493
rect 105 435 171 527
rect 19 206 60 417
rect 295 401 361 493
rect 395 435 433 527
rect 467 401 533 493
rect 295 365 533 401
rect 19 156 229 206
rect 19 56 76 156
rect 110 17 229 122
rect 467 17 533 119
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 356 153 434 323 6 A1
port 1 nsew signal input
rlabel locali s 468 153 523 287 6 A2
port 2 nsew signal input
rlabel locali s 94 240 179 391 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 551 157 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 263 51 322 240 6 Y
port 8 nsew signal output
rlabel locali s 213 240 322 331 6 Y
port 8 nsew signal output
rlabel locali s 213 331 261 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4003510
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3998334
<< end >>
