magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1563 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 687 47 717 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1194 47 1224 177
rect 1278 47 1308 177
rect 1371 47 1401 177
rect 1455 47 1485 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 687 297 717 497
rect 771 297 801 497
rect 855 297 885 497
rect 939 297 969 497
rect 1203 297 1233 497
rect 1287 297 1317 497
rect 1371 297 1401 497
rect 1455 297 1485 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 101 163 177
rect 109 67 119 101
rect 153 67 163 101
rect 109 47 163 67
rect 193 93 247 177
rect 193 59 203 93
rect 237 59 247 93
rect 193 47 247 59
rect 277 101 331 177
rect 277 67 287 101
rect 321 67 331 101
rect 277 47 331 67
rect 361 93 415 177
rect 361 59 371 93
rect 405 59 415 93
rect 361 47 415 59
rect 445 101 499 177
rect 445 67 455 101
rect 489 67 499 101
rect 445 47 499 67
rect 529 93 581 177
rect 529 59 539 93
rect 573 59 581 93
rect 529 47 581 59
rect 635 93 687 177
rect 635 59 643 93
rect 677 59 687 93
rect 635 47 687 59
rect 717 165 771 177
rect 717 131 727 165
rect 761 131 771 165
rect 717 47 771 131
rect 801 93 855 177
rect 801 59 811 93
rect 845 59 855 93
rect 801 47 855 59
rect 885 161 939 177
rect 885 127 895 161
rect 929 127 939 161
rect 885 47 939 127
rect 969 93 1021 177
rect 969 59 979 93
rect 1013 59 1021 93
rect 969 47 1021 59
rect 1142 93 1194 177
rect 1142 59 1150 93
rect 1184 59 1194 93
rect 1142 47 1194 59
rect 1224 161 1278 177
rect 1224 127 1234 161
rect 1268 127 1278 161
rect 1224 47 1278 127
rect 1308 101 1371 177
rect 1308 67 1327 101
rect 1361 67 1371 101
rect 1308 47 1371 67
rect 1401 93 1455 177
rect 1401 59 1411 93
rect 1445 59 1455 93
rect 1401 47 1455 59
rect 1485 101 1537 177
rect 1485 67 1495 101
rect 1529 67 1537 101
rect 1485 47 1537 67
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 297 79 383
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 477 331 497
rect 277 443 287 477
rect 321 443 331 477
rect 277 409 331 443
rect 277 375 287 409
rect 321 375 331 409
rect 277 297 331 375
rect 361 485 415 497
rect 361 451 371 485
rect 405 451 415 485
rect 361 417 415 451
rect 361 383 371 417
rect 405 383 415 417
rect 361 297 415 383
rect 445 477 499 497
rect 445 443 455 477
rect 489 443 499 477
rect 445 297 499 443
rect 529 485 581 497
rect 529 451 539 485
rect 573 451 581 485
rect 529 297 581 451
rect 635 477 687 497
rect 635 443 643 477
rect 677 443 687 477
rect 635 297 687 443
rect 717 485 771 497
rect 717 451 727 485
rect 761 451 771 485
rect 717 297 771 451
rect 801 477 855 497
rect 801 443 811 477
rect 845 443 855 477
rect 801 297 855 443
rect 885 485 939 497
rect 885 451 895 485
rect 929 451 939 485
rect 885 297 939 451
rect 969 485 1203 497
rect 969 451 1159 485
rect 1193 451 1203 485
rect 969 297 1203 451
rect 1233 417 1287 497
rect 1233 383 1243 417
rect 1277 383 1287 417
rect 1233 297 1287 383
rect 1317 485 1371 497
rect 1317 451 1327 485
rect 1361 451 1371 485
rect 1317 297 1371 451
rect 1401 417 1455 497
rect 1401 383 1411 417
rect 1445 383 1455 417
rect 1401 297 1455 383
rect 1485 485 1537 497
rect 1485 451 1495 485
rect 1529 451 1537 485
rect 1485 401 1537 451
rect 1485 367 1495 401
rect 1529 367 1537 401
rect 1485 297 1537 367
<< ndiffc >>
rect 35 59 69 93
rect 119 67 153 101
rect 203 59 237 93
rect 287 67 321 101
rect 371 59 405 93
rect 455 67 489 101
rect 539 59 573 93
rect 643 59 677 93
rect 727 131 761 165
rect 811 59 845 93
rect 895 127 929 161
rect 979 59 1013 93
rect 1150 59 1184 93
rect 1234 127 1268 161
rect 1327 67 1361 101
rect 1411 59 1445 93
rect 1495 67 1529 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 119 443 153 477
rect 119 375 153 409
rect 203 451 237 485
rect 203 383 237 417
rect 287 443 321 477
rect 287 375 321 409
rect 371 451 405 485
rect 371 383 405 417
rect 455 443 489 477
rect 539 451 573 485
rect 643 443 677 477
rect 727 451 761 485
rect 811 443 845 477
rect 895 451 929 485
rect 1159 451 1193 485
rect 1243 383 1277 417
rect 1327 451 1361 485
rect 1411 383 1445 417
rect 1495 451 1529 485
rect 1495 367 1529 401
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 687 497 717 523
rect 771 497 801 523
rect 855 497 885 523
rect 939 497 969 523
rect 1203 497 1233 523
rect 1287 497 1317 523
rect 1371 497 1401 523
rect 1455 497 1485 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 79 249 361 265
rect 79 215 114 249
rect 148 215 188 249
rect 222 215 262 249
rect 296 215 361 249
rect 79 199 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 687 269 717 297
rect 771 269 801 297
rect 415 261 542 265
rect 415 249 576 261
rect 687 259 801 269
rect 415 215 458 249
rect 492 215 526 249
rect 560 215 576 249
rect 415 203 576 215
rect 667 249 801 259
rect 667 215 683 249
rect 717 215 751 249
rect 785 215 801 249
rect 667 205 801 215
rect 415 199 542 203
rect 687 199 801 205
rect 415 177 445 199
rect 499 177 529 199
rect 687 177 717 199
rect 771 177 801 199
rect 855 269 885 297
rect 939 269 969 297
rect 855 261 969 269
rect 1203 265 1233 297
rect 1287 265 1317 297
rect 855 249 1015 261
rect 1203 259 1317 265
rect 855 215 897 249
rect 931 215 965 249
rect 999 215 1015 249
rect 855 205 1015 215
rect 1183 249 1317 259
rect 1183 215 1199 249
rect 1233 215 1267 249
rect 1301 215 1317 249
rect 1183 205 1317 215
rect 1371 265 1401 297
rect 1455 265 1485 297
rect 1371 261 1485 265
rect 1371 249 1542 261
rect 1371 215 1424 249
rect 1458 215 1492 249
rect 1526 215 1542 249
rect 1371 205 1542 215
rect 855 177 885 205
rect 939 203 1015 205
rect 939 177 969 203
rect 1194 177 1224 205
rect 1278 177 1308 205
rect 1371 177 1401 205
rect 1455 203 1542 205
rect 1455 177 1485 203
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 687 21 717 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1194 21 1224 47
rect 1278 21 1308 47
rect 1371 21 1401 47
rect 1455 21 1485 47
<< polycont >>
rect 114 215 148 249
rect 188 215 222 249
rect 262 215 296 249
rect 458 215 492 249
rect 526 215 560 249
rect 683 215 717 249
rect 751 215 785 249
rect 897 215 931 249
rect 965 215 999 249
rect 1199 215 1233 249
rect 1267 215 1301 249
rect 1424 215 1458 249
rect 1492 215 1526 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 19 485 85 527
rect 19 451 35 485
rect 69 451 85 485
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 119 477 153 493
rect 119 409 153 443
rect 187 485 253 527
rect 187 451 203 485
rect 237 451 253 485
rect 187 417 253 451
rect 187 383 203 417
rect 237 383 253 417
rect 287 477 321 493
rect 287 409 321 443
rect 119 333 153 375
rect 355 485 421 527
rect 355 451 371 485
rect 405 451 421 485
rect 355 417 421 451
rect 355 383 371 417
rect 405 383 421 417
rect 455 477 489 493
rect 523 485 589 527
rect 523 451 539 485
rect 573 451 589 485
rect 643 477 677 493
rect 455 417 489 443
rect 711 485 777 527
rect 711 451 727 485
rect 761 451 777 485
rect 811 477 845 493
rect 643 417 677 443
rect 879 485 945 527
rect 879 451 895 485
rect 929 451 945 485
rect 979 451 1159 485
rect 1193 451 1327 485
rect 1361 451 1495 485
rect 1529 451 1545 485
rect 811 417 845 443
rect 979 417 1013 451
rect 455 383 1013 417
rect 1227 415 1243 417
rect 1056 383 1243 415
rect 1277 383 1411 417
rect 1445 383 1461 417
rect 1495 401 1545 451
rect 287 333 321 375
rect 1056 381 1240 383
rect 1056 333 1090 381
rect 1529 367 1545 401
rect 1495 351 1545 367
rect 24 299 321 333
rect 360 299 1090 333
rect 24 161 68 299
rect 360 265 394 299
rect 114 249 394 265
rect 148 215 188 249
rect 222 215 262 249
rect 296 215 394 249
rect 442 249 621 259
rect 442 215 458 249
rect 492 215 526 249
rect 560 215 621 249
rect 667 249 806 265
rect 667 215 683 249
rect 717 215 751 249
rect 785 215 806 249
rect 856 249 1015 265
rect 856 215 897 249
rect 931 215 965 249
rect 999 215 1015 249
rect 114 199 394 215
rect 24 127 321 161
rect 119 101 153 127
rect 19 59 35 93
rect 69 59 85 93
rect 19 17 85 59
rect 287 101 321 127
rect 119 51 153 67
rect 187 59 203 93
rect 237 59 253 93
rect 187 17 253 59
rect 455 131 727 165
rect 761 131 777 165
rect 1056 161 1090 299
rect 1126 249 1356 325
rect 1126 215 1199 249
rect 1233 215 1267 249
rect 1301 215 1356 249
rect 1406 259 1445 327
rect 1406 249 1542 259
rect 1406 215 1424 249
rect 1458 215 1492 249
rect 1526 215 1542 249
rect 455 101 489 131
rect 879 127 895 161
rect 929 127 1234 161
rect 1268 127 1285 161
rect 1327 129 1529 163
rect 287 51 321 67
rect 355 59 371 93
rect 405 59 421 93
rect 355 17 421 59
rect 1327 101 1361 129
rect 455 51 489 67
rect 523 59 539 93
rect 573 59 589 93
rect 627 59 643 93
rect 677 59 811 93
rect 845 59 979 93
rect 1013 59 1029 93
rect 1134 59 1150 93
rect 1184 67 1327 93
rect 1495 101 1529 129
rect 1184 59 1361 67
rect 523 17 589 59
rect 1327 51 1361 59
rect 1395 59 1411 93
rect 1445 59 1461 93
rect 1395 17 1461 59
rect 1495 51 1529 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 678 221 712 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 30 153 64 187 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 1224 289 1258 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1132 289 1166 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1132 221 1166 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1500 221 1534 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 1316 289 1350 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 1316 221 1350 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1224 221 1258 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1408 289 1442 323 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 1408 221 1442 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a32o_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 3479836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3467700
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 39.100 0.000 
<< end >>
