* NGSPICE file created from brbufhalf_lvs_flat.ext - technology: sky130A

.subckt brbufhalf_lvs_flat OUT RESET1 RESET2 IN VSS VDD
X0 VSS a_6572_3230# a_7497_3153# VSS sky130_fd_pr__nfet_01v8 ad=2.49028e+13p pd=2.6672e+08u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1 a_17894_3230# a_17400_3147# a_17455_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2 a_8460_3230# a_8192_3293# a_8021_4451# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X3 a_21231_4451# a_21226_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X4 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X5 a_3891_3153# a_3721_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=3.92256e+13p ps=3.6968e+08u w=790000u l=150000u
X6 a_8556_3230# a_8558_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X7 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X8 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VSS a_n3183_4389# a_10444_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X10 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X11 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_2894_4286# a_2528_3293# a_908_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X13 a_23654_3230# a_23290_3293# a_23558_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X14 a_8192_3293# a_7966_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_6572_3230# a_6078_3147# a_6133_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X16 a_4780_3230# a_4190_3147# a_4684_3230# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X17 a_n2868_3230# a_n1248_3293# a_n1424_4353# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X18 VSS a_11915_4389# a_14214_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X19 a_24653_3153# a_24483_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X20 a_11443_3153# a_11273_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X21 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X23 a_11962_3293# a_11736_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X24 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_n3362_3147# a_n3448_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X26 a_n980_3230# a_n1248_3293# a_n1419_4451# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X27 a_10446_4286# a_10080_3293# a_8460_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X28 VDD a_15738_3293# a_15562_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X29 VSS a_n3183_4389# a_6668_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X30 a_2892_3230# a_2528_3293# a_2796_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X31 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_19288_3147# a_19202_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X33 VSS a_n3183_4389# a_2892_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X34 a_23558_3230# a_24952_3147# a_25002_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X35 a_n2868_3230# a_n1474_3147# a_n1424_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X36 a_21766_3230# a_21768_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X37 a_n2770_4286# a_n3136_3293# IN VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X38 VSS a_11915_4389# a_25007_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X39 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 a_3891_3153# a_3721_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X41 a_14118_3230# a_15512_3147# a_15562_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X42 a_22765_3153# a_22595_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X43 VDD a_4416_3293# a_4240_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X44 a_n3136_3293# a_n3362_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X45 a_n980_3230# a_640_3293# a_464_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X46 a_n980_3230# a_n1474_3147# a_n1419_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X47 VDD a_11915_4389# a_19425_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X48 VSS a_11915_4389# a_11791_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X49 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X52 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X53 a_10444_3230# a_10080_3293# a_10348_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X54 a_n2772_3230# a_n3136_3293# a_n2868_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X55 a_21768_4286# a_21402_3293# a_19782_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X56 a_6215_4451# a_6128_4353# a_6133_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X57 a_2796_3230# a_4190_3147# a_4240_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_2439_4451# a_2352_4353# a_2357_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X59 a_25446_3230# a_24952_3147# a_25007_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=3.3e+11p pd=2.66e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X60 a_25544_4286# a_24952_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X61 a_17455_4451# a_17450_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X62 VSS a_n3183_4389# a_4245_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X63 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 a_11443_3153# a_11273_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X65 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 VDD a_n3183_4389# a_8103_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X67 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X68 a_17626_3293# a_17400_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X69 a_16006_3230# a_15512_3147# a_15567_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X70 a_6572_3230# a_6304_3293# a_6133_4451# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X71 a_2003_3153# a_1833_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X72 a_6668_3230# a_6670_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X73 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X74 a_908_3230# a_640_3293# a_469_4451# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X75 VDD a_n3183_4389# a_n3225_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X76 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 VDD a_17894_3230# a_18819_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X78 a_21766_3230# a_21402_3293# a_21670_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X79 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X80 a_6304_3293# a_6078_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X81 a_4684_3230# a_4190_3147# a_4245_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X82 a_469_4451# a_464_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X83 a_23290_3293# a_23064_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X84 a_18351_4451# a_17992_4286# a_17990_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X85 a_17400_3147# a_17314_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X86 a_2892_3230# a_2302_3147# a_2796_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X87 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X88 a_22765_3153# a_22595_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X89 a_13850_3293# a_13624_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X90 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X91 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X92 VDD a_23290_3293# a_23114_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X93 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_17101_3153# a_16931_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X95 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X96 a_17894_3230# a_19514_3293# a_19338_4353# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X97 a_25903_4451# a_25544_4286# a_25542_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X98 VDD a_13850_3293# a_13674_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X99 VSS a_n3183_4389# a_4780_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X100 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 VSS a_n3183_4389# a_1004_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X102 a_25089_4451# a_25002_4353# a_25007_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X103 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X104 a_16104_4286# a_15738_3293# a_14118_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X105 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 VSS a_11915_4389# a_23119_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X107 a_n2411_4451# a_n2770_4286# a_n2772_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X108 a_2003_3153# a_1833_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X109 a_25544_4286# a_24952_3147# a_23558_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X110 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X111 a_20877_3153# a_20707_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X112 VDD a_2528_3293# a_2352_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X113 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 a_16104_4286# a_15512_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 VDD a_11915_4389# a_17537_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X117 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X118 a_6078_3147# a_5992_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X119 VSS a_17894_3230# a_18819_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X120 a_24952_3147# a_24866_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X121 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X122 a_414_3147# a_328_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X123 a_4327_4451# a_4240_4353# a_4245_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X124 a_10080_3293# a_9854_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X125 a_908_3230# a_2302_3147# a_2352_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 VSS a_n3183_4389# a_n3307_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X127 a_25178_3293# a_24952_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X128 a_19343_4451# a_19338_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X129 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 a_23558_3230# a_23064_3147# a_23119_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X131 a_n882_4286# a_n1474_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X132 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X133 VSS a_n3183_4389# a_2357_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X134 a_23656_4286# a_23064_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X135 a_16102_3230# a_15738_3293# a_16006_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X136 a_15567_4451# a_15562_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X137 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X138 a_n1248_3293# a_n1474_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X139 VDD a_n3183_4389# a_6215_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 a_15738_3293# a_15512_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X141 a_n882_4286# a_n1474_3147# a_n2868_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X142 VDD a_n3183_4389# a_551_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X143 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X144 a_17101_3153# a_16931_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X145 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X146 VDD a_25446_3230# a_26371_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X147 VDD a_n3183_4389# a_n1337_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X148 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X149 a_8021_4451# a_8016_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X150 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X151 a_n884_3230# a_n1474_3147# a_n980_3230# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X152 VSS a_11915_4389# a_23654_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X153 VDD a_16006_3230# a_16931_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X154 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 a_n3225_4451# a_n3312_4353# a_n3307_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X156 a_4416_3293# a_4190_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X157 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X158 a_2796_3230# a_2302_3147# a_2357_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 VSS a_n3183_4389# a_9909_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X160 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X161 a_21402_3293# a_21176_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X162 a_16463_4451# a_16104_4286# a_16102_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X163 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X164 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X165 a_15512_3147# a_15426_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X166 a_20877_3153# a_20707_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X167 a_11736_3147# a_11650_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X168 VDD a_25178_3293# a_25002_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X169 VDD a_4684_3230# a_5609_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X170 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X171 a_15213_3153# a_15043_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X172 VDD a_11915_4389# a_20239_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X173 a_16006_3230# a_17626_3293# a_17450_4353# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X174 a_24015_4451# a_23656_4286# a_23654_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X175 a_5141_4451# a_4782_4286# a_4780_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X176 VSS a_n3183_4389# a_n884_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 a_4190_3147# a_4104_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X178 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X179 a_10348_3230# a_9854_3147# a_9909_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X180 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X181 a_10446_4286# a_9854_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 a_640_3293# a_414_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X183 VDD a_11915_4389# a_25903_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X184 a_14216_4286# a_13850_3293# a_12230_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X185 VSS a_11915_4389# a_21231_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X186 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X187 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X188 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X189 a_9854_3147# a_9768_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X190 a_23656_4286# a_23064_3147# a_21670_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X191 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 a_17992_4286# a_17400_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X193 a_4684_3230# a_6304_3293# a_6128_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X194 VSS a_25446_3230# a_26371_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X195 a_13761_4451# a_13674_4353# a_13679_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X196 a_16102_3230# a_15512_3147# a_16006_3230# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X197 a_14216_4286# a_13624_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X198 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X199 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X200 VSS a_16006_3230# a_16931_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X201 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X202 a_17894_3230# a_17626_3293# a_17455_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X203 a_9555_3153# a_9385_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X204 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X205 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 VSS a_n3183_4389# a_n1419_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X207 IN a_n3136_3293# a_n3312_4353# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X208 a_14214_3230# a_13850_3293# a_14118_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X209 a_8558_4286# a_8192_3293# a_6572_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X210 a_2894_4286# a_2302_3147# a_908_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X211 VDD a_n3183_4389# a_4327_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X212 a_23654_3230# a_23064_3147# a_23558_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X213 VSS a_4684_3230# a_5609_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X214 a_19878_3230# a_19514_3293# a_19782_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X215 a_15213_3153# a_15043_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X216 VDD a_23558_3230# a_24483_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X217 a_10805_4451# a_10446_4286# a_10444_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X218 a_6133_4451# a_6128_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X219 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X220 a_2357_4451# a_2352_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X221 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X222 a_23064_3147# a_22978_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X223 a_n1337_4451# a_n1424_4353# a_n1419_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 a_2528_3293# a_2302_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X225 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X226 a_19514_3293# a_19288_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X227 a_14575_4451# a_14216_4286# a_14214_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X228 a_10446_4286# a_9854_3147# a_8460_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X229 a_13624_3147# a_13538_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X230 a_8556_3230# a_8192_3293# a_8460_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X231 VSS a_11915_4389# a_12326_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X232 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 a_23558_3230# a_25178_3293# a_25002_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X234 VDD a_11915_4389# a_16463_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X235 VDD a_2796_3230# a_3721_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X236 a_9555_3153# a_9385_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X237 a_14216_4286# a_13624_3147# a_12230_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X238 a_13325_3153# a_13155_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X239 a_14118_3230# a_15738_3293# a_15562_4353# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X240 a_3253_4451# a_2894_4286# a_2892_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X241 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 a_2302_3147# a_2216_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X243 a_17990_3230# a_17992_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X244 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X245 a_17400_3147# a_17314_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X246 a_18989_3153# a_18819_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X247 a_21670_3230# a_23064_3147# a_23114_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X248 a_12328_4286# a_11962_3293# a_10348_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X249 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X250 a_10444_3230# a_9854_3147# a_10348_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X251 a_21768_4286# a_21176_3147# a_19782_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X252 a_7966_3147# a_7880_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X253 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X254 VSS a_23558_3230# a_24483_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X255 a_2796_3230# a_4416_3293# a_4240_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X256 a_11873_4451# a_11786_4353# a_11791_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X257 a_25446_3230# a_25178_3293# a_25007_4451# VSS sky130_fd_pr__nfet_01v8 ad=2.145e+11p pd=1.96e+06u as=0p ps=0u w=650000u l=150000u
X258 VDD a_10348_3230# a_11273_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X259 a_12328_4286# a_11736_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X260 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X261 VDD a_n3183_4389# a_n523_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X262 a_25542_3230# a_25544_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X263 a_14214_3230# a_13624_3147# a_14118_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X264 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X265 a_25007_4451# a_25002_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X266 a_16006_3230# a_15738_3293# a_15567_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X267 a_7667_3153# a_7497_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X268 VDD a_11915_4389# a_13761_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X269 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X270 VSS a_n3183_4389# a_469_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X271 a_n882_4286# a_n1248_3293# a_n2868_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_4782_4286# a_4190_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X273 a_n2772_3230# a_n2770_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X274 a_12326_3230# a_11962_3293# a_12230_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X275 a_1006_4286# a_414_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X276 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X278 VDD a_10080_3293# a_9904_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X279 a_21766_3230# a_21176_3147# a_21670_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X280 VSS a_2796_3230# a_3721_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X281 a_9991_4451# a_9904_4353# a_9909_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X282 a_1006_4286# a_640_3293# a_n980_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X283 a_4684_3230# a_4416_3293# a_4245_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X284 a_n884_3230# a_n1248_3293# a_n980_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X285 a_13325_3153# a_13155_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X286 a_11962_3293# a_11736_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X287 VDD a_21670_3230# a_22595_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X288 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X289 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X290 a_4245_4451# a_4240_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X291 VDD a_n2868_3230# a_n1943_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X292 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X293 a_18989_3153# a_18819_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X294 a_21176_3147# a_21090_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X295 a_8460_3230# a_9854_3147# a_9904_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 VDD a_n3183_4389# a_10805_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X297 a_12687_4451# a_12328_4286# a_12326_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X298 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X299 a_6668_3230# a_6304_3293# a_6572_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X300 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X301 VSS a_10348_3230# a_11273_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X302 VDD a_11915_4389# a_18351_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X303 a_8192_3293# a_7966_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X304 a_1004_3230# a_640_3293# a_908_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X305 a_21670_3230# a_23290_3293# a_23114_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X306 VDD a_11915_4389# a_14575_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X307 a_16104_4286# a_15512_3147# a_14118_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X308 VDD a_908_3230# a_1833_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X309 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X310 VDD a_21402_3293# a_21226_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X311 a_7667_3153# a_7497_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X312 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X313 a_12328_4286# a_11736_3147# a_10348_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X314 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X315 a_n3307_4451# a_n3312_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X316 a_1365_4451# a_1006_4286# a_1004_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X317 VSS a_11915_4389# a_19343_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X318 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X319 VDD a_11962_3293# a_11786_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X320 a_16102_3230# a_16104_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X321 a_15512_3147# a_15426_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X322 a_23201_4451# a_23114_4353# a_23119_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X323 VDD a_n3183_4389# a_7029_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X324 a_19782_3230# a_21176_3147# a_21226_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X325 a_11736_3147# a_11650_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X326 a_14118_3230# a_13624_3147# a_13679_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X327 VSS a_n3183_4389# a_8556_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X328 VDD a_11915_4389# a_25089_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X329 a_908_3230# a_2528_3293# a_2352_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X330 VSS a_21670_3230# a_22595_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X331 a_23558_3230# a_23290_3293# a_23119_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X332 VSS a_n3183_4389# a_8021_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X333 a_23654_3230# a_23656_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X334 a_19880_4286# a_19514_3293# a_17894_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X335 a_4780_3230# a_4782_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X336 a_12326_3230# a_11736_3147# a_12230_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X337 VDD a_11915_4389# a_15649_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X338 a_4190_3147# a_4104_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X339 VSS a_n2868_3230# a_n1943_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X340 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X341 VDD a_11915_4389# a_11873_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X342 a_5779_3153# a_5609_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X343 a_n523_4451# a_n882_4286# a_n884_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X344 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X345 VDD a_12230_3230# a_13155_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X346 a_n3136_3293# a_n3362_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X347 a_2894_4286# a_2302_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X348 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X349 a_115_3153# a_n55_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X350 a_21670_3230# a_21176_3147# a_21231_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X351 a_23290_3293# a_23064_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X352 a_9854_3147# a_9768_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X353 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X354 a_13679_4451# a_13674_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X355 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X356 a_8460_3230# a_10080_3293# a_9904_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X357 a_13850_3293# a_13624_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X358 VSS a_908_3230# a_1833_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X359 a_n1474_3147# a_n1560_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X360 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X361 a_2796_3230# a_2528_3293# a_2357_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 a_8558_4286# a_7966_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X363 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X364 a_n2868_3230# a_n3136_3293# a_n3307_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X365 VDD a_19782_3230# a_20707_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X366 a_17626_3293# a_17400_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X367 a_12230_3230# a_13850_3293# a_13674_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X368 a_20239_4451# a_19880_4286# a_19878_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X369 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X370 VSS a_11915_4389# a_21766_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X371 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X372 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X373 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X374 a_10348_3230# a_10080_3293# a_9909_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X375 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X376 a_6304_3293# a_6078_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X377 VDD a_n980_3230# a_n55_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X378 a_19782_3230# a_21402_3293# a_21226_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X379 VDD a_11915_4389# a_12687_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X380 a_10348_3230# a_11736_3147# a_11786_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X381 a_10444_3230# a_10446_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X382 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X383 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X385 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X386 a_5779_3153# a_5609_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X387 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X388 a_23064_3147# a_22978_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X389 a_n1419_4451# a_n1424_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X390 VSS a_12230_3230# a_13155_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X391 a_14118_3230# a_13850_3293# a_13679_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X392 a_115_3153# a_n55_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X393 a_14214_3230# a_14216_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X394 a_19880_4286# a_19288_3147# a_17894_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X395 a_10080_3293# a_9854_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X396 a_21313_4451# a_21226_4353# a_21231_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X397 VDD RESET2 a_11915_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 a_13624_3147# a_13538_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X399 VDD a_640_3293# a_464_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X400 VDD a_n3183_4389# a_5141_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X401 a_21768_4286# a_21176_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X402 a_8917_4451# a_8558_4286# a_8556_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X403 VDD a_n3183_4389# a_1365_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X404 a_n1773_3153# a_n1943_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X405 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X406 VDD a_11915_4389# a_23201_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X407 VSS a_19782_3230# a_20707_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X408 a_12230_3230# a_11736_3147# a_11791_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X409 VSS a_n3183_4389# a_6133_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X410 a_21670_3230# a_21402_3293# a_21231_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X411 VDD a_n3136_3293# a_n3312_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X412 a_8558_4286# a_7966_3147# a_6572_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X413 a_17992_4286# a_17626_3293# a_16006_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X414 a_2892_3230# a_2894_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X415 a_2302_3147# a_2216_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X416 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X417 VDD a_14118_3230# a_15043_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X418 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X419 a_19878_3230# a_19288_3147# a_19782_3230# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X420 a_21402_3293# a_21176_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X421 a_7966_3147# a_7880_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X422 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 a_11791_4451# a_11786_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X424 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X425 VSS a_n980_3230# a_n55_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X426 a_n3362_3147# a_n3448_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X427 a_6670_4286# a_6304_3293# a_4684_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X428 VDD a_n3183_4389# a_2439_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X429 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X430 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X431 a_25178_3293# a_24952_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X432 a_6670_4286# a_6078_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X433 a_17990_3230# a_17626_3293# a_17894_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X434 a_19288_3147# a_19202_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X435 a_908_3230# a_414_3147# a_469_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X436 a_8556_3230# a_7966_3147# a_8460_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X437 a_n1248_3293# a_n1474_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X438 VSS a_11915_4389# a_17990_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X439 a_15738_3293# a_15512_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X440 a_22127_4451# a_21768_4286# a_21766_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X441 a_10348_3230# a_11962_3293# a_11786_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X442 VDD a_8460_3230# a_9385_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X443 VSS a_11915_4389# a_19878_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X444 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X445 a_n1773_3153# a_n1943_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X446 a_640_3293# a_414_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X447 VDD a_11915_4389# a_24015_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X448 a_9909_4451# a_9904_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X449 VDD a_19514_3293# a_19338_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X450 VDD a_n3183_4389# a_9991_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X451 VDD a_n3183_4389# a_n2411_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X452 VSS a_11915_4389# a_25542_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X453 a_12230_3230# a_13624_3147# a_13674_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X454 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X455 a_4416_3293# a_4190_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X456 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X457 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X458 VSS a_14118_3230# a_15043_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X459 a_21176_3147# a_21090_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X460 a_17894_3230# a_19288_3147# a_19338_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X461 a_17537_4451# a_17450_4353# a_17455_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X462 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X463 a_12230_3230# a_11962_3293# a_11791_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X464 OUT a_26371_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X465 VDD a_8192_3293# a_8016_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X466 a_n2770_4286# a_n3362_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X467 a_17992_4286# a_17400_3147# a_16006_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X468 a_12326_3230# a_12328_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X469 a_11915_4389# RESET2 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X470 VSS a_11915_4389# a_15567_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X471 VDD a_n3183_4389# a_3253_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X472 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X473 a_19880_4286# a_19288_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X474 a_7029_4451# a_6670_4286# a_6668_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X475 a_n2770_4286# a_n3362_3147# IN VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X476 a_25544_4286# a_25178_3293# a_23558_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X477 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X478 VDD a_11915_4389# a_21313_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X479 a_6572_3230# a_7966_3147# a_8016_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X480 IN a_n3362_3147# a_n3312_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X481 VDD a_n3183_4389# a_8917_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X482 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X483 VDD a_n1248_3293# a_n1424_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X484 a_1004_3230# a_1006_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X485 a_6670_4286# a_6078_3147# a_4684_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X486 a_551_4451# a_464_4353# a_469_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X487 a_n2772_3230# a_n3362_3147# a_n2868_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X488 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X489 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X490 a_19782_3230# a_19288_3147# a_19343_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X491 VSS a_8460_3230# a_9385_3153# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X492 a_23119_4451# a_23114_4353# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X493 a_1006_4286# a_414_3147# a_n980_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X494 a_n2868_3230# a_n3362_3147# a_n3307_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X495 a_17990_3230# a_17400_3147# a_17894_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X496 VSS RESET1 a_n3183_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X497 a_19514_3293# a_19288_3147# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X498 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X499 a_4782_4286# a_4416_3293# a_2796_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X500 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X501 a_25542_3230# a_25178_3293# a_25446_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X502 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X503 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X504 a_8460_3230# a_7966_3147# a_8021_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X505 VSS a_n3183_4389# a_n2772_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X506 a_n884_3230# a_n882_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X507 a_6668_3230# a_6078_3147# a_6572_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X508 OUT a_26371_3153# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X509 VSS a_11915_4389# a_16102_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X510 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X511 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X512 a_1004_3230# a_414_3147# a_908_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X513 VDD a_6572_3230# a_7497_3153# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X514 a_n3183_4389# RESET1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X515 VDD a_11915_4389# a_22127_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X516 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X517 a_n1474_3147# a_n1560_3299# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X518 VDD a_17626_3293# a_17450_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X519 a_6078_3147# a_5992_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X520 a_4780_3230# a_4416_3293# a_4684_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X521 a_11915_4389# RESET2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X522 a_2528_3293# a_2302_3147# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X523 a_24952_3147# a_24866_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X524 a_414_3147# a_328_3299# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X525 a_19878_3230# a_19880_4286# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X526 a_19425_4451# a_19338_4353# a_19343_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X527 a_16006_3230# a_17400_3147# a_17450_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X528 a_6572_3230# a_8192_3293# a_8016_4353# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X529 a_15649_4451# a_15562_4353# a_15567_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X530 VSS a_11915_4389# a_17455_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X531 a_24653_3153# a_24483_3153# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X532 VDD a_6304_3293# a_6128_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X533 VSS a_11915_4389# a_13679_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X534 a_19782_3230# a_19514_3293# a_19343_4451# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X535 a_n3183_4389# RESET1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X536 a_23656_4286# a_23290_3293# a_21670_3230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X537 a_8103_4451# a_8016_4353# a_8021_4451# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X538 a_4684_3230# a_6078_3147# a_6128_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X539 VSS RESET2 a_11915_4389# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X540 a_n980_3230# a_414_3147# a_464_4353# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X541 a_4782_4286# a_4190_3147# a_2796_3230# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X542 VDD RESET1 a_n3183_4389# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X543 a_25542_3230# a_24952_3147# a_25446_3230# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

