magic
tech sky130A
magscale 1 2
timestamp 1654151355
<< nwell >>
rect -3374 4412 -2206 4746
rect -1486 4412 -318 4746
rect 402 4412 1570 4746
rect 2074 4740 3622 5061
rect 2290 4412 3458 4740
rect 3956 4738 5504 5059
rect 4178 4412 5346 4738
rect 6066 4412 7234 4746
rect 7954 4412 9122 4746
rect 9842 4412 11010 4746
rect 11724 4412 12892 4746
rect 13612 4412 14780 4746
rect 15500 4412 16668 4746
rect 17172 4740 18720 5061
rect 17388 4412 18556 4740
rect 19054 4738 20602 5059
rect 19276 4412 20444 4738
rect 21164 4412 22332 4746
rect 23052 4412 24220 4746
rect 24940 4412 26108 4746
rect -2994 4224 -2672 4412
rect -2994 4186 -2768 4224
rect -1106 4224 -784 4412
rect -1106 4186 -880 4224
rect 782 4224 1104 4412
rect 782 4186 1008 4224
rect 2670 4224 2992 4412
rect 2670 4186 2896 4224
rect 4558 4224 4880 4412
rect 4558 4186 4784 4224
rect 6446 4224 6768 4412
rect 6446 4186 6672 4224
rect 8334 4224 8656 4412
rect 8334 4186 8560 4224
rect 10222 4224 10544 4412
rect 10222 4186 10448 4224
rect 12104 4224 12426 4412
rect 12104 4186 12330 4224
rect 13992 4224 14314 4412
rect 13992 4186 14218 4224
rect 15880 4224 16202 4412
rect 15880 4186 16106 4224
rect 17768 4224 18090 4412
rect 17768 4186 17994 4224
rect 19656 4224 19978 4412
rect 19656 4186 19882 4224
rect 21544 4224 21866 4412
rect 21544 4186 21770 4224
rect 23432 4224 23754 4412
rect 23432 4186 23658 4224
rect 25320 4224 25642 4412
rect 25320 4186 25546 4224
rect -3212 3688 -2002 3690
rect -1324 3688 -114 3690
rect 564 3688 1774 3690
rect 2452 3688 3662 3690
rect 4340 3688 5550 3690
rect 6228 3688 7438 3690
rect 8116 3688 9326 3690
rect 10004 3688 11214 3690
rect 11886 3688 13096 3690
rect 13774 3688 14984 3690
rect 15662 3688 16872 3690
rect 17550 3688 18760 3690
rect 19438 3688 20648 3690
rect 21326 3688 22536 3690
rect 23214 3688 24424 3690
rect 25102 3688 26312 3690
rect -3212 3682 -1656 3688
rect -1324 3682 232 3688
rect 564 3682 2120 3688
rect 2452 3682 4008 3688
rect 4340 3682 5896 3688
rect 6228 3682 7784 3688
rect 8116 3682 9672 3688
rect 10004 3682 11560 3688
rect 11886 3682 13442 3688
rect 13774 3682 15330 3688
rect 15662 3682 17218 3688
rect 17550 3682 19106 3688
rect 19438 3682 20994 3688
rect 21326 3682 22882 3688
rect 23214 3682 24770 3688
rect 25102 3682 26658 3688
rect -3550 3369 26658 3682
rect -3550 3361 -2348 3369
rect -2008 3367 -460 3369
rect -120 3367 1428 3369
rect 1768 3367 3316 3369
rect 3656 3367 5204 3369
rect 5544 3367 7092 3369
rect 7432 3367 8980 3369
rect 9320 3367 10868 3369
rect 11208 3367 12750 3369
rect 13090 3367 14638 3369
rect 14978 3367 16526 3369
rect 16866 3367 18414 3369
rect 18754 3367 20302 3369
rect 20642 3367 22190 3369
rect 22530 3367 24078 3369
rect 24418 3367 25966 3369
rect 26306 3367 26658 3369
rect -1662 3361 -460 3367
rect 226 3361 1428 3367
rect 2114 3361 3316 3367
rect 4002 3361 5204 3367
rect 5890 3361 7092 3367
rect 7778 3361 8980 3367
rect 9666 3361 10868 3367
rect 11548 3361 12750 3367
rect 13436 3361 14638 3367
rect 15324 3361 16526 3367
rect 17212 3361 18414 3367
rect 19100 3361 20302 3367
rect 20988 3361 22190 3367
rect 22876 3361 24078 3367
rect 24764 3361 25966 3367
rect -3212 3290 -2348 3361
rect -2996 3168 -2674 3290
rect -2996 3130 -2770 3168
rect -1324 3290 -460 3361
rect -1108 3168 -786 3290
rect -1108 3130 -882 3168
rect 564 3290 1428 3361
rect 780 3168 1102 3290
rect 780 3130 1006 3168
rect 2452 3290 3316 3361
rect 2668 3168 2990 3290
rect 2668 3130 2894 3168
rect 4340 3290 5204 3361
rect 4556 3168 4878 3290
rect 4556 3130 4782 3168
rect 6228 3290 7092 3361
rect 6444 3168 6766 3290
rect 6444 3130 6670 3168
rect 8116 3290 8980 3361
rect 8332 3168 8654 3290
rect 8332 3130 8558 3168
rect 10004 3290 10868 3361
rect 10220 3168 10542 3290
rect 10220 3130 10446 3168
rect 11886 3290 12750 3361
rect 12102 3168 12424 3290
rect 12102 3130 12328 3168
rect 13774 3290 14638 3361
rect 13990 3168 14312 3290
rect 13990 3130 14216 3168
rect 15662 3290 16526 3361
rect 15878 3168 16200 3290
rect 15878 3130 16104 3168
rect 17550 3290 18414 3361
rect 17766 3168 18088 3290
rect 17766 3130 17992 3168
rect 19438 3290 20302 3361
rect 19654 3168 19976 3290
rect 19654 3130 19880 3168
rect 21326 3290 22190 3361
rect 21542 3168 21864 3290
rect 21542 3130 21768 3168
rect 23214 3290 24078 3361
rect 23430 3168 23752 3290
rect 23430 3130 23656 3168
rect 25102 3290 25966 3361
rect 25318 3168 25640 3290
rect 25318 3130 25544 3168
<< pwell >>
rect 2126 5119 3572 5301
rect 4008 5117 5454 5299
rect 17224 5119 18670 5301
rect 19106 5117 20552 5299
rect -3333 4175 -3063 4357
rect -2519 4175 -2249 4357
rect -1445 4175 -1175 4357
rect -631 4175 -361 4357
rect 443 4175 713 4357
rect 1257 4175 1527 4357
rect 2331 4175 2601 4357
rect 3145 4175 3415 4357
rect 4219 4175 4489 4357
rect 5033 4175 5303 4357
rect 6107 4175 6377 4357
rect 6921 4175 7191 4357
rect 7995 4175 8265 4357
rect 8809 4175 9079 4357
rect 9883 4175 10153 4357
rect 10697 4175 10967 4357
rect 11765 4175 12035 4357
rect 12579 4175 12849 4357
rect 13653 4175 13923 4357
rect 14467 4175 14737 4357
rect 15541 4175 15811 4357
rect 16355 4175 16625 4357
rect 17429 4175 17699 4357
rect 18243 4175 18513 4357
rect 19317 4175 19587 4357
rect 20131 4175 20401 4357
rect 21205 4175 21475 4357
rect 22019 4175 22289 4357
rect 23093 4175 23363 4357
rect 23907 4175 24177 4357
rect 24981 4175 25251 4357
rect 25795 4175 26065 4357
rect -2968 3930 -2666 4112
rect -1080 3930 -778 4112
rect 808 3930 1110 4112
rect 2696 3930 2998 4112
rect 4584 3930 4886 4112
rect 6472 3930 6774 4112
rect 8360 3930 8662 4112
rect 10248 3930 10550 4112
rect 12130 3930 12432 4112
rect 14018 3930 14320 4112
rect 15906 3930 16208 4112
rect 17794 3930 18096 4112
rect 19682 3930 19984 4112
rect 21570 3930 21872 4112
rect 23458 3930 23760 4112
rect 25346 3930 25648 4112
rect -2924 3746 -2712 3846
rect -1036 3746 -824 3846
rect 852 3746 1064 3846
rect 2740 3746 2952 3846
rect 4628 3746 4840 3846
rect 6516 3746 6728 3846
rect 8404 3746 8616 3846
rect 10292 3746 10504 3846
rect 12174 3746 12386 3846
rect 14062 3746 14274 3846
rect 15950 3746 16162 3846
rect 17838 3746 18050 3846
rect 19726 3746 19938 3846
rect 21614 3746 21826 3846
rect 23502 3746 23714 3846
rect 25390 3746 25602 3846
rect -3470 3121 -3284 3303
rect -2274 3129 -2088 3311
rect -1969 3127 -1695 3283
rect -1582 3121 -1396 3303
rect -386 3129 -200 3311
rect -81 3127 193 3283
rect 306 3121 492 3303
rect 1502 3129 1688 3311
rect 1807 3127 2081 3283
rect 2194 3121 2380 3303
rect 3390 3129 3576 3311
rect 3695 3127 3969 3283
rect 4082 3121 4268 3303
rect 5278 3129 5464 3311
rect 5583 3127 5857 3283
rect 5970 3121 6156 3303
rect 7166 3129 7352 3311
rect 7471 3127 7745 3283
rect 7858 3121 8044 3303
rect 9054 3129 9240 3311
rect 9359 3127 9633 3283
rect 9746 3121 9932 3303
rect 10942 3129 11128 3311
rect 11247 3127 11521 3283
rect 11628 3121 11814 3303
rect 12824 3129 13010 3311
rect 13129 3127 13403 3283
rect 13516 3121 13702 3303
rect 14712 3129 14898 3311
rect 15017 3127 15291 3283
rect 15404 3121 15590 3303
rect 16600 3129 16786 3311
rect 16905 3127 17179 3283
rect 17292 3121 17478 3303
rect 18488 3129 18674 3311
rect 18793 3127 19067 3283
rect 19180 3121 19366 3303
rect 20376 3129 20562 3311
rect 20681 3127 20955 3283
rect 21068 3121 21254 3303
rect 22264 3129 22450 3311
rect 22569 3127 22843 3283
rect 22956 3121 23142 3303
rect 24152 3129 24338 3311
rect 24457 3127 24731 3283
rect 24844 3121 25030 3303
rect 26040 3129 26226 3311
rect 26345 3127 26619 3283
rect -2970 2874 -2668 3056
rect -1082 2874 -780 3056
rect 806 2874 1108 3056
rect 2694 2874 2996 3056
rect 4582 2874 4884 3056
rect 6470 2874 6772 3056
rect 8358 2874 8660 3056
rect 10246 2874 10548 3056
rect 12128 2874 12430 3056
rect 14016 2874 14318 3056
rect 15904 2874 16206 3056
rect 17792 2874 18094 3056
rect 19680 2874 19982 3056
rect 21568 2874 21870 3056
rect 23456 2874 23758 3056
rect 25344 2874 25646 3056
rect -2926 2690 -2714 2790
rect -1038 2690 -826 2790
rect 850 2690 1062 2790
rect 2738 2690 2950 2790
rect 4626 2690 4838 2790
rect 6514 2690 6726 2790
rect 8402 2690 8614 2790
rect 10290 2690 10502 2790
rect 12172 2690 12384 2790
rect 14060 2690 14272 2790
rect 15948 2690 16160 2790
rect 17836 2690 18048 2790
rect 19724 2690 19936 2790
rect 21612 2690 21824 2790
rect 23500 2690 23712 2790
rect 25388 2690 25600 2790
<< nmos >>
rect -2880 3956 -2850 4086
rect -2784 3956 -2754 4086
rect -992 3956 -962 4086
rect -896 3956 -866 4086
rect 896 3956 926 4086
rect 992 3956 1022 4086
rect 2784 3956 2814 4086
rect 2880 3956 2910 4086
rect 4672 3956 4702 4086
rect 4768 3956 4798 4086
rect 6560 3956 6590 4086
rect 6656 3956 6686 4086
rect 8448 3956 8478 4086
rect 8544 3956 8574 4086
rect 10336 3956 10366 4086
rect 10432 3956 10462 4086
rect 12218 3956 12248 4086
rect 12314 3956 12344 4086
rect 14106 3956 14136 4086
rect 14202 3956 14232 4086
rect 15994 3956 16024 4086
rect 16090 3956 16120 4086
rect 17882 3956 17912 4086
rect 17978 3956 18008 4086
rect 19770 3956 19800 4086
rect 19866 3956 19896 4086
rect 21658 3956 21688 4086
rect 21754 3956 21784 4086
rect 23546 3956 23576 4086
rect 23642 3956 23672 4086
rect 25434 3956 25464 4086
rect 25530 3956 25560 4086
rect -2882 2900 -2852 3030
rect -2786 2900 -2756 3030
rect -994 2900 -964 3030
rect -898 2900 -868 3030
rect 894 2900 924 3030
rect 990 2900 1020 3030
rect 2782 2900 2812 3030
rect 2878 2900 2908 3030
rect 4670 2900 4700 3030
rect 4766 2900 4796 3030
rect 6558 2900 6588 3030
rect 6654 2900 6684 3030
rect 8446 2900 8476 3030
rect 8542 2900 8572 3030
rect 10334 2900 10364 3030
rect 10430 2900 10460 3030
rect 12216 2900 12246 3030
rect 12312 2900 12342 3030
rect 14104 2900 14134 3030
rect 14200 2900 14230 3030
rect 15992 2900 16022 3030
rect 16088 2900 16118 3030
rect 17880 2900 17910 3030
rect 17976 2900 18006 3030
rect 19768 2900 19798 3030
rect 19864 2900 19894 3030
rect 21656 2900 21686 3030
rect 21752 2900 21782 3030
rect 23544 2900 23574 3030
rect 23640 2900 23670 3030
rect 25432 2900 25462 3030
rect 25528 2900 25558 3030
<< scnmos >>
rect 2204 5145 2234 5275
rect 2288 5145 2318 5275
rect 2372 5145 2402 5275
rect 2456 5145 2486 5275
rect 2540 5145 2570 5275
rect 2624 5145 2654 5275
rect 2708 5145 2738 5275
rect 2792 5145 2822 5275
rect 2876 5145 2906 5275
rect 2960 5145 2990 5275
rect 3044 5145 3074 5275
rect 3128 5145 3158 5275
rect 3212 5145 3242 5275
rect 3296 5145 3326 5275
rect 3380 5145 3410 5275
rect 3464 5145 3494 5275
rect 4086 5143 4116 5273
rect 4170 5143 4200 5273
rect 4254 5143 4284 5273
rect 4338 5143 4368 5273
rect 4422 5143 4452 5273
rect 4506 5143 4536 5273
rect 4590 5143 4620 5273
rect 4674 5143 4704 5273
rect 4758 5143 4788 5273
rect 4842 5143 4872 5273
rect 4926 5143 4956 5273
rect 5010 5143 5040 5273
rect 5094 5143 5124 5273
rect 5178 5143 5208 5273
rect 5262 5143 5292 5273
rect 5346 5143 5376 5273
rect 17302 5145 17332 5275
rect 17386 5145 17416 5275
rect 17470 5145 17500 5275
rect 17554 5145 17584 5275
rect 17638 5145 17668 5275
rect 17722 5145 17752 5275
rect 17806 5145 17836 5275
rect 17890 5145 17920 5275
rect 17974 5145 18004 5275
rect 18058 5145 18088 5275
rect 18142 5145 18172 5275
rect 18226 5145 18256 5275
rect 18310 5145 18340 5275
rect 18394 5145 18424 5275
rect 18478 5145 18508 5275
rect 18562 5145 18592 5275
rect 19184 5143 19214 5273
rect 19268 5143 19298 5273
rect 19352 5143 19382 5273
rect 19436 5143 19466 5273
rect 19520 5143 19550 5273
rect 19604 5143 19634 5273
rect 19688 5143 19718 5273
rect 19772 5143 19802 5273
rect 19856 5143 19886 5273
rect 19940 5143 19970 5273
rect 20024 5143 20054 5273
rect 20108 5143 20138 5273
rect 20192 5143 20222 5273
rect 20276 5143 20306 5273
rect 20360 5143 20390 5273
rect 20444 5143 20474 5273
rect -3255 4201 -3225 4331
rect -3171 4201 -3141 4331
rect -2441 4201 -2411 4331
rect -2357 4201 -2327 4331
rect -1367 4201 -1337 4331
rect -1283 4201 -1253 4331
rect -553 4201 -523 4331
rect -469 4201 -439 4331
rect 521 4201 551 4331
rect 605 4201 635 4331
rect 1335 4201 1365 4331
rect 1419 4201 1449 4331
rect 2409 4201 2439 4331
rect 2493 4201 2523 4331
rect 3223 4201 3253 4331
rect 3307 4201 3337 4331
rect 4297 4201 4327 4331
rect 4381 4201 4411 4331
rect 5111 4201 5141 4331
rect 5195 4201 5225 4331
rect 6185 4201 6215 4331
rect 6269 4201 6299 4331
rect 6999 4201 7029 4331
rect 7083 4201 7113 4331
rect 8073 4201 8103 4331
rect 8157 4201 8187 4331
rect 8887 4201 8917 4331
rect 8971 4201 9001 4331
rect 9961 4201 9991 4331
rect 10045 4201 10075 4331
rect 10775 4201 10805 4331
rect 10859 4201 10889 4331
rect 11843 4201 11873 4331
rect 11927 4201 11957 4331
rect 12657 4201 12687 4331
rect 12741 4201 12771 4331
rect 13731 4201 13761 4331
rect 13815 4201 13845 4331
rect 14545 4201 14575 4331
rect 14629 4201 14659 4331
rect 15619 4201 15649 4331
rect 15703 4201 15733 4331
rect 16433 4201 16463 4331
rect 16517 4201 16547 4331
rect 17507 4201 17537 4331
rect 17591 4201 17621 4331
rect 18321 4201 18351 4331
rect 18405 4201 18435 4331
rect 19395 4201 19425 4331
rect 19479 4201 19509 4331
rect 20209 4201 20239 4331
rect 20293 4201 20323 4331
rect 21283 4201 21313 4331
rect 21367 4201 21397 4331
rect 22097 4201 22127 4331
rect 22181 4201 22211 4331
rect 23171 4201 23201 4331
rect 23255 4201 23285 4331
rect 23985 4201 24015 4331
rect 24069 4201 24099 4331
rect 25059 4201 25089 4331
rect 25143 4201 25173 4331
rect 25873 4201 25903 4331
rect 25957 4201 25987 4331
rect -3392 3147 -3362 3277
rect -2196 3155 -2166 3285
rect -1891 3153 -1861 3257
rect -1803 3153 -1773 3257
rect -1504 3147 -1474 3277
rect -308 3155 -278 3285
rect -3 3153 27 3257
rect 85 3153 115 3257
rect 384 3147 414 3277
rect 1580 3155 1610 3285
rect 1885 3153 1915 3257
rect 1973 3153 2003 3257
rect 2272 3147 2302 3277
rect 3468 3155 3498 3285
rect 3773 3153 3803 3257
rect 3861 3153 3891 3257
rect 4160 3147 4190 3277
rect 5356 3155 5386 3285
rect 5661 3153 5691 3257
rect 5749 3153 5779 3257
rect 6048 3147 6078 3277
rect 7244 3155 7274 3285
rect 7549 3153 7579 3257
rect 7637 3153 7667 3257
rect 7936 3147 7966 3277
rect 9132 3155 9162 3285
rect 9437 3153 9467 3257
rect 9525 3153 9555 3257
rect 9824 3147 9854 3277
rect 11020 3155 11050 3285
rect 11325 3153 11355 3257
rect 11413 3153 11443 3257
rect 11706 3147 11736 3277
rect 12902 3155 12932 3285
rect 13207 3153 13237 3257
rect 13295 3153 13325 3257
rect 13594 3147 13624 3277
rect 14790 3155 14820 3285
rect 15095 3153 15125 3257
rect 15183 3153 15213 3257
rect 15482 3147 15512 3277
rect 16678 3155 16708 3285
rect 16983 3153 17013 3257
rect 17071 3153 17101 3257
rect 17370 3147 17400 3277
rect 18566 3155 18596 3285
rect 18871 3153 18901 3257
rect 18959 3153 18989 3257
rect 19258 3147 19288 3277
rect 20454 3155 20484 3285
rect 20759 3153 20789 3257
rect 20847 3153 20877 3257
rect 21146 3147 21176 3277
rect 22342 3155 22372 3285
rect 22647 3153 22677 3257
rect 22735 3153 22765 3257
rect 23034 3147 23064 3277
rect 24230 3155 24260 3285
rect 24535 3153 24565 3257
rect 24623 3153 24653 3257
rect 24922 3147 24952 3277
rect 26118 3155 26148 3285
rect 26423 3153 26453 3257
rect 26511 3153 26541 3257
<< scpmoshvt >>
rect 2204 4825 2234 5025
rect 2288 4825 2318 5025
rect 2372 4825 2402 5025
rect 2456 4825 2486 5025
rect 2540 4825 2570 5025
rect 2624 4825 2654 5025
rect 2708 4825 2738 5025
rect 2792 4825 2822 5025
rect 2876 4825 2906 5025
rect 2960 4825 2990 5025
rect 3044 4825 3074 5025
rect 3128 4825 3158 5025
rect 3212 4825 3242 5025
rect 3296 4825 3326 5025
rect 3380 4825 3410 5025
rect 3464 4825 3494 5025
rect 4086 4823 4116 5023
rect 4170 4823 4200 5023
rect 4254 4823 4284 5023
rect 4338 4823 4368 5023
rect 4422 4823 4452 5023
rect 4506 4823 4536 5023
rect 4590 4823 4620 5023
rect 4674 4823 4704 5023
rect 4758 4823 4788 5023
rect 4842 4823 4872 5023
rect 4926 4823 4956 5023
rect 5010 4823 5040 5023
rect 5094 4823 5124 5023
rect 5178 4823 5208 5023
rect 5262 4823 5292 5023
rect 5346 4823 5376 5023
rect 17302 4825 17332 5025
rect 17386 4825 17416 5025
rect 17470 4825 17500 5025
rect 17554 4825 17584 5025
rect 17638 4825 17668 5025
rect 17722 4825 17752 5025
rect 17806 4825 17836 5025
rect 17890 4825 17920 5025
rect 17974 4825 18004 5025
rect 18058 4825 18088 5025
rect 18142 4825 18172 5025
rect 18226 4825 18256 5025
rect 18310 4825 18340 5025
rect 18394 4825 18424 5025
rect 18478 4825 18508 5025
rect 18562 4825 18592 5025
rect 19184 4823 19214 5023
rect 19268 4823 19298 5023
rect 19352 4823 19382 5023
rect 19436 4823 19466 5023
rect 19520 4823 19550 5023
rect 19604 4823 19634 5023
rect 19688 4823 19718 5023
rect 19772 4823 19802 5023
rect 19856 4823 19886 5023
rect 19940 4823 19970 5023
rect 20024 4823 20054 5023
rect 20108 4823 20138 5023
rect 20192 4823 20222 5023
rect 20276 4823 20306 5023
rect 20360 4823 20390 5023
rect 20444 4823 20474 5023
rect -3255 4451 -3225 4651
rect -3183 4451 -3153 4651
rect -2441 4451 -2411 4651
rect -2369 4451 -2339 4651
rect -1367 4451 -1337 4651
rect -1295 4451 -1265 4651
rect -553 4451 -523 4651
rect -481 4451 -451 4651
rect 521 4451 551 4651
rect 593 4451 623 4651
rect 1335 4451 1365 4651
rect 1407 4451 1437 4651
rect 2409 4451 2439 4651
rect 2481 4451 2511 4651
rect 3223 4451 3253 4651
rect 3295 4451 3325 4651
rect 4297 4451 4327 4651
rect 4369 4451 4399 4651
rect 5111 4451 5141 4651
rect 5183 4451 5213 4651
rect 6185 4451 6215 4651
rect 6257 4451 6287 4651
rect 6999 4451 7029 4651
rect 7071 4451 7101 4651
rect 8073 4451 8103 4651
rect 8145 4451 8175 4651
rect 8887 4451 8917 4651
rect 8959 4451 8989 4651
rect 9961 4451 9991 4651
rect 10033 4451 10063 4651
rect 10775 4451 10805 4651
rect 10847 4451 10877 4651
rect 11843 4451 11873 4651
rect 11915 4451 11945 4651
rect 12657 4451 12687 4651
rect 12729 4451 12759 4651
rect 13731 4451 13761 4651
rect 13803 4451 13833 4651
rect 14545 4451 14575 4651
rect 14617 4451 14647 4651
rect 15619 4451 15649 4651
rect 15691 4451 15721 4651
rect 16433 4451 16463 4651
rect 16505 4451 16535 4651
rect 17507 4451 17537 4651
rect 17579 4451 17609 4651
rect 18321 4451 18351 4651
rect 18393 4451 18423 4651
rect 19395 4451 19425 4651
rect 19467 4451 19497 4651
rect 20209 4451 20239 4651
rect 20281 4451 20311 4651
rect 21283 4451 21313 4651
rect 21355 4451 21385 4651
rect 22097 4451 22127 4651
rect 22169 4451 22199 4651
rect 23171 4451 23201 4651
rect 23243 4451 23273 4651
rect 23985 4451 24015 4651
rect 24057 4451 24087 4651
rect 25059 4451 25089 4651
rect 25131 4451 25161 4651
rect 25873 4451 25903 4651
rect 25945 4451 25975 4651
rect -3392 3397 -3362 3597
rect -2196 3405 -2166 3605
rect -1891 3445 -1861 3603
rect -1803 3445 -1773 3603
rect -1504 3397 -1474 3597
rect -308 3405 -278 3605
rect -3 3445 27 3603
rect 85 3445 115 3603
rect 384 3397 414 3597
rect 1580 3405 1610 3605
rect 1885 3445 1915 3603
rect 1973 3445 2003 3603
rect 2272 3397 2302 3597
rect 3468 3405 3498 3605
rect 3773 3445 3803 3603
rect 3861 3445 3891 3603
rect 4160 3397 4190 3597
rect 5356 3405 5386 3605
rect 5661 3445 5691 3603
rect 5749 3445 5779 3603
rect 6048 3397 6078 3597
rect 7244 3405 7274 3605
rect 7549 3445 7579 3603
rect 7637 3445 7667 3603
rect 7936 3397 7966 3597
rect 9132 3405 9162 3605
rect 9437 3445 9467 3603
rect 9525 3445 9555 3603
rect 9824 3397 9854 3597
rect 11020 3405 11050 3605
rect 11325 3445 11355 3603
rect 11413 3445 11443 3603
rect 11706 3397 11736 3597
rect 12902 3405 12932 3605
rect 13207 3445 13237 3603
rect 13295 3445 13325 3603
rect 13594 3397 13624 3597
rect 14790 3405 14820 3605
rect 15095 3445 15125 3603
rect 15183 3445 15213 3603
rect 15482 3397 15512 3597
rect 16678 3405 16708 3605
rect 16983 3445 17013 3603
rect 17071 3445 17101 3603
rect 17370 3397 17400 3597
rect 18566 3405 18596 3605
rect 18871 3445 18901 3603
rect 18959 3445 18989 3603
rect 19258 3397 19288 3597
rect 20454 3405 20484 3605
rect 20759 3445 20789 3603
rect 20847 3445 20877 3603
rect 21146 3397 21176 3597
rect 22342 3405 22372 3605
rect 22647 3445 22677 3603
rect 22735 3445 22765 3603
rect 23034 3397 23064 3597
rect 24230 3405 24260 3605
rect 24535 3445 24565 3603
rect 24623 3445 24653 3603
rect 24922 3397 24952 3597
rect 26118 3405 26148 3605
rect 26423 3445 26453 3603
rect 26511 3445 26541 3603
<< pmoshvt >>
rect -2896 4286 -2866 4486
rect -2800 4286 -2770 4486
rect -1008 4286 -978 4486
rect -912 4286 -882 4486
rect 880 4286 910 4486
rect 976 4286 1006 4486
rect 2768 4286 2798 4486
rect 2864 4286 2894 4486
rect 4656 4286 4686 4486
rect 4752 4286 4782 4486
rect 6544 4286 6574 4486
rect 6640 4286 6670 4486
rect 8432 4286 8462 4486
rect 8528 4286 8558 4486
rect 10320 4286 10350 4486
rect 10416 4286 10446 4486
rect 12202 4286 12232 4486
rect 12298 4286 12328 4486
rect 14090 4286 14120 4486
rect 14186 4286 14216 4486
rect 15978 4286 16008 4486
rect 16074 4286 16104 4486
rect 17866 4286 17896 4486
rect 17962 4286 17992 4486
rect 19754 4286 19784 4486
rect 19850 4286 19880 4486
rect 21642 4286 21672 4486
rect 21738 4286 21768 4486
rect 23530 4286 23560 4486
rect 23626 4286 23656 4486
rect 25418 4286 25448 4486
rect 25514 4286 25544 4486
rect -3118 3390 -3088 3590
rect -2898 3230 -2868 3430
rect -2802 3230 -2772 3430
rect -2472 3390 -2442 3590
rect -1230 3390 -1200 3590
rect -1010 3230 -980 3430
rect -914 3230 -884 3430
rect -584 3390 -554 3590
rect 658 3390 688 3590
rect 878 3230 908 3430
rect 974 3230 1004 3430
rect 1304 3390 1334 3590
rect 2546 3390 2576 3590
rect 2766 3230 2796 3430
rect 2862 3230 2892 3430
rect 3192 3390 3222 3590
rect 4434 3390 4464 3590
rect 4654 3230 4684 3430
rect 4750 3230 4780 3430
rect 5080 3390 5110 3590
rect 6322 3390 6352 3590
rect 6542 3230 6572 3430
rect 6638 3230 6668 3430
rect 6968 3390 6998 3590
rect 8210 3390 8240 3590
rect 8430 3230 8460 3430
rect 8526 3230 8556 3430
rect 8856 3390 8886 3590
rect 10098 3390 10128 3590
rect 10318 3230 10348 3430
rect 10414 3230 10444 3430
rect 10744 3390 10774 3590
rect 11980 3390 12010 3590
rect 12200 3230 12230 3430
rect 12296 3230 12326 3430
rect 12626 3390 12656 3590
rect 13868 3390 13898 3590
rect 14088 3230 14118 3430
rect 14184 3230 14214 3430
rect 14514 3390 14544 3590
rect 15756 3390 15786 3590
rect 15976 3230 16006 3430
rect 16072 3230 16102 3430
rect 16402 3390 16432 3590
rect 17644 3390 17674 3590
rect 17864 3230 17894 3430
rect 17960 3230 17990 3430
rect 18290 3390 18320 3590
rect 19532 3390 19562 3590
rect 19752 3230 19782 3430
rect 19848 3230 19878 3430
rect 20178 3390 20208 3590
rect 21420 3390 21450 3590
rect 21640 3230 21670 3430
rect 21736 3230 21766 3430
rect 22066 3390 22096 3590
rect 23308 3390 23338 3590
rect 23528 3230 23558 3430
rect 23624 3230 23654 3430
rect 23954 3390 23984 3590
rect 25196 3390 25226 3590
rect 25416 3230 25446 3430
rect 25512 3230 25542 3430
rect 25842 3390 25872 3590
<< ndiff >>
rect 2152 5263 2204 5275
rect 2152 5229 2160 5263
rect 2194 5229 2204 5263
rect 2152 5195 2204 5229
rect 2152 5161 2160 5195
rect 2194 5161 2204 5195
rect 2152 5145 2204 5161
rect 2234 5263 2288 5275
rect 2234 5229 2244 5263
rect 2278 5229 2288 5263
rect 2234 5195 2288 5229
rect 2234 5161 2244 5195
rect 2278 5161 2288 5195
rect 2234 5145 2288 5161
rect 2318 5263 2372 5275
rect 2318 5229 2328 5263
rect 2362 5229 2372 5263
rect 2318 5145 2372 5229
rect 2402 5263 2456 5275
rect 2402 5229 2412 5263
rect 2446 5229 2456 5263
rect 2402 5195 2456 5229
rect 2402 5161 2412 5195
rect 2446 5161 2456 5195
rect 2402 5145 2456 5161
rect 2486 5263 2540 5275
rect 2486 5229 2496 5263
rect 2530 5229 2540 5263
rect 2486 5145 2540 5229
rect 2570 5263 2624 5275
rect 2570 5229 2580 5263
rect 2614 5229 2624 5263
rect 2570 5195 2624 5229
rect 2570 5161 2580 5195
rect 2614 5161 2624 5195
rect 2570 5145 2624 5161
rect 2654 5263 2708 5275
rect 2654 5229 2664 5263
rect 2698 5229 2708 5263
rect 2654 5145 2708 5229
rect 2738 5263 2792 5275
rect 2738 5229 2748 5263
rect 2782 5229 2792 5263
rect 2738 5195 2792 5229
rect 2738 5161 2748 5195
rect 2782 5161 2792 5195
rect 2738 5145 2792 5161
rect 2822 5263 2876 5275
rect 2822 5229 2832 5263
rect 2866 5229 2876 5263
rect 2822 5145 2876 5229
rect 2906 5263 2960 5275
rect 2906 5229 2916 5263
rect 2950 5229 2960 5263
rect 2906 5195 2960 5229
rect 2906 5161 2916 5195
rect 2950 5161 2960 5195
rect 2906 5145 2960 5161
rect 2990 5263 3044 5275
rect 2990 5229 3000 5263
rect 3034 5229 3044 5263
rect 2990 5145 3044 5229
rect 3074 5263 3128 5275
rect 3074 5229 3084 5263
rect 3118 5229 3128 5263
rect 3074 5195 3128 5229
rect 3074 5161 3084 5195
rect 3118 5161 3128 5195
rect 3074 5145 3128 5161
rect 3158 5263 3212 5275
rect 3158 5229 3168 5263
rect 3202 5229 3212 5263
rect 3158 5145 3212 5229
rect 3242 5263 3296 5275
rect 3242 5229 3252 5263
rect 3286 5229 3296 5263
rect 3242 5195 3296 5229
rect 3242 5161 3252 5195
rect 3286 5161 3296 5195
rect 3242 5145 3296 5161
rect 3326 5263 3380 5275
rect 3326 5229 3336 5263
rect 3370 5229 3380 5263
rect 3326 5145 3380 5229
rect 3410 5263 3464 5275
rect 3410 5229 3420 5263
rect 3454 5229 3464 5263
rect 3410 5195 3464 5229
rect 3410 5161 3420 5195
rect 3454 5161 3464 5195
rect 3410 5145 3464 5161
rect 3494 5263 3546 5275
rect 3494 5229 3504 5263
rect 3538 5229 3546 5263
rect 3494 5195 3546 5229
rect 3494 5161 3504 5195
rect 3538 5161 3546 5195
rect 3494 5145 3546 5161
rect 4034 5261 4086 5273
rect 4034 5227 4042 5261
rect 4076 5227 4086 5261
rect 4034 5193 4086 5227
rect 4034 5159 4042 5193
rect 4076 5159 4086 5193
rect 4034 5143 4086 5159
rect 4116 5261 4170 5273
rect 4116 5227 4126 5261
rect 4160 5227 4170 5261
rect 4116 5193 4170 5227
rect 4116 5159 4126 5193
rect 4160 5159 4170 5193
rect 4116 5143 4170 5159
rect 4200 5261 4254 5273
rect 4200 5227 4210 5261
rect 4244 5227 4254 5261
rect 4200 5143 4254 5227
rect 4284 5261 4338 5273
rect 4284 5227 4294 5261
rect 4328 5227 4338 5261
rect 4284 5193 4338 5227
rect 4284 5159 4294 5193
rect 4328 5159 4338 5193
rect 4284 5143 4338 5159
rect 4368 5261 4422 5273
rect 4368 5227 4378 5261
rect 4412 5227 4422 5261
rect 4368 5143 4422 5227
rect 4452 5261 4506 5273
rect 4452 5227 4462 5261
rect 4496 5227 4506 5261
rect 4452 5193 4506 5227
rect 4452 5159 4462 5193
rect 4496 5159 4506 5193
rect 4452 5143 4506 5159
rect 4536 5261 4590 5273
rect 4536 5227 4546 5261
rect 4580 5227 4590 5261
rect 4536 5143 4590 5227
rect 4620 5261 4674 5273
rect 4620 5227 4630 5261
rect 4664 5227 4674 5261
rect 4620 5193 4674 5227
rect 4620 5159 4630 5193
rect 4664 5159 4674 5193
rect 4620 5143 4674 5159
rect 4704 5261 4758 5273
rect 4704 5227 4714 5261
rect 4748 5227 4758 5261
rect 4704 5143 4758 5227
rect 4788 5261 4842 5273
rect 4788 5227 4798 5261
rect 4832 5227 4842 5261
rect 4788 5193 4842 5227
rect 4788 5159 4798 5193
rect 4832 5159 4842 5193
rect 4788 5143 4842 5159
rect 4872 5261 4926 5273
rect 4872 5227 4882 5261
rect 4916 5227 4926 5261
rect 4872 5143 4926 5227
rect 4956 5261 5010 5273
rect 4956 5227 4966 5261
rect 5000 5227 5010 5261
rect 4956 5193 5010 5227
rect 4956 5159 4966 5193
rect 5000 5159 5010 5193
rect 4956 5143 5010 5159
rect 5040 5261 5094 5273
rect 5040 5227 5050 5261
rect 5084 5227 5094 5261
rect 5040 5143 5094 5227
rect 5124 5261 5178 5273
rect 5124 5227 5134 5261
rect 5168 5227 5178 5261
rect 5124 5193 5178 5227
rect 5124 5159 5134 5193
rect 5168 5159 5178 5193
rect 5124 5143 5178 5159
rect 5208 5261 5262 5273
rect 5208 5227 5218 5261
rect 5252 5227 5262 5261
rect 5208 5143 5262 5227
rect 5292 5261 5346 5273
rect 5292 5227 5302 5261
rect 5336 5227 5346 5261
rect 5292 5193 5346 5227
rect 5292 5159 5302 5193
rect 5336 5159 5346 5193
rect 5292 5143 5346 5159
rect 5376 5261 5428 5273
rect 5376 5227 5386 5261
rect 5420 5227 5428 5261
rect 5376 5193 5428 5227
rect 5376 5159 5386 5193
rect 5420 5159 5428 5193
rect 5376 5143 5428 5159
rect 17250 5263 17302 5275
rect 17250 5229 17258 5263
rect 17292 5229 17302 5263
rect 17250 5195 17302 5229
rect 17250 5161 17258 5195
rect 17292 5161 17302 5195
rect 17250 5145 17302 5161
rect 17332 5263 17386 5275
rect 17332 5229 17342 5263
rect 17376 5229 17386 5263
rect 17332 5195 17386 5229
rect 17332 5161 17342 5195
rect 17376 5161 17386 5195
rect 17332 5145 17386 5161
rect 17416 5263 17470 5275
rect 17416 5229 17426 5263
rect 17460 5229 17470 5263
rect 17416 5145 17470 5229
rect 17500 5263 17554 5275
rect 17500 5229 17510 5263
rect 17544 5229 17554 5263
rect 17500 5195 17554 5229
rect 17500 5161 17510 5195
rect 17544 5161 17554 5195
rect 17500 5145 17554 5161
rect 17584 5263 17638 5275
rect 17584 5229 17594 5263
rect 17628 5229 17638 5263
rect 17584 5145 17638 5229
rect 17668 5263 17722 5275
rect 17668 5229 17678 5263
rect 17712 5229 17722 5263
rect 17668 5195 17722 5229
rect 17668 5161 17678 5195
rect 17712 5161 17722 5195
rect 17668 5145 17722 5161
rect 17752 5263 17806 5275
rect 17752 5229 17762 5263
rect 17796 5229 17806 5263
rect 17752 5145 17806 5229
rect 17836 5263 17890 5275
rect 17836 5229 17846 5263
rect 17880 5229 17890 5263
rect 17836 5195 17890 5229
rect 17836 5161 17846 5195
rect 17880 5161 17890 5195
rect 17836 5145 17890 5161
rect 17920 5263 17974 5275
rect 17920 5229 17930 5263
rect 17964 5229 17974 5263
rect 17920 5145 17974 5229
rect 18004 5263 18058 5275
rect 18004 5229 18014 5263
rect 18048 5229 18058 5263
rect 18004 5195 18058 5229
rect 18004 5161 18014 5195
rect 18048 5161 18058 5195
rect 18004 5145 18058 5161
rect 18088 5263 18142 5275
rect 18088 5229 18098 5263
rect 18132 5229 18142 5263
rect 18088 5145 18142 5229
rect 18172 5263 18226 5275
rect 18172 5229 18182 5263
rect 18216 5229 18226 5263
rect 18172 5195 18226 5229
rect 18172 5161 18182 5195
rect 18216 5161 18226 5195
rect 18172 5145 18226 5161
rect 18256 5263 18310 5275
rect 18256 5229 18266 5263
rect 18300 5229 18310 5263
rect 18256 5145 18310 5229
rect 18340 5263 18394 5275
rect 18340 5229 18350 5263
rect 18384 5229 18394 5263
rect 18340 5195 18394 5229
rect 18340 5161 18350 5195
rect 18384 5161 18394 5195
rect 18340 5145 18394 5161
rect 18424 5263 18478 5275
rect 18424 5229 18434 5263
rect 18468 5229 18478 5263
rect 18424 5145 18478 5229
rect 18508 5263 18562 5275
rect 18508 5229 18518 5263
rect 18552 5229 18562 5263
rect 18508 5195 18562 5229
rect 18508 5161 18518 5195
rect 18552 5161 18562 5195
rect 18508 5145 18562 5161
rect 18592 5263 18644 5275
rect 18592 5229 18602 5263
rect 18636 5229 18644 5263
rect 18592 5195 18644 5229
rect 18592 5161 18602 5195
rect 18636 5161 18644 5195
rect 18592 5145 18644 5161
rect 19132 5261 19184 5273
rect 19132 5227 19140 5261
rect 19174 5227 19184 5261
rect 19132 5193 19184 5227
rect 19132 5159 19140 5193
rect 19174 5159 19184 5193
rect 19132 5143 19184 5159
rect 19214 5261 19268 5273
rect 19214 5227 19224 5261
rect 19258 5227 19268 5261
rect 19214 5193 19268 5227
rect 19214 5159 19224 5193
rect 19258 5159 19268 5193
rect 19214 5143 19268 5159
rect 19298 5261 19352 5273
rect 19298 5227 19308 5261
rect 19342 5227 19352 5261
rect 19298 5143 19352 5227
rect 19382 5261 19436 5273
rect 19382 5227 19392 5261
rect 19426 5227 19436 5261
rect 19382 5193 19436 5227
rect 19382 5159 19392 5193
rect 19426 5159 19436 5193
rect 19382 5143 19436 5159
rect 19466 5261 19520 5273
rect 19466 5227 19476 5261
rect 19510 5227 19520 5261
rect 19466 5143 19520 5227
rect 19550 5261 19604 5273
rect 19550 5227 19560 5261
rect 19594 5227 19604 5261
rect 19550 5193 19604 5227
rect 19550 5159 19560 5193
rect 19594 5159 19604 5193
rect 19550 5143 19604 5159
rect 19634 5261 19688 5273
rect 19634 5227 19644 5261
rect 19678 5227 19688 5261
rect 19634 5143 19688 5227
rect 19718 5261 19772 5273
rect 19718 5227 19728 5261
rect 19762 5227 19772 5261
rect 19718 5193 19772 5227
rect 19718 5159 19728 5193
rect 19762 5159 19772 5193
rect 19718 5143 19772 5159
rect 19802 5261 19856 5273
rect 19802 5227 19812 5261
rect 19846 5227 19856 5261
rect 19802 5143 19856 5227
rect 19886 5261 19940 5273
rect 19886 5227 19896 5261
rect 19930 5227 19940 5261
rect 19886 5193 19940 5227
rect 19886 5159 19896 5193
rect 19930 5159 19940 5193
rect 19886 5143 19940 5159
rect 19970 5261 20024 5273
rect 19970 5227 19980 5261
rect 20014 5227 20024 5261
rect 19970 5143 20024 5227
rect 20054 5261 20108 5273
rect 20054 5227 20064 5261
rect 20098 5227 20108 5261
rect 20054 5193 20108 5227
rect 20054 5159 20064 5193
rect 20098 5159 20108 5193
rect 20054 5143 20108 5159
rect 20138 5261 20192 5273
rect 20138 5227 20148 5261
rect 20182 5227 20192 5261
rect 20138 5143 20192 5227
rect 20222 5261 20276 5273
rect 20222 5227 20232 5261
rect 20266 5227 20276 5261
rect 20222 5193 20276 5227
rect 20222 5159 20232 5193
rect 20266 5159 20276 5193
rect 20222 5143 20276 5159
rect 20306 5261 20360 5273
rect 20306 5227 20316 5261
rect 20350 5227 20360 5261
rect 20306 5143 20360 5227
rect 20390 5261 20444 5273
rect 20390 5227 20400 5261
rect 20434 5227 20444 5261
rect 20390 5193 20444 5227
rect 20390 5159 20400 5193
rect 20434 5159 20444 5193
rect 20390 5143 20444 5159
rect 20474 5261 20526 5273
rect 20474 5227 20484 5261
rect 20518 5227 20526 5261
rect 20474 5193 20526 5227
rect 20474 5159 20484 5193
rect 20518 5159 20526 5193
rect 20474 5143 20526 5159
rect -3307 4317 -3255 4331
rect -3307 4283 -3299 4317
rect -3265 4283 -3255 4317
rect -3307 4249 -3255 4283
rect -3307 4215 -3299 4249
rect -3265 4215 -3255 4249
rect -3307 4201 -3255 4215
rect -3225 4317 -3171 4331
rect -3225 4283 -3215 4317
rect -3181 4283 -3171 4317
rect -3225 4249 -3171 4283
rect -3225 4215 -3215 4249
rect -3181 4215 -3171 4249
rect -3225 4201 -3171 4215
rect -3141 4317 -3089 4331
rect -3141 4283 -3131 4317
rect -3097 4283 -3089 4317
rect -2493 4317 -2441 4331
rect -3141 4249 -3089 4283
rect -2493 4283 -2485 4317
rect -2451 4283 -2441 4317
rect -3141 4215 -3131 4249
rect -3097 4215 -3089 4249
rect -3141 4201 -3089 4215
rect -2493 4249 -2441 4283
rect -2493 4215 -2485 4249
rect -2451 4215 -2441 4249
rect -2493 4201 -2441 4215
rect -2411 4317 -2357 4331
rect -2411 4283 -2401 4317
rect -2367 4283 -2357 4317
rect -2411 4249 -2357 4283
rect -2411 4215 -2401 4249
rect -2367 4215 -2357 4249
rect -2411 4201 -2357 4215
rect -2327 4317 -2275 4331
rect -2327 4283 -2317 4317
rect -2283 4283 -2275 4317
rect -2327 4249 -2275 4283
rect -2327 4215 -2317 4249
rect -2283 4215 -2275 4249
rect -2327 4201 -2275 4215
rect -1419 4317 -1367 4331
rect -1419 4283 -1411 4317
rect -1377 4283 -1367 4317
rect -1419 4249 -1367 4283
rect -1419 4215 -1411 4249
rect -1377 4215 -1367 4249
rect -1419 4201 -1367 4215
rect -1337 4317 -1283 4331
rect -1337 4283 -1327 4317
rect -1293 4283 -1283 4317
rect -1337 4249 -1283 4283
rect -1337 4215 -1327 4249
rect -1293 4215 -1283 4249
rect -1337 4201 -1283 4215
rect -1253 4317 -1201 4331
rect -1253 4283 -1243 4317
rect -1209 4283 -1201 4317
rect -605 4317 -553 4331
rect -1253 4249 -1201 4283
rect -605 4283 -597 4317
rect -563 4283 -553 4317
rect -1253 4215 -1243 4249
rect -1209 4215 -1201 4249
rect -1253 4201 -1201 4215
rect -605 4249 -553 4283
rect -605 4215 -597 4249
rect -563 4215 -553 4249
rect -605 4201 -553 4215
rect -523 4317 -469 4331
rect -523 4283 -513 4317
rect -479 4283 -469 4317
rect -523 4249 -469 4283
rect -523 4215 -513 4249
rect -479 4215 -469 4249
rect -523 4201 -469 4215
rect -439 4317 -387 4331
rect -439 4283 -429 4317
rect -395 4283 -387 4317
rect -439 4249 -387 4283
rect -439 4215 -429 4249
rect -395 4215 -387 4249
rect -439 4201 -387 4215
rect 469 4317 521 4331
rect 469 4283 477 4317
rect 511 4283 521 4317
rect 469 4249 521 4283
rect 469 4215 477 4249
rect 511 4215 521 4249
rect 469 4201 521 4215
rect 551 4317 605 4331
rect 551 4283 561 4317
rect 595 4283 605 4317
rect 551 4249 605 4283
rect 551 4215 561 4249
rect 595 4215 605 4249
rect 551 4201 605 4215
rect 635 4317 687 4331
rect 635 4283 645 4317
rect 679 4283 687 4317
rect 1283 4317 1335 4331
rect 635 4249 687 4283
rect 1283 4283 1291 4317
rect 1325 4283 1335 4317
rect 635 4215 645 4249
rect 679 4215 687 4249
rect 635 4201 687 4215
rect 1283 4249 1335 4283
rect 1283 4215 1291 4249
rect 1325 4215 1335 4249
rect 1283 4201 1335 4215
rect 1365 4317 1419 4331
rect 1365 4283 1375 4317
rect 1409 4283 1419 4317
rect 1365 4249 1419 4283
rect 1365 4215 1375 4249
rect 1409 4215 1419 4249
rect 1365 4201 1419 4215
rect 1449 4317 1501 4331
rect 1449 4283 1459 4317
rect 1493 4283 1501 4317
rect 1449 4249 1501 4283
rect 1449 4215 1459 4249
rect 1493 4215 1501 4249
rect 1449 4201 1501 4215
rect 2357 4317 2409 4331
rect 2357 4283 2365 4317
rect 2399 4283 2409 4317
rect 2357 4249 2409 4283
rect 2357 4215 2365 4249
rect 2399 4215 2409 4249
rect 2357 4201 2409 4215
rect 2439 4317 2493 4331
rect 2439 4283 2449 4317
rect 2483 4283 2493 4317
rect 2439 4249 2493 4283
rect 2439 4215 2449 4249
rect 2483 4215 2493 4249
rect 2439 4201 2493 4215
rect 2523 4317 2575 4331
rect 2523 4283 2533 4317
rect 2567 4283 2575 4317
rect 3171 4317 3223 4331
rect 2523 4249 2575 4283
rect 3171 4283 3179 4317
rect 3213 4283 3223 4317
rect 2523 4215 2533 4249
rect 2567 4215 2575 4249
rect 2523 4201 2575 4215
rect 3171 4249 3223 4283
rect 3171 4215 3179 4249
rect 3213 4215 3223 4249
rect 3171 4201 3223 4215
rect 3253 4317 3307 4331
rect 3253 4283 3263 4317
rect 3297 4283 3307 4317
rect 3253 4249 3307 4283
rect 3253 4215 3263 4249
rect 3297 4215 3307 4249
rect 3253 4201 3307 4215
rect 3337 4317 3389 4331
rect 3337 4283 3347 4317
rect 3381 4283 3389 4317
rect 3337 4249 3389 4283
rect 3337 4215 3347 4249
rect 3381 4215 3389 4249
rect 3337 4201 3389 4215
rect 4245 4317 4297 4331
rect 4245 4283 4253 4317
rect 4287 4283 4297 4317
rect 4245 4249 4297 4283
rect 4245 4215 4253 4249
rect 4287 4215 4297 4249
rect 4245 4201 4297 4215
rect 4327 4317 4381 4331
rect 4327 4283 4337 4317
rect 4371 4283 4381 4317
rect 4327 4249 4381 4283
rect 4327 4215 4337 4249
rect 4371 4215 4381 4249
rect 4327 4201 4381 4215
rect 4411 4317 4463 4331
rect 4411 4283 4421 4317
rect 4455 4283 4463 4317
rect 5059 4317 5111 4331
rect 4411 4249 4463 4283
rect 5059 4283 5067 4317
rect 5101 4283 5111 4317
rect 4411 4215 4421 4249
rect 4455 4215 4463 4249
rect 4411 4201 4463 4215
rect 5059 4249 5111 4283
rect 5059 4215 5067 4249
rect 5101 4215 5111 4249
rect 5059 4201 5111 4215
rect 5141 4317 5195 4331
rect 5141 4283 5151 4317
rect 5185 4283 5195 4317
rect 5141 4249 5195 4283
rect 5141 4215 5151 4249
rect 5185 4215 5195 4249
rect 5141 4201 5195 4215
rect 5225 4317 5277 4331
rect 5225 4283 5235 4317
rect 5269 4283 5277 4317
rect 5225 4249 5277 4283
rect 5225 4215 5235 4249
rect 5269 4215 5277 4249
rect 5225 4201 5277 4215
rect 6133 4317 6185 4331
rect 6133 4283 6141 4317
rect 6175 4283 6185 4317
rect 6133 4249 6185 4283
rect 6133 4215 6141 4249
rect 6175 4215 6185 4249
rect 6133 4201 6185 4215
rect 6215 4317 6269 4331
rect 6215 4283 6225 4317
rect 6259 4283 6269 4317
rect 6215 4249 6269 4283
rect 6215 4215 6225 4249
rect 6259 4215 6269 4249
rect 6215 4201 6269 4215
rect 6299 4317 6351 4331
rect 6299 4283 6309 4317
rect 6343 4283 6351 4317
rect 6947 4317 6999 4331
rect 6299 4249 6351 4283
rect 6947 4283 6955 4317
rect 6989 4283 6999 4317
rect 6299 4215 6309 4249
rect 6343 4215 6351 4249
rect 6299 4201 6351 4215
rect 6947 4249 6999 4283
rect 6947 4215 6955 4249
rect 6989 4215 6999 4249
rect 6947 4201 6999 4215
rect 7029 4317 7083 4331
rect 7029 4283 7039 4317
rect 7073 4283 7083 4317
rect 7029 4249 7083 4283
rect 7029 4215 7039 4249
rect 7073 4215 7083 4249
rect 7029 4201 7083 4215
rect 7113 4317 7165 4331
rect 7113 4283 7123 4317
rect 7157 4283 7165 4317
rect 7113 4249 7165 4283
rect 7113 4215 7123 4249
rect 7157 4215 7165 4249
rect 7113 4201 7165 4215
rect 8021 4317 8073 4331
rect 8021 4283 8029 4317
rect 8063 4283 8073 4317
rect 8021 4249 8073 4283
rect 8021 4215 8029 4249
rect 8063 4215 8073 4249
rect 8021 4201 8073 4215
rect 8103 4317 8157 4331
rect 8103 4283 8113 4317
rect 8147 4283 8157 4317
rect 8103 4249 8157 4283
rect 8103 4215 8113 4249
rect 8147 4215 8157 4249
rect 8103 4201 8157 4215
rect 8187 4317 8239 4331
rect 8187 4283 8197 4317
rect 8231 4283 8239 4317
rect 8835 4317 8887 4331
rect 8187 4249 8239 4283
rect 8835 4283 8843 4317
rect 8877 4283 8887 4317
rect 8187 4215 8197 4249
rect 8231 4215 8239 4249
rect 8187 4201 8239 4215
rect 8835 4249 8887 4283
rect 8835 4215 8843 4249
rect 8877 4215 8887 4249
rect 8835 4201 8887 4215
rect 8917 4317 8971 4331
rect 8917 4283 8927 4317
rect 8961 4283 8971 4317
rect 8917 4249 8971 4283
rect 8917 4215 8927 4249
rect 8961 4215 8971 4249
rect 8917 4201 8971 4215
rect 9001 4317 9053 4331
rect 9001 4283 9011 4317
rect 9045 4283 9053 4317
rect 9001 4249 9053 4283
rect 9001 4215 9011 4249
rect 9045 4215 9053 4249
rect 9001 4201 9053 4215
rect 9909 4317 9961 4331
rect 9909 4283 9917 4317
rect 9951 4283 9961 4317
rect 9909 4249 9961 4283
rect 9909 4215 9917 4249
rect 9951 4215 9961 4249
rect 9909 4201 9961 4215
rect 9991 4317 10045 4331
rect 9991 4283 10001 4317
rect 10035 4283 10045 4317
rect 9991 4249 10045 4283
rect 9991 4215 10001 4249
rect 10035 4215 10045 4249
rect 9991 4201 10045 4215
rect 10075 4317 10127 4331
rect 10075 4283 10085 4317
rect 10119 4283 10127 4317
rect 10723 4317 10775 4331
rect 10075 4249 10127 4283
rect 10723 4283 10731 4317
rect 10765 4283 10775 4317
rect 10075 4215 10085 4249
rect 10119 4215 10127 4249
rect 10075 4201 10127 4215
rect 10723 4249 10775 4283
rect 10723 4215 10731 4249
rect 10765 4215 10775 4249
rect 10723 4201 10775 4215
rect 10805 4317 10859 4331
rect 10805 4283 10815 4317
rect 10849 4283 10859 4317
rect 10805 4249 10859 4283
rect 10805 4215 10815 4249
rect 10849 4215 10859 4249
rect 10805 4201 10859 4215
rect 10889 4317 10941 4331
rect 10889 4283 10899 4317
rect 10933 4283 10941 4317
rect 10889 4249 10941 4283
rect 10889 4215 10899 4249
rect 10933 4215 10941 4249
rect 10889 4201 10941 4215
rect 11791 4317 11843 4331
rect 11791 4283 11799 4317
rect 11833 4283 11843 4317
rect 11791 4249 11843 4283
rect 11791 4215 11799 4249
rect 11833 4215 11843 4249
rect 11791 4201 11843 4215
rect 11873 4317 11927 4331
rect 11873 4283 11883 4317
rect 11917 4283 11927 4317
rect 11873 4249 11927 4283
rect 11873 4215 11883 4249
rect 11917 4215 11927 4249
rect 11873 4201 11927 4215
rect 11957 4317 12009 4331
rect 11957 4283 11967 4317
rect 12001 4283 12009 4317
rect 12605 4317 12657 4331
rect 11957 4249 12009 4283
rect 12605 4283 12613 4317
rect 12647 4283 12657 4317
rect 11957 4215 11967 4249
rect 12001 4215 12009 4249
rect 11957 4201 12009 4215
rect 12605 4249 12657 4283
rect 12605 4215 12613 4249
rect 12647 4215 12657 4249
rect 12605 4201 12657 4215
rect 12687 4317 12741 4331
rect 12687 4283 12697 4317
rect 12731 4283 12741 4317
rect 12687 4249 12741 4283
rect 12687 4215 12697 4249
rect 12731 4215 12741 4249
rect 12687 4201 12741 4215
rect 12771 4317 12823 4331
rect 12771 4283 12781 4317
rect 12815 4283 12823 4317
rect 12771 4249 12823 4283
rect 12771 4215 12781 4249
rect 12815 4215 12823 4249
rect 12771 4201 12823 4215
rect 13679 4317 13731 4331
rect 13679 4283 13687 4317
rect 13721 4283 13731 4317
rect 13679 4249 13731 4283
rect 13679 4215 13687 4249
rect 13721 4215 13731 4249
rect 13679 4201 13731 4215
rect 13761 4317 13815 4331
rect 13761 4283 13771 4317
rect 13805 4283 13815 4317
rect 13761 4249 13815 4283
rect 13761 4215 13771 4249
rect 13805 4215 13815 4249
rect 13761 4201 13815 4215
rect 13845 4317 13897 4331
rect 13845 4283 13855 4317
rect 13889 4283 13897 4317
rect 14493 4317 14545 4331
rect 13845 4249 13897 4283
rect 14493 4283 14501 4317
rect 14535 4283 14545 4317
rect 13845 4215 13855 4249
rect 13889 4215 13897 4249
rect 13845 4201 13897 4215
rect 14493 4249 14545 4283
rect 14493 4215 14501 4249
rect 14535 4215 14545 4249
rect 14493 4201 14545 4215
rect 14575 4317 14629 4331
rect 14575 4283 14585 4317
rect 14619 4283 14629 4317
rect 14575 4249 14629 4283
rect 14575 4215 14585 4249
rect 14619 4215 14629 4249
rect 14575 4201 14629 4215
rect 14659 4317 14711 4331
rect 14659 4283 14669 4317
rect 14703 4283 14711 4317
rect 14659 4249 14711 4283
rect 14659 4215 14669 4249
rect 14703 4215 14711 4249
rect 14659 4201 14711 4215
rect 15567 4317 15619 4331
rect 15567 4283 15575 4317
rect 15609 4283 15619 4317
rect 15567 4249 15619 4283
rect 15567 4215 15575 4249
rect 15609 4215 15619 4249
rect 15567 4201 15619 4215
rect 15649 4317 15703 4331
rect 15649 4283 15659 4317
rect 15693 4283 15703 4317
rect 15649 4249 15703 4283
rect 15649 4215 15659 4249
rect 15693 4215 15703 4249
rect 15649 4201 15703 4215
rect 15733 4317 15785 4331
rect 15733 4283 15743 4317
rect 15777 4283 15785 4317
rect 16381 4317 16433 4331
rect 15733 4249 15785 4283
rect 16381 4283 16389 4317
rect 16423 4283 16433 4317
rect 15733 4215 15743 4249
rect 15777 4215 15785 4249
rect 15733 4201 15785 4215
rect 16381 4249 16433 4283
rect 16381 4215 16389 4249
rect 16423 4215 16433 4249
rect 16381 4201 16433 4215
rect 16463 4317 16517 4331
rect 16463 4283 16473 4317
rect 16507 4283 16517 4317
rect 16463 4249 16517 4283
rect 16463 4215 16473 4249
rect 16507 4215 16517 4249
rect 16463 4201 16517 4215
rect 16547 4317 16599 4331
rect 16547 4283 16557 4317
rect 16591 4283 16599 4317
rect 16547 4249 16599 4283
rect 16547 4215 16557 4249
rect 16591 4215 16599 4249
rect 16547 4201 16599 4215
rect 17455 4317 17507 4331
rect 17455 4283 17463 4317
rect 17497 4283 17507 4317
rect 17455 4249 17507 4283
rect 17455 4215 17463 4249
rect 17497 4215 17507 4249
rect 17455 4201 17507 4215
rect 17537 4317 17591 4331
rect 17537 4283 17547 4317
rect 17581 4283 17591 4317
rect 17537 4249 17591 4283
rect 17537 4215 17547 4249
rect 17581 4215 17591 4249
rect 17537 4201 17591 4215
rect 17621 4317 17673 4331
rect 17621 4283 17631 4317
rect 17665 4283 17673 4317
rect 18269 4317 18321 4331
rect 17621 4249 17673 4283
rect 18269 4283 18277 4317
rect 18311 4283 18321 4317
rect 17621 4215 17631 4249
rect 17665 4215 17673 4249
rect 17621 4201 17673 4215
rect 18269 4249 18321 4283
rect 18269 4215 18277 4249
rect 18311 4215 18321 4249
rect 18269 4201 18321 4215
rect 18351 4317 18405 4331
rect 18351 4283 18361 4317
rect 18395 4283 18405 4317
rect 18351 4249 18405 4283
rect 18351 4215 18361 4249
rect 18395 4215 18405 4249
rect 18351 4201 18405 4215
rect 18435 4317 18487 4331
rect 18435 4283 18445 4317
rect 18479 4283 18487 4317
rect 18435 4249 18487 4283
rect 18435 4215 18445 4249
rect 18479 4215 18487 4249
rect 18435 4201 18487 4215
rect 19343 4317 19395 4331
rect 19343 4283 19351 4317
rect 19385 4283 19395 4317
rect 19343 4249 19395 4283
rect 19343 4215 19351 4249
rect 19385 4215 19395 4249
rect 19343 4201 19395 4215
rect 19425 4317 19479 4331
rect 19425 4283 19435 4317
rect 19469 4283 19479 4317
rect 19425 4249 19479 4283
rect 19425 4215 19435 4249
rect 19469 4215 19479 4249
rect 19425 4201 19479 4215
rect 19509 4317 19561 4331
rect 19509 4283 19519 4317
rect 19553 4283 19561 4317
rect 20157 4317 20209 4331
rect 19509 4249 19561 4283
rect 20157 4283 20165 4317
rect 20199 4283 20209 4317
rect 19509 4215 19519 4249
rect 19553 4215 19561 4249
rect 19509 4201 19561 4215
rect 20157 4249 20209 4283
rect 20157 4215 20165 4249
rect 20199 4215 20209 4249
rect 20157 4201 20209 4215
rect 20239 4317 20293 4331
rect 20239 4283 20249 4317
rect 20283 4283 20293 4317
rect 20239 4249 20293 4283
rect 20239 4215 20249 4249
rect 20283 4215 20293 4249
rect 20239 4201 20293 4215
rect 20323 4317 20375 4331
rect 20323 4283 20333 4317
rect 20367 4283 20375 4317
rect 20323 4249 20375 4283
rect 20323 4215 20333 4249
rect 20367 4215 20375 4249
rect 20323 4201 20375 4215
rect 21231 4317 21283 4331
rect 21231 4283 21239 4317
rect 21273 4283 21283 4317
rect 21231 4249 21283 4283
rect 21231 4215 21239 4249
rect 21273 4215 21283 4249
rect 21231 4201 21283 4215
rect 21313 4317 21367 4331
rect 21313 4283 21323 4317
rect 21357 4283 21367 4317
rect 21313 4249 21367 4283
rect 21313 4215 21323 4249
rect 21357 4215 21367 4249
rect 21313 4201 21367 4215
rect 21397 4317 21449 4331
rect 21397 4283 21407 4317
rect 21441 4283 21449 4317
rect 22045 4317 22097 4331
rect 21397 4249 21449 4283
rect 22045 4283 22053 4317
rect 22087 4283 22097 4317
rect 21397 4215 21407 4249
rect 21441 4215 21449 4249
rect 21397 4201 21449 4215
rect 22045 4249 22097 4283
rect 22045 4215 22053 4249
rect 22087 4215 22097 4249
rect 22045 4201 22097 4215
rect 22127 4317 22181 4331
rect 22127 4283 22137 4317
rect 22171 4283 22181 4317
rect 22127 4249 22181 4283
rect 22127 4215 22137 4249
rect 22171 4215 22181 4249
rect 22127 4201 22181 4215
rect 22211 4317 22263 4331
rect 22211 4283 22221 4317
rect 22255 4283 22263 4317
rect 22211 4249 22263 4283
rect 22211 4215 22221 4249
rect 22255 4215 22263 4249
rect 22211 4201 22263 4215
rect 23119 4317 23171 4331
rect 23119 4283 23127 4317
rect 23161 4283 23171 4317
rect 23119 4249 23171 4283
rect 23119 4215 23127 4249
rect 23161 4215 23171 4249
rect 23119 4201 23171 4215
rect 23201 4317 23255 4331
rect 23201 4283 23211 4317
rect 23245 4283 23255 4317
rect 23201 4249 23255 4283
rect 23201 4215 23211 4249
rect 23245 4215 23255 4249
rect 23201 4201 23255 4215
rect 23285 4317 23337 4331
rect 23285 4283 23295 4317
rect 23329 4283 23337 4317
rect 23933 4317 23985 4331
rect 23285 4249 23337 4283
rect 23933 4283 23941 4317
rect 23975 4283 23985 4317
rect 23285 4215 23295 4249
rect 23329 4215 23337 4249
rect 23285 4201 23337 4215
rect 23933 4249 23985 4283
rect 23933 4215 23941 4249
rect 23975 4215 23985 4249
rect 23933 4201 23985 4215
rect 24015 4317 24069 4331
rect 24015 4283 24025 4317
rect 24059 4283 24069 4317
rect 24015 4249 24069 4283
rect 24015 4215 24025 4249
rect 24059 4215 24069 4249
rect 24015 4201 24069 4215
rect 24099 4317 24151 4331
rect 24099 4283 24109 4317
rect 24143 4283 24151 4317
rect 24099 4249 24151 4283
rect 24099 4215 24109 4249
rect 24143 4215 24151 4249
rect 24099 4201 24151 4215
rect 25007 4317 25059 4331
rect 25007 4283 25015 4317
rect 25049 4283 25059 4317
rect 25007 4249 25059 4283
rect 25007 4215 25015 4249
rect 25049 4215 25059 4249
rect 25007 4201 25059 4215
rect 25089 4317 25143 4331
rect 25089 4283 25099 4317
rect 25133 4283 25143 4317
rect 25089 4249 25143 4283
rect 25089 4215 25099 4249
rect 25133 4215 25143 4249
rect 25089 4201 25143 4215
rect 25173 4317 25225 4331
rect 25173 4283 25183 4317
rect 25217 4283 25225 4317
rect 25821 4317 25873 4331
rect 25173 4249 25225 4283
rect 25821 4283 25829 4317
rect 25863 4283 25873 4317
rect 25173 4215 25183 4249
rect 25217 4215 25225 4249
rect 25173 4201 25225 4215
rect 25821 4249 25873 4283
rect 25821 4215 25829 4249
rect 25863 4215 25873 4249
rect 25821 4201 25873 4215
rect 25903 4317 25957 4331
rect 25903 4283 25913 4317
rect 25947 4283 25957 4317
rect 25903 4249 25957 4283
rect 25903 4215 25913 4249
rect 25947 4215 25957 4249
rect 25903 4201 25957 4215
rect 25987 4317 26039 4331
rect 25987 4283 25997 4317
rect 26031 4283 26039 4317
rect 25987 4249 26039 4283
rect 25987 4215 25997 4249
rect 26031 4215 26039 4249
rect 25987 4201 26039 4215
rect -2942 4072 -2880 4086
rect -2942 4038 -2930 4072
rect -2896 4038 -2880 4072
rect -2942 4004 -2880 4038
rect -2942 3970 -2930 4004
rect -2896 3970 -2880 4004
rect -2942 3956 -2880 3970
rect -2850 4072 -2784 4086
rect -2850 4038 -2834 4072
rect -2800 4038 -2784 4072
rect -2850 4004 -2784 4038
rect -2850 3970 -2834 4004
rect -2800 3970 -2784 4004
rect -2850 3956 -2784 3970
rect -2754 4072 -2692 4086
rect -2754 4038 -2738 4072
rect -2704 4038 -2692 4072
rect -2754 4004 -2692 4038
rect -2754 3970 -2738 4004
rect -2704 3970 -2692 4004
rect -2754 3956 -2692 3970
rect -1054 4072 -992 4086
rect -1054 4038 -1042 4072
rect -1008 4038 -992 4072
rect -1054 4004 -992 4038
rect -1054 3970 -1042 4004
rect -1008 3970 -992 4004
rect -1054 3956 -992 3970
rect -962 4072 -896 4086
rect -962 4038 -946 4072
rect -912 4038 -896 4072
rect -962 4004 -896 4038
rect -962 3970 -946 4004
rect -912 3970 -896 4004
rect -962 3956 -896 3970
rect -866 4072 -804 4086
rect -866 4038 -850 4072
rect -816 4038 -804 4072
rect -866 4004 -804 4038
rect -866 3970 -850 4004
rect -816 3970 -804 4004
rect -866 3956 -804 3970
rect 834 4072 896 4086
rect 834 4038 846 4072
rect 880 4038 896 4072
rect 834 4004 896 4038
rect 834 3970 846 4004
rect 880 3970 896 4004
rect 834 3956 896 3970
rect 926 4072 992 4086
rect 926 4038 942 4072
rect 976 4038 992 4072
rect 926 4004 992 4038
rect 926 3970 942 4004
rect 976 3970 992 4004
rect 926 3956 992 3970
rect 1022 4072 1084 4086
rect 1022 4038 1038 4072
rect 1072 4038 1084 4072
rect 1022 4004 1084 4038
rect 1022 3970 1038 4004
rect 1072 3970 1084 4004
rect 1022 3956 1084 3970
rect 2722 4072 2784 4086
rect 2722 4038 2734 4072
rect 2768 4038 2784 4072
rect 2722 4004 2784 4038
rect 2722 3970 2734 4004
rect 2768 3970 2784 4004
rect 2722 3956 2784 3970
rect 2814 4072 2880 4086
rect 2814 4038 2830 4072
rect 2864 4038 2880 4072
rect 2814 4004 2880 4038
rect 2814 3970 2830 4004
rect 2864 3970 2880 4004
rect 2814 3956 2880 3970
rect 2910 4072 2972 4086
rect 2910 4038 2926 4072
rect 2960 4038 2972 4072
rect 2910 4004 2972 4038
rect 2910 3970 2926 4004
rect 2960 3970 2972 4004
rect 2910 3956 2972 3970
rect 4610 4072 4672 4086
rect 4610 4038 4622 4072
rect 4656 4038 4672 4072
rect 4610 4004 4672 4038
rect 4610 3970 4622 4004
rect 4656 3970 4672 4004
rect 4610 3956 4672 3970
rect 4702 4072 4768 4086
rect 4702 4038 4718 4072
rect 4752 4038 4768 4072
rect 4702 4004 4768 4038
rect 4702 3970 4718 4004
rect 4752 3970 4768 4004
rect 4702 3956 4768 3970
rect 4798 4072 4860 4086
rect 4798 4038 4814 4072
rect 4848 4038 4860 4072
rect 4798 4004 4860 4038
rect 4798 3970 4814 4004
rect 4848 3970 4860 4004
rect 4798 3956 4860 3970
rect 6498 4072 6560 4086
rect 6498 4038 6510 4072
rect 6544 4038 6560 4072
rect 6498 4004 6560 4038
rect 6498 3970 6510 4004
rect 6544 3970 6560 4004
rect 6498 3956 6560 3970
rect 6590 4072 6656 4086
rect 6590 4038 6606 4072
rect 6640 4038 6656 4072
rect 6590 4004 6656 4038
rect 6590 3970 6606 4004
rect 6640 3970 6656 4004
rect 6590 3956 6656 3970
rect 6686 4072 6748 4086
rect 6686 4038 6702 4072
rect 6736 4038 6748 4072
rect 6686 4004 6748 4038
rect 6686 3970 6702 4004
rect 6736 3970 6748 4004
rect 6686 3956 6748 3970
rect 8386 4072 8448 4086
rect 8386 4038 8398 4072
rect 8432 4038 8448 4072
rect 8386 4004 8448 4038
rect 8386 3970 8398 4004
rect 8432 3970 8448 4004
rect 8386 3956 8448 3970
rect 8478 4072 8544 4086
rect 8478 4038 8494 4072
rect 8528 4038 8544 4072
rect 8478 4004 8544 4038
rect 8478 3970 8494 4004
rect 8528 3970 8544 4004
rect 8478 3956 8544 3970
rect 8574 4072 8636 4086
rect 8574 4038 8590 4072
rect 8624 4038 8636 4072
rect 8574 4004 8636 4038
rect 8574 3970 8590 4004
rect 8624 3970 8636 4004
rect 8574 3956 8636 3970
rect 10274 4072 10336 4086
rect 10274 4038 10286 4072
rect 10320 4038 10336 4072
rect 10274 4004 10336 4038
rect 10274 3970 10286 4004
rect 10320 3970 10336 4004
rect 10274 3956 10336 3970
rect 10366 4072 10432 4086
rect 10366 4038 10382 4072
rect 10416 4038 10432 4072
rect 10366 4004 10432 4038
rect 10366 3970 10382 4004
rect 10416 3970 10432 4004
rect 10366 3956 10432 3970
rect 10462 4072 10524 4086
rect 10462 4038 10478 4072
rect 10512 4038 10524 4072
rect 10462 4004 10524 4038
rect 10462 3970 10478 4004
rect 10512 3970 10524 4004
rect 10462 3956 10524 3970
rect 12156 4072 12218 4086
rect 12156 4038 12168 4072
rect 12202 4038 12218 4072
rect 12156 4004 12218 4038
rect 12156 3970 12168 4004
rect 12202 3970 12218 4004
rect 12156 3956 12218 3970
rect 12248 4072 12314 4086
rect 12248 4038 12264 4072
rect 12298 4038 12314 4072
rect 12248 4004 12314 4038
rect 12248 3970 12264 4004
rect 12298 3970 12314 4004
rect 12248 3956 12314 3970
rect 12344 4072 12406 4086
rect 12344 4038 12360 4072
rect 12394 4038 12406 4072
rect 12344 4004 12406 4038
rect 12344 3970 12360 4004
rect 12394 3970 12406 4004
rect 12344 3956 12406 3970
rect 14044 4072 14106 4086
rect 14044 4038 14056 4072
rect 14090 4038 14106 4072
rect 14044 4004 14106 4038
rect 14044 3970 14056 4004
rect 14090 3970 14106 4004
rect 14044 3956 14106 3970
rect 14136 4072 14202 4086
rect 14136 4038 14152 4072
rect 14186 4038 14202 4072
rect 14136 4004 14202 4038
rect 14136 3970 14152 4004
rect 14186 3970 14202 4004
rect 14136 3956 14202 3970
rect 14232 4072 14294 4086
rect 14232 4038 14248 4072
rect 14282 4038 14294 4072
rect 14232 4004 14294 4038
rect 14232 3970 14248 4004
rect 14282 3970 14294 4004
rect 14232 3956 14294 3970
rect 15932 4072 15994 4086
rect 15932 4038 15944 4072
rect 15978 4038 15994 4072
rect 15932 4004 15994 4038
rect 15932 3970 15944 4004
rect 15978 3970 15994 4004
rect 15932 3956 15994 3970
rect 16024 4072 16090 4086
rect 16024 4038 16040 4072
rect 16074 4038 16090 4072
rect 16024 4004 16090 4038
rect 16024 3970 16040 4004
rect 16074 3970 16090 4004
rect 16024 3956 16090 3970
rect 16120 4072 16182 4086
rect 16120 4038 16136 4072
rect 16170 4038 16182 4072
rect 16120 4004 16182 4038
rect 16120 3970 16136 4004
rect 16170 3970 16182 4004
rect 16120 3956 16182 3970
rect 17820 4072 17882 4086
rect 17820 4038 17832 4072
rect 17866 4038 17882 4072
rect 17820 4004 17882 4038
rect 17820 3970 17832 4004
rect 17866 3970 17882 4004
rect 17820 3956 17882 3970
rect 17912 4072 17978 4086
rect 17912 4038 17928 4072
rect 17962 4038 17978 4072
rect 17912 4004 17978 4038
rect 17912 3970 17928 4004
rect 17962 3970 17978 4004
rect 17912 3956 17978 3970
rect 18008 4072 18070 4086
rect 18008 4038 18024 4072
rect 18058 4038 18070 4072
rect 18008 4004 18070 4038
rect 18008 3970 18024 4004
rect 18058 3970 18070 4004
rect 18008 3956 18070 3970
rect 19708 4072 19770 4086
rect 19708 4038 19720 4072
rect 19754 4038 19770 4072
rect 19708 4004 19770 4038
rect 19708 3970 19720 4004
rect 19754 3970 19770 4004
rect 19708 3956 19770 3970
rect 19800 4072 19866 4086
rect 19800 4038 19816 4072
rect 19850 4038 19866 4072
rect 19800 4004 19866 4038
rect 19800 3970 19816 4004
rect 19850 3970 19866 4004
rect 19800 3956 19866 3970
rect 19896 4072 19958 4086
rect 19896 4038 19912 4072
rect 19946 4038 19958 4072
rect 19896 4004 19958 4038
rect 19896 3970 19912 4004
rect 19946 3970 19958 4004
rect 19896 3956 19958 3970
rect 21596 4072 21658 4086
rect 21596 4038 21608 4072
rect 21642 4038 21658 4072
rect 21596 4004 21658 4038
rect 21596 3970 21608 4004
rect 21642 3970 21658 4004
rect 21596 3956 21658 3970
rect 21688 4072 21754 4086
rect 21688 4038 21704 4072
rect 21738 4038 21754 4072
rect 21688 4004 21754 4038
rect 21688 3970 21704 4004
rect 21738 3970 21754 4004
rect 21688 3956 21754 3970
rect 21784 4072 21846 4086
rect 21784 4038 21800 4072
rect 21834 4038 21846 4072
rect 21784 4004 21846 4038
rect 21784 3970 21800 4004
rect 21834 3970 21846 4004
rect 21784 3956 21846 3970
rect 23484 4072 23546 4086
rect 23484 4038 23496 4072
rect 23530 4038 23546 4072
rect 23484 4004 23546 4038
rect 23484 3970 23496 4004
rect 23530 3970 23546 4004
rect 23484 3956 23546 3970
rect 23576 4072 23642 4086
rect 23576 4038 23592 4072
rect 23626 4038 23642 4072
rect 23576 4004 23642 4038
rect 23576 3970 23592 4004
rect 23626 3970 23642 4004
rect 23576 3956 23642 3970
rect 23672 4072 23734 4086
rect 23672 4038 23688 4072
rect 23722 4038 23734 4072
rect 23672 4004 23734 4038
rect 23672 3970 23688 4004
rect 23722 3970 23734 4004
rect 23672 3956 23734 3970
rect 25372 4072 25434 4086
rect 25372 4038 25384 4072
rect 25418 4038 25434 4072
rect 25372 4004 25434 4038
rect 25372 3970 25384 4004
rect 25418 3970 25434 4004
rect 25372 3956 25434 3970
rect 25464 4072 25530 4086
rect 25464 4038 25480 4072
rect 25514 4038 25530 4072
rect 25464 4004 25530 4038
rect 25464 3970 25480 4004
rect 25514 3970 25530 4004
rect 25464 3956 25530 3970
rect 25560 4072 25622 4086
rect 25560 4038 25576 4072
rect 25610 4038 25622 4072
rect 25560 4004 25622 4038
rect 25560 3970 25576 4004
rect 25610 3970 25622 4004
rect 25560 3956 25622 3970
rect -3444 3265 -3392 3277
rect -3444 3231 -3436 3265
rect -3402 3231 -3392 3265
rect -3444 3197 -3392 3231
rect -3444 3163 -3436 3197
rect -3402 3163 -3392 3197
rect -3444 3147 -3392 3163
rect -3362 3265 -3310 3277
rect -3362 3231 -3352 3265
rect -3318 3231 -3310 3265
rect -3362 3197 -3310 3231
rect -2248 3273 -2196 3285
rect -2248 3239 -2240 3273
rect -2206 3239 -2196 3273
rect -2248 3205 -2196 3239
rect -3362 3163 -3352 3197
rect -3318 3163 -3310 3197
rect -3362 3147 -3310 3163
rect -2248 3171 -2240 3205
rect -2206 3171 -2196 3205
rect -2248 3155 -2196 3171
rect -2166 3273 -2114 3285
rect -2166 3239 -2156 3273
rect -2122 3239 -2114 3273
rect -1556 3265 -1504 3277
rect -2166 3205 -2114 3239
rect -2166 3171 -2156 3205
rect -2122 3171 -2114 3205
rect -2166 3155 -2114 3171
rect -1943 3212 -1891 3257
rect -1943 3178 -1935 3212
rect -1901 3178 -1891 3212
rect -1943 3153 -1891 3178
rect -1861 3199 -1803 3257
rect -1861 3165 -1849 3199
rect -1815 3165 -1803 3199
rect -1861 3153 -1803 3165
rect -1773 3229 -1721 3257
rect -1773 3195 -1763 3229
rect -1729 3195 -1721 3229
rect -1773 3153 -1721 3195
rect -1556 3231 -1548 3265
rect -1514 3231 -1504 3265
rect -1556 3197 -1504 3231
rect -1556 3163 -1548 3197
rect -1514 3163 -1504 3197
rect -1556 3147 -1504 3163
rect -1474 3265 -1422 3277
rect -1474 3231 -1464 3265
rect -1430 3231 -1422 3265
rect -1474 3197 -1422 3231
rect -360 3273 -308 3285
rect -360 3239 -352 3273
rect -318 3239 -308 3273
rect -360 3205 -308 3239
rect -1474 3163 -1464 3197
rect -1430 3163 -1422 3197
rect -1474 3147 -1422 3163
rect -360 3171 -352 3205
rect -318 3171 -308 3205
rect -360 3155 -308 3171
rect -278 3273 -226 3285
rect -278 3239 -268 3273
rect -234 3239 -226 3273
rect 332 3265 384 3277
rect -278 3205 -226 3239
rect -278 3171 -268 3205
rect -234 3171 -226 3205
rect -278 3155 -226 3171
rect -55 3212 -3 3257
rect -55 3178 -47 3212
rect -13 3178 -3 3212
rect -55 3153 -3 3178
rect 27 3199 85 3257
rect 27 3165 39 3199
rect 73 3165 85 3199
rect 27 3153 85 3165
rect 115 3229 167 3257
rect 115 3195 125 3229
rect 159 3195 167 3229
rect 115 3153 167 3195
rect 332 3231 340 3265
rect 374 3231 384 3265
rect 332 3197 384 3231
rect 332 3163 340 3197
rect 374 3163 384 3197
rect 332 3147 384 3163
rect 414 3265 466 3277
rect 414 3231 424 3265
rect 458 3231 466 3265
rect 414 3197 466 3231
rect 1528 3273 1580 3285
rect 1528 3239 1536 3273
rect 1570 3239 1580 3273
rect 1528 3205 1580 3239
rect 414 3163 424 3197
rect 458 3163 466 3197
rect 414 3147 466 3163
rect 1528 3171 1536 3205
rect 1570 3171 1580 3205
rect 1528 3155 1580 3171
rect 1610 3273 1662 3285
rect 1610 3239 1620 3273
rect 1654 3239 1662 3273
rect 2220 3265 2272 3277
rect 1610 3205 1662 3239
rect 1610 3171 1620 3205
rect 1654 3171 1662 3205
rect 1610 3155 1662 3171
rect 1833 3212 1885 3257
rect 1833 3178 1841 3212
rect 1875 3178 1885 3212
rect 1833 3153 1885 3178
rect 1915 3199 1973 3257
rect 1915 3165 1927 3199
rect 1961 3165 1973 3199
rect 1915 3153 1973 3165
rect 2003 3229 2055 3257
rect 2003 3195 2013 3229
rect 2047 3195 2055 3229
rect 2003 3153 2055 3195
rect 2220 3231 2228 3265
rect 2262 3231 2272 3265
rect 2220 3197 2272 3231
rect 2220 3163 2228 3197
rect 2262 3163 2272 3197
rect 2220 3147 2272 3163
rect 2302 3265 2354 3277
rect 2302 3231 2312 3265
rect 2346 3231 2354 3265
rect 2302 3197 2354 3231
rect 3416 3273 3468 3285
rect 3416 3239 3424 3273
rect 3458 3239 3468 3273
rect 3416 3205 3468 3239
rect 2302 3163 2312 3197
rect 2346 3163 2354 3197
rect 2302 3147 2354 3163
rect 3416 3171 3424 3205
rect 3458 3171 3468 3205
rect 3416 3155 3468 3171
rect 3498 3273 3550 3285
rect 3498 3239 3508 3273
rect 3542 3239 3550 3273
rect 4108 3265 4160 3277
rect 3498 3205 3550 3239
rect 3498 3171 3508 3205
rect 3542 3171 3550 3205
rect 3498 3155 3550 3171
rect 3721 3212 3773 3257
rect 3721 3178 3729 3212
rect 3763 3178 3773 3212
rect 3721 3153 3773 3178
rect 3803 3199 3861 3257
rect 3803 3165 3815 3199
rect 3849 3165 3861 3199
rect 3803 3153 3861 3165
rect 3891 3229 3943 3257
rect 3891 3195 3901 3229
rect 3935 3195 3943 3229
rect 3891 3153 3943 3195
rect 4108 3231 4116 3265
rect 4150 3231 4160 3265
rect 4108 3197 4160 3231
rect 4108 3163 4116 3197
rect 4150 3163 4160 3197
rect 4108 3147 4160 3163
rect 4190 3265 4242 3277
rect 4190 3231 4200 3265
rect 4234 3231 4242 3265
rect 4190 3197 4242 3231
rect 5304 3273 5356 3285
rect 5304 3239 5312 3273
rect 5346 3239 5356 3273
rect 5304 3205 5356 3239
rect 4190 3163 4200 3197
rect 4234 3163 4242 3197
rect 4190 3147 4242 3163
rect 5304 3171 5312 3205
rect 5346 3171 5356 3205
rect 5304 3155 5356 3171
rect 5386 3273 5438 3285
rect 5386 3239 5396 3273
rect 5430 3239 5438 3273
rect 5996 3265 6048 3277
rect 5386 3205 5438 3239
rect 5386 3171 5396 3205
rect 5430 3171 5438 3205
rect 5386 3155 5438 3171
rect 5609 3212 5661 3257
rect 5609 3178 5617 3212
rect 5651 3178 5661 3212
rect 5609 3153 5661 3178
rect 5691 3199 5749 3257
rect 5691 3165 5703 3199
rect 5737 3165 5749 3199
rect 5691 3153 5749 3165
rect 5779 3229 5831 3257
rect 5779 3195 5789 3229
rect 5823 3195 5831 3229
rect 5779 3153 5831 3195
rect 5996 3231 6004 3265
rect 6038 3231 6048 3265
rect 5996 3197 6048 3231
rect 5996 3163 6004 3197
rect 6038 3163 6048 3197
rect 5996 3147 6048 3163
rect 6078 3265 6130 3277
rect 6078 3231 6088 3265
rect 6122 3231 6130 3265
rect 6078 3197 6130 3231
rect 7192 3273 7244 3285
rect 7192 3239 7200 3273
rect 7234 3239 7244 3273
rect 7192 3205 7244 3239
rect 6078 3163 6088 3197
rect 6122 3163 6130 3197
rect 6078 3147 6130 3163
rect 7192 3171 7200 3205
rect 7234 3171 7244 3205
rect 7192 3155 7244 3171
rect 7274 3273 7326 3285
rect 7274 3239 7284 3273
rect 7318 3239 7326 3273
rect 7884 3265 7936 3277
rect 7274 3205 7326 3239
rect 7274 3171 7284 3205
rect 7318 3171 7326 3205
rect 7274 3155 7326 3171
rect 7497 3212 7549 3257
rect 7497 3178 7505 3212
rect 7539 3178 7549 3212
rect 7497 3153 7549 3178
rect 7579 3199 7637 3257
rect 7579 3165 7591 3199
rect 7625 3165 7637 3199
rect 7579 3153 7637 3165
rect 7667 3229 7719 3257
rect 7667 3195 7677 3229
rect 7711 3195 7719 3229
rect 7667 3153 7719 3195
rect 7884 3231 7892 3265
rect 7926 3231 7936 3265
rect 7884 3197 7936 3231
rect 7884 3163 7892 3197
rect 7926 3163 7936 3197
rect 7884 3147 7936 3163
rect 7966 3265 8018 3277
rect 7966 3231 7976 3265
rect 8010 3231 8018 3265
rect 7966 3197 8018 3231
rect 9080 3273 9132 3285
rect 9080 3239 9088 3273
rect 9122 3239 9132 3273
rect 9080 3205 9132 3239
rect 7966 3163 7976 3197
rect 8010 3163 8018 3197
rect 7966 3147 8018 3163
rect 9080 3171 9088 3205
rect 9122 3171 9132 3205
rect 9080 3155 9132 3171
rect 9162 3273 9214 3285
rect 9162 3239 9172 3273
rect 9206 3239 9214 3273
rect 9772 3265 9824 3277
rect 9162 3205 9214 3239
rect 9162 3171 9172 3205
rect 9206 3171 9214 3205
rect 9162 3155 9214 3171
rect 9385 3212 9437 3257
rect 9385 3178 9393 3212
rect 9427 3178 9437 3212
rect 9385 3153 9437 3178
rect 9467 3199 9525 3257
rect 9467 3165 9479 3199
rect 9513 3165 9525 3199
rect 9467 3153 9525 3165
rect 9555 3229 9607 3257
rect 9555 3195 9565 3229
rect 9599 3195 9607 3229
rect 9555 3153 9607 3195
rect 9772 3231 9780 3265
rect 9814 3231 9824 3265
rect 9772 3197 9824 3231
rect 9772 3163 9780 3197
rect 9814 3163 9824 3197
rect 9772 3147 9824 3163
rect 9854 3265 9906 3277
rect 9854 3231 9864 3265
rect 9898 3231 9906 3265
rect 9854 3197 9906 3231
rect 10968 3273 11020 3285
rect 10968 3239 10976 3273
rect 11010 3239 11020 3273
rect 10968 3205 11020 3239
rect 9854 3163 9864 3197
rect 9898 3163 9906 3197
rect 9854 3147 9906 3163
rect 10968 3171 10976 3205
rect 11010 3171 11020 3205
rect 10968 3155 11020 3171
rect 11050 3273 11102 3285
rect 11050 3239 11060 3273
rect 11094 3239 11102 3273
rect 11654 3265 11706 3277
rect 11050 3205 11102 3239
rect 11050 3171 11060 3205
rect 11094 3171 11102 3205
rect 11050 3155 11102 3171
rect 11273 3212 11325 3257
rect 11273 3178 11281 3212
rect 11315 3178 11325 3212
rect 11273 3153 11325 3178
rect 11355 3199 11413 3257
rect 11355 3165 11367 3199
rect 11401 3165 11413 3199
rect 11355 3153 11413 3165
rect 11443 3229 11495 3257
rect 11443 3195 11453 3229
rect 11487 3195 11495 3229
rect 11443 3153 11495 3195
rect 11654 3231 11662 3265
rect 11696 3231 11706 3265
rect 11654 3197 11706 3231
rect 11654 3163 11662 3197
rect 11696 3163 11706 3197
rect 11654 3147 11706 3163
rect 11736 3265 11788 3277
rect 11736 3231 11746 3265
rect 11780 3231 11788 3265
rect 11736 3197 11788 3231
rect 12850 3273 12902 3285
rect 12850 3239 12858 3273
rect 12892 3239 12902 3273
rect 12850 3205 12902 3239
rect 11736 3163 11746 3197
rect 11780 3163 11788 3197
rect 11736 3147 11788 3163
rect 12850 3171 12858 3205
rect 12892 3171 12902 3205
rect 12850 3155 12902 3171
rect 12932 3273 12984 3285
rect 12932 3239 12942 3273
rect 12976 3239 12984 3273
rect 13542 3265 13594 3277
rect 12932 3205 12984 3239
rect 12932 3171 12942 3205
rect 12976 3171 12984 3205
rect 12932 3155 12984 3171
rect 13155 3212 13207 3257
rect 13155 3178 13163 3212
rect 13197 3178 13207 3212
rect 13155 3153 13207 3178
rect 13237 3199 13295 3257
rect 13237 3165 13249 3199
rect 13283 3165 13295 3199
rect 13237 3153 13295 3165
rect 13325 3229 13377 3257
rect 13325 3195 13335 3229
rect 13369 3195 13377 3229
rect 13325 3153 13377 3195
rect 13542 3231 13550 3265
rect 13584 3231 13594 3265
rect 13542 3197 13594 3231
rect 13542 3163 13550 3197
rect 13584 3163 13594 3197
rect 13542 3147 13594 3163
rect 13624 3265 13676 3277
rect 13624 3231 13634 3265
rect 13668 3231 13676 3265
rect 13624 3197 13676 3231
rect 14738 3273 14790 3285
rect 14738 3239 14746 3273
rect 14780 3239 14790 3273
rect 14738 3205 14790 3239
rect 13624 3163 13634 3197
rect 13668 3163 13676 3197
rect 13624 3147 13676 3163
rect 14738 3171 14746 3205
rect 14780 3171 14790 3205
rect 14738 3155 14790 3171
rect 14820 3273 14872 3285
rect 14820 3239 14830 3273
rect 14864 3239 14872 3273
rect 15430 3265 15482 3277
rect 14820 3205 14872 3239
rect 14820 3171 14830 3205
rect 14864 3171 14872 3205
rect 14820 3155 14872 3171
rect 15043 3212 15095 3257
rect 15043 3178 15051 3212
rect 15085 3178 15095 3212
rect 15043 3153 15095 3178
rect 15125 3199 15183 3257
rect 15125 3165 15137 3199
rect 15171 3165 15183 3199
rect 15125 3153 15183 3165
rect 15213 3229 15265 3257
rect 15213 3195 15223 3229
rect 15257 3195 15265 3229
rect 15213 3153 15265 3195
rect 15430 3231 15438 3265
rect 15472 3231 15482 3265
rect 15430 3197 15482 3231
rect 15430 3163 15438 3197
rect 15472 3163 15482 3197
rect 15430 3147 15482 3163
rect 15512 3265 15564 3277
rect 15512 3231 15522 3265
rect 15556 3231 15564 3265
rect 15512 3197 15564 3231
rect 16626 3273 16678 3285
rect 16626 3239 16634 3273
rect 16668 3239 16678 3273
rect 16626 3205 16678 3239
rect 15512 3163 15522 3197
rect 15556 3163 15564 3197
rect 15512 3147 15564 3163
rect 16626 3171 16634 3205
rect 16668 3171 16678 3205
rect 16626 3155 16678 3171
rect 16708 3273 16760 3285
rect 16708 3239 16718 3273
rect 16752 3239 16760 3273
rect 17318 3265 17370 3277
rect 16708 3205 16760 3239
rect 16708 3171 16718 3205
rect 16752 3171 16760 3205
rect 16708 3155 16760 3171
rect 16931 3212 16983 3257
rect 16931 3178 16939 3212
rect 16973 3178 16983 3212
rect 16931 3153 16983 3178
rect 17013 3199 17071 3257
rect 17013 3165 17025 3199
rect 17059 3165 17071 3199
rect 17013 3153 17071 3165
rect 17101 3229 17153 3257
rect 17101 3195 17111 3229
rect 17145 3195 17153 3229
rect 17101 3153 17153 3195
rect 17318 3231 17326 3265
rect 17360 3231 17370 3265
rect 17318 3197 17370 3231
rect 17318 3163 17326 3197
rect 17360 3163 17370 3197
rect 17318 3147 17370 3163
rect 17400 3265 17452 3277
rect 17400 3231 17410 3265
rect 17444 3231 17452 3265
rect 17400 3197 17452 3231
rect 18514 3273 18566 3285
rect 18514 3239 18522 3273
rect 18556 3239 18566 3273
rect 18514 3205 18566 3239
rect 17400 3163 17410 3197
rect 17444 3163 17452 3197
rect 17400 3147 17452 3163
rect 18514 3171 18522 3205
rect 18556 3171 18566 3205
rect 18514 3155 18566 3171
rect 18596 3273 18648 3285
rect 18596 3239 18606 3273
rect 18640 3239 18648 3273
rect 19206 3265 19258 3277
rect 18596 3205 18648 3239
rect 18596 3171 18606 3205
rect 18640 3171 18648 3205
rect 18596 3155 18648 3171
rect 18819 3212 18871 3257
rect 18819 3178 18827 3212
rect 18861 3178 18871 3212
rect 18819 3153 18871 3178
rect 18901 3199 18959 3257
rect 18901 3165 18913 3199
rect 18947 3165 18959 3199
rect 18901 3153 18959 3165
rect 18989 3229 19041 3257
rect 18989 3195 18999 3229
rect 19033 3195 19041 3229
rect 18989 3153 19041 3195
rect 19206 3231 19214 3265
rect 19248 3231 19258 3265
rect 19206 3197 19258 3231
rect 19206 3163 19214 3197
rect 19248 3163 19258 3197
rect 19206 3147 19258 3163
rect 19288 3265 19340 3277
rect 19288 3231 19298 3265
rect 19332 3231 19340 3265
rect 19288 3197 19340 3231
rect 20402 3273 20454 3285
rect 20402 3239 20410 3273
rect 20444 3239 20454 3273
rect 20402 3205 20454 3239
rect 19288 3163 19298 3197
rect 19332 3163 19340 3197
rect 19288 3147 19340 3163
rect 20402 3171 20410 3205
rect 20444 3171 20454 3205
rect 20402 3155 20454 3171
rect 20484 3273 20536 3285
rect 20484 3239 20494 3273
rect 20528 3239 20536 3273
rect 21094 3265 21146 3277
rect 20484 3205 20536 3239
rect 20484 3171 20494 3205
rect 20528 3171 20536 3205
rect 20484 3155 20536 3171
rect 20707 3212 20759 3257
rect 20707 3178 20715 3212
rect 20749 3178 20759 3212
rect 20707 3153 20759 3178
rect 20789 3199 20847 3257
rect 20789 3165 20801 3199
rect 20835 3165 20847 3199
rect 20789 3153 20847 3165
rect 20877 3229 20929 3257
rect 20877 3195 20887 3229
rect 20921 3195 20929 3229
rect 20877 3153 20929 3195
rect 21094 3231 21102 3265
rect 21136 3231 21146 3265
rect 21094 3197 21146 3231
rect 21094 3163 21102 3197
rect 21136 3163 21146 3197
rect 21094 3147 21146 3163
rect 21176 3265 21228 3277
rect 21176 3231 21186 3265
rect 21220 3231 21228 3265
rect 21176 3197 21228 3231
rect 22290 3273 22342 3285
rect 22290 3239 22298 3273
rect 22332 3239 22342 3273
rect 22290 3205 22342 3239
rect 21176 3163 21186 3197
rect 21220 3163 21228 3197
rect 21176 3147 21228 3163
rect 22290 3171 22298 3205
rect 22332 3171 22342 3205
rect 22290 3155 22342 3171
rect 22372 3273 22424 3285
rect 22372 3239 22382 3273
rect 22416 3239 22424 3273
rect 22982 3265 23034 3277
rect 22372 3205 22424 3239
rect 22372 3171 22382 3205
rect 22416 3171 22424 3205
rect 22372 3155 22424 3171
rect 22595 3212 22647 3257
rect 22595 3178 22603 3212
rect 22637 3178 22647 3212
rect 22595 3153 22647 3178
rect 22677 3199 22735 3257
rect 22677 3165 22689 3199
rect 22723 3165 22735 3199
rect 22677 3153 22735 3165
rect 22765 3229 22817 3257
rect 22765 3195 22775 3229
rect 22809 3195 22817 3229
rect 22765 3153 22817 3195
rect 22982 3231 22990 3265
rect 23024 3231 23034 3265
rect 22982 3197 23034 3231
rect 22982 3163 22990 3197
rect 23024 3163 23034 3197
rect 22982 3147 23034 3163
rect 23064 3265 23116 3277
rect 23064 3231 23074 3265
rect 23108 3231 23116 3265
rect 23064 3197 23116 3231
rect 24178 3273 24230 3285
rect 24178 3239 24186 3273
rect 24220 3239 24230 3273
rect 24178 3205 24230 3239
rect 23064 3163 23074 3197
rect 23108 3163 23116 3197
rect 23064 3147 23116 3163
rect 24178 3171 24186 3205
rect 24220 3171 24230 3205
rect 24178 3155 24230 3171
rect 24260 3273 24312 3285
rect 24260 3239 24270 3273
rect 24304 3239 24312 3273
rect 24870 3265 24922 3277
rect 24260 3205 24312 3239
rect 24260 3171 24270 3205
rect 24304 3171 24312 3205
rect 24260 3155 24312 3171
rect 24483 3212 24535 3257
rect 24483 3178 24491 3212
rect 24525 3178 24535 3212
rect 24483 3153 24535 3178
rect 24565 3199 24623 3257
rect 24565 3165 24577 3199
rect 24611 3165 24623 3199
rect 24565 3153 24623 3165
rect 24653 3229 24705 3257
rect 24653 3195 24663 3229
rect 24697 3195 24705 3229
rect 24653 3153 24705 3195
rect 24870 3231 24878 3265
rect 24912 3231 24922 3265
rect 24870 3197 24922 3231
rect 24870 3163 24878 3197
rect 24912 3163 24922 3197
rect 24870 3147 24922 3163
rect 24952 3265 25004 3277
rect 24952 3231 24962 3265
rect 24996 3231 25004 3265
rect 24952 3197 25004 3231
rect 26066 3273 26118 3285
rect 26066 3239 26074 3273
rect 26108 3239 26118 3273
rect 26066 3205 26118 3239
rect 24952 3163 24962 3197
rect 24996 3163 25004 3197
rect 24952 3147 25004 3163
rect 26066 3171 26074 3205
rect 26108 3171 26118 3205
rect 26066 3155 26118 3171
rect 26148 3273 26200 3285
rect 26148 3239 26158 3273
rect 26192 3239 26200 3273
rect 26148 3205 26200 3239
rect 26148 3171 26158 3205
rect 26192 3171 26200 3205
rect 26148 3155 26200 3171
rect 26371 3212 26423 3257
rect 26371 3178 26379 3212
rect 26413 3178 26423 3212
rect 26371 3153 26423 3178
rect 26453 3199 26511 3257
rect 26453 3165 26465 3199
rect 26499 3165 26511 3199
rect 26453 3153 26511 3165
rect 26541 3229 26593 3257
rect 26541 3195 26551 3229
rect 26585 3195 26593 3229
rect 26541 3153 26593 3195
rect -2944 3016 -2882 3030
rect -2944 2982 -2932 3016
rect -2898 2982 -2882 3016
rect -2944 2948 -2882 2982
rect -2944 2914 -2932 2948
rect -2898 2914 -2882 2948
rect -2944 2900 -2882 2914
rect -2852 3016 -2786 3030
rect -2852 2982 -2836 3016
rect -2802 2982 -2786 3016
rect -2852 2948 -2786 2982
rect -2852 2914 -2836 2948
rect -2802 2914 -2786 2948
rect -2852 2900 -2786 2914
rect -2756 3016 -2694 3030
rect -2756 2982 -2740 3016
rect -2706 2982 -2694 3016
rect -2756 2948 -2694 2982
rect -2756 2914 -2740 2948
rect -2706 2914 -2694 2948
rect -2756 2900 -2694 2914
rect -1056 3016 -994 3030
rect -1056 2982 -1044 3016
rect -1010 2982 -994 3016
rect -1056 2948 -994 2982
rect -1056 2914 -1044 2948
rect -1010 2914 -994 2948
rect -1056 2900 -994 2914
rect -964 3016 -898 3030
rect -964 2982 -948 3016
rect -914 2982 -898 3016
rect -964 2948 -898 2982
rect -964 2914 -948 2948
rect -914 2914 -898 2948
rect -964 2900 -898 2914
rect -868 3016 -806 3030
rect -868 2982 -852 3016
rect -818 2982 -806 3016
rect -868 2948 -806 2982
rect -868 2914 -852 2948
rect -818 2914 -806 2948
rect -868 2900 -806 2914
rect 832 3016 894 3030
rect 832 2982 844 3016
rect 878 2982 894 3016
rect 832 2948 894 2982
rect 832 2914 844 2948
rect 878 2914 894 2948
rect 832 2900 894 2914
rect 924 3016 990 3030
rect 924 2982 940 3016
rect 974 2982 990 3016
rect 924 2948 990 2982
rect 924 2914 940 2948
rect 974 2914 990 2948
rect 924 2900 990 2914
rect 1020 3016 1082 3030
rect 1020 2982 1036 3016
rect 1070 2982 1082 3016
rect 1020 2948 1082 2982
rect 1020 2914 1036 2948
rect 1070 2914 1082 2948
rect 1020 2900 1082 2914
rect 2720 3016 2782 3030
rect 2720 2982 2732 3016
rect 2766 2982 2782 3016
rect 2720 2948 2782 2982
rect 2720 2914 2732 2948
rect 2766 2914 2782 2948
rect 2720 2900 2782 2914
rect 2812 3016 2878 3030
rect 2812 2982 2828 3016
rect 2862 2982 2878 3016
rect 2812 2948 2878 2982
rect 2812 2914 2828 2948
rect 2862 2914 2878 2948
rect 2812 2900 2878 2914
rect 2908 3016 2970 3030
rect 2908 2982 2924 3016
rect 2958 2982 2970 3016
rect 2908 2948 2970 2982
rect 2908 2914 2924 2948
rect 2958 2914 2970 2948
rect 2908 2900 2970 2914
rect 4608 3016 4670 3030
rect 4608 2982 4620 3016
rect 4654 2982 4670 3016
rect 4608 2948 4670 2982
rect 4608 2914 4620 2948
rect 4654 2914 4670 2948
rect 4608 2900 4670 2914
rect 4700 3016 4766 3030
rect 4700 2982 4716 3016
rect 4750 2982 4766 3016
rect 4700 2948 4766 2982
rect 4700 2914 4716 2948
rect 4750 2914 4766 2948
rect 4700 2900 4766 2914
rect 4796 3016 4858 3030
rect 4796 2982 4812 3016
rect 4846 2982 4858 3016
rect 4796 2948 4858 2982
rect 4796 2914 4812 2948
rect 4846 2914 4858 2948
rect 4796 2900 4858 2914
rect 6496 3016 6558 3030
rect 6496 2982 6508 3016
rect 6542 2982 6558 3016
rect 6496 2948 6558 2982
rect 6496 2914 6508 2948
rect 6542 2914 6558 2948
rect 6496 2900 6558 2914
rect 6588 3016 6654 3030
rect 6588 2982 6604 3016
rect 6638 2982 6654 3016
rect 6588 2948 6654 2982
rect 6588 2914 6604 2948
rect 6638 2914 6654 2948
rect 6588 2900 6654 2914
rect 6684 3016 6746 3030
rect 6684 2982 6700 3016
rect 6734 2982 6746 3016
rect 6684 2948 6746 2982
rect 6684 2914 6700 2948
rect 6734 2914 6746 2948
rect 6684 2900 6746 2914
rect 8384 3016 8446 3030
rect 8384 2982 8396 3016
rect 8430 2982 8446 3016
rect 8384 2948 8446 2982
rect 8384 2914 8396 2948
rect 8430 2914 8446 2948
rect 8384 2900 8446 2914
rect 8476 3016 8542 3030
rect 8476 2982 8492 3016
rect 8526 2982 8542 3016
rect 8476 2948 8542 2982
rect 8476 2914 8492 2948
rect 8526 2914 8542 2948
rect 8476 2900 8542 2914
rect 8572 3016 8634 3030
rect 8572 2982 8588 3016
rect 8622 2982 8634 3016
rect 8572 2948 8634 2982
rect 8572 2914 8588 2948
rect 8622 2914 8634 2948
rect 8572 2900 8634 2914
rect 10272 3016 10334 3030
rect 10272 2982 10284 3016
rect 10318 2982 10334 3016
rect 10272 2948 10334 2982
rect 10272 2914 10284 2948
rect 10318 2914 10334 2948
rect 10272 2900 10334 2914
rect 10364 3016 10430 3030
rect 10364 2982 10380 3016
rect 10414 2982 10430 3016
rect 10364 2948 10430 2982
rect 10364 2914 10380 2948
rect 10414 2914 10430 2948
rect 10364 2900 10430 2914
rect 10460 3016 10522 3030
rect 10460 2982 10476 3016
rect 10510 2982 10522 3016
rect 10460 2948 10522 2982
rect 10460 2914 10476 2948
rect 10510 2914 10522 2948
rect 10460 2900 10522 2914
rect 12154 3016 12216 3030
rect 12154 2982 12166 3016
rect 12200 2982 12216 3016
rect 12154 2948 12216 2982
rect 12154 2914 12166 2948
rect 12200 2914 12216 2948
rect 12154 2900 12216 2914
rect 12246 3016 12312 3030
rect 12246 2982 12262 3016
rect 12296 2982 12312 3016
rect 12246 2948 12312 2982
rect 12246 2914 12262 2948
rect 12296 2914 12312 2948
rect 12246 2900 12312 2914
rect 12342 3016 12404 3030
rect 12342 2982 12358 3016
rect 12392 2982 12404 3016
rect 12342 2948 12404 2982
rect 12342 2914 12358 2948
rect 12392 2914 12404 2948
rect 12342 2900 12404 2914
rect 14042 3016 14104 3030
rect 14042 2982 14054 3016
rect 14088 2982 14104 3016
rect 14042 2948 14104 2982
rect 14042 2914 14054 2948
rect 14088 2914 14104 2948
rect 14042 2900 14104 2914
rect 14134 3016 14200 3030
rect 14134 2982 14150 3016
rect 14184 2982 14200 3016
rect 14134 2948 14200 2982
rect 14134 2914 14150 2948
rect 14184 2914 14200 2948
rect 14134 2900 14200 2914
rect 14230 3016 14292 3030
rect 14230 2982 14246 3016
rect 14280 2982 14292 3016
rect 14230 2948 14292 2982
rect 14230 2914 14246 2948
rect 14280 2914 14292 2948
rect 14230 2900 14292 2914
rect 15930 3016 15992 3030
rect 15930 2982 15942 3016
rect 15976 2982 15992 3016
rect 15930 2948 15992 2982
rect 15930 2914 15942 2948
rect 15976 2914 15992 2948
rect 15930 2900 15992 2914
rect 16022 3016 16088 3030
rect 16022 2982 16038 3016
rect 16072 2982 16088 3016
rect 16022 2948 16088 2982
rect 16022 2914 16038 2948
rect 16072 2914 16088 2948
rect 16022 2900 16088 2914
rect 16118 3016 16180 3030
rect 16118 2982 16134 3016
rect 16168 2982 16180 3016
rect 16118 2948 16180 2982
rect 16118 2914 16134 2948
rect 16168 2914 16180 2948
rect 16118 2900 16180 2914
rect 17818 3016 17880 3030
rect 17818 2982 17830 3016
rect 17864 2982 17880 3016
rect 17818 2948 17880 2982
rect 17818 2914 17830 2948
rect 17864 2914 17880 2948
rect 17818 2900 17880 2914
rect 17910 3016 17976 3030
rect 17910 2982 17926 3016
rect 17960 2982 17976 3016
rect 17910 2948 17976 2982
rect 17910 2914 17926 2948
rect 17960 2914 17976 2948
rect 17910 2900 17976 2914
rect 18006 3016 18068 3030
rect 18006 2982 18022 3016
rect 18056 2982 18068 3016
rect 18006 2948 18068 2982
rect 18006 2914 18022 2948
rect 18056 2914 18068 2948
rect 18006 2900 18068 2914
rect 19706 3016 19768 3030
rect 19706 2982 19718 3016
rect 19752 2982 19768 3016
rect 19706 2948 19768 2982
rect 19706 2914 19718 2948
rect 19752 2914 19768 2948
rect 19706 2900 19768 2914
rect 19798 3016 19864 3030
rect 19798 2982 19814 3016
rect 19848 2982 19864 3016
rect 19798 2948 19864 2982
rect 19798 2914 19814 2948
rect 19848 2914 19864 2948
rect 19798 2900 19864 2914
rect 19894 3016 19956 3030
rect 19894 2982 19910 3016
rect 19944 2982 19956 3016
rect 19894 2948 19956 2982
rect 19894 2914 19910 2948
rect 19944 2914 19956 2948
rect 19894 2900 19956 2914
rect 21594 3016 21656 3030
rect 21594 2982 21606 3016
rect 21640 2982 21656 3016
rect 21594 2948 21656 2982
rect 21594 2914 21606 2948
rect 21640 2914 21656 2948
rect 21594 2900 21656 2914
rect 21686 3016 21752 3030
rect 21686 2982 21702 3016
rect 21736 2982 21752 3016
rect 21686 2948 21752 2982
rect 21686 2914 21702 2948
rect 21736 2914 21752 2948
rect 21686 2900 21752 2914
rect 21782 3016 21844 3030
rect 21782 2982 21798 3016
rect 21832 2982 21844 3016
rect 21782 2948 21844 2982
rect 21782 2914 21798 2948
rect 21832 2914 21844 2948
rect 21782 2900 21844 2914
rect 23482 3016 23544 3030
rect 23482 2982 23494 3016
rect 23528 2982 23544 3016
rect 23482 2948 23544 2982
rect 23482 2914 23494 2948
rect 23528 2914 23544 2948
rect 23482 2900 23544 2914
rect 23574 3016 23640 3030
rect 23574 2982 23590 3016
rect 23624 2982 23640 3016
rect 23574 2948 23640 2982
rect 23574 2914 23590 2948
rect 23624 2914 23640 2948
rect 23574 2900 23640 2914
rect 23670 3016 23732 3030
rect 23670 2982 23686 3016
rect 23720 2982 23732 3016
rect 23670 2948 23732 2982
rect 23670 2914 23686 2948
rect 23720 2914 23732 2948
rect 23670 2900 23732 2914
rect 25370 3016 25432 3030
rect 25370 2982 25382 3016
rect 25416 2982 25432 3016
rect 25370 2948 25432 2982
rect 25370 2914 25382 2948
rect 25416 2914 25432 2948
rect 25370 2900 25432 2914
rect 25462 3016 25528 3030
rect 25462 2982 25478 3016
rect 25512 2982 25528 3016
rect 25462 2948 25528 2982
rect 25462 2914 25478 2948
rect 25512 2914 25528 2948
rect 25462 2900 25528 2914
rect 25558 3016 25620 3030
rect 25558 2982 25574 3016
rect 25608 2982 25620 3016
rect 25558 2948 25620 2982
rect 25558 2914 25574 2948
rect 25608 2914 25620 2948
rect 25558 2900 25620 2914
<< pdiff >>
rect 2152 5009 2204 5025
rect 2152 4975 2160 5009
rect 2194 4975 2204 5009
rect 2152 4939 2204 4975
rect 2152 4905 2160 4939
rect 2194 4905 2204 4939
rect 2152 4871 2204 4905
rect 2152 4837 2160 4871
rect 2194 4837 2204 4871
rect 2152 4825 2204 4837
rect 2234 5009 2288 5025
rect 2234 4975 2244 5009
rect 2278 4975 2288 5009
rect 2234 4939 2288 4975
rect 2234 4905 2244 4939
rect 2278 4905 2288 4939
rect 2234 4871 2288 4905
rect 2234 4837 2244 4871
rect 2278 4837 2288 4871
rect 2234 4825 2288 4837
rect 2318 4939 2372 5025
rect 2318 4905 2328 4939
rect 2362 4905 2372 4939
rect 2318 4871 2372 4905
rect 2318 4837 2328 4871
rect 2362 4837 2372 4871
rect 2318 4825 2372 4837
rect 2402 5009 2456 5025
rect 2402 4975 2412 5009
rect 2446 4975 2456 5009
rect 2402 4939 2456 4975
rect 2402 4905 2412 4939
rect 2446 4905 2456 4939
rect 2402 4871 2456 4905
rect 2402 4837 2412 4871
rect 2446 4837 2456 4871
rect 2402 4825 2456 4837
rect 2486 4939 2540 5025
rect 2486 4905 2496 4939
rect 2530 4905 2540 4939
rect 2486 4871 2540 4905
rect 2486 4837 2496 4871
rect 2530 4837 2540 4871
rect 2486 4825 2540 4837
rect 2570 5009 2624 5025
rect 2570 4975 2580 5009
rect 2614 4975 2624 5009
rect 2570 4939 2624 4975
rect 2570 4905 2580 4939
rect 2614 4905 2624 4939
rect 2570 4871 2624 4905
rect 2570 4837 2580 4871
rect 2614 4837 2624 4871
rect 2570 4825 2624 4837
rect 2654 4939 2708 5025
rect 2654 4905 2664 4939
rect 2698 4905 2708 4939
rect 2654 4871 2708 4905
rect 2654 4837 2664 4871
rect 2698 4837 2708 4871
rect 2654 4825 2708 4837
rect 2738 5009 2792 5025
rect 2738 4975 2748 5009
rect 2782 4975 2792 5009
rect 2738 4939 2792 4975
rect 2738 4905 2748 4939
rect 2782 4905 2792 4939
rect 2738 4871 2792 4905
rect 2738 4837 2748 4871
rect 2782 4837 2792 4871
rect 2738 4825 2792 4837
rect 2822 4939 2876 5025
rect 2822 4905 2832 4939
rect 2866 4905 2876 4939
rect 2822 4871 2876 4905
rect 2822 4837 2832 4871
rect 2866 4837 2876 4871
rect 2822 4825 2876 4837
rect 2906 5009 2960 5025
rect 2906 4975 2916 5009
rect 2950 4975 2960 5009
rect 2906 4939 2960 4975
rect 2906 4905 2916 4939
rect 2950 4905 2960 4939
rect 2906 4871 2960 4905
rect 2906 4837 2916 4871
rect 2950 4837 2960 4871
rect 2906 4825 2960 4837
rect 2990 4939 3044 5025
rect 2990 4905 3000 4939
rect 3034 4905 3044 4939
rect 2990 4871 3044 4905
rect 2990 4837 3000 4871
rect 3034 4837 3044 4871
rect 2990 4825 3044 4837
rect 3074 5009 3128 5025
rect 3074 4975 3084 5009
rect 3118 4975 3128 5009
rect 3074 4939 3128 4975
rect 3074 4905 3084 4939
rect 3118 4905 3128 4939
rect 3074 4871 3128 4905
rect 3074 4837 3084 4871
rect 3118 4837 3128 4871
rect 3074 4825 3128 4837
rect 3158 4939 3212 5025
rect 3158 4905 3168 4939
rect 3202 4905 3212 4939
rect 3158 4871 3212 4905
rect 3158 4837 3168 4871
rect 3202 4837 3212 4871
rect 3158 4825 3212 4837
rect 3242 5009 3296 5025
rect 3242 4975 3252 5009
rect 3286 4975 3296 5009
rect 3242 4939 3296 4975
rect 3242 4905 3252 4939
rect 3286 4905 3296 4939
rect 3242 4871 3296 4905
rect 3242 4837 3252 4871
rect 3286 4837 3296 4871
rect 3242 4825 3296 4837
rect 3326 4939 3380 5025
rect 3326 4905 3336 4939
rect 3370 4905 3380 4939
rect 3326 4871 3380 4905
rect 3326 4837 3336 4871
rect 3370 4837 3380 4871
rect 3326 4825 3380 4837
rect 3410 5009 3464 5025
rect 3410 4975 3420 5009
rect 3454 4975 3464 5009
rect 3410 4939 3464 4975
rect 3410 4905 3420 4939
rect 3454 4905 3464 4939
rect 3410 4871 3464 4905
rect 3410 4837 3420 4871
rect 3454 4837 3464 4871
rect 3410 4825 3464 4837
rect 3494 4939 3546 5025
rect 3494 4905 3504 4939
rect 3538 4905 3546 4939
rect 3494 4871 3546 4905
rect 3494 4837 3504 4871
rect 3538 4837 3546 4871
rect 3494 4825 3546 4837
rect 4034 5007 4086 5023
rect 4034 4973 4042 5007
rect 4076 4973 4086 5007
rect 4034 4937 4086 4973
rect 4034 4903 4042 4937
rect 4076 4903 4086 4937
rect 4034 4869 4086 4903
rect 4034 4835 4042 4869
rect 4076 4835 4086 4869
rect 4034 4823 4086 4835
rect 4116 5007 4170 5023
rect 4116 4973 4126 5007
rect 4160 4973 4170 5007
rect 4116 4937 4170 4973
rect 4116 4903 4126 4937
rect 4160 4903 4170 4937
rect 4116 4869 4170 4903
rect 4116 4835 4126 4869
rect 4160 4835 4170 4869
rect 4116 4823 4170 4835
rect 4200 4937 4254 5023
rect 4200 4903 4210 4937
rect 4244 4903 4254 4937
rect 4200 4869 4254 4903
rect 4200 4835 4210 4869
rect 4244 4835 4254 4869
rect 4200 4823 4254 4835
rect 4284 5007 4338 5023
rect 4284 4973 4294 5007
rect 4328 4973 4338 5007
rect 4284 4937 4338 4973
rect 4284 4903 4294 4937
rect 4328 4903 4338 4937
rect 4284 4869 4338 4903
rect 4284 4835 4294 4869
rect 4328 4835 4338 4869
rect 4284 4823 4338 4835
rect 4368 4937 4422 5023
rect 4368 4903 4378 4937
rect 4412 4903 4422 4937
rect 4368 4869 4422 4903
rect 4368 4835 4378 4869
rect 4412 4835 4422 4869
rect 4368 4823 4422 4835
rect 4452 5007 4506 5023
rect 4452 4973 4462 5007
rect 4496 4973 4506 5007
rect 4452 4937 4506 4973
rect 4452 4903 4462 4937
rect 4496 4903 4506 4937
rect 4452 4869 4506 4903
rect 4452 4835 4462 4869
rect 4496 4835 4506 4869
rect 4452 4823 4506 4835
rect 4536 4937 4590 5023
rect 4536 4903 4546 4937
rect 4580 4903 4590 4937
rect 4536 4869 4590 4903
rect 4536 4835 4546 4869
rect 4580 4835 4590 4869
rect 4536 4823 4590 4835
rect 4620 5007 4674 5023
rect 4620 4973 4630 5007
rect 4664 4973 4674 5007
rect 4620 4937 4674 4973
rect 4620 4903 4630 4937
rect 4664 4903 4674 4937
rect 4620 4869 4674 4903
rect 4620 4835 4630 4869
rect 4664 4835 4674 4869
rect 4620 4823 4674 4835
rect 4704 4937 4758 5023
rect 4704 4903 4714 4937
rect 4748 4903 4758 4937
rect 4704 4869 4758 4903
rect 4704 4835 4714 4869
rect 4748 4835 4758 4869
rect 4704 4823 4758 4835
rect 4788 5007 4842 5023
rect 4788 4973 4798 5007
rect 4832 4973 4842 5007
rect 4788 4937 4842 4973
rect 4788 4903 4798 4937
rect 4832 4903 4842 4937
rect 4788 4869 4842 4903
rect 4788 4835 4798 4869
rect 4832 4835 4842 4869
rect 4788 4823 4842 4835
rect 4872 4937 4926 5023
rect 4872 4903 4882 4937
rect 4916 4903 4926 4937
rect 4872 4869 4926 4903
rect 4872 4835 4882 4869
rect 4916 4835 4926 4869
rect 4872 4823 4926 4835
rect 4956 5007 5010 5023
rect 4956 4973 4966 5007
rect 5000 4973 5010 5007
rect 4956 4937 5010 4973
rect 4956 4903 4966 4937
rect 5000 4903 5010 4937
rect 4956 4869 5010 4903
rect 4956 4835 4966 4869
rect 5000 4835 5010 4869
rect 4956 4823 5010 4835
rect 5040 4937 5094 5023
rect 5040 4903 5050 4937
rect 5084 4903 5094 4937
rect 5040 4869 5094 4903
rect 5040 4835 5050 4869
rect 5084 4835 5094 4869
rect 5040 4823 5094 4835
rect 5124 5007 5178 5023
rect 5124 4973 5134 5007
rect 5168 4973 5178 5007
rect 5124 4937 5178 4973
rect 5124 4903 5134 4937
rect 5168 4903 5178 4937
rect 5124 4869 5178 4903
rect 5124 4835 5134 4869
rect 5168 4835 5178 4869
rect 5124 4823 5178 4835
rect 5208 4937 5262 5023
rect 5208 4903 5218 4937
rect 5252 4903 5262 4937
rect 5208 4869 5262 4903
rect 5208 4835 5218 4869
rect 5252 4835 5262 4869
rect 5208 4823 5262 4835
rect 5292 5007 5346 5023
rect 5292 4973 5302 5007
rect 5336 4973 5346 5007
rect 5292 4937 5346 4973
rect 5292 4903 5302 4937
rect 5336 4903 5346 4937
rect 5292 4869 5346 4903
rect 5292 4835 5302 4869
rect 5336 4835 5346 4869
rect 5292 4823 5346 4835
rect 5376 4937 5428 5023
rect 5376 4903 5386 4937
rect 5420 4903 5428 4937
rect 5376 4869 5428 4903
rect 5376 4835 5386 4869
rect 5420 4835 5428 4869
rect 5376 4823 5428 4835
rect 17250 5009 17302 5025
rect 17250 4975 17258 5009
rect 17292 4975 17302 5009
rect 17250 4939 17302 4975
rect 17250 4905 17258 4939
rect 17292 4905 17302 4939
rect 17250 4871 17302 4905
rect 17250 4837 17258 4871
rect 17292 4837 17302 4871
rect 17250 4825 17302 4837
rect 17332 5009 17386 5025
rect 17332 4975 17342 5009
rect 17376 4975 17386 5009
rect 17332 4939 17386 4975
rect 17332 4905 17342 4939
rect 17376 4905 17386 4939
rect 17332 4871 17386 4905
rect 17332 4837 17342 4871
rect 17376 4837 17386 4871
rect 17332 4825 17386 4837
rect 17416 4939 17470 5025
rect 17416 4905 17426 4939
rect 17460 4905 17470 4939
rect 17416 4871 17470 4905
rect 17416 4837 17426 4871
rect 17460 4837 17470 4871
rect 17416 4825 17470 4837
rect 17500 5009 17554 5025
rect 17500 4975 17510 5009
rect 17544 4975 17554 5009
rect 17500 4939 17554 4975
rect 17500 4905 17510 4939
rect 17544 4905 17554 4939
rect 17500 4871 17554 4905
rect 17500 4837 17510 4871
rect 17544 4837 17554 4871
rect 17500 4825 17554 4837
rect 17584 4939 17638 5025
rect 17584 4905 17594 4939
rect 17628 4905 17638 4939
rect 17584 4871 17638 4905
rect 17584 4837 17594 4871
rect 17628 4837 17638 4871
rect 17584 4825 17638 4837
rect 17668 5009 17722 5025
rect 17668 4975 17678 5009
rect 17712 4975 17722 5009
rect 17668 4939 17722 4975
rect 17668 4905 17678 4939
rect 17712 4905 17722 4939
rect 17668 4871 17722 4905
rect 17668 4837 17678 4871
rect 17712 4837 17722 4871
rect 17668 4825 17722 4837
rect 17752 4939 17806 5025
rect 17752 4905 17762 4939
rect 17796 4905 17806 4939
rect 17752 4871 17806 4905
rect 17752 4837 17762 4871
rect 17796 4837 17806 4871
rect 17752 4825 17806 4837
rect 17836 5009 17890 5025
rect 17836 4975 17846 5009
rect 17880 4975 17890 5009
rect 17836 4939 17890 4975
rect 17836 4905 17846 4939
rect 17880 4905 17890 4939
rect 17836 4871 17890 4905
rect 17836 4837 17846 4871
rect 17880 4837 17890 4871
rect 17836 4825 17890 4837
rect 17920 4939 17974 5025
rect 17920 4905 17930 4939
rect 17964 4905 17974 4939
rect 17920 4871 17974 4905
rect 17920 4837 17930 4871
rect 17964 4837 17974 4871
rect 17920 4825 17974 4837
rect 18004 5009 18058 5025
rect 18004 4975 18014 5009
rect 18048 4975 18058 5009
rect 18004 4939 18058 4975
rect 18004 4905 18014 4939
rect 18048 4905 18058 4939
rect 18004 4871 18058 4905
rect 18004 4837 18014 4871
rect 18048 4837 18058 4871
rect 18004 4825 18058 4837
rect 18088 4939 18142 5025
rect 18088 4905 18098 4939
rect 18132 4905 18142 4939
rect 18088 4871 18142 4905
rect 18088 4837 18098 4871
rect 18132 4837 18142 4871
rect 18088 4825 18142 4837
rect 18172 5009 18226 5025
rect 18172 4975 18182 5009
rect 18216 4975 18226 5009
rect 18172 4939 18226 4975
rect 18172 4905 18182 4939
rect 18216 4905 18226 4939
rect 18172 4871 18226 4905
rect 18172 4837 18182 4871
rect 18216 4837 18226 4871
rect 18172 4825 18226 4837
rect 18256 4939 18310 5025
rect 18256 4905 18266 4939
rect 18300 4905 18310 4939
rect 18256 4871 18310 4905
rect 18256 4837 18266 4871
rect 18300 4837 18310 4871
rect 18256 4825 18310 4837
rect 18340 5009 18394 5025
rect 18340 4975 18350 5009
rect 18384 4975 18394 5009
rect 18340 4939 18394 4975
rect 18340 4905 18350 4939
rect 18384 4905 18394 4939
rect 18340 4871 18394 4905
rect 18340 4837 18350 4871
rect 18384 4837 18394 4871
rect 18340 4825 18394 4837
rect 18424 4939 18478 5025
rect 18424 4905 18434 4939
rect 18468 4905 18478 4939
rect 18424 4871 18478 4905
rect 18424 4837 18434 4871
rect 18468 4837 18478 4871
rect 18424 4825 18478 4837
rect 18508 5009 18562 5025
rect 18508 4975 18518 5009
rect 18552 4975 18562 5009
rect 18508 4939 18562 4975
rect 18508 4905 18518 4939
rect 18552 4905 18562 4939
rect 18508 4871 18562 4905
rect 18508 4837 18518 4871
rect 18552 4837 18562 4871
rect 18508 4825 18562 4837
rect 18592 4939 18644 5025
rect 18592 4905 18602 4939
rect 18636 4905 18644 4939
rect 18592 4871 18644 4905
rect 18592 4837 18602 4871
rect 18636 4837 18644 4871
rect 18592 4825 18644 4837
rect 19132 5007 19184 5023
rect 19132 4973 19140 5007
rect 19174 4973 19184 5007
rect 19132 4937 19184 4973
rect 19132 4903 19140 4937
rect 19174 4903 19184 4937
rect 19132 4869 19184 4903
rect 19132 4835 19140 4869
rect 19174 4835 19184 4869
rect 19132 4823 19184 4835
rect 19214 5007 19268 5023
rect 19214 4973 19224 5007
rect 19258 4973 19268 5007
rect 19214 4937 19268 4973
rect 19214 4903 19224 4937
rect 19258 4903 19268 4937
rect 19214 4869 19268 4903
rect 19214 4835 19224 4869
rect 19258 4835 19268 4869
rect 19214 4823 19268 4835
rect 19298 4937 19352 5023
rect 19298 4903 19308 4937
rect 19342 4903 19352 4937
rect 19298 4869 19352 4903
rect 19298 4835 19308 4869
rect 19342 4835 19352 4869
rect 19298 4823 19352 4835
rect 19382 5007 19436 5023
rect 19382 4973 19392 5007
rect 19426 4973 19436 5007
rect 19382 4937 19436 4973
rect 19382 4903 19392 4937
rect 19426 4903 19436 4937
rect 19382 4869 19436 4903
rect 19382 4835 19392 4869
rect 19426 4835 19436 4869
rect 19382 4823 19436 4835
rect 19466 4937 19520 5023
rect 19466 4903 19476 4937
rect 19510 4903 19520 4937
rect 19466 4869 19520 4903
rect 19466 4835 19476 4869
rect 19510 4835 19520 4869
rect 19466 4823 19520 4835
rect 19550 5007 19604 5023
rect 19550 4973 19560 5007
rect 19594 4973 19604 5007
rect 19550 4937 19604 4973
rect 19550 4903 19560 4937
rect 19594 4903 19604 4937
rect 19550 4869 19604 4903
rect 19550 4835 19560 4869
rect 19594 4835 19604 4869
rect 19550 4823 19604 4835
rect 19634 4937 19688 5023
rect 19634 4903 19644 4937
rect 19678 4903 19688 4937
rect 19634 4869 19688 4903
rect 19634 4835 19644 4869
rect 19678 4835 19688 4869
rect 19634 4823 19688 4835
rect 19718 5007 19772 5023
rect 19718 4973 19728 5007
rect 19762 4973 19772 5007
rect 19718 4937 19772 4973
rect 19718 4903 19728 4937
rect 19762 4903 19772 4937
rect 19718 4869 19772 4903
rect 19718 4835 19728 4869
rect 19762 4835 19772 4869
rect 19718 4823 19772 4835
rect 19802 4937 19856 5023
rect 19802 4903 19812 4937
rect 19846 4903 19856 4937
rect 19802 4869 19856 4903
rect 19802 4835 19812 4869
rect 19846 4835 19856 4869
rect 19802 4823 19856 4835
rect 19886 5007 19940 5023
rect 19886 4973 19896 5007
rect 19930 4973 19940 5007
rect 19886 4937 19940 4973
rect 19886 4903 19896 4937
rect 19930 4903 19940 4937
rect 19886 4869 19940 4903
rect 19886 4835 19896 4869
rect 19930 4835 19940 4869
rect 19886 4823 19940 4835
rect 19970 4937 20024 5023
rect 19970 4903 19980 4937
rect 20014 4903 20024 4937
rect 19970 4869 20024 4903
rect 19970 4835 19980 4869
rect 20014 4835 20024 4869
rect 19970 4823 20024 4835
rect 20054 5007 20108 5023
rect 20054 4973 20064 5007
rect 20098 4973 20108 5007
rect 20054 4937 20108 4973
rect 20054 4903 20064 4937
rect 20098 4903 20108 4937
rect 20054 4869 20108 4903
rect 20054 4835 20064 4869
rect 20098 4835 20108 4869
rect 20054 4823 20108 4835
rect 20138 4937 20192 5023
rect 20138 4903 20148 4937
rect 20182 4903 20192 4937
rect 20138 4869 20192 4903
rect 20138 4835 20148 4869
rect 20182 4835 20192 4869
rect 20138 4823 20192 4835
rect 20222 5007 20276 5023
rect 20222 4973 20232 5007
rect 20266 4973 20276 5007
rect 20222 4937 20276 4973
rect 20222 4903 20232 4937
rect 20266 4903 20276 4937
rect 20222 4869 20276 4903
rect 20222 4835 20232 4869
rect 20266 4835 20276 4869
rect 20222 4823 20276 4835
rect 20306 4937 20360 5023
rect 20306 4903 20316 4937
rect 20350 4903 20360 4937
rect 20306 4869 20360 4903
rect 20306 4835 20316 4869
rect 20350 4835 20360 4869
rect 20306 4823 20360 4835
rect 20390 5007 20444 5023
rect 20390 4973 20400 5007
rect 20434 4973 20444 5007
rect 20390 4937 20444 4973
rect 20390 4903 20400 4937
rect 20434 4903 20444 4937
rect 20390 4869 20444 4903
rect 20390 4835 20400 4869
rect 20434 4835 20444 4869
rect 20390 4823 20444 4835
rect 20474 4937 20526 5023
rect 20474 4903 20484 4937
rect 20518 4903 20526 4937
rect 20474 4869 20526 4903
rect 20474 4835 20484 4869
rect 20518 4835 20526 4869
rect 20474 4823 20526 4835
rect -3307 4639 -3255 4651
rect -3307 4605 -3299 4639
rect -3265 4605 -3255 4639
rect -3307 4571 -3255 4605
rect -3307 4537 -3299 4571
rect -3265 4537 -3255 4571
rect -3307 4503 -3255 4537
rect -3307 4469 -3299 4503
rect -3265 4469 -3255 4503
rect -3307 4451 -3255 4469
rect -3225 4451 -3183 4651
rect -3153 4639 -3101 4651
rect -3153 4605 -3143 4639
rect -3109 4605 -3101 4639
rect -2493 4639 -2441 4651
rect -3153 4571 -3101 4605
rect -2493 4605 -2485 4639
rect -2451 4605 -2441 4639
rect -3153 4537 -3143 4571
rect -3109 4537 -3101 4571
rect -3153 4503 -3101 4537
rect -2493 4571 -2441 4605
rect -2493 4537 -2485 4571
rect -2451 4537 -2441 4571
rect -3153 4469 -3143 4503
rect -3109 4469 -3101 4503
rect -2493 4503 -2441 4537
rect -3153 4451 -3101 4469
rect -2958 4471 -2896 4486
rect -2958 4437 -2946 4471
rect -2912 4437 -2896 4471
rect -2958 4403 -2896 4437
rect -2958 4369 -2946 4403
rect -2912 4369 -2896 4403
rect -2958 4335 -2896 4369
rect -2958 4301 -2946 4335
rect -2912 4301 -2896 4335
rect -2958 4286 -2896 4301
rect -2866 4471 -2800 4486
rect -2866 4437 -2850 4471
rect -2816 4437 -2800 4471
rect -2866 4403 -2800 4437
rect -2866 4369 -2850 4403
rect -2816 4369 -2800 4403
rect -2866 4335 -2800 4369
rect -2866 4301 -2850 4335
rect -2816 4301 -2800 4335
rect -2866 4286 -2800 4301
rect -2770 4471 -2708 4486
rect -2770 4437 -2754 4471
rect -2720 4437 -2708 4471
rect -2493 4469 -2485 4503
rect -2451 4469 -2441 4503
rect -2493 4451 -2441 4469
rect -2411 4451 -2369 4651
rect -2339 4639 -2287 4651
rect -2339 4605 -2329 4639
rect -2295 4605 -2287 4639
rect -2339 4571 -2287 4605
rect -2339 4537 -2329 4571
rect -2295 4537 -2287 4571
rect -2339 4503 -2287 4537
rect -2339 4469 -2329 4503
rect -2295 4469 -2287 4503
rect -2339 4451 -2287 4469
rect -1419 4639 -1367 4651
rect -1419 4605 -1411 4639
rect -1377 4605 -1367 4639
rect -1419 4571 -1367 4605
rect -1419 4537 -1411 4571
rect -1377 4537 -1367 4571
rect -1419 4503 -1367 4537
rect -1419 4469 -1411 4503
rect -1377 4469 -1367 4503
rect -1419 4451 -1367 4469
rect -1337 4451 -1295 4651
rect -1265 4639 -1213 4651
rect -1265 4605 -1255 4639
rect -1221 4605 -1213 4639
rect -605 4639 -553 4651
rect -1265 4571 -1213 4605
rect -605 4605 -597 4639
rect -563 4605 -553 4639
rect -1265 4537 -1255 4571
rect -1221 4537 -1213 4571
rect -1265 4503 -1213 4537
rect -605 4571 -553 4605
rect -605 4537 -597 4571
rect -563 4537 -553 4571
rect -1265 4469 -1255 4503
rect -1221 4469 -1213 4503
rect -605 4503 -553 4537
rect -1265 4451 -1213 4469
rect -1070 4471 -1008 4486
rect -2770 4403 -2708 4437
rect -2770 4369 -2754 4403
rect -2720 4369 -2708 4403
rect -2770 4335 -2708 4369
rect -2770 4301 -2754 4335
rect -2720 4301 -2708 4335
rect -1070 4437 -1058 4471
rect -1024 4437 -1008 4471
rect -1070 4403 -1008 4437
rect -1070 4369 -1058 4403
rect -1024 4369 -1008 4403
rect -1070 4335 -1008 4369
rect -2770 4286 -2708 4301
rect -1070 4301 -1058 4335
rect -1024 4301 -1008 4335
rect -1070 4286 -1008 4301
rect -978 4471 -912 4486
rect -978 4437 -962 4471
rect -928 4437 -912 4471
rect -978 4403 -912 4437
rect -978 4369 -962 4403
rect -928 4369 -912 4403
rect -978 4335 -912 4369
rect -978 4301 -962 4335
rect -928 4301 -912 4335
rect -978 4286 -912 4301
rect -882 4471 -820 4486
rect -882 4437 -866 4471
rect -832 4437 -820 4471
rect -605 4469 -597 4503
rect -563 4469 -553 4503
rect -605 4451 -553 4469
rect -523 4451 -481 4651
rect -451 4639 -399 4651
rect -451 4605 -441 4639
rect -407 4605 -399 4639
rect -451 4571 -399 4605
rect -451 4537 -441 4571
rect -407 4537 -399 4571
rect -451 4503 -399 4537
rect -451 4469 -441 4503
rect -407 4469 -399 4503
rect -451 4451 -399 4469
rect 469 4639 521 4651
rect 469 4605 477 4639
rect 511 4605 521 4639
rect 469 4571 521 4605
rect 469 4537 477 4571
rect 511 4537 521 4571
rect 469 4503 521 4537
rect 469 4469 477 4503
rect 511 4469 521 4503
rect 469 4451 521 4469
rect 551 4451 593 4651
rect 623 4639 675 4651
rect 623 4605 633 4639
rect 667 4605 675 4639
rect 1283 4639 1335 4651
rect 623 4571 675 4605
rect 1283 4605 1291 4639
rect 1325 4605 1335 4639
rect 623 4537 633 4571
rect 667 4537 675 4571
rect 623 4503 675 4537
rect 1283 4571 1335 4605
rect 1283 4537 1291 4571
rect 1325 4537 1335 4571
rect 623 4469 633 4503
rect 667 4469 675 4503
rect 1283 4503 1335 4537
rect 623 4451 675 4469
rect 818 4471 880 4486
rect -882 4403 -820 4437
rect -882 4369 -866 4403
rect -832 4369 -820 4403
rect -882 4335 -820 4369
rect -882 4301 -866 4335
rect -832 4301 -820 4335
rect 818 4437 830 4471
rect 864 4437 880 4471
rect 818 4403 880 4437
rect 818 4369 830 4403
rect 864 4369 880 4403
rect 818 4335 880 4369
rect -882 4286 -820 4301
rect 818 4301 830 4335
rect 864 4301 880 4335
rect 818 4286 880 4301
rect 910 4471 976 4486
rect 910 4437 926 4471
rect 960 4437 976 4471
rect 910 4403 976 4437
rect 910 4369 926 4403
rect 960 4369 976 4403
rect 910 4335 976 4369
rect 910 4301 926 4335
rect 960 4301 976 4335
rect 910 4286 976 4301
rect 1006 4471 1068 4486
rect 1006 4437 1022 4471
rect 1056 4437 1068 4471
rect 1283 4469 1291 4503
rect 1325 4469 1335 4503
rect 1283 4451 1335 4469
rect 1365 4451 1407 4651
rect 1437 4639 1489 4651
rect 1437 4605 1447 4639
rect 1481 4605 1489 4639
rect 1437 4571 1489 4605
rect 1437 4537 1447 4571
rect 1481 4537 1489 4571
rect 1437 4503 1489 4537
rect 1437 4469 1447 4503
rect 1481 4469 1489 4503
rect 1437 4451 1489 4469
rect 2357 4639 2409 4651
rect 2357 4605 2365 4639
rect 2399 4605 2409 4639
rect 2357 4571 2409 4605
rect 2357 4537 2365 4571
rect 2399 4537 2409 4571
rect 2357 4503 2409 4537
rect 2357 4469 2365 4503
rect 2399 4469 2409 4503
rect 2357 4451 2409 4469
rect 2439 4451 2481 4651
rect 2511 4639 2563 4651
rect 2511 4605 2521 4639
rect 2555 4605 2563 4639
rect 3171 4639 3223 4651
rect 2511 4571 2563 4605
rect 3171 4605 3179 4639
rect 3213 4605 3223 4639
rect 2511 4537 2521 4571
rect 2555 4537 2563 4571
rect 2511 4503 2563 4537
rect 3171 4571 3223 4605
rect 3171 4537 3179 4571
rect 3213 4537 3223 4571
rect 2511 4469 2521 4503
rect 2555 4469 2563 4503
rect 3171 4503 3223 4537
rect 2511 4451 2563 4469
rect 2706 4471 2768 4486
rect 1006 4403 1068 4437
rect 1006 4369 1022 4403
rect 1056 4369 1068 4403
rect 1006 4335 1068 4369
rect 1006 4301 1022 4335
rect 1056 4301 1068 4335
rect 2706 4437 2718 4471
rect 2752 4437 2768 4471
rect 2706 4403 2768 4437
rect 2706 4369 2718 4403
rect 2752 4369 2768 4403
rect 2706 4335 2768 4369
rect 1006 4286 1068 4301
rect 2706 4301 2718 4335
rect 2752 4301 2768 4335
rect 2706 4286 2768 4301
rect 2798 4471 2864 4486
rect 2798 4437 2814 4471
rect 2848 4437 2864 4471
rect 2798 4403 2864 4437
rect 2798 4369 2814 4403
rect 2848 4369 2864 4403
rect 2798 4335 2864 4369
rect 2798 4301 2814 4335
rect 2848 4301 2864 4335
rect 2798 4286 2864 4301
rect 2894 4471 2956 4486
rect 2894 4437 2910 4471
rect 2944 4437 2956 4471
rect 3171 4469 3179 4503
rect 3213 4469 3223 4503
rect 3171 4451 3223 4469
rect 3253 4451 3295 4651
rect 3325 4639 3377 4651
rect 3325 4605 3335 4639
rect 3369 4605 3377 4639
rect 3325 4571 3377 4605
rect 3325 4537 3335 4571
rect 3369 4537 3377 4571
rect 3325 4503 3377 4537
rect 3325 4469 3335 4503
rect 3369 4469 3377 4503
rect 3325 4451 3377 4469
rect 4245 4639 4297 4651
rect 4245 4605 4253 4639
rect 4287 4605 4297 4639
rect 4245 4571 4297 4605
rect 4245 4537 4253 4571
rect 4287 4537 4297 4571
rect 4245 4503 4297 4537
rect 4245 4469 4253 4503
rect 4287 4469 4297 4503
rect 4245 4451 4297 4469
rect 4327 4451 4369 4651
rect 4399 4639 4451 4651
rect 4399 4605 4409 4639
rect 4443 4605 4451 4639
rect 5059 4639 5111 4651
rect 4399 4571 4451 4605
rect 5059 4605 5067 4639
rect 5101 4605 5111 4639
rect 4399 4537 4409 4571
rect 4443 4537 4451 4571
rect 4399 4503 4451 4537
rect 5059 4571 5111 4605
rect 5059 4537 5067 4571
rect 5101 4537 5111 4571
rect 4399 4469 4409 4503
rect 4443 4469 4451 4503
rect 5059 4503 5111 4537
rect 4399 4451 4451 4469
rect 4594 4471 4656 4486
rect 2894 4403 2956 4437
rect 2894 4369 2910 4403
rect 2944 4369 2956 4403
rect 2894 4335 2956 4369
rect 2894 4301 2910 4335
rect 2944 4301 2956 4335
rect 4594 4437 4606 4471
rect 4640 4437 4656 4471
rect 4594 4403 4656 4437
rect 4594 4369 4606 4403
rect 4640 4369 4656 4403
rect 4594 4335 4656 4369
rect 2894 4286 2956 4301
rect 4594 4301 4606 4335
rect 4640 4301 4656 4335
rect 4594 4286 4656 4301
rect 4686 4471 4752 4486
rect 4686 4437 4702 4471
rect 4736 4437 4752 4471
rect 4686 4403 4752 4437
rect 4686 4369 4702 4403
rect 4736 4369 4752 4403
rect 4686 4335 4752 4369
rect 4686 4301 4702 4335
rect 4736 4301 4752 4335
rect 4686 4286 4752 4301
rect 4782 4471 4844 4486
rect 4782 4437 4798 4471
rect 4832 4437 4844 4471
rect 5059 4469 5067 4503
rect 5101 4469 5111 4503
rect 5059 4451 5111 4469
rect 5141 4451 5183 4651
rect 5213 4639 5265 4651
rect 5213 4605 5223 4639
rect 5257 4605 5265 4639
rect 5213 4571 5265 4605
rect 5213 4537 5223 4571
rect 5257 4537 5265 4571
rect 5213 4503 5265 4537
rect 5213 4469 5223 4503
rect 5257 4469 5265 4503
rect 5213 4451 5265 4469
rect 6133 4639 6185 4651
rect 6133 4605 6141 4639
rect 6175 4605 6185 4639
rect 6133 4571 6185 4605
rect 6133 4537 6141 4571
rect 6175 4537 6185 4571
rect 6133 4503 6185 4537
rect 6133 4469 6141 4503
rect 6175 4469 6185 4503
rect 6133 4451 6185 4469
rect 6215 4451 6257 4651
rect 6287 4639 6339 4651
rect 6287 4605 6297 4639
rect 6331 4605 6339 4639
rect 6947 4639 6999 4651
rect 6287 4571 6339 4605
rect 6947 4605 6955 4639
rect 6989 4605 6999 4639
rect 6287 4537 6297 4571
rect 6331 4537 6339 4571
rect 6287 4503 6339 4537
rect 6947 4571 6999 4605
rect 6947 4537 6955 4571
rect 6989 4537 6999 4571
rect 6287 4469 6297 4503
rect 6331 4469 6339 4503
rect 6947 4503 6999 4537
rect 6287 4451 6339 4469
rect 6482 4471 6544 4486
rect 4782 4403 4844 4437
rect 4782 4369 4798 4403
rect 4832 4369 4844 4403
rect 4782 4335 4844 4369
rect 4782 4301 4798 4335
rect 4832 4301 4844 4335
rect 6482 4437 6494 4471
rect 6528 4437 6544 4471
rect 6482 4403 6544 4437
rect 6482 4369 6494 4403
rect 6528 4369 6544 4403
rect 6482 4335 6544 4369
rect 4782 4286 4844 4301
rect 6482 4301 6494 4335
rect 6528 4301 6544 4335
rect 6482 4286 6544 4301
rect 6574 4471 6640 4486
rect 6574 4437 6590 4471
rect 6624 4437 6640 4471
rect 6574 4403 6640 4437
rect 6574 4369 6590 4403
rect 6624 4369 6640 4403
rect 6574 4335 6640 4369
rect 6574 4301 6590 4335
rect 6624 4301 6640 4335
rect 6574 4286 6640 4301
rect 6670 4471 6732 4486
rect 6670 4437 6686 4471
rect 6720 4437 6732 4471
rect 6947 4469 6955 4503
rect 6989 4469 6999 4503
rect 6947 4451 6999 4469
rect 7029 4451 7071 4651
rect 7101 4639 7153 4651
rect 7101 4605 7111 4639
rect 7145 4605 7153 4639
rect 7101 4571 7153 4605
rect 7101 4537 7111 4571
rect 7145 4537 7153 4571
rect 7101 4503 7153 4537
rect 7101 4469 7111 4503
rect 7145 4469 7153 4503
rect 7101 4451 7153 4469
rect 8021 4639 8073 4651
rect 8021 4605 8029 4639
rect 8063 4605 8073 4639
rect 8021 4571 8073 4605
rect 8021 4537 8029 4571
rect 8063 4537 8073 4571
rect 8021 4503 8073 4537
rect 8021 4469 8029 4503
rect 8063 4469 8073 4503
rect 8021 4451 8073 4469
rect 8103 4451 8145 4651
rect 8175 4639 8227 4651
rect 8175 4605 8185 4639
rect 8219 4605 8227 4639
rect 8835 4639 8887 4651
rect 8175 4571 8227 4605
rect 8835 4605 8843 4639
rect 8877 4605 8887 4639
rect 8175 4537 8185 4571
rect 8219 4537 8227 4571
rect 8175 4503 8227 4537
rect 8835 4571 8887 4605
rect 8835 4537 8843 4571
rect 8877 4537 8887 4571
rect 8175 4469 8185 4503
rect 8219 4469 8227 4503
rect 8835 4503 8887 4537
rect 8175 4451 8227 4469
rect 8370 4471 8432 4486
rect 6670 4403 6732 4437
rect 6670 4369 6686 4403
rect 6720 4369 6732 4403
rect 6670 4335 6732 4369
rect 6670 4301 6686 4335
rect 6720 4301 6732 4335
rect 8370 4437 8382 4471
rect 8416 4437 8432 4471
rect 8370 4403 8432 4437
rect 8370 4369 8382 4403
rect 8416 4369 8432 4403
rect 8370 4335 8432 4369
rect 6670 4286 6732 4301
rect 8370 4301 8382 4335
rect 8416 4301 8432 4335
rect 8370 4286 8432 4301
rect 8462 4471 8528 4486
rect 8462 4437 8478 4471
rect 8512 4437 8528 4471
rect 8462 4403 8528 4437
rect 8462 4369 8478 4403
rect 8512 4369 8528 4403
rect 8462 4335 8528 4369
rect 8462 4301 8478 4335
rect 8512 4301 8528 4335
rect 8462 4286 8528 4301
rect 8558 4471 8620 4486
rect 8558 4437 8574 4471
rect 8608 4437 8620 4471
rect 8835 4469 8843 4503
rect 8877 4469 8887 4503
rect 8835 4451 8887 4469
rect 8917 4451 8959 4651
rect 8989 4639 9041 4651
rect 8989 4605 8999 4639
rect 9033 4605 9041 4639
rect 8989 4571 9041 4605
rect 8989 4537 8999 4571
rect 9033 4537 9041 4571
rect 8989 4503 9041 4537
rect 8989 4469 8999 4503
rect 9033 4469 9041 4503
rect 8989 4451 9041 4469
rect 9909 4639 9961 4651
rect 9909 4605 9917 4639
rect 9951 4605 9961 4639
rect 9909 4571 9961 4605
rect 9909 4537 9917 4571
rect 9951 4537 9961 4571
rect 9909 4503 9961 4537
rect 9909 4469 9917 4503
rect 9951 4469 9961 4503
rect 9909 4451 9961 4469
rect 9991 4451 10033 4651
rect 10063 4639 10115 4651
rect 10063 4605 10073 4639
rect 10107 4605 10115 4639
rect 10723 4639 10775 4651
rect 10063 4571 10115 4605
rect 10723 4605 10731 4639
rect 10765 4605 10775 4639
rect 10063 4537 10073 4571
rect 10107 4537 10115 4571
rect 10063 4503 10115 4537
rect 10723 4571 10775 4605
rect 10723 4537 10731 4571
rect 10765 4537 10775 4571
rect 10063 4469 10073 4503
rect 10107 4469 10115 4503
rect 10723 4503 10775 4537
rect 10063 4451 10115 4469
rect 10258 4471 10320 4486
rect 8558 4403 8620 4437
rect 8558 4369 8574 4403
rect 8608 4369 8620 4403
rect 8558 4335 8620 4369
rect 8558 4301 8574 4335
rect 8608 4301 8620 4335
rect 10258 4437 10270 4471
rect 10304 4437 10320 4471
rect 10258 4403 10320 4437
rect 10258 4369 10270 4403
rect 10304 4369 10320 4403
rect 10258 4335 10320 4369
rect 8558 4286 8620 4301
rect 10258 4301 10270 4335
rect 10304 4301 10320 4335
rect 10258 4286 10320 4301
rect 10350 4471 10416 4486
rect 10350 4437 10366 4471
rect 10400 4437 10416 4471
rect 10350 4403 10416 4437
rect 10350 4369 10366 4403
rect 10400 4369 10416 4403
rect 10350 4335 10416 4369
rect 10350 4301 10366 4335
rect 10400 4301 10416 4335
rect 10350 4286 10416 4301
rect 10446 4471 10508 4486
rect 10446 4437 10462 4471
rect 10496 4437 10508 4471
rect 10723 4469 10731 4503
rect 10765 4469 10775 4503
rect 10723 4451 10775 4469
rect 10805 4451 10847 4651
rect 10877 4639 10929 4651
rect 10877 4605 10887 4639
rect 10921 4605 10929 4639
rect 10877 4571 10929 4605
rect 10877 4537 10887 4571
rect 10921 4537 10929 4571
rect 10877 4503 10929 4537
rect 10877 4469 10887 4503
rect 10921 4469 10929 4503
rect 10877 4451 10929 4469
rect 11791 4639 11843 4651
rect 11791 4605 11799 4639
rect 11833 4605 11843 4639
rect 11791 4571 11843 4605
rect 11791 4537 11799 4571
rect 11833 4537 11843 4571
rect 11791 4503 11843 4537
rect 11791 4469 11799 4503
rect 11833 4469 11843 4503
rect 11791 4451 11843 4469
rect 11873 4451 11915 4651
rect 11945 4639 11997 4651
rect 11945 4605 11955 4639
rect 11989 4605 11997 4639
rect 12605 4639 12657 4651
rect 11945 4571 11997 4605
rect 12605 4605 12613 4639
rect 12647 4605 12657 4639
rect 11945 4537 11955 4571
rect 11989 4537 11997 4571
rect 11945 4503 11997 4537
rect 12605 4571 12657 4605
rect 12605 4537 12613 4571
rect 12647 4537 12657 4571
rect 11945 4469 11955 4503
rect 11989 4469 11997 4503
rect 12605 4503 12657 4537
rect 11945 4451 11997 4469
rect 12140 4471 12202 4486
rect 10446 4403 10508 4437
rect 10446 4369 10462 4403
rect 10496 4369 10508 4403
rect 10446 4335 10508 4369
rect 10446 4301 10462 4335
rect 10496 4301 10508 4335
rect 12140 4437 12152 4471
rect 12186 4437 12202 4471
rect 12140 4403 12202 4437
rect 12140 4369 12152 4403
rect 12186 4369 12202 4403
rect 12140 4335 12202 4369
rect 10446 4286 10508 4301
rect 12140 4301 12152 4335
rect 12186 4301 12202 4335
rect 12140 4286 12202 4301
rect 12232 4471 12298 4486
rect 12232 4437 12248 4471
rect 12282 4437 12298 4471
rect 12232 4403 12298 4437
rect 12232 4369 12248 4403
rect 12282 4369 12298 4403
rect 12232 4335 12298 4369
rect 12232 4301 12248 4335
rect 12282 4301 12298 4335
rect 12232 4286 12298 4301
rect 12328 4471 12390 4486
rect 12328 4437 12344 4471
rect 12378 4437 12390 4471
rect 12605 4469 12613 4503
rect 12647 4469 12657 4503
rect 12605 4451 12657 4469
rect 12687 4451 12729 4651
rect 12759 4639 12811 4651
rect 12759 4605 12769 4639
rect 12803 4605 12811 4639
rect 12759 4571 12811 4605
rect 12759 4537 12769 4571
rect 12803 4537 12811 4571
rect 12759 4503 12811 4537
rect 12759 4469 12769 4503
rect 12803 4469 12811 4503
rect 12759 4451 12811 4469
rect 13679 4639 13731 4651
rect 13679 4605 13687 4639
rect 13721 4605 13731 4639
rect 13679 4571 13731 4605
rect 13679 4537 13687 4571
rect 13721 4537 13731 4571
rect 13679 4503 13731 4537
rect 13679 4469 13687 4503
rect 13721 4469 13731 4503
rect 13679 4451 13731 4469
rect 13761 4451 13803 4651
rect 13833 4639 13885 4651
rect 13833 4605 13843 4639
rect 13877 4605 13885 4639
rect 14493 4639 14545 4651
rect 13833 4571 13885 4605
rect 14493 4605 14501 4639
rect 14535 4605 14545 4639
rect 13833 4537 13843 4571
rect 13877 4537 13885 4571
rect 13833 4503 13885 4537
rect 14493 4571 14545 4605
rect 14493 4537 14501 4571
rect 14535 4537 14545 4571
rect 13833 4469 13843 4503
rect 13877 4469 13885 4503
rect 14493 4503 14545 4537
rect 13833 4451 13885 4469
rect 14028 4471 14090 4486
rect 12328 4403 12390 4437
rect 12328 4369 12344 4403
rect 12378 4369 12390 4403
rect 12328 4335 12390 4369
rect 12328 4301 12344 4335
rect 12378 4301 12390 4335
rect 14028 4437 14040 4471
rect 14074 4437 14090 4471
rect 14028 4403 14090 4437
rect 14028 4369 14040 4403
rect 14074 4369 14090 4403
rect 14028 4335 14090 4369
rect 12328 4286 12390 4301
rect 14028 4301 14040 4335
rect 14074 4301 14090 4335
rect 14028 4286 14090 4301
rect 14120 4471 14186 4486
rect 14120 4437 14136 4471
rect 14170 4437 14186 4471
rect 14120 4403 14186 4437
rect 14120 4369 14136 4403
rect 14170 4369 14186 4403
rect 14120 4335 14186 4369
rect 14120 4301 14136 4335
rect 14170 4301 14186 4335
rect 14120 4286 14186 4301
rect 14216 4471 14278 4486
rect 14216 4437 14232 4471
rect 14266 4437 14278 4471
rect 14493 4469 14501 4503
rect 14535 4469 14545 4503
rect 14493 4451 14545 4469
rect 14575 4451 14617 4651
rect 14647 4639 14699 4651
rect 14647 4605 14657 4639
rect 14691 4605 14699 4639
rect 14647 4571 14699 4605
rect 14647 4537 14657 4571
rect 14691 4537 14699 4571
rect 14647 4503 14699 4537
rect 14647 4469 14657 4503
rect 14691 4469 14699 4503
rect 14647 4451 14699 4469
rect 15567 4639 15619 4651
rect 15567 4605 15575 4639
rect 15609 4605 15619 4639
rect 15567 4571 15619 4605
rect 15567 4537 15575 4571
rect 15609 4537 15619 4571
rect 15567 4503 15619 4537
rect 15567 4469 15575 4503
rect 15609 4469 15619 4503
rect 15567 4451 15619 4469
rect 15649 4451 15691 4651
rect 15721 4639 15773 4651
rect 15721 4605 15731 4639
rect 15765 4605 15773 4639
rect 16381 4639 16433 4651
rect 15721 4571 15773 4605
rect 16381 4605 16389 4639
rect 16423 4605 16433 4639
rect 15721 4537 15731 4571
rect 15765 4537 15773 4571
rect 15721 4503 15773 4537
rect 16381 4571 16433 4605
rect 16381 4537 16389 4571
rect 16423 4537 16433 4571
rect 15721 4469 15731 4503
rect 15765 4469 15773 4503
rect 16381 4503 16433 4537
rect 15721 4451 15773 4469
rect 15916 4471 15978 4486
rect 14216 4403 14278 4437
rect 14216 4369 14232 4403
rect 14266 4369 14278 4403
rect 14216 4335 14278 4369
rect 14216 4301 14232 4335
rect 14266 4301 14278 4335
rect 15916 4437 15928 4471
rect 15962 4437 15978 4471
rect 15916 4403 15978 4437
rect 15916 4369 15928 4403
rect 15962 4369 15978 4403
rect 15916 4335 15978 4369
rect 14216 4286 14278 4301
rect 15916 4301 15928 4335
rect 15962 4301 15978 4335
rect 15916 4286 15978 4301
rect 16008 4471 16074 4486
rect 16008 4437 16024 4471
rect 16058 4437 16074 4471
rect 16008 4403 16074 4437
rect 16008 4369 16024 4403
rect 16058 4369 16074 4403
rect 16008 4335 16074 4369
rect 16008 4301 16024 4335
rect 16058 4301 16074 4335
rect 16008 4286 16074 4301
rect 16104 4471 16166 4486
rect 16104 4437 16120 4471
rect 16154 4437 16166 4471
rect 16381 4469 16389 4503
rect 16423 4469 16433 4503
rect 16381 4451 16433 4469
rect 16463 4451 16505 4651
rect 16535 4639 16587 4651
rect 16535 4605 16545 4639
rect 16579 4605 16587 4639
rect 16535 4571 16587 4605
rect 16535 4537 16545 4571
rect 16579 4537 16587 4571
rect 16535 4503 16587 4537
rect 16535 4469 16545 4503
rect 16579 4469 16587 4503
rect 16535 4451 16587 4469
rect 17455 4639 17507 4651
rect 17455 4605 17463 4639
rect 17497 4605 17507 4639
rect 17455 4571 17507 4605
rect 17455 4537 17463 4571
rect 17497 4537 17507 4571
rect 17455 4503 17507 4537
rect 17455 4469 17463 4503
rect 17497 4469 17507 4503
rect 17455 4451 17507 4469
rect 17537 4451 17579 4651
rect 17609 4639 17661 4651
rect 17609 4605 17619 4639
rect 17653 4605 17661 4639
rect 18269 4639 18321 4651
rect 17609 4571 17661 4605
rect 18269 4605 18277 4639
rect 18311 4605 18321 4639
rect 17609 4537 17619 4571
rect 17653 4537 17661 4571
rect 17609 4503 17661 4537
rect 18269 4571 18321 4605
rect 18269 4537 18277 4571
rect 18311 4537 18321 4571
rect 17609 4469 17619 4503
rect 17653 4469 17661 4503
rect 18269 4503 18321 4537
rect 17609 4451 17661 4469
rect 17804 4471 17866 4486
rect 16104 4403 16166 4437
rect 16104 4369 16120 4403
rect 16154 4369 16166 4403
rect 16104 4335 16166 4369
rect 16104 4301 16120 4335
rect 16154 4301 16166 4335
rect 17804 4437 17816 4471
rect 17850 4437 17866 4471
rect 17804 4403 17866 4437
rect 17804 4369 17816 4403
rect 17850 4369 17866 4403
rect 17804 4335 17866 4369
rect 16104 4286 16166 4301
rect 17804 4301 17816 4335
rect 17850 4301 17866 4335
rect 17804 4286 17866 4301
rect 17896 4471 17962 4486
rect 17896 4437 17912 4471
rect 17946 4437 17962 4471
rect 17896 4403 17962 4437
rect 17896 4369 17912 4403
rect 17946 4369 17962 4403
rect 17896 4335 17962 4369
rect 17896 4301 17912 4335
rect 17946 4301 17962 4335
rect 17896 4286 17962 4301
rect 17992 4471 18054 4486
rect 17992 4437 18008 4471
rect 18042 4437 18054 4471
rect 18269 4469 18277 4503
rect 18311 4469 18321 4503
rect 18269 4451 18321 4469
rect 18351 4451 18393 4651
rect 18423 4639 18475 4651
rect 18423 4605 18433 4639
rect 18467 4605 18475 4639
rect 18423 4571 18475 4605
rect 18423 4537 18433 4571
rect 18467 4537 18475 4571
rect 18423 4503 18475 4537
rect 18423 4469 18433 4503
rect 18467 4469 18475 4503
rect 18423 4451 18475 4469
rect 19343 4639 19395 4651
rect 19343 4605 19351 4639
rect 19385 4605 19395 4639
rect 19343 4571 19395 4605
rect 19343 4537 19351 4571
rect 19385 4537 19395 4571
rect 19343 4503 19395 4537
rect 19343 4469 19351 4503
rect 19385 4469 19395 4503
rect 19343 4451 19395 4469
rect 19425 4451 19467 4651
rect 19497 4639 19549 4651
rect 19497 4605 19507 4639
rect 19541 4605 19549 4639
rect 20157 4639 20209 4651
rect 19497 4571 19549 4605
rect 20157 4605 20165 4639
rect 20199 4605 20209 4639
rect 19497 4537 19507 4571
rect 19541 4537 19549 4571
rect 19497 4503 19549 4537
rect 20157 4571 20209 4605
rect 20157 4537 20165 4571
rect 20199 4537 20209 4571
rect 19497 4469 19507 4503
rect 19541 4469 19549 4503
rect 20157 4503 20209 4537
rect 19497 4451 19549 4469
rect 19692 4471 19754 4486
rect 17992 4403 18054 4437
rect 17992 4369 18008 4403
rect 18042 4369 18054 4403
rect 17992 4335 18054 4369
rect 17992 4301 18008 4335
rect 18042 4301 18054 4335
rect 19692 4437 19704 4471
rect 19738 4437 19754 4471
rect 19692 4403 19754 4437
rect 19692 4369 19704 4403
rect 19738 4369 19754 4403
rect 19692 4335 19754 4369
rect 17992 4286 18054 4301
rect 19692 4301 19704 4335
rect 19738 4301 19754 4335
rect 19692 4286 19754 4301
rect 19784 4471 19850 4486
rect 19784 4437 19800 4471
rect 19834 4437 19850 4471
rect 19784 4403 19850 4437
rect 19784 4369 19800 4403
rect 19834 4369 19850 4403
rect 19784 4335 19850 4369
rect 19784 4301 19800 4335
rect 19834 4301 19850 4335
rect 19784 4286 19850 4301
rect 19880 4471 19942 4486
rect 19880 4437 19896 4471
rect 19930 4437 19942 4471
rect 20157 4469 20165 4503
rect 20199 4469 20209 4503
rect 20157 4451 20209 4469
rect 20239 4451 20281 4651
rect 20311 4639 20363 4651
rect 20311 4605 20321 4639
rect 20355 4605 20363 4639
rect 20311 4571 20363 4605
rect 20311 4537 20321 4571
rect 20355 4537 20363 4571
rect 20311 4503 20363 4537
rect 20311 4469 20321 4503
rect 20355 4469 20363 4503
rect 20311 4451 20363 4469
rect 21231 4639 21283 4651
rect 21231 4605 21239 4639
rect 21273 4605 21283 4639
rect 21231 4571 21283 4605
rect 21231 4537 21239 4571
rect 21273 4537 21283 4571
rect 21231 4503 21283 4537
rect 21231 4469 21239 4503
rect 21273 4469 21283 4503
rect 21231 4451 21283 4469
rect 21313 4451 21355 4651
rect 21385 4639 21437 4651
rect 21385 4605 21395 4639
rect 21429 4605 21437 4639
rect 22045 4639 22097 4651
rect 21385 4571 21437 4605
rect 22045 4605 22053 4639
rect 22087 4605 22097 4639
rect 21385 4537 21395 4571
rect 21429 4537 21437 4571
rect 21385 4503 21437 4537
rect 22045 4571 22097 4605
rect 22045 4537 22053 4571
rect 22087 4537 22097 4571
rect 21385 4469 21395 4503
rect 21429 4469 21437 4503
rect 22045 4503 22097 4537
rect 21385 4451 21437 4469
rect 21580 4471 21642 4486
rect 19880 4403 19942 4437
rect 19880 4369 19896 4403
rect 19930 4369 19942 4403
rect 19880 4335 19942 4369
rect 19880 4301 19896 4335
rect 19930 4301 19942 4335
rect 21580 4437 21592 4471
rect 21626 4437 21642 4471
rect 21580 4403 21642 4437
rect 21580 4369 21592 4403
rect 21626 4369 21642 4403
rect 21580 4335 21642 4369
rect 19880 4286 19942 4301
rect 21580 4301 21592 4335
rect 21626 4301 21642 4335
rect 21580 4286 21642 4301
rect 21672 4471 21738 4486
rect 21672 4437 21688 4471
rect 21722 4437 21738 4471
rect 21672 4403 21738 4437
rect 21672 4369 21688 4403
rect 21722 4369 21738 4403
rect 21672 4335 21738 4369
rect 21672 4301 21688 4335
rect 21722 4301 21738 4335
rect 21672 4286 21738 4301
rect 21768 4471 21830 4486
rect 21768 4437 21784 4471
rect 21818 4437 21830 4471
rect 22045 4469 22053 4503
rect 22087 4469 22097 4503
rect 22045 4451 22097 4469
rect 22127 4451 22169 4651
rect 22199 4639 22251 4651
rect 22199 4605 22209 4639
rect 22243 4605 22251 4639
rect 22199 4571 22251 4605
rect 22199 4537 22209 4571
rect 22243 4537 22251 4571
rect 22199 4503 22251 4537
rect 22199 4469 22209 4503
rect 22243 4469 22251 4503
rect 22199 4451 22251 4469
rect 23119 4639 23171 4651
rect 23119 4605 23127 4639
rect 23161 4605 23171 4639
rect 23119 4571 23171 4605
rect 23119 4537 23127 4571
rect 23161 4537 23171 4571
rect 23119 4503 23171 4537
rect 23119 4469 23127 4503
rect 23161 4469 23171 4503
rect 23119 4451 23171 4469
rect 23201 4451 23243 4651
rect 23273 4639 23325 4651
rect 23273 4605 23283 4639
rect 23317 4605 23325 4639
rect 23933 4639 23985 4651
rect 23273 4571 23325 4605
rect 23933 4605 23941 4639
rect 23975 4605 23985 4639
rect 23273 4537 23283 4571
rect 23317 4537 23325 4571
rect 23273 4503 23325 4537
rect 23933 4571 23985 4605
rect 23933 4537 23941 4571
rect 23975 4537 23985 4571
rect 23273 4469 23283 4503
rect 23317 4469 23325 4503
rect 23933 4503 23985 4537
rect 23273 4451 23325 4469
rect 23468 4471 23530 4486
rect 21768 4403 21830 4437
rect 21768 4369 21784 4403
rect 21818 4369 21830 4403
rect 21768 4335 21830 4369
rect 21768 4301 21784 4335
rect 21818 4301 21830 4335
rect 23468 4437 23480 4471
rect 23514 4437 23530 4471
rect 23468 4403 23530 4437
rect 23468 4369 23480 4403
rect 23514 4369 23530 4403
rect 23468 4335 23530 4369
rect 21768 4286 21830 4301
rect 23468 4301 23480 4335
rect 23514 4301 23530 4335
rect 23468 4286 23530 4301
rect 23560 4471 23626 4486
rect 23560 4437 23576 4471
rect 23610 4437 23626 4471
rect 23560 4403 23626 4437
rect 23560 4369 23576 4403
rect 23610 4369 23626 4403
rect 23560 4335 23626 4369
rect 23560 4301 23576 4335
rect 23610 4301 23626 4335
rect 23560 4286 23626 4301
rect 23656 4471 23718 4486
rect 23656 4437 23672 4471
rect 23706 4437 23718 4471
rect 23933 4469 23941 4503
rect 23975 4469 23985 4503
rect 23933 4451 23985 4469
rect 24015 4451 24057 4651
rect 24087 4639 24139 4651
rect 24087 4605 24097 4639
rect 24131 4605 24139 4639
rect 24087 4571 24139 4605
rect 24087 4537 24097 4571
rect 24131 4537 24139 4571
rect 24087 4503 24139 4537
rect 24087 4469 24097 4503
rect 24131 4469 24139 4503
rect 24087 4451 24139 4469
rect 25007 4639 25059 4651
rect 25007 4605 25015 4639
rect 25049 4605 25059 4639
rect 25007 4571 25059 4605
rect 25007 4537 25015 4571
rect 25049 4537 25059 4571
rect 25007 4503 25059 4537
rect 25007 4469 25015 4503
rect 25049 4469 25059 4503
rect 25007 4451 25059 4469
rect 25089 4451 25131 4651
rect 25161 4639 25213 4651
rect 25161 4605 25171 4639
rect 25205 4605 25213 4639
rect 25821 4639 25873 4651
rect 25161 4571 25213 4605
rect 25821 4605 25829 4639
rect 25863 4605 25873 4639
rect 25161 4537 25171 4571
rect 25205 4537 25213 4571
rect 25161 4503 25213 4537
rect 25821 4571 25873 4605
rect 25821 4537 25829 4571
rect 25863 4537 25873 4571
rect 25161 4469 25171 4503
rect 25205 4469 25213 4503
rect 25821 4503 25873 4537
rect 25161 4451 25213 4469
rect 25356 4471 25418 4486
rect 23656 4403 23718 4437
rect 23656 4369 23672 4403
rect 23706 4369 23718 4403
rect 23656 4335 23718 4369
rect 23656 4301 23672 4335
rect 23706 4301 23718 4335
rect 25356 4437 25368 4471
rect 25402 4437 25418 4471
rect 25356 4403 25418 4437
rect 25356 4369 25368 4403
rect 25402 4369 25418 4403
rect 25356 4335 25418 4369
rect 23656 4286 23718 4301
rect 25356 4301 25368 4335
rect 25402 4301 25418 4335
rect 25356 4286 25418 4301
rect 25448 4471 25514 4486
rect 25448 4437 25464 4471
rect 25498 4437 25514 4471
rect 25448 4403 25514 4437
rect 25448 4369 25464 4403
rect 25498 4369 25514 4403
rect 25448 4335 25514 4369
rect 25448 4301 25464 4335
rect 25498 4301 25514 4335
rect 25448 4286 25514 4301
rect 25544 4471 25606 4486
rect 25544 4437 25560 4471
rect 25594 4437 25606 4471
rect 25821 4469 25829 4503
rect 25863 4469 25873 4503
rect 25821 4451 25873 4469
rect 25903 4451 25945 4651
rect 25975 4639 26027 4651
rect 25975 4605 25985 4639
rect 26019 4605 26027 4639
rect 25975 4571 26027 4605
rect 25975 4537 25985 4571
rect 26019 4537 26027 4571
rect 25975 4503 26027 4537
rect 25975 4469 25985 4503
rect 26019 4469 26027 4503
rect 25975 4451 26027 4469
rect 25544 4403 25606 4437
rect 25544 4369 25560 4403
rect 25594 4369 25606 4403
rect 25544 4335 25606 4369
rect 25544 4301 25560 4335
rect 25594 4301 25606 4335
rect 25544 4286 25606 4301
rect -3444 3585 -3392 3597
rect -3444 3551 -3436 3585
rect -3402 3551 -3392 3585
rect -3444 3517 -3392 3551
rect -3444 3483 -3436 3517
rect -3402 3483 -3392 3517
rect -3444 3449 -3392 3483
rect -3444 3415 -3436 3449
rect -3402 3415 -3392 3449
rect -3444 3397 -3392 3415
rect -3362 3585 -3310 3597
rect -3362 3551 -3352 3585
rect -3318 3551 -3310 3585
rect -3362 3517 -3310 3551
rect -3362 3483 -3352 3517
rect -3318 3483 -3310 3517
rect -3362 3449 -3310 3483
rect -3362 3415 -3352 3449
rect -3318 3415 -3310 3449
rect -3362 3397 -3310 3415
rect -3176 3575 -3118 3590
rect -3176 3541 -3164 3575
rect -3130 3541 -3118 3575
rect -3176 3507 -3118 3541
rect -3176 3473 -3164 3507
rect -3130 3473 -3118 3507
rect -3176 3439 -3118 3473
rect -3176 3405 -3164 3439
rect -3130 3405 -3118 3439
rect -3176 3390 -3118 3405
rect -3088 3575 -3030 3590
rect -3088 3541 -3076 3575
rect -3042 3541 -3030 3575
rect -3088 3507 -3030 3541
rect -2248 3593 -2196 3605
rect -2530 3575 -2472 3590
rect -2530 3541 -2518 3575
rect -2484 3541 -2472 3575
rect -3088 3473 -3076 3507
rect -3042 3473 -3030 3507
rect -3088 3439 -3030 3473
rect -3088 3405 -3076 3439
rect -3042 3405 -3030 3439
rect -2530 3507 -2472 3541
rect -2530 3473 -2518 3507
rect -2484 3473 -2472 3507
rect -2530 3439 -2472 3473
rect -3088 3390 -3030 3405
rect -2960 3415 -2898 3430
rect -2960 3381 -2948 3415
rect -2914 3381 -2898 3415
rect -2960 3347 -2898 3381
rect -2960 3313 -2948 3347
rect -2914 3313 -2898 3347
rect -2960 3279 -2898 3313
rect -2960 3245 -2948 3279
rect -2914 3245 -2898 3279
rect -2960 3230 -2898 3245
rect -2868 3415 -2802 3430
rect -2868 3381 -2852 3415
rect -2818 3381 -2802 3415
rect -2868 3347 -2802 3381
rect -2868 3313 -2852 3347
rect -2818 3313 -2802 3347
rect -2868 3279 -2802 3313
rect -2868 3245 -2852 3279
rect -2818 3245 -2802 3279
rect -2868 3230 -2802 3245
rect -2772 3415 -2710 3430
rect -2772 3381 -2756 3415
rect -2722 3381 -2710 3415
rect -2530 3405 -2518 3439
rect -2484 3405 -2472 3439
rect -2530 3390 -2472 3405
rect -2442 3575 -2384 3590
rect -2442 3541 -2430 3575
rect -2396 3541 -2384 3575
rect -2442 3507 -2384 3541
rect -2442 3473 -2430 3507
rect -2396 3473 -2384 3507
rect -2442 3439 -2384 3473
rect -2442 3405 -2430 3439
rect -2396 3405 -2384 3439
rect -2248 3559 -2240 3593
rect -2206 3559 -2196 3593
rect -2248 3525 -2196 3559
rect -2248 3491 -2240 3525
rect -2206 3491 -2196 3525
rect -2248 3457 -2196 3491
rect -2248 3423 -2240 3457
rect -2206 3423 -2196 3457
rect -2248 3405 -2196 3423
rect -2166 3593 -2114 3605
rect -2166 3559 -2156 3593
rect -2122 3559 -2114 3593
rect -2166 3525 -2114 3559
rect -2166 3491 -2156 3525
rect -2122 3491 -2114 3525
rect -2166 3457 -2114 3491
rect -2166 3423 -2156 3457
rect -2122 3423 -2114 3457
rect -1943 3583 -1891 3603
rect -1943 3549 -1935 3583
rect -1901 3549 -1891 3583
rect -1943 3515 -1891 3549
rect -1943 3481 -1935 3515
rect -1901 3481 -1891 3515
rect -1943 3445 -1891 3481
rect -1861 3583 -1803 3603
rect -1861 3549 -1849 3583
rect -1815 3549 -1803 3583
rect -1861 3515 -1803 3549
rect -1861 3481 -1849 3515
rect -1815 3481 -1803 3515
rect -1861 3445 -1803 3481
rect -1773 3583 -1721 3603
rect -1773 3549 -1763 3583
rect -1729 3549 -1721 3583
rect -1773 3502 -1721 3549
rect -1773 3468 -1763 3502
rect -1729 3468 -1721 3502
rect -1773 3445 -1721 3468
rect -1556 3585 -1504 3597
rect -1556 3551 -1548 3585
rect -1514 3551 -1504 3585
rect -1556 3517 -1504 3551
rect -1556 3483 -1548 3517
rect -1514 3483 -1504 3517
rect -1556 3449 -1504 3483
rect -2166 3405 -2114 3423
rect -2442 3390 -2384 3405
rect -2772 3347 -2710 3381
rect -2772 3313 -2756 3347
rect -2722 3313 -2710 3347
rect -2772 3279 -2710 3313
rect -1556 3415 -1548 3449
rect -1514 3415 -1504 3449
rect -1556 3397 -1504 3415
rect -1474 3585 -1422 3597
rect -1474 3551 -1464 3585
rect -1430 3551 -1422 3585
rect -1474 3517 -1422 3551
rect -1474 3483 -1464 3517
rect -1430 3483 -1422 3517
rect -1474 3449 -1422 3483
rect -1474 3415 -1464 3449
rect -1430 3415 -1422 3449
rect -1474 3397 -1422 3415
rect -1288 3575 -1230 3590
rect -1288 3541 -1276 3575
rect -1242 3541 -1230 3575
rect -1288 3507 -1230 3541
rect -1288 3473 -1276 3507
rect -1242 3473 -1230 3507
rect -1288 3439 -1230 3473
rect -1288 3405 -1276 3439
rect -1242 3405 -1230 3439
rect -1288 3390 -1230 3405
rect -1200 3575 -1142 3590
rect -1200 3541 -1188 3575
rect -1154 3541 -1142 3575
rect -1200 3507 -1142 3541
rect -360 3593 -308 3605
rect -642 3575 -584 3590
rect -642 3541 -630 3575
rect -596 3541 -584 3575
rect -1200 3473 -1188 3507
rect -1154 3473 -1142 3507
rect -1200 3439 -1142 3473
rect -1200 3405 -1188 3439
rect -1154 3405 -1142 3439
rect -642 3507 -584 3541
rect -642 3473 -630 3507
rect -596 3473 -584 3507
rect -642 3439 -584 3473
rect -1200 3390 -1142 3405
rect -1072 3415 -1010 3430
rect -1072 3381 -1060 3415
rect -1026 3381 -1010 3415
rect -2772 3245 -2756 3279
rect -2722 3245 -2710 3279
rect -2772 3230 -2710 3245
rect -1072 3347 -1010 3381
rect -1072 3313 -1060 3347
rect -1026 3313 -1010 3347
rect -1072 3279 -1010 3313
rect -1072 3245 -1060 3279
rect -1026 3245 -1010 3279
rect -1072 3230 -1010 3245
rect -980 3415 -914 3430
rect -980 3381 -964 3415
rect -930 3381 -914 3415
rect -980 3347 -914 3381
rect -980 3313 -964 3347
rect -930 3313 -914 3347
rect -980 3279 -914 3313
rect -980 3245 -964 3279
rect -930 3245 -914 3279
rect -980 3230 -914 3245
rect -884 3415 -822 3430
rect -884 3381 -868 3415
rect -834 3381 -822 3415
rect -642 3405 -630 3439
rect -596 3405 -584 3439
rect -642 3390 -584 3405
rect -554 3575 -496 3590
rect -554 3541 -542 3575
rect -508 3541 -496 3575
rect -554 3507 -496 3541
rect -554 3473 -542 3507
rect -508 3473 -496 3507
rect -554 3439 -496 3473
rect -554 3405 -542 3439
rect -508 3405 -496 3439
rect -360 3559 -352 3593
rect -318 3559 -308 3593
rect -360 3525 -308 3559
rect -360 3491 -352 3525
rect -318 3491 -308 3525
rect -360 3457 -308 3491
rect -360 3423 -352 3457
rect -318 3423 -308 3457
rect -360 3405 -308 3423
rect -278 3593 -226 3605
rect -278 3559 -268 3593
rect -234 3559 -226 3593
rect -278 3525 -226 3559
rect -278 3491 -268 3525
rect -234 3491 -226 3525
rect -278 3457 -226 3491
rect -278 3423 -268 3457
rect -234 3423 -226 3457
rect -55 3583 -3 3603
rect -55 3549 -47 3583
rect -13 3549 -3 3583
rect -55 3515 -3 3549
rect -55 3481 -47 3515
rect -13 3481 -3 3515
rect -55 3445 -3 3481
rect 27 3583 85 3603
rect 27 3549 39 3583
rect 73 3549 85 3583
rect 27 3515 85 3549
rect 27 3481 39 3515
rect 73 3481 85 3515
rect 27 3445 85 3481
rect 115 3583 167 3603
rect 115 3549 125 3583
rect 159 3549 167 3583
rect 115 3502 167 3549
rect 115 3468 125 3502
rect 159 3468 167 3502
rect 115 3445 167 3468
rect 332 3585 384 3597
rect 332 3551 340 3585
rect 374 3551 384 3585
rect 332 3517 384 3551
rect 332 3483 340 3517
rect 374 3483 384 3517
rect 332 3449 384 3483
rect -278 3405 -226 3423
rect -554 3390 -496 3405
rect -884 3347 -822 3381
rect -884 3313 -868 3347
rect -834 3313 -822 3347
rect -884 3279 -822 3313
rect 332 3415 340 3449
rect 374 3415 384 3449
rect 332 3397 384 3415
rect 414 3585 466 3597
rect 414 3551 424 3585
rect 458 3551 466 3585
rect 414 3517 466 3551
rect 414 3483 424 3517
rect 458 3483 466 3517
rect 414 3449 466 3483
rect 414 3415 424 3449
rect 458 3415 466 3449
rect 414 3397 466 3415
rect 600 3575 658 3590
rect 600 3541 612 3575
rect 646 3541 658 3575
rect 600 3507 658 3541
rect 600 3473 612 3507
rect 646 3473 658 3507
rect 600 3439 658 3473
rect 600 3405 612 3439
rect 646 3405 658 3439
rect 600 3390 658 3405
rect 688 3575 746 3590
rect 688 3541 700 3575
rect 734 3541 746 3575
rect 688 3507 746 3541
rect 1528 3593 1580 3605
rect 1246 3575 1304 3590
rect 1246 3541 1258 3575
rect 1292 3541 1304 3575
rect 688 3473 700 3507
rect 734 3473 746 3507
rect 688 3439 746 3473
rect 688 3405 700 3439
rect 734 3405 746 3439
rect 1246 3507 1304 3541
rect 1246 3473 1258 3507
rect 1292 3473 1304 3507
rect 1246 3439 1304 3473
rect 688 3390 746 3405
rect 816 3415 878 3430
rect 816 3381 828 3415
rect 862 3381 878 3415
rect -884 3245 -868 3279
rect -834 3245 -822 3279
rect -884 3230 -822 3245
rect 816 3347 878 3381
rect 816 3313 828 3347
rect 862 3313 878 3347
rect 816 3279 878 3313
rect 816 3245 828 3279
rect 862 3245 878 3279
rect 816 3230 878 3245
rect 908 3415 974 3430
rect 908 3381 924 3415
rect 958 3381 974 3415
rect 908 3347 974 3381
rect 908 3313 924 3347
rect 958 3313 974 3347
rect 908 3279 974 3313
rect 908 3245 924 3279
rect 958 3245 974 3279
rect 908 3230 974 3245
rect 1004 3415 1066 3430
rect 1004 3381 1020 3415
rect 1054 3381 1066 3415
rect 1246 3405 1258 3439
rect 1292 3405 1304 3439
rect 1246 3390 1304 3405
rect 1334 3575 1392 3590
rect 1334 3541 1346 3575
rect 1380 3541 1392 3575
rect 1334 3507 1392 3541
rect 1334 3473 1346 3507
rect 1380 3473 1392 3507
rect 1334 3439 1392 3473
rect 1334 3405 1346 3439
rect 1380 3405 1392 3439
rect 1528 3559 1536 3593
rect 1570 3559 1580 3593
rect 1528 3525 1580 3559
rect 1528 3491 1536 3525
rect 1570 3491 1580 3525
rect 1528 3457 1580 3491
rect 1528 3423 1536 3457
rect 1570 3423 1580 3457
rect 1528 3405 1580 3423
rect 1610 3593 1662 3605
rect 1610 3559 1620 3593
rect 1654 3559 1662 3593
rect 1610 3525 1662 3559
rect 1610 3491 1620 3525
rect 1654 3491 1662 3525
rect 1610 3457 1662 3491
rect 1610 3423 1620 3457
rect 1654 3423 1662 3457
rect 1833 3583 1885 3603
rect 1833 3549 1841 3583
rect 1875 3549 1885 3583
rect 1833 3515 1885 3549
rect 1833 3481 1841 3515
rect 1875 3481 1885 3515
rect 1833 3445 1885 3481
rect 1915 3583 1973 3603
rect 1915 3549 1927 3583
rect 1961 3549 1973 3583
rect 1915 3515 1973 3549
rect 1915 3481 1927 3515
rect 1961 3481 1973 3515
rect 1915 3445 1973 3481
rect 2003 3583 2055 3603
rect 2003 3549 2013 3583
rect 2047 3549 2055 3583
rect 2003 3502 2055 3549
rect 2003 3468 2013 3502
rect 2047 3468 2055 3502
rect 2003 3445 2055 3468
rect 2220 3585 2272 3597
rect 2220 3551 2228 3585
rect 2262 3551 2272 3585
rect 2220 3517 2272 3551
rect 2220 3483 2228 3517
rect 2262 3483 2272 3517
rect 2220 3449 2272 3483
rect 1610 3405 1662 3423
rect 1334 3390 1392 3405
rect 1004 3347 1066 3381
rect 1004 3313 1020 3347
rect 1054 3313 1066 3347
rect 1004 3279 1066 3313
rect 2220 3415 2228 3449
rect 2262 3415 2272 3449
rect 2220 3397 2272 3415
rect 2302 3585 2354 3597
rect 2302 3551 2312 3585
rect 2346 3551 2354 3585
rect 2302 3517 2354 3551
rect 2302 3483 2312 3517
rect 2346 3483 2354 3517
rect 2302 3449 2354 3483
rect 2302 3415 2312 3449
rect 2346 3415 2354 3449
rect 2302 3397 2354 3415
rect 2488 3575 2546 3590
rect 2488 3541 2500 3575
rect 2534 3541 2546 3575
rect 2488 3507 2546 3541
rect 2488 3473 2500 3507
rect 2534 3473 2546 3507
rect 2488 3439 2546 3473
rect 2488 3405 2500 3439
rect 2534 3405 2546 3439
rect 2488 3390 2546 3405
rect 2576 3575 2634 3590
rect 2576 3541 2588 3575
rect 2622 3541 2634 3575
rect 2576 3507 2634 3541
rect 3416 3593 3468 3605
rect 3134 3575 3192 3590
rect 3134 3541 3146 3575
rect 3180 3541 3192 3575
rect 2576 3473 2588 3507
rect 2622 3473 2634 3507
rect 2576 3439 2634 3473
rect 2576 3405 2588 3439
rect 2622 3405 2634 3439
rect 3134 3507 3192 3541
rect 3134 3473 3146 3507
rect 3180 3473 3192 3507
rect 3134 3439 3192 3473
rect 2576 3390 2634 3405
rect 2704 3415 2766 3430
rect 2704 3381 2716 3415
rect 2750 3381 2766 3415
rect 1004 3245 1020 3279
rect 1054 3245 1066 3279
rect 1004 3230 1066 3245
rect 2704 3347 2766 3381
rect 2704 3313 2716 3347
rect 2750 3313 2766 3347
rect 2704 3279 2766 3313
rect 2704 3245 2716 3279
rect 2750 3245 2766 3279
rect 2704 3230 2766 3245
rect 2796 3415 2862 3430
rect 2796 3381 2812 3415
rect 2846 3381 2862 3415
rect 2796 3347 2862 3381
rect 2796 3313 2812 3347
rect 2846 3313 2862 3347
rect 2796 3279 2862 3313
rect 2796 3245 2812 3279
rect 2846 3245 2862 3279
rect 2796 3230 2862 3245
rect 2892 3415 2954 3430
rect 2892 3381 2908 3415
rect 2942 3381 2954 3415
rect 3134 3405 3146 3439
rect 3180 3405 3192 3439
rect 3134 3390 3192 3405
rect 3222 3575 3280 3590
rect 3222 3541 3234 3575
rect 3268 3541 3280 3575
rect 3222 3507 3280 3541
rect 3222 3473 3234 3507
rect 3268 3473 3280 3507
rect 3222 3439 3280 3473
rect 3222 3405 3234 3439
rect 3268 3405 3280 3439
rect 3416 3559 3424 3593
rect 3458 3559 3468 3593
rect 3416 3525 3468 3559
rect 3416 3491 3424 3525
rect 3458 3491 3468 3525
rect 3416 3457 3468 3491
rect 3416 3423 3424 3457
rect 3458 3423 3468 3457
rect 3416 3405 3468 3423
rect 3498 3593 3550 3605
rect 3498 3559 3508 3593
rect 3542 3559 3550 3593
rect 3498 3525 3550 3559
rect 3498 3491 3508 3525
rect 3542 3491 3550 3525
rect 3498 3457 3550 3491
rect 3498 3423 3508 3457
rect 3542 3423 3550 3457
rect 3721 3583 3773 3603
rect 3721 3549 3729 3583
rect 3763 3549 3773 3583
rect 3721 3515 3773 3549
rect 3721 3481 3729 3515
rect 3763 3481 3773 3515
rect 3721 3445 3773 3481
rect 3803 3583 3861 3603
rect 3803 3549 3815 3583
rect 3849 3549 3861 3583
rect 3803 3515 3861 3549
rect 3803 3481 3815 3515
rect 3849 3481 3861 3515
rect 3803 3445 3861 3481
rect 3891 3583 3943 3603
rect 3891 3549 3901 3583
rect 3935 3549 3943 3583
rect 3891 3502 3943 3549
rect 3891 3468 3901 3502
rect 3935 3468 3943 3502
rect 3891 3445 3943 3468
rect 4108 3585 4160 3597
rect 4108 3551 4116 3585
rect 4150 3551 4160 3585
rect 4108 3517 4160 3551
rect 4108 3483 4116 3517
rect 4150 3483 4160 3517
rect 4108 3449 4160 3483
rect 3498 3405 3550 3423
rect 3222 3390 3280 3405
rect 2892 3347 2954 3381
rect 2892 3313 2908 3347
rect 2942 3313 2954 3347
rect 2892 3279 2954 3313
rect 4108 3415 4116 3449
rect 4150 3415 4160 3449
rect 4108 3397 4160 3415
rect 4190 3585 4242 3597
rect 4190 3551 4200 3585
rect 4234 3551 4242 3585
rect 4190 3517 4242 3551
rect 4190 3483 4200 3517
rect 4234 3483 4242 3517
rect 4190 3449 4242 3483
rect 4190 3415 4200 3449
rect 4234 3415 4242 3449
rect 4190 3397 4242 3415
rect 4376 3575 4434 3590
rect 4376 3541 4388 3575
rect 4422 3541 4434 3575
rect 4376 3507 4434 3541
rect 4376 3473 4388 3507
rect 4422 3473 4434 3507
rect 4376 3439 4434 3473
rect 4376 3405 4388 3439
rect 4422 3405 4434 3439
rect 4376 3390 4434 3405
rect 4464 3575 4522 3590
rect 4464 3541 4476 3575
rect 4510 3541 4522 3575
rect 4464 3507 4522 3541
rect 5304 3593 5356 3605
rect 5022 3575 5080 3590
rect 5022 3541 5034 3575
rect 5068 3541 5080 3575
rect 4464 3473 4476 3507
rect 4510 3473 4522 3507
rect 4464 3439 4522 3473
rect 4464 3405 4476 3439
rect 4510 3405 4522 3439
rect 5022 3507 5080 3541
rect 5022 3473 5034 3507
rect 5068 3473 5080 3507
rect 5022 3439 5080 3473
rect 4464 3390 4522 3405
rect 4592 3415 4654 3430
rect 4592 3381 4604 3415
rect 4638 3381 4654 3415
rect 2892 3245 2908 3279
rect 2942 3245 2954 3279
rect 2892 3230 2954 3245
rect 4592 3347 4654 3381
rect 4592 3313 4604 3347
rect 4638 3313 4654 3347
rect 4592 3279 4654 3313
rect 4592 3245 4604 3279
rect 4638 3245 4654 3279
rect 4592 3230 4654 3245
rect 4684 3415 4750 3430
rect 4684 3381 4700 3415
rect 4734 3381 4750 3415
rect 4684 3347 4750 3381
rect 4684 3313 4700 3347
rect 4734 3313 4750 3347
rect 4684 3279 4750 3313
rect 4684 3245 4700 3279
rect 4734 3245 4750 3279
rect 4684 3230 4750 3245
rect 4780 3415 4842 3430
rect 4780 3381 4796 3415
rect 4830 3381 4842 3415
rect 5022 3405 5034 3439
rect 5068 3405 5080 3439
rect 5022 3390 5080 3405
rect 5110 3575 5168 3590
rect 5110 3541 5122 3575
rect 5156 3541 5168 3575
rect 5110 3507 5168 3541
rect 5110 3473 5122 3507
rect 5156 3473 5168 3507
rect 5110 3439 5168 3473
rect 5110 3405 5122 3439
rect 5156 3405 5168 3439
rect 5304 3559 5312 3593
rect 5346 3559 5356 3593
rect 5304 3525 5356 3559
rect 5304 3491 5312 3525
rect 5346 3491 5356 3525
rect 5304 3457 5356 3491
rect 5304 3423 5312 3457
rect 5346 3423 5356 3457
rect 5304 3405 5356 3423
rect 5386 3593 5438 3605
rect 5386 3559 5396 3593
rect 5430 3559 5438 3593
rect 5386 3525 5438 3559
rect 5386 3491 5396 3525
rect 5430 3491 5438 3525
rect 5386 3457 5438 3491
rect 5386 3423 5396 3457
rect 5430 3423 5438 3457
rect 5609 3583 5661 3603
rect 5609 3549 5617 3583
rect 5651 3549 5661 3583
rect 5609 3515 5661 3549
rect 5609 3481 5617 3515
rect 5651 3481 5661 3515
rect 5609 3445 5661 3481
rect 5691 3583 5749 3603
rect 5691 3549 5703 3583
rect 5737 3549 5749 3583
rect 5691 3515 5749 3549
rect 5691 3481 5703 3515
rect 5737 3481 5749 3515
rect 5691 3445 5749 3481
rect 5779 3583 5831 3603
rect 5779 3549 5789 3583
rect 5823 3549 5831 3583
rect 5779 3502 5831 3549
rect 5779 3468 5789 3502
rect 5823 3468 5831 3502
rect 5779 3445 5831 3468
rect 5996 3585 6048 3597
rect 5996 3551 6004 3585
rect 6038 3551 6048 3585
rect 5996 3517 6048 3551
rect 5996 3483 6004 3517
rect 6038 3483 6048 3517
rect 5996 3449 6048 3483
rect 5386 3405 5438 3423
rect 5110 3390 5168 3405
rect 4780 3347 4842 3381
rect 4780 3313 4796 3347
rect 4830 3313 4842 3347
rect 4780 3279 4842 3313
rect 5996 3415 6004 3449
rect 6038 3415 6048 3449
rect 5996 3397 6048 3415
rect 6078 3585 6130 3597
rect 6078 3551 6088 3585
rect 6122 3551 6130 3585
rect 6078 3517 6130 3551
rect 6078 3483 6088 3517
rect 6122 3483 6130 3517
rect 6078 3449 6130 3483
rect 6078 3415 6088 3449
rect 6122 3415 6130 3449
rect 6078 3397 6130 3415
rect 6264 3575 6322 3590
rect 6264 3541 6276 3575
rect 6310 3541 6322 3575
rect 6264 3507 6322 3541
rect 6264 3473 6276 3507
rect 6310 3473 6322 3507
rect 6264 3439 6322 3473
rect 6264 3405 6276 3439
rect 6310 3405 6322 3439
rect 6264 3390 6322 3405
rect 6352 3575 6410 3590
rect 6352 3541 6364 3575
rect 6398 3541 6410 3575
rect 6352 3507 6410 3541
rect 7192 3593 7244 3605
rect 6910 3575 6968 3590
rect 6910 3541 6922 3575
rect 6956 3541 6968 3575
rect 6352 3473 6364 3507
rect 6398 3473 6410 3507
rect 6352 3439 6410 3473
rect 6352 3405 6364 3439
rect 6398 3405 6410 3439
rect 6910 3507 6968 3541
rect 6910 3473 6922 3507
rect 6956 3473 6968 3507
rect 6910 3439 6968 3473
rect 6352 3390 6410 3405
rect 6480 3415 6542 3430
rect 6480 3381 6492 3415
rect 6526 3381 6542 3415
rect 4780 3245 4796 3279
rect 4830 3245 4842 3279
rect 4780 3230 4842 3245
rect 6480 3347 6542 3381
rect 6480 3313 6492 3347
rect 6526 3313 6542 3347
rect 6480 3279 6542 3313
rect 6480 3245 6492 3279
rect 6526 3245 6542 3279
rect 6480 3230 6542 3245
rect 6572 3415 6638 3430
rect 6572 3381 6588 3415
rect 6622 3381 6638 3415
rect 6572 3347 6638 3381
rect 6572 3313 6588 3347
rect 6622 3313 6638 3347
rect 6572 3279 6638 3313
rect 6572 3245 6588 3279
rect 6622 3245 6638 3279
rect 6572 3230 6638 3245
rect 6668 3415 6730 3430
rect 6668 3381 6684 3415
rect 6718 3381 6730 3415
rect 6910 3405 6922 3439
rect 6956 3405 6968 3439
rect 6910 3390 6968 3405
rect 6998 3575 7056 3590
rect 6998 3541 7010 3575
rect 7044 3541 7056 3575
rect 6998 3507 7056 3541
rect 6998 3473 7010 3507
rect 7044 3473 7056 3507
rect 6998 3439 7056 3473
rect 6998 3405 7010 3439
rect 7044 3405 7056 3439
rect 7192 3559 7200 3593
rect 7234 3559 7244 3593
rect 7192 3525 7244 3559
rect 7192 3491 7200 3525
rect 7234 3491 7244 3525
rect 7192 3457 7244 3491
rect 7192 3423 7200 3457
rect 7234 3423 7244 3457
rect 7192 3405 7244 3423
rect 7274 3593 7326 3605
rect 7274 3559 7284 3593
rect 7318 3559 7326 3593
rect 7274 3525 7326 3559
rect 7274 3491 7284 3525
rect 7318 3491 7326 3525
rect 7274 3457 7326 3491
rect 7274 3423 7284 3457
rect 7318 3423 7326 3457
rect 7497 3583 7549 3603
rect 7497 3549 7505 3583
rect 7539 3549 7549 3583
rect 7497 3515 7549 3549
rect 7497 3481 7505 3515
rect 7539 3481 7549 3515
rect 7497 3445 7549 3481
rect 7579 3583 7637 3603
rect 7579 3549 7591 3583
rect 7625 3549 7637 3583
rect 7579 3515 7637 3549
rect 7579 3481 7591 3515
rect 7625 3481 7637 3515
rect 7579 3445 7637 3481
rect 7667 3583 7719 3603
rect 7667 3549 7677 3583
rect 7711 3549 7719 3583
rect 7667 3502 7719 3549
rect 7667 3468 7677 3502
rect 7711 3468 7719 3502
rect 7667 3445 7719 3468
rect 7884 3585 7936 3597
rect 7884 3551 7892 3585
rect 7926 3551 7936 3585
rect 7884 3517 7936 3551
rect 7884 3483 7892 3517
rect 7926 3483 7936 3517
rect 7884 3449 7936 3483
rect 7274 3405 7326 3423
rect 6998 3390 7056 3405
rect 6668 3347 6730 3381
rect 6668 3313 6684 3347
rect 6718 3313 6730 3347
rect 6668 3279 6730 3313
rect 7884 3415 7892 3449
rect 7926 3415 7936 3449
rect 7884 3397 7936 3415
rect 7966 3585 8018 3597
rect 7966 3551 7976 3585
rect 8010 3551 8018 3585
rect 7966 3517 8018 3551
rect 7966 3483 7976 3517
rect 8010 3483 8018 3517
rect 7966 3449 8018 3483
rect 7966 3415 7976 3449
rect 8010 3415 8018 3449
rect 7966 3397 8018 3415
rect 8152 3575 8210 3590
rect 8152 3541 8164 3575
rect 8198 3541 8210 3575
rect 8152 3507 8210 3541
rect 8152 3473 8164 3507
rect 8198 3473 8210 3507
rect 8152 3439 8210 3473
rect 8152 3405 8164 3439
rect 8198 3405 8210 3439
rect 8152 3390 8210 3405
rect 8240 3575 8298 3590
rect 8240 3541 8252 3575
rect 8286 3541 8298 3575
rect 8240 3507 8298 3541
rect 9080 3593 9132 3605
rect 8798 3575 8856 3590
rect 8798 3541 8810 3575
rect 8844 3541 8856 3575
rect 8240 3473 8252 3507
rect 8286 3473 8298 3507
rect 8240 3439 8298 3473
rect 8240 3405 8252 3439
rect 8286 3405 8298 3439
rect 8798 3507 8856 3541
rect 8798 3473 8810 3507
rect 8844 3473 8856 3507
rect 8798 3439 8856 3473
rect 8240 3390 8298 3405
rect 8368 3415 8430 3430
rect 8368 3381 8380 3415
rect 8414 3381 8430 3415
rect 6668 3245 6684 3279
rect 6718 3245 6730 3279
rect 6668 3230 6730 3245
rect 8368 3347 8430 3381
rect 8368 3313 8380 3347
rect 8414 3313 8430 3347
rect 8368 3279 8430 3313
rect 8368 3245 8380 3279
rect 8414 3245 8430 3279
rect 8368 3230 8430 3245
rect 8460 3415 8526 3430
rect 8460 3381 8476 3415
rect 8510 3381 8526 3415
rect 8460 3347 8526 3381
rect 8460 3313 8476 3347
rect 8510 3313 8526 3347
rect 8460 3279 8526 3313
rect 8460 3245 8476 3279
rect 8510 3245 8526 3279
rect 8460 3230 8526 3245
rect 8556 3415 8618 3430
rect 8556 3381 8572 3415
rect 8606 3381 8618 3415
rect 8798 3405 8810 3439
rect 8844 3405 8856 3439
rect 8798 3390 8856 3405
rect 8886 3575 8944 3590
rect 8886 3541 8898 3575
rect 8932 3541 8944 3575
rect 8886 3507 8944 3541
rect 8886 3473 8898 3507
rect 8932 3473 8944 3507
rect 8886 3439 8944 3473
rect 8886 3405 8898 3439
rect 8932 3405 8944 3439
rect 9080 3559 9088 3593
rect 9122 3559 9132 3593
rect 9080 3525 9132 3559
rect 9080 3491 9088 3525
rect 9122 3491 9132 3525
rect 9080 3457 9132 3491
rect 9080 3423 9088 3457
rect 9122 3423 9132 3457
rect 9080 3405 9132 3423
rect 9162 3593 9214 3605
rect 9162 3559 9172 3593
rect 9206 3559 9214 3593
rect 9162 3525 9214 3559
rect 9162 3491 9172 3525
rect 9206 3491 9214 3525
rect 9162 3457 9214 3491
rect 9162 3423 9172 3457
rect 9206 3423 9214 3457
rect 9385 3583 9437 3603
rect 9385 3549 9393 3583
rect 9427 3549 9437 3583
rect 9385 3515 9437 3549
rect 9385 3481 9393 3515
rect 9427 3481 9437 3515
rect 9385 3445 9437 3481
rect 9467 3583 9525 3603
rect 9467 3549 9479 3583
rect 9513 3549 9525 3583
rect 9467 3515 9525 3549
rect 9467 3481 9479 3515
rect 9513 3481 9525 3515
rect 9467 3445 9525 3481
rect 9555 3583 9607 3603
rect 9555 3549 9565 3583
rect 9599 3549 9607 3583
rect 9555 3502 9607 3549
rect 9555 3468 9565 3502
rect 9599 3468 9607 3502
rect 9555 3445 9607 3468
rect 9772 3585 9824 3597
rect 9772 3551 9780 3585
rect 9814 3551 9824 3585
rect 9772 3517 9824 3551
rect 9772 3483 9780 3517
rect 9814 3483 9824 3517
rect 9772 3449 9824 3483
rect 9162 3405 9214 3423
rect 8886 3390 8944 3405
rect 8556 3347 8618 3381
rect 8556 3313 8572 3347
rect 8606 3313 8618 3347
rect 8556 3279 8618 3313
rect 9772 3415 9780 3449
rect 9814 3415 9824 3449
rect 9772 3397 9824 3415
rect 9854 3585 9906 3597
rect 9854 3551 9864 3585
rect 9898 3551 9906 3585
rect 9854 3517 9906 3551
rect 9854 3483 9864 3517
rect 9898 3483 9906 3517
rect 9854 3449 9906 3483
rect 9854 3415 9864 3449
rect 9898 3415 9906 3449
rect 9854 3397 9906 3415
rect 10040 3575 10098 3590
rect 10040 3541 10052 3575
rect 10086 3541 10098 3575
rect 10040 3507 10098 3541
rect 10040 3473 10052 3507
rect 10086 3473 10098 3507
rect 10040 3439 10098 3473
rect 10040 3405 10052 3439
rect 10086 3405 10098 3439
rect 10040 3390 10098 3405
rect 10128 3575 10186 3590
rect 10128 3541 10140 3575
rect 10174 3541 10186 3575
rect 10128 3507 10186 3541
rect 10968 3593 11020 3605
rect 10686 3575 10744 3590
rect 10686 3541 10698 3575
rect 10732 3541 10744 3575
rect 10128 3473 10140 3507
rect 10174 3473 10186 3507
rect 10128 3439 10186 3473
rect 10128 3405 10140 3439
rect 10174 3405 10186 3439
rect 10686 3507 10744 3541
rect 10686 3473 10698 3507
rect 10732 3473 10744 3507
rect 10686 3439 10744 3473
rect 10128 3390 10186 3405
rect 10256 3415 10318 3430
rect 10256 3381 10268 3415
rect 10302 3381 10318 3415
rect 8556 3245 8572 3279
rect 8606 3245 8618 3279
rect 8556 3230 8618 3245
rect 10256 3347 10318 3381
rect 10256 3313 10268 3347
rect 10302 3313 10318 3347
rect 10256 3279 10318 3313
rect 10256 3245 10268 3279
rect 10302 3245 10318 3279
rect 10256 3230 10318 3245
rect 10348 3415 10414 3430
rect 10348 3381 10364 3415
rect 10398 3381 10414 3415
rect 10348 3347 10414 3381
rect 10348 3313 10364 3347
rect 10398 3313 10414 3347
rect 10348 3279 10414 3313
rect 10348 3245 10364 3279
rect 10398 3245 10414 3279
rect 10348 3230 10414 3245
rect 10444 3415 10506 3430
rect 10444 3381 10460 3415
rect 10494 3381 10506 3415
rect 10686 3405 10698 3439
rect 10732 3405 10744 3439
rect 10686 3390 10744 3405
rect 10774 3575 10832 3590
rect 10774 3541 10786 3575
rect 10820 3541 10832 3575
rect 10774 3507 10832 3541
rect 10774 3473 10786 3507
rect 10820 3473 10832 3507
rect 10774 3439 10832 3473
rect 10774 3405 10786 3439
rect 10820 3405 10832 3439
rect 10968 3559 10976 3593
rect 11010 3559 11020 3593
rect 10968 3525 11020 3559
rect 10968 3491 10976 3525
rect 11010 3491 11020 3525
rect 10968 3457 11020 3491
rect 10968 3423 10976 3457
rect 11010 3423 11020 3457
rect 10968 3405 11020 3423
rect 11050 3593 11102 3605
rect 11050 3559 11060 3593
rect 11094 3559 11102 3593
rect 11050 3525 11102 3559
rect 11050 3491 11060 3525
rect 11094 3491 11102 3525
rect 11050 3457 11102 3491
rect 11050 3423 11060 3457
rect 11094 3423 11102 3457
rect 11273 3583 11325 3603
rect 11273 3549 11281 3583
rect 11315 3549 11325 3583
rect 11273 3515 11325 3549
rect 11273 3481 11281 3515
rect 11315 3481 11325 3515
rect 11273 3445 11325 3481
rect 11355 3583 11413 3603
rect 11355 3549 11367 3583
rect 11401 3549 11413 3583
rect 11355 3515 11413 3549
rect 11355 3481 11367 3515
rect 11401 3481 11413 3515
rect 11355 3445 11413 3481
rect 11443 3583 11495 3603
rect 11443 3549 11453 3583
rect 11487 3549 11495 3583
rect 11443 3502 11495 3549
rect 11443 3468 11453 3502
rect 11487 3468 11495 3502
rect 11443 3445 11495 3468
rect 11654 3585 11706 3597
rect 11654 3551 11662 3585
rect 11696 3551 11706 3585
rect 11654 3517 11706 3551
rect 11654 3483 11662 3517
rect 11696 3483 11706 3517
rect 11654 3449 11706 3483
rect 11050 3405 11102 3423
rect 10774 3390 10832 3405
rect 10444 3347 10506 3381
rect 10444 3313 10460 3347
rect 10494 3313 10506 3347
rect 10444 3279 10506 3313
rect 11654 3415 11662 3449
rect 11696 3415 11706 3449
rect 11654 3397 11706 3415
rect 11736 3585 11788 3597
rect 11736 3551 11746 3585
rect 11780 3551 11788 3585
rect 11736 3517 11788 3551
rect 11736 3483 11746 3517
rect 11780 3483 11788 3517
rect 11736 3449 11788 3483
rect 11736 3415 11746 3449
rect 11780 3415 11788 3449
rect 11736 3397 11788 3415
rect 11922 3575 11980 3590
rect 11922 3541 11934 3575
rect 11968 3541 11980 3575
rect 11922 3507 11980 3541
rect 11922 3473 11934 3507
rect 11968 3473 11980 3507
rect 11922 3439 11980 3473
rect 11922 3405 11934 3439
rect 11968 3405 11980 3439
rect 11922 3390 11980 3405
rect 12010 3575 12068 3590
rect 12010 3541 12022 3575
rect 12056 3541 12068 3575
rect 12010 3507 12068 3541
rect 12850 3593 12902 3605
rect 12568 3575 12626 3590
rect 12568 3541 12580 3575
rect 12614 3541 12626 3575
rect 12010 3473 12022 3507
rect 12056 3473 12068 3507
rect 12010 3439 12068 3473
rect 12010 3405 12022 3439
rect 12056 3405 12068 3439
rect 12568 3507 12626 3541
rect 12568 3473 12580 3507
rect 12614 3473 12626 3507
rect 12568 3439 12626 3473
rect 12010 3390 12068 3405
rect 12138 3415 12200 3430
rect 12138 3381 12150 3415
rect 12184 3381 12200 3415
rect 10444 3245 10460 3279
rect 10494 3245 10506 3279
rect 10444 3230 10506 3245
rect 12138 3347 12200 3381
rect 12138 3313 12150 3347
rect 12184 3313 12200 3347
rect 12138 3279 12200 3313
rect 12138 3245 12150 3279
rect 12184 3245 12200 3279
rect 12138 3230 12200 3245
rect 12230 3415 12296 3430
rect 12230 3381 12246 3415
rect 12280 3381 12296 3415
rect 12230 3347 12296 3381
rect 12230 3313 12246 3347
rect 12280 3313 12296 3347
rect 12230 3279 12296 3313
rect 12230 3245 12246 3279
rect 12280 3245 12296 3279
rect 12230 3230 12296 3245
rect 12326 3415 12388 3430
rect 12326 3381 12342 3415
rect 12376 3381 12388 3415
rect 12568 3405 12580 3439
rect 12614 3405 12626 3439
rect 12568 3390 12626 3405
rect 12656 3575 12714 3590
rect 12656 3541 12668 3575
rect 12702 3541 12714 3575
rect 12656 3507 12714 3541
rect 12656 3473 12668 3507
rect 12702 3473 12714 3507
rect 12656 3439 12714 3473
rect 12656 3405 12668 3439
rect 12702 3405 12714 3439
rect 12850 3559 12858 3593
rect 12892 3559 12902 3593
rect 12850 3525 12902 3559
rect 12850 3491 12858 3525
rect 12892 3491 12902 3525
rect 12850 3457 12902 3491
rect 12850 3423 12858 3457
rect 12892 3423 12902 3457
rect 12850 3405 12902 3423
rect 12932 3593 12984 3605
rect 12932 3559 12942 3593
rect 12976 3559 12984 3593
rect 12932 3525 12984 3559
rect 12932 3491 12942 3525
rect 12976 3491 12984 3525
rect 12932 3457 12984 3491
rect 12932 3423 12942 3457
rect 12976 3423 12984 3457
rect 13155 3583 13207 3603
rect 13155 3549 13163 3583
rect 13197 3549 13207 3583
rect 13155 3515 13207 3549
rect 13155 3481 13163 3515
rect 13197 3481 13207 3515
rect 13155 3445 13207 3481
rect 13237 3583 13295 3603
rect 13237 3549 13249 3583
rect 13283 3549 13295 3583
rect 13237 3515 13295 3549
rect 13237 3481 13249 3515
rect 13283 3481 13295 3515
rect 13237 3445 13295 3481
rect 13325 3583 13377 3603
rect 13325 3549 13335 3583
rect 13369 3549 13377 3583
rect 13325 3502 13377 3549
rect 13325 3468 13335 3502
rect 13369 3468 13377 3502
rect 13325 3445 13377 3468
rect 13542 3585 13594 3597
rect 13542 3551 13550 3585
rect 13584 3551 13594 3585
rect 13542 3517 13594 3551
rect 13542 3483 13550 3517
rect 13584 3483 13594 3517
rect 13542 3449 13594 3483
rect 12932 3405 12984 3423
rect 12656 3390 12714 3405
rect 12326 3347 12388 3381
rect 12326 3313 12342 3347
rect 12376 3313 12388 3347
rect 12326 3279 12388 3313
rect 13542 3415 13550 3449
rect 13584 3415 13594 3449
rect 13542 3397 13594 3415
rect 13624 3585 13676 3597
rect 13624 3551 13634 3585
rect 13668 3551 13676 3585
rect 13624 3517 13676 3551
rect 13624 3483 13634 3517
rect 13668 3483 13676 3517
rect 13624 3449 13676 3483
rect 13624 3415 13634 3449
rect 13668 3415 13676 3449
rect 13624 3397 13676 3415
rect 13810 3575 13868 3590
rect 13810 3541 13822 3575
rect 13856 3541 13868 3575
rect 13810 3507 13868 3541
rect 13810 3473 13822 3507
rect 13856 3473 13868 3507
rect 13810 3439 13868 3473
rect 13810 3405 13822 3439
rect 13856 3405 13868 3439
rect 13810 3390 13868 3405
rect 13898 3575 13956 3590
rect 13898 3541 13910 3575
rect 13944 3541 13956 3575
rect 13898 3507 13956 3541
rect 14738 3593 14790 3605
rect 14456 3575 14514 3590
rect 14456 3541 14468 3575
rect 14502 3541 14514 3575
rect 13898 3473 13910 3507
rect 13944 3473 13956 3507
rect 13898 3439 13956 3473
rect 13898 3405 13910 3439
rect 13944 3405 13956 3439
rect 14456 3507 14514 3541
rect 14456 3473 14468 3507
rect 14502 3473 14514 3507
rect 14456 3439 14514 3473
rect 13898 3390 13956 3405
rect 14026 3415 14088 3430
rect 14026 3381 14038 3415
rect 14072 3381 14088 3415
rect 12326 3245 12342 3279
rect 12376 3245 12388 3279
rect 12326 3230 12388 3245
rect 14026 3347 14088 3381
rect 14026 3313 14038 3347
rect 14072 3313 14088 3347
rect 14026 3279 14088 3313
rect 14026 3245 14038 3279
rect 14072 3245 14088 3279
rect 14026 3230 14088 3245
rect 14118 3415 14184 3430
rect 14118 3381 14134 3415
rect 14168 3381 14184 3415
rect 14118 3347 14184 3381
rect 14118 3313 14134 3347
rect 14168 3313 14184 3347
rect 14118 3279 14184 3313
rect 14118 3245 14134 3279
rect 14168 3245 14184 3279
rect 14118 3230 14184 3245
rect 14214 3415 14276 3430
rect 14214 3381 14230 3415
rect 14264 3381 14276 3415
rect 14456 3405 14468 3439
rect 14502 3405 14514 3439
rect 14456 3390 14514 3405
rect 14544 3575 14602 3590
rect 14544 3541 14556 3575
rect 14590 3541 14602 3575
rect 14544 3507 14602 3541
rect 14544 3473 14556 3507
rect 14590 3473 14602 3507
rect 14544 3439 14602 3473
rect 14544 3405 14556 3439
rect 14590 3405 14602 3439
rect 14738 3559 14746 3593
rect 14780 3559 14790 3593
rect 14738 3525 14790 3559
rect 14738 3491 14746 3525
rect 14780 3491 14790 3525
rect 14738 3457 14790 3491
rect 14738 3423 14746 3457
rect 14780 3423 14790 3457
rect 14738 3405 14790 3423
rect 14820 3593 14872 3605
rect 14820 3559 14830 3593
rect 14864 3559 14872 3593
rect 14820 3525 14872 3559
rect 14820 3491 14830 3525
rect 14864 3491 14872 3525
rect 14820 3457 14872 3491
rect 14820 3423 14830 3457
rect 14864 3423 14872 3457
rect 15043 3583 15095 3603
rect 15043 3549 15051 3583
rect 15085 3549 15095 3583
rect 15043 3515 15095 3549
rect 15043 3481 15051 3515
rect 15085 3481 15095 3515
rect 15043 3445 15095 3481
rect 15125 3583 15183 3603
rect 15125 3549 15137 3583
rect 15171 3549 15183 3583
rect 15125 3515 15183 3549
rect 15125 3481 15137 3515
rect 15171 3481 15183 3515
rect 15125 3445 15183 3481
rect 15213 3583 15265 3603
rect 15213 3549 15223 3583
rect 15257 3549 15265 3583
rect 15213 3502 15265 3549
rect 15213 3468 15223 3502
rect 15257 3468 15265 3502
rect 15213 3445 15265 3468
rect 15430 3585 15482 3597
rect 15430 3551 15438 3585
rect 15472 3551 15482 3585
rect 15430 3517 15482 3551
rect 15430 3483 15438 3517
rect 15472 3483 15482 3517
rect 15430 3449 15482 3483
rect 14820 3405 14872 3423
rect 14544 3390 14602 3405
rect 14214 3347 14276 3381
rect 14214 3313 14230 3347
rect 14264 3313 14276 3347
rect 14214 3279 14276 3313
rect 15430 3415 15438 3449
rect 15472 3415 15482 3449
rect 15430 3397 15482 3415
rect 15512 3585 15564 3597
rect 15512 3551 15522 3585
rect 15556 3551 15564 3585
rect 15512 3517 15564 3551
rect 15512 3483 15522 3517
rect 15556 3483 15564 3517
rect 15512 3449 15564 3483
rect 15512 3415 15522 3449
rect 15556 3415 15564 3449
rect 15512 3397 15564 3415
rect 15698 3575 15756 3590
rect 15698 3541 15710 3575
rect 15744 3541 15756 3575
rect 15698 3507 15756 3541
rect 15698 3473 15710 3507
rect 15744 3473 15756 3507
rect 15698 3439 15756 3473
rect 15698 3405 15710 3439
rect 15744 3405 15756 3439
rect 15698 3390 15756 3405
rect 15786 3575 15844 3590
rect 15786 3541 15798 3575
rect 15832 3541 15844 3575
rect 15786 3507 15844 3541
rect 16626 3593 16678 3605
rect 16344 3575 16402 3590
rect 16344 3541 16356 3575
rect 16390 3541 16402 3575
rect 15786 3473 15798 3507
rect 15832 3473 15844 3507
rect 15786 3439 15844 3473
rect 15786 3405 15798 3439
rect 15832 3405 15844 3439
rect 16344 3507 16402 3541
rect 16344 3473 16356 3507
rect 16390 3473 16402 3507
rect 16344 3439 16402 3473
rect 15786 3390 15844 3405
rect 15914 3415 15976 3430
rect 15914 3381 15926 3415
rect 15960 3381 15976 3415
rect 14214 3245 14230 3279
rect 14264 3245 14276 3279
rect 14214 3230 14276 3245
rect 15914 3347 15976 3381
rect 15914 3313 15926 3347
rect 15960 3313 15976 3347
rect 15914 3279 15976 3313
rect 15914 3245 15926 3279
rect 15960 3245 15976 3279
rect 15914 3230 15976 3245
rect 16006 3415 16072 3430
rect 16006 3381 16022 3415
rect 16056 3381 16072 3415
rect 16006 3347 16072 3381
rect 16006 3313 16022 3347
rect 16056 3313 16072 3347
rect 16006 3279 16072 3313
rect 16006 3245 16022 3279
rect 16056 3245 16072 3279
rect 16006 3230 16072 3245
rect 16102 3415 16164 3430
rect 16102 3381 16118 3415
rect 16152 3381 16164 3415
rect 16344 3405 16356 3439
rect 16390 3405 16402 3439
rect 16344 3390 16402 3405
rect 16432 3575 16490 3590
rect 16432 3541 16444 3575
rect 16478 3541 16490 3575
rect 16432 3507 16490 3541
rect 16432 3473 16444 3507
rect 16478 3473 16490 3507
rect 16432 3439 16490 3473
rect 16432 3405 16444 3439
rect 16478 3405 16490 3439
rect 16626 3559 16634 3593
rect 16668 3559 16678 3593
rect 16626 3525 16678 3559
rect 16626 3491 16634 3525
rect 16668 3491 16678 3525
rect 16626 3457 16678 3491
rect 16626 3423 16634 3457
rect 16668 3423 16678 3457
rect 16626 3405 16678 3423
rect 16708 3593 16760 3605
rect 16708 3559 16718 3593
rect 16752 3559 16760 3593
rect 16708 3525 16760 3559
rect 16708 3491 16718 3525
rect 16752 3491 16760 3525
rect 16708 3457 16760 3491
rect 16708 3423 16718 3457
rect 16752 3423 16760 3457
rect 16931 3583 16983 3603
rect 16931 3549 16939 3583
rect 16973 3549 16983 3583
rect 16931 3515 16983 3549
rect 16931 3481 16939 3515
rect 16973 3481 16983 3515
rect 16931 3445 16983 3481
rect 17013 3583 17071 3603
rect 17013 3549 17025 3583
rect 17059 3549 17071 3583
rect 17013 3515 17071 3549
rect 17013 3481 17025 3515
rect 17059 3481 17071 3515
rect 17013 3445 17071 3481
rect 17101 3583 17153 3603
rect 17101 3549 17111 3583
rect 17145 3549 17153 3583
rect 17101 3502 17153 3549
rect 17101 3468 17111 3502
rect 17145 3468 17153 3502
rect 17101 3445 17153 3468
rect 17318 3585 17370 3597
rect 17318 3551 17326 3585
rect 17360 3551 17370 3585
rect 17318 3517 17370 3551
rect 17318 3483 17326 3517
rect 17360 3483 17370 3517
rect 17318 3449 17370 3483
rect 16708 3405 16760 3423
rect 16432 3390 16490 3405
rect 16102 3347 16164 3381
rect 16102 3313 16118 3347
rect 16152 3313 16164 3347
rect 16102 3279 16164 3313
rect 17318 3415 17326 3449
rect 17360 3415 17370 3449
rect 17318 3397 17370 3415
rect 17400 3585 17452 3597
rect 17400 3551 17410 3585
rect 17444 3551 17452 3585
rect 17400 3517 17452 3551
rect 17400 3483 17410 3517
rect 17444 3483 17452 3517
rect 17400 3449 17452 3483
rect 17400 3415 17410 3449
rect 17444 3415 17452 3449
rect 17400 3397 17452 3415
rect 17586 3575 17644 3590
rect 17586 3541 17598 3575
rect 17632 3541 17644 3575
rect 17586 3507 17644 3541
rect 17586 3473 17598 3507
rect 17632 3473 17644 3507
rect 17586 3439 17644 3473
rect 17586 3405 17598 3439
rect 17632 3405 17644 3439
rect 17586 3390 17644 3405
rect 17674 3575 17732 3590
rect 17674 3541 17686 3575
rect 17720 3541 17732 3575
rect 17674 3507 17732 3541
rect 18514 3593 18566 3605
rect 18232 3575 18290 3590
rect 18232 3541 18244 3575
rect 18278 3541 18290 3575
rect 17674 3473 17686 3507
rect 17720 3473 17732 3507
rect 17674 3439 17732 3473
rect 17674 3405 17686 3439
rect 17720 3405 17732 3439
rect 18232 3507 18290 3541
rect 18232 3473 18244 3507
rect 18278 3473 18290 3507
rect 18232 3439 18290 3473
rect 17674 3390 17732 3405
rect 17802 3415 17864 3430
rect 17802 3381 17814 3415
rect 17848 3381 17864 3415
rect 16102 3245 16118 3279
rect 16152 3245 16164 3279
rect 16102 3230 16164 3245
rect 17802 3347 17864 3381
rect 17802 3313 17814 3347
rect 17848 3313 17864 3347
rect 17802 3279 17864 3313
rect 17802 3245 17814 3279
rect 17848 3245 17864 3279
rect 17802 3230 17864 3245
rect 17894 3415 17960 3430
rect 17894 3381 17910 3415
rect 17944 3381 17960 3415
rect 17894 3347 17960 3381
rect 17894 3313 17910 3347
rect 17944 3313 17960 3347
rect 17894 3279 17960 3313
rect 17894 3245 17910 3279
rect 17944 3245 17960 3279
rect 17894 3230 17960 3245
rect 17990 3415 18052 3430
rect 17990 3381 18006 3415
rect 18040 3381 18052 3415
rect 18232 3405 18244 3439
rect 18278 3405 18290 3439
rect 18232 3390 18290 3405
rect 18320 3575 18378 3590
rect 18320 3541 18332 3575
rect 18366 3541 18378 3575
rect 18320 3507 18378 3541
rect 18320 3473 18332 3507
rect 18366 3473 18378 3507
rect 18320 3439 18378 3473
rect 18320 3405 18332 3439
rect 18366 3405 18378 3439
rect 18514 3559 18522 3593
rect 18556 3559 18566 3593
rect 18514 3525 18566 3559
rect 18514 3491 18522 3525
rect 18556 3491 18566 3525
rect 18514 3457 18566 3491
rect 18514 3423 18522 3457
rect 18556 3423 18566 3457
rect 18514 3405 18566 3423
rect 18596 3593 18648 3605
rect 18596 3559 18606 3593
rect 18640 3559 18648 3593
rect 18596 3525 18648 3559
rect 18596 3491 18606 3525
rect 18640 3491 18648 3525
rect 18596 3457 18648 3491
rect 18596 3423 18606 3457
rect 18640 3423 18648 3457
rect 18819 3583 18871 3603
rect 18819 3549 18827 3583
rect 18861 3549 18871 3583
rect 18819 3515 18871 3549
rect 18819 3481 18827 3515
rect 18861 3481 18871 3515
rect 18819 3445 18871 3481
rect 18901 3583 18959 3603
rect 18901 3549 18913 3583
rect 18947 3549 18959 3583
rect 18901 3515 18959 3549
rect 18901 3481 18913 3515
rect 18947 3481 18959 3515
rect 18901 3445 18959 3481
rect 18989 3583 19041 3603
rect 18989 3549 18999 3583
rect 19033 3549 19041 3583
rect 18989 3502 19041 3549
rect 18989 3468 18999 3502
rect 19033 3468 19041 3502
rect 18989 3445 19041 3468
rect 19206 3585 19258 3597
rect 19206 3551 19214 3585
rect 19248 3551 19258 3585
rect 19206 3517 19258 3551
rect 19206 3483 19214 3517
rect 19248 3483 19258 3517
rect 19206 3449 19258 3483
rect 18596 3405 18648 3423
rect 18320 3390 18378 3405
rect 17990 3347 18052 3381
rect 17990 3313 18006 3347
rect 18040 3313 18052 3347
rect 17990 3279 18052 3313
rect 19206 3415 19214 3449
rect 19248 3415 19258 3449
rect 19206 3397 19258 3415
rect 19288 3585 19340 3597
rect 19288 3551 19298 3585
rect 19332 3551 19340 3585
rect 19288 3517 19340 3551
rect 19288 3483 19298 3517
rect 19332 3483 19340 3517
rect 19288 3449 19340 3483
rect 19288 3415 19298 3449
rect 19332 3415 19340 3449
rect 19288 3397 19340 3415
rect 19474 3575 19532 3590
rect 19474 3541 19486 3575
rect 19520 3541 19532 3575
rect 19474 3507 19532 3541
rect 19474 3473 19486 3507
rect 19520 3473 19532 3507
rect 19474 3439 19532 3473
rect 19474 3405 19486 3439
rect 19520 3405 19532 3439
rect 19474 3390 19532 3405
rect 19562 3575 19620 3590
rect 19562 3541 19574 3575
rect 19608 3541 19620 3575
rect 19562 3507 19620 3541
rect 20402 3593 20454 3605
rect 20120 3575 20178 3590
rect 20120 3541 20132 3575
rect 20166 3541 20178 3575
rect 19562 3473 19574 3507
rect 19608 3473 19620 3507
rect 19562 3439 19620 3473
rect 19562 3405 19574 3439
rect 19608 3405 19620 3439
rect 20120 3507 20178 3541
rect 20120 3473 20132 3507
rect 20166 3473 20178 3507
rect 20120 3439 20178 3473
rect 19562 3390 19620 3405
rect 19690 3415 19752 3430
rect 19690 3381 19702 3415
rect 19736 3381 19752 3415
rect 17990 3245 18006 3279
rect 18040 3245 18052 3279
rect 17990 3230 18052 3245
rect 19690 3347 19752 3381
rect 19690 3313 19702 3347
rect 19736 3313 19752 3347
rect 19690 3279 19752 3313
rect 19690 3245 19702 3279
rect 19736 3245 19752 3279
rect 19690 3230 19752 3245
rect 19782 3415 19848 3430
rect 19782 3381 19798 3415
rect 19832 3381 19848 3415
rect 19782 3347 19848 3381
rect 19782 3313 19798 3347
rect 19832 3313 19848 3347
rect 19782 3279 19848 3313
rect 19782 3245 19798 3279
rect 19832 3245 19848 3279
rect 19782 3230 19848 3245
rect 19878 3415 19940 3430
rect 19878 3381 19894 3415
rect 19928 3381 19940 3415
rect 20120 3405 20132 3439
rect 20166 3405 20178 3439
rect 20120 3390 20178 3405
rect 20208 3575 20266 3590
rect 20208 3541 20220 3575
rect 20254 3541 20266 3575
rect 20208 3507 20266 3541
rect 20208 3473 20220 3507
rect 20254 3473 20266 3507
rect 20208 3439 20266 3473
rect 20208 3405 20220 3439
rect 20254 3405 20266 3439
rect 20402 3559 20410 3593
rect 20444 3559 20454 3593
rect 20402 3525 20454 3559
rect 20402 3491 20410 3525
rect 20444 3491 20454 3525
rect 20402 3457 20454 3491
rect 20402 3423 20410 3457
rect 20444 3423 20454 3457
rect 20402 3405 20454 3423
rect 20484 3593 20536 3605
rect 20484 3559 20494 3593
rect 20528 3559 20536 3593
rect 20484 3525 20536 3559
rect 20484 3491 20494 3525
rect 20528 3491 20536 3525
rect 20484 3457 20536 3491
rect 20484 3423 20494 3457
rect 20528 3423 20536 3457
rect 20707 3583 20759 3603
rect 20707 3549 20715 3583
rect 20749 3549 20759 3583
rect 20707 3515 20759 3549
rect 20707 3481 20715 3515
rect 20749 3481 20759 3515
rect 20707 3445 20759 3481
rect 20789 3583 20847 3603
rect 20789 3549 20801 3583
rect 20835 3549 20847 3583
rect 20789 3515 20847 3549
rect 20789 3481 20801 3515
rect 20835 3481 20847 3515
rect 20789 3445 20847 3481
rect 20877 3583 20929 3603
rect 20877 3549 20887 3583
rect 20921 3549 20929 3583
rect 20877 3502 20929 3549
rect 20877 3468 20887 3502
rect 20921 3468 20929 3502
rect 20877 3445 20929 3468
rect 21094 3585 21146 3597
rect 21094 3551 21102 3585
rect 21136 3551 21146 3585
rect 21094 3517 21146 3551
rect 21094 3483 21102 3517
rect 21136 3483 21146 3517
rect 21094 3449 21146 3483
rect 20484 3405 20536 3423
rect 20208 3390 20266 3405
rect 19878 3347 19940 3381
rect 19878 3313 19894 3347
rect 19928 3313 19940 3347
rect 19878 3279 19940 3313
rect 21094 3415 21102 3449
rect 21136 3415 21146 3449
rect 21094 3397 21146 3415
rect 21176 3585 21228 3597
rect 21176 3551 21186 3585
rect 21220 3551 21228 3585
rect 21176 3517 21228 3551
rect 21176 3483 21186 3517
rect 21220 3483 21228 3517
rect 21176 3449 21228 3483
rect 21176 3415 21186 3449
rect 21220 3415 21228 3449
rect 21176 3397 21228 3415
rect 21362 3575 21420 3590
rect 21362 3541 21374 3575
rect 21408 3541 21420 3575
rect 21362 3507 21420 3541
rect 21362 3473 21374 3507
rect 21408 3473 21420 3507
rect 21362 3439 21420 3473
rect 21362 3405 21374 3439
rect 21408 3405 21420 3439
rect 21362 3390 21420 3405
rect 21450 3575 21508 3590
rect 21450 3541 21462 3575
rect 21496 3541 21508 3575
rect 21450 3507 21508 3541
rect 22290 3593 22342 3605
rect 22008 3575 22066 3590
rect 22008 3541 22020 3575
rect 22054 3541 22066 3575
rect 21450 3473 21462 3507
rect 21496 3473 21508 3507
rect 21450 3439 21508 3473
rect 21450 3405 21462 3439
rect 21496 3405 21508 3439
rect 22008 3507 22066 3541
rect 22008 3473 22020 3507
rect 22054 3473 22066 3507
rect 22008 3439 22066 3473
rect 21450 3390 21508 3405
rect 21578 3415 21640 3430
rect 21578 3381 21590 3415
rect 21624 3381 21640 3415
rect 19878 3245 19894 3279
rect 19928 3245 19940 3279
rect 19878 3230 19940 3245
rect 21578 3347 21640 3381
rect 21578 3313 21590 3347
rect 21624 3313 21640 3347
rect 21578 3279 21640 3313
rect 21578 3245 21590 3279
rect 21624 3245 21640 3279
rect 21578 3230 21640 3245
rect 21670 3415 21736 3430
rect 21670 3381 21686 3415
rect 21720 3381 21736 3415
rect 21670 3347 21736 3381
rect 21670 3313 21686 3347
rect 21720 3313 21736 3347
rect 21670 3279 21736 3313
rect 21670 3245 21686 3279
rect 21720 3245 21736 3279
rect 21670 3230 21736 3245
rect 21766 3415 21828 3430
rect 21766 3381 21782 3415
rect 21816 3381 21828 3415
rect 22008 3405 22020 3439
rect 22054 3405 22066 3439
rect 22008 3390 22066 3405
rect 22096 3575 22154 3590
rect 22096 3541 22108 3575
rect 22142 3541 22154 3575
rect 22096 3507 22154 3541
rect 22096 3473 22108 3507
rect 22142 3473 22154 3507
rect 22096 3439 22154 3473
rect 22096 3405 22108 3439
rect 22142 3405 22154 3439
rect 22290 3559 22298 3593
rect 22332 3559 22342 3593
rect 22290 3525 22342 3559
rect 22290 3491 22298 3525
rect 22332 3491 22342 3525
rect 22290 3457 22342 3491
rect 22290 3423 22298 3457
rect 22332 3423 22342 3457
rect 22290 3405 22342 3423
rect 22372 3593 22424 3605
rect 22372 3559 22382 3593
rect 22416 3559 22424 3593
rect 22372 3525 22424 3559
rect 22372 3491 22382 3525
rect 22416 3491 22424 3525
rect 22372 3457 22424 3491
rect 22372 3423 22382 3457
rect 22416 3423 22424 3457
rect 22595 3583 22647 3603
rect 22595 3549 22603 3583
rect 22637 3549 22647 3583
rect 22595 3515 22647 3549
rect 22595 3481 22603 3515
rect 22637 3481 22647 3515
rect 22595 3445 22647 3481
rect 22677 3583 22735 3603
rect 22677 3549 22689 3583
rect 22723 3549 22735 3583
rect 22677 3515 22735 3549
rect 22677 3481 22689 3515
rect 22723 3481 22735 3515
rect 22677 3445 22735 3481
rect 22765 3583 22817 3603
rect 22765 3549 22775 3583
rect 22809 3549 22817 3583
rect 22765 3502 22817 3549
rect 22765 3468 22775 3502
rect 22809 3468 22817 3502
rect 22765 3445 22817 3468
rect 22982 3585 23034 3597
rect 22982 3551 22990 3585
rect 23024 3551 23034 3585
rect 22982 3517 23034 3551
rect 22982 3483 22990 3517
rect 23024 3483 23034 3517
rect 22982 3449 23034 3483
rect 22372 3405 22424 3423
rect 22096 3390 22154 3405
rect 21766 3347 21828 3381
rect 21766 3313 21782 3347
rect 21816 3313 21828 3347
rect 21766 3279 21828 3313
rect 22982 3415 22990 3449
rect 23024 3415 23034 3449
rect 22982 3397 23034 3415
rect 23064 3585 23116 3597
rect 23064 3551 23074 3585
rect 23108 3551 23116 3585
rect 23064 3517 23116 3551
rect 23064 3483 23074 3517
rect 23108 3483 23116 3517
rect 23064 3449 23116 3483
rect 23064 3415 23074 3449
rect 23108 3415 23116 3449
rect 23064 3397 23116 3415
rect 23250 3575 23308 3590
rect 23250 3541 23262 3575
rect 23296 3541 23308 3575
rect 23250 3507 23308 3541
rect 23250 3473 23262 3507
rect 23296 3473 23308 3507
rect 23250 3439 23308 3473
rect 23250 3405 23262 3439
rect 23296 3405 23308 3439
rect 23250 3390 23308 3405
rect 23338 3575 23396 3590
rect 23338 3541 23350 3575
rect 23384 3541 23396 3575
rect 23338 3507 23396 3541
rect 24178 3593 24230 3605
rect 23896 3575 23954 3590
rect 23896 3541 23908 3575
rect 23942 3541 23954 3575
rect 23338 3473 23350 3507
rect 23384 3473 23396 3507
rect 23338 3439 23396 3473
rect 23338 3405 23350 3439
rect 23384 3405 23396 3439
rect 23896 3507 23954 3541
rect 23896 3473 23908 3507
rect 23942 3473 23954 3507
rect 23896 3439 23954 3473
rect 23338 3390 23396 3405
rect 23466 3415 23528 3430
rect 23466 3381 23478 3415
rect 23512 3381 23528 3415
rect 21766 3245 21782 3279
rect 21816 3245 21828 3279
rect 21766 3230 21828 3245
rect 23466 3347 23528 3381
rect 23466 3313 23478 3347
rect 23512 3313 23528 3347
rect 23466 3279 23528 3313
rect 23466 3245 23478 3279
rect 23512 3245 23528 3279
rect 23466 3230 23528 3245
rect 23558 3415 23624 3430
rect 23558 3381 23574 3415
rect 23608 3381 23624 3415
rect 23558 3347 23624 3381
rect 23558 3313 23574 3347
rect 23608 3313 23624 3347
rect 23558 3279 23624 3313
rect 23558 3245 23574 3279
rect 23608 3245 23624 3279
rect 23558 3230 23624 3245
rect 23654 3415 23716 3430
rect 23654 3381 23670 3415
rect 23704 3381 23716 3415
rect 23896 3405 23908 3439
rect 23942 3405 23954 3439
rect 23896 3390 23954 3405
rect 23984 3575 24042 3590
rect 23984 3541 23996 3575
rect 24030 3541 24042 3575
rect 23984 3507 24042 3541
rect 23984 3473 23996 3507
rect 24030 3473 24042 3507
rect 23984 3439 24042 3473
rect 23984 3405 23996 3439
rect 24030 3405 24042 3439
rect 24178 3559 24186 3593
rect 24220 3559 24230 3593
rect 24178 3525 24230 3559
rect 24178 3491 24186 3525
rect 24220 3491 24230 3525
rect 24178 3457 24230 3491
rect 24178 3423 24186 3457
rect 24220 3423 24230 3457
rect 24178 3405 24230 3423
rect 24260 3593 24312 3605
rect 24260 3559 24270 3593
rect 24304 3559 24312 3593
rect 24260 3525 24312 3559
rect 24260 3491 24270 3525
rect 24304 3491 24312 3525
rect 24260 3457 24312 3491
rect 24260 3423 24270 3457
rect 24304 3423 24312 3457
rect 24483 3583 24535 3603
rect 24483 3549 24491 3583
rect 24525 3549 24535 3583
rect 24483 3515 24535 3549
rect 24483 3481 24491 3515
rect 24525 3481 24535 3515
rect 24483 3445 24535 3481
rect 24565 3583 24623 3603
rect 24565 3549 24577 3583
rect 24611 3549 24623 3583
rect 24565 3515 24623 3549
rect 24565 3481 24577 3515
rect 24611 3481 24623 3515
rect 24565 3445 24623 3481
rect 24653 3583 24705 3603
rect 24653 3549 24663 3583
rect 24697 3549 24705 3583
rect 24653 3502 24705 3549
rect 24653 3468 24663 3502
rect 24697 3468 24705 3502
rect 24653 3445 24705 3468
rect 24870 3585 24922 3597
rect 24870 3551 24878 3585
rect 24912 3551 24922 3585
rect 24870 3517 24922 3551
rect 24870 3483 24878 3517
rect 24912 3483 24922 3517
rect 24870 3449 24922 3483
rect 24260 3405 24312 3423
rect 23984 3390 24042 3405
rect 23654 3347 23716 3381
rect 23654 3313 23670 3347
rect 23704 3313 23716 3347
rect 23654 3279 23716 3313
rect 24870 3415 24878 3449
rect 24912 3415 24922 3449
rect 24870 3397 24922 3415
rect 24952 3585 25004 3597
rect 24952 3551 24962 3585
rect 24996 3551 25004 3585
rect 24952 3517 25004 3551
rect 24952 3483 24962 3517
rect 24996 3483 25004 3517
rect 24952 3449 25004 3483
rect 24952 3415 24962 3449
rect 24996 3415 25004 3449
rect 24952 3397 25004 3415
rect 25138 3575 25196 3590
rect 25138 3541 25150 3575
rect 25184 3541 25196 3575
rect 25138 3507 25196 3541
rect 25138 3473 25150 3507
rect 25184 3473 25196 3507
rect 25138 3439 25196 3473
rect 25138 3405 25150 3439
rect 25184 3405 25196 3439
rect 25138 3390 25196 3405
rect 25226 3575 25284 3590
rect 25226 3541 25238 3575
rect 25272 3541 25284 3575
rect 25226 3507 25284 3541
rect 26066 3593 26118 3605
rect 25784 3575 25842 3590
rect 25784 3541 25796 3575
rect 25830 3541 25842 3575
rect 25226 3473 25238 3507
rect 25272 3473 25284 3507
rect 25226 3439 25284 3473
rect 25226 3405 25238 3439
rect 25272 3405 25284 3439
rect 25784 3507 25842 3541
rect 25784 3473 25796 3507
rect 25830 3473 25842 3507
rect 25784 3439 25842 3473
rect 25226 3390 25284 3405
rect 25354 3415 25416 3430
rect 25354 3381 25366 3415
rect 25400 3381 25416 3415
rect 23654 3245 23670 3279
rect 23704 3245 23716 3279
rect 23654 3230 23716 3245
rect 25354 3347 25416 3381
rect 25354 3313 25366 3347
rect 25400 3313 25416 3347
rect 25354 3279 25416 3313
rect 25354 3245 25366 3279
rect 25400 3245 25416 3279
rect 25354 3230 25416 3245
rect 25446 3415 25512 3430
rect 25446 3381 25462 3415
rect 25496 3381 25512 3415
rect 25446 3347 25512 3381
rect 25446 3313 25462 3347
rect 25496 3313 25512 3347
rect 25446 3279 25512 3313
rect 25446 3245 25462 3279
rect 25496 3245 25512 3279
rect 25446 3230 25512 3245
rect 25542 3415 25604 3430
rect 25542 3381 25558 3415
rect 25592 3381 25604 3415
rect 25784 3405 25796 3439
rect 25830 3405 25842 3439
rect 25784 3390 25842 3405
rect 25872 3575 25930 3590
rect 25872 3541 25884 3575
rect 25918 3541 25930 3575
rect 25872 3507 25930 3541
rect 25872 3473 25884 3507
rect 25918 3473 25930 3507
rect 25872 3439 25930 3473
rect 25872 3405 25884 3439
rect 25918 3405 25930 3439
rect 26066 3559 26074 3593
rect 26108 3559 26118 3593
rect 26066 3525 26118 3559
rect 26066 3491 26074 3525
rect 26108 3491 26118 3525
rect 26066 3457 26118 3491
rect 26066 3423 26074 3457
rect 26108 3423 26118 3457
rect 26066 3405 26118 3423
rect 26148 3593 26200 3605
rect 26148 3559 26158 3593
rect 26192 3559 26200 3593
rect 26148 3525 26200 3559
rect 26148 3491 26158 3525
rect 26192 3491 26200 3525
rect 26148 3457 26200 3491
rect 26148 3423 26158 3457
rect 26192 3423 26200 3457
rect 26371 3583 26423 3603
rect 26371 3549 26379 3583
rect 26413 3549 26423 3583
rect 26371 3515 26423 3549
rect 26371 3481 26379 3515
rect 26413 3481 26423 3515
rect 26371 3445 26423 3481
rect 26453 3583 26511 3603
rect 26453 3549 26465 3583
rect 26499 3549 26511 3583
rect 26453 3515 26511 3549
rect 26453 3481 26465 3515
rect 26499 3481 26511 3515
rect 26453 3445 26511 3481
rect 26541 3583 26593 3603
rect 26541 3549 26551 3583
rect 26585 3549 26593 3583
rect 26541 3502 26593 3549
rect 26541 3468 26551 3502
rect 26585 3468 26593 3502
rect 26541 3445 26593 3468
rect 26148 3405 26200 3423
rect 25872 3390 25930 3405
rect 25542 3347 25604 3381
rect 25542 3313 25558 3347
rect 25592 3313 25604 3347
rect 25542 3279 25604 3313
rect 25542 3245 25558 3279
rect 25592 3245 25604 3279
rect 25542 3230 25604 3245
<< ndiffc >>
rect 2160 5229 2194 5263
rect 2160 5161 2194 5195
rect 2244 5229 2278 5263
rect 2244 5161 2278 5195
rect 2328 5229 2362 5263
rect 2412 5229 2446 5263
rect 2412 5161 2446 5195
rect 2496 5229 2530 5263
rect 2580 5229 2614 5263
rect 2580 5161 2614 5195
rect 2664 5229 2698 5263
rect 2748 5229 2782 5263
rect 2748 5161 2782 5195
rect 2832 5229 2866 5263
rect 2916 5229 2950 5263
rect 2916 5161 2950 5195
rect 3000 5229 3034 5263
rect 3084 5229 3118 5263
rect 3084 5161 3118 5195
rect 3168 5229 3202 5263
rect 3252 5229 3286 5263
rect 3252 5161 3286 5195
rect 3336 5229 3370 5263
rect 3420 5229 3454 5263
rect 3420 5161 3454 5195
rect 3504 5229 3538 5263
rect 3504 5161 3538 5195
rect 4042 5227 4076 5261
rect 4042 5159 4076 5193
rect 4126 5227 4160 5261
rect 4126 5159 4160 5193
rect 4210 5227 4244 5261
rect 4294 5227 4328 5261
rect 4294 5159 4328 5193
rect 4378 5227 4412 5261
rect 4462 5227 4496 5261
rect 4462 5159 4496 5193
rect 4546 5227 4580 5261
rect 4630 5227 4664 5261
rect 4630 5159 4664 5193
rect 4714 5227 4748 5261
rect 4798 5227 4832 5261
rect 4798 5159 4832 5193
rect 4882 5227 4916 5261
rect 4966 5227 5000 5261
rect 4966 5159 5000 5193
rect 5050 5227 5084 5261
rect 5134 5227 5168 5261
rect 5134 5159 5168 5193
rect 5218 5227 5252 5261
rect 5302 5227 5336 5261
rect 5302 5159 5336 5193
rect 5386 5227 5420 5261
rect 5386 5159 5420 5193
rect 17258 5229 17292 5263
rect 17258 5161 17292 5195
rect 17342 5229 17376 5263
rect 17342 5161 17376 5195
rect 17426 5229 17460 5263
rect 17510 5229 17544 5263
rect 17510 5161 17544 5195
rect 17594 5229 17628 5263
rect 17678 5229 17712 5263
rect 17678 5161 17712 5195
rect 17762 5229 17796 5263
rect 17846 5229 17880 5263
rect 17846 5161 17880 5195
rect 17930 5229 17964 5263
rect 18014 5229 18048 5263
rect 18014 5161 18048 5195
rect 18098 5229 18132 5263
rect 18182 5229 18216 5263
rect 18182 5161 18216 5195
rect 18266 5229 18300 5263
rect 18350 5229 18384 5263
rect 18350 5161 18384 5195
rect 18434 5229 18468 5263
rect 18518 5229 18552 5263
rect 18518 5161 18552 5195
rect 18602 5229 18636 5263
rect 18602 5161 18636 5195
rect 19140 5227 19174 5261
rect 19140 5159 19174 5193
rect 19224 5227 19258 5261
rect 19224 5159 19258 5193
rect 19308 5227 19342 5261
rect 19392 5227 19426 5261
rect 19392 5159 19426 5193
rect 19476 5227 19510 5261
rect 19560 5227 19594 5261
rect 19560 5159 19594 5193
rect 19644 5227 19678 5261
rect 19728 5227 19762 5261
rect 19728 5159 19762 5193
rect 19812 5227 19846 5261
rect 19896 5227 19930 5261
rect 19896 5159 19930 5193
rect 19980 5227 20014 5261
rect 20064 5227 20098 5261
rect 20064 5159 20098 5193
rect 20148 5227 20182 5261
rect 20232 5227 20266 5261
rect 20232 5159 20266 5193
rect 20316 5227 20350 5261
rect 20400 5227 20434 5261
rect 20400 5159 20434 5193
rect 20484 5227 20518 5261
rect 20484 5159 20518 5193
rect -3299 4283 -3265 4317
rect -3299 4215 -3265 4249
rect -3215 4283 -3181 4317
rect -3215 4215 -3181 4249
rect -3131 4283 -3097 4317
rect -2485 4283 -2451 4317
rect -3131 4215 -3097 4249
rect -2485 4215 -2451 4249
rect -2401 4283 -2367 4317
rect -2401 4215 -2367 4249
rect -2317 4283 -2283 4317
rect -2317 4215 -2283 4249
rect -1411 4283 -1377 4317
rect -1411 4215 -1377 4249
rect -1327 4283 -1293 4317
rect -1327 4215 -1293 4249
rect -1243 4283 -1209 4317
rect -597 4283 -563 4317
rect -1243 4215 -1209 4249
rect -597 4215 -563 4249
rect -513 4283 -479 4317
rect -513 4215 -479 4249
rect -429 4283 -395 4317
rect -429 4215 -395 4249
rect 477 4283 511 4317
rect 477 4215 511 4249
rect 561 4283 595 4317
rect 561 4215 595 4249
rect 645 4283 679 4317
rect 1291 4283 1325 4317
rect 645 4215 679 4249
rect 1291 4215 1325 4249
rect 1375 4283 1409 4317
rect 1375 4215 1409 4249
rect 1459 4283 1493 4317
rect 1459 4215 1493 4249
rect 2365 4283 2399 4317
rect 2365 4215 2399 4249
rect 2449 4283 2483 4317
rect 2449 4215 2483 4249
rect 2533 4283 2567 4317
rect 3179 4283 3213 4317
rect 2533 4215 2567 4249
rect 3179 4215 3213 4249
rect 3263 4283 3297 4317
rect 3263 4215 3297 4249
rect 3347 4283 3381 4317
rect 3347 4215 3381 4249
rect 4253 4283 4287 4317
rect 4253 4215 4287 4249
rect 4337 4283 4371 4317
rect 4337 4215 4371 4249
rect 4421 4283 4455 4317
rect 5067 4283 5101 4317
rect 4421 4215 4455 4249
rect 5067 4215 5101 4249
rect 5151 4283 5185 4317
rect 5151 4215 5185 4249
rect 5235 4283 5269 4317
rect 5235 4215 5269 4249
rect 6141 4283 6175 4317
rect 6141 4215 6175 4249
rect 6225 4283 6259 4317
rect 6225 4215 6259 4249
rect 6309 4283 6343 4317
rect 6955 4283 6989 4317
rect 6309 4215 6343 4249
rect 6955 4215 6989 4249
rect 7039 4283 7073 4317
rect 7039 4215 7073 4249
rect 7123 4283 7157 4317
rect 7123 4215 7157 4249
rect 8029 4283 8063 4317
rect 8029 4215 8063 4249
rect 8113 4283 8147 4317
rect 8113 4215 8147 4249
rect 8197 4283 8231 4317
rect 8843 4283 8877 4317
rect 8197 4215 8231 4249
rect 8843 4215 8877 4249
rect 8927 4283 8961 4317
rect 8927 4215 8961 4249
rect 9011 4283 9045 4317
rect 9011 4215 9045 4249
rect 9917 4283 9951 4317
rect 9917 4215 9951 4249
rect 10001 4283 10035 4317
rect 10001 4215 10035 4249
rect 10085 4283 10119 4317
rect 10731 4283 10765 4317
rect 10085 4215 10119 4249
rect 10731 4215 10765 4249
rect 10815 4283 10849 4317
rect 10815 4215 10849 4249
rect 10899 4283 10933 4317
rect 10899 4215 10933 4249
rect 11799 4283 11833 4317
rect 11799 4215 11833 4249
rect 11883 4283 11917 4317
rect 11883 4215 11917 4249
rect 11967 4283 12001 4317
rect 12613 4283 12647 4317
rect 11967 4215 12001 4249
rect 12613 4215 12647 4249
rect 12697 4283 12731 4317
rect 12697 4215 12731 4249
rect 12781 4283 12815 4317
rect 12781 4215 12815 4249
rect 13687 4283 13721 4317
rect 13687 4215 13721 4249
rect 13771 4283 13805 4317
rect 13771 4215 13805 4249
rect 13855 4283 13889 4317
rect 14501 4283 14535 4317
rect 13855 4215 13889 4249
rect 14501 4215 14535 4249
rect 14585 4283 14619 4317
rect 14585 4215 14619 4249
rect 14669 4283 14703 4317
rect 14669 4215 14703 4249
rect 15575 4283 15609 4317
rect 15575 4215 15609 4249
rect 15659 4283 15693 4317
rect 15659 4215 15693 4249
rect 15743 4283 15777 4317
rect 16389 4283 16423 4317
rect 15743 4215 15777 4249
rect 16389 4215 16423 4249
rect 16473 4283 16507 4317
rect 16473 4215 16507 4249
rect 16557 4283 16591 4317
rect 16557 4215 16591 4249
rect 17463 4283 17497 4317
rect 17463 4215 17497 4249
rect 17547 4283 17581 4317
rect 17547 4215 17581 4249
rect 17631 4283 17665 4317
rect 18277 4283 18311 4317
rect 17631 4215 17665 4249
rect 18277 4215 18311 4249
rect 18361 4283 18395 4317
rect 18361 4215 18395 4249
rect 18445 4283 18479 4317
rect 18445 4215 18479 4249
rect 19351 4283 19385 4317
rect 19351 4215 19385 4249
rect 19435 4283 19469 4317
rect 19435 4215 19469 4249
rect 19519 4283 19553 4317
rect 20165 4283 20199 4317
rect 19519 4215 19553 4249
rect 20165 4215 20199 4249
rect 20249 4283 20283 4317
rect 20249 4215 20283 4249
rect 20333 4283 20367 4317
rect 20333 4215 20367 4249
rect 21239 4283 21273 4317
rect 21239 4215 21273 4249
rect 21323 4283 21357 4317
rect 21323 4215 21357 4249
rect 21407 4283 21441 4317
rect 22053 4283 22087 4317
rect 21407 4215 21441 4249
rect 22053 4215 22087 4249
rect 22137 4283 22171 4317
rect 22137 4215 22171 4249
rect 22221 4283 22255 4317
rect 22221 4215 22255 4249
rect 23127 4283 23161 4317
rect 23127 4215 23161 4249
rect 23211 4283 23245 4317
rect 23211 4215 23245 4249
rect 23295 4283 23329 4317
rect 23941 4283 23975 4317
rect 23295 4215 23329 4249
rect 23941 4215 23975 4249
rect 24025 4283 24059 4317
rect 24025 4215 24059 4249
rect 24109 4283 24143 4317
rect 24109 4215 24143 4249
rect 25015 4283 25049 4317
rect 25015 4215 25049 4249
rect 25099 4283 25133 4317
rect 25099 4215 25133 4249
rect 25183 4283 25217 4317
rect 25829 4283 25863 4317
rect 25183 4215 25217 4249
rect 25829 4215 25863 4249
rect 25913 4283 25947 4317
rect 25913 4215 25947 4249
rect 25997 4283 26031 4317
rect 25997 4215 26031 4249
rect -2930 4038 -2896 4072
rect -2930 3970 -2896 4004
rect -2834 4038 -2800 4072
rect -2834 3970 -2800 4004
rect -2738 4038 -2704 4072
rect -2738 3970 -2704 4004
rect -1042 4038 -1008 4072
rect -1042 3970 -1008 4004
rect -946 4038 -912 4072
rect -946 3970 -912 4004
rect -850 4038 -816 4072
rect -850 3970 -816 4004
rect 846 4038 880 4072
rect 846 3970 880 4004
rect 942 4038 976 4072
rect 942 3970 976 4004
rect 1038 4038 1072 4072
rect 1038 3970 1072 4004
rect 2734 4038 2768 4072
rect 2734 3970 2768 4004
rect 2830 4038 2864 4072
rect 2830 3970 2864 4004
rect 2926 4038 2960 4072
rect 2926 3970 2960 4004
rect 4622 4038 4656 4072
rect 4622 3970 4656 4004
rect 4718 4038 4752 4072
rect 4718 3970 4752 4004
rect 4814 4038 4848 4072
rect 4814 3970 4848 4004
rect 6510 4038 6544 4072
rect 6510 3970 6544 4004
rect 6606 4038 6640 4072
rect 6606 3970 6640 4004
rect 6702 4038 6736 4072
rect 6702 3970 6736 4004
rect 8398 4038 8432 4072
rect 8398 3970 8432 4004
rect 8494 4038 8528 4072
rect 8494 3970 8528 4004
rect 8590 4038 8624 4072
rect 8590 3970 8624 4004
rect 10286 4038 10320 4072
rect 10286 3970 10320 4004
rect 10382 4038 10416 4072
rect 10382 3970 10416 4004
rect 10478 4038 10512 4072
rect 10478 3970 10512 4004
rect 12168 4038 12202 4072
rect 12168 3970 12202 4004
rect 12264 4038 12298 4072
rect 12264 3970 12298 4004
rect 12360 4038 12394 4072
rect 12360 3970 12394 4004
rect 14056 4038 14090 4072
rect 14056 3970 14090 4004
rect 14152 4038 14186 4072
rect 14152 3970 14186 4004
rect 14248 4038 14282 4072
rect 14248 3970 14282 4004
rect 15944 4038 15978 4072
rect 15944 3970 15978 4004
rect 16040 4038 16074 4072
rect 16040 3970 16074 4004
rect 16136 4038 16170 4072
rect 16136 3970 16170 4004
rect 17832 4038 17866 4072
rect 17832 3970 17866 4004
rect 17928 4038 17962 4072
rect 17928 3970 17962 4004
rect 18024 4038 18058 4072
rect 18024 3970 18058 4004
rect 19720 4038 19754 4072
rect 19720 3970 19754 4004
rect 19816 4038 19850 4072
rect 19816 3970 19850 4004
rect 19912 4038 19946 4072
rect 19912 3970 19946 4004
rect 21608 4038 21642 4072
rect 21608 3970 21642 4004
rect 21704 4038 21738 4072
rect 21704 3970 21738 4004
rect 21800 4038 21834 4072
rect 21800 3970 21834 4004
rect 23496 4038 23530 4072
rect 23496 3970 23530 4004
rect 23592 4038 23626 4072
rect 23592 3970 23626 4004
rect 23688 4038 23722 4072
rect 23688 3970 23722 4004
rect 25384 4038 25418 4072
rect 25384 3970 25418 4004
rect 25480 4038 25514 4072
rect 25480 3970 25514 4004
rect 25576 4038 25610 4072
rect 25576 3970 25610 4004
rect -3436 3231 -3402 3265
rect -3436 3163 -3402 3197
rect -3352 3231 -3318 3265
rect -2240 3239 -2206 3273
rect -3352 3163 -3318 3197
rect -2240 3171 -2206 3205
rect -2156 3239 -2122 3273
rect -2156 3171 -2122 3205
rect -1935 3178 -1901 3212
rect -1849 3165 -1815 3199
rect -1763 3195 -1729 3229
rect -1548 3231 -1514 3265
rect -1548 3163 -1514 3197
rect -1464 3231 -1430 3265
rect -352 3239 -318 3273
rect -1464 3163 -1430 3197
rect -352 3171 -318 3205
rect -268 3239 -234 3273
rect -268 3171 -234 3205
rect -47 3178 -13 3212
rect 39 3165 73 3199
rect 125 3195 159 3229
rect 340 3231 374 3265
rect 340 3163 374 3197
rect 424 3231 458 3265
rect 1536 3239 1570 3273
rect 424 3163 458 3197
rect 1536 3171 1570 3205
rect 1620 3239 1654 3273
rect 1620 3171 1654 3205
rect 1841 3178 1875 3212
rect 1927 3165 1961 3199
rect 2013 3195 2047 3229
rect 2228 3231 2262 3265
rect 2228 3163 2262 3197
rect 2312 3231 2346 3265
rect 3424 3239 3458 3273
rect 2312 3163 2346 3197
rect 3424 3171 3458 3205
rect 3508 3239 3542 3273
rect 3508 3171 3542 3205
rect 3729 3178 3763 3212
rect 3815 3165 3849 3199
rect 3901 3195 3935 3229
rect 4116 3231 4150 3265
rect 4116 3163 4150 3197
rect 4200 3231 4234 3265
rect 5312 3239 5346 3273
rect 4200 3163 4234 3197
rect 5312 3171 5346 3205
rect 5396 3239 5430 3273
rect 5396 3171 5430 3205
rect 5617 3178 5651 3212
rect 5703 3165 5737 3199
rect 5789 3195 5823 3229
rect 6004 3231 6038 3265
rect 6004 3163 6038 3197
rect 6088 3231 6122 3265
rect 7200 3239 7234 3273
rect 6088 3163 6122 3197
rect 7200 3171 7234 3205
rect 7284 3239 7318 3273
rect 7284 3171 7318 3205
rect 7505 3178 7539 3212
rect 7591 3165 7625 3199
rect 7677 3195 7711 3229
rect 7892 3231 7926 3265
rect 7892 3163 7926 3197
rect 7976 3231 8010 3265
rect 9088 3239 9122 3273
rect 7976 3163 8010 3197
rect 9088 3171 9122 3205
rect 9172 3239 9206 3273
rect 9172 3171 9206 3205
rect 9393 3178 9427 3212
rect 9479 3165 9513 3199
rect 9565 3195 9599 3229
rect 9780 3231 9814 3265
rect 9780 3163 9814 3197
rect 9864 3231 9898 3265
rect 10976 3239 11010 3273
rect 9864 3163 9898 3197
rect 10976 3171 11010 3205
rect 11060 3239 11094 3273
rect 11060 3171 11094 3205
rect 11281 3178 11315 3212
rect 11367 3165 11401 3199
rect 11453 3195 11487 3229
rect 11662 3231 11696 3265
rect 11662 3163 11696 3197
rect 11746 3231 11780 3265
rect 12858 3239 12892 3273
rect 11746 3163 11780 3197
rect 12858 3171 12892 3205
rect 12942 3239 12976 3273
rect 12942 3171 12976 3205
rect 13163 3178 13197 3212
rect 13249 3165 13283 3199
rect 13335 3195 13369 3229
rect 13550 3231 13584 3265
rect 13550 3163 13584 3197
rect 13634 3231 13668 3265
rect 14746 3239 14780 3273
rect 13634 3163 13668 3197
rect 14746 3171 14780 3205
rect 14830 3239 14864 3273
rect 14830 3171 14864 3205
rect 15051 3178 15085 3212
rect 15137 3165 15171 3199
rect 15223 3195 15257 3229
rect 15438 3231 15472 3265
rect 15438 3163 15472 3197
rect 15522 3231 15556 3265
rect 16634 3239 16668 3273
rect 15522 3163 15556 3197
rect 16634 3171 16668 3205
rect 16718 3239 16752 3273
rect 16718 3171 16752 3205
rect 16939 3178 16973 3212
rect 17025 3165 17059 3199
rect 17111 3195 17145 3229
rect 17326 3231 17360 3265
rect 17326 3163 17360 3197
rect 17410 3231 17444 3265
rect 18522 3239 18556 3273
rect 17410 3163 17444 3197
rect 18522 3171 18556 3205
rect 18606 3239 18640 3273
rect 18606 3171 18640 3205
rect 18827 3178 18861 3212
rect 18913 3165 18947 3199
rect 18999 3195 19033 3229
rect 19214 3231 19248 3265
rect 19214 3163 19248 3197
rect 19298 3231 19332 3265
rect 20410 3239 20444 3273
rect 19298 3163 19332 3197
rect 20410 3171 20444 3205
rect 20494 3239 20528 3273
rect 20494 3171 20528 3205
rect 20715 3178 20749 3212
rect 20801 3165 20835 3199
rect 20887 3195 20921 3229
rect 21102 3231 21136 3265
rect 21102 3163 21136 3197
rect 21186 3231 21220 3265
rect 22298 3239 22332 3273
rect 21186 3163 21220 3197
rect 22298 3171 22332 3205
rect 22382 3239 22416 3273
rect 22382 3171 22416 3205
rect 22603 3178 22637 3212
rect 22689 3165 22723 3199
rect 22775 3195 22809 3229
rect 22990 3231 23024 3265
rect 22990 3163 23024 3197
rect 23074 3231 23108 3265
rect 24186 3239 24220 3273
rect 23074 3163 23108 3197
rect 24186 3171 24220 3205
rect 24270 3239 24304 3273
rect 24270 3171 24304 3205
rect 24491 3178 24525 3212
rect 24577 3165 24611 3199
rect 24663 3195 24697 3229
rect 24878 3231 24912 3265
rect 24878 3163 24912 3197
rect 24962 3231 24996 3265
rect 26074 3239 26108 3273
rect 24962 3163 24996 3197
rect 26074 3171 26108 3205
rect 26158 3239 26192 3273
rect 26158 3171 26192 3205
rect 26379 3178 26413 3212
rect 26465 3165 26499 3199
rect 26551 3195 26585 3229
rect -2932 2982 -2898 3016
rect -2932 2914 -2898 2948
rect -2836 2982 -2802 3016
rect -2836 2914 -2802 2948
rect -2740 2982 -2706 3016
rect -2740 2914 -2706 2948
rect -1044 2982 -1010 3016
rect -1044 2914 -1010 2948
rect -948 2982 -914 3016
rect -948 2914 -914 2948
rect -852 2982 -818 3016
rect -852 2914 -818 2948
rect 844 2982 878 3016
rect 844 2914 878 2948
rect 940 2982 974 3016
rect 940 2914 974 2948
rect 1036 2982 1070 3016
rect 1036 2914 1070 2948
rect 2732 2982 2766 3016
rect 2732 2914 2766 2948
rect 2828 2982 2862 3016
rect 2828 2914 2862 2948
rect 2924 2982 2958 3016
rect 2924 2914 2958 2948
rect 4620 2982 4654 3016
rect 4620 2914 4654 2948
rect 4716 2982 4750 3016
rect 4716 2914 4750 2948
rect 4812 2982 4846 3016
rect 4812 2914 4846 2948
rect 6508 2982 6542 3016
rect 6508 2914 6542 2948
rect 6604 2982 6638 3016
rect 6604 2914 6638 2948
rect 6700 2982 6734 3016
rect 6700 2914 6734 2948
rect 8396 2982 8430 3016
rect 8396 2914 8430 2948
rect 8492 2982 8526 3016
rect 8492 2914 8526 2948
rect 8588 2982 8622 3016
rect 8588 2914 8622 2948
rect 10284 2982 10318 3016
rect 10284 2914 10318 2948
rect 10380 2982 10414 3016
rect 10380 2914 10414 2948
rect 10476 2982 10510 3016
rect 10476 2914 10510 2948
rect 12166 2982 12200 3016
rect 12166 2914 12200 2948
rect 12262 2982 12296 3016
rect 12262 2914 12296 2948
rect 12358 2982 12392 3016
rect 12358 2914 12392 2948
rect 14054 2982 14088 3016
rect 14054 2914 14088 2948
rect 14150 2982 14184 3016
rect 14150 2914 14184 2948
rect 14246 2982 14280 3016
rect 14246 2914 14280 2948
rect 15942 2982 15976 3016
rect 15942 2914 15976 2948
rect 16038 2982 16072 3016
rect 16038 2914 16072 2948
rect 16134 2982 16168 3016
rect 16134 2914 16168 2948
rect 17830 2982 17864 3016
rect 17830 2914 17864 2948
rect 17926 2982 17960 3016
rect 17926 2914 17960 2948
rect 18022 2982 18056 3016
rect 18022 2914 18056 2948
rect 19718 2982 19752 3016
rect 19718 2914 19752 2948
rect 19814 2982 19848 3016
rect 19814 2914 19848 2948
rect 19910 2982 19944 3016
rect 19910 2914 19944 2948
rect 21606 2982 21640 3016
rect 21606 2914 21640 2948
rect 21702 2982 21736 3016
rect 21702 2914 21736 2948
rect 21798 2982 21832 3016
rect 21798 2914 21832 2948
rect 23494 2982 23528 3016
rect 23494 2914 23528 2948
rect 23590 2982 23624 3016
rect 23590 2914 23624 2948
rect 23686 2982 23720 3016
rect 23686 2914 23720 2948
rect 25382 2982 25416 3016
rect 25382 2914 25416 2948
rect 25478 2982 25512 3016
rect 25478 2914 25512 2948
rect 25574 2982 25608 3016
rect 25574 2914 25608 2948
<< pdiffc >>
rect 2160 4975 2194 5009
rect 2160 4905 2194 4939
rect 2160 4837 2194 4871
rect 2244 4975 2278 5009
rect 2244 4905 2278 4939
rect 2244 4837 2278 4871
rect 2328 4905 2362 4939
rect 2328 4837 2362 4871
rect 2412 4975 2446 5009
rect 2412 4905 2446 4939
rect 2412 4837 2446 4871
rect 2496 4905 2530 4939
rect 2496 4837 2530 4871
rect 2580 4975 2614 5009
rect 2580 4905 2614 4939
rect 2580 4837 2614 4871
rect 2664 4905 2698 4939
rect 2664 4837 2698 4871
rect 2748 4975 2782 5009
rect 2748 4905 2782 4939
rect 2748 4837 2782 4871
rect 2832 4905 2866 4939
rect 2832 4837 2866 4871
rect 2916 4975 2950 5009
rect 2916 4905 2950 4939
rect 2916 4837 2950 4871
rect 3000 4905 3034 4939
rect 3000 4837 3034 4871
rect 3084 4975 3118 5009
rect 3084 4905 3118 4939
rect 3084 4837 3118 4871
rect 3168 4905 3202 4939
rect 3168 4837 3202 4871
rect 3252 4975 3286 5009
rect 3252 4905 3286 4939
rect 3252 4837 3286 4871
rect 3336 4905 3370 4939
rect 3336 4837 3370 4871
rect 3420 4975 3454 5009
rect 3420 4905 3454 4939
rect 3420 4837 3454 4871
rect 3504 4905 3538 4939
rect 3504 4837 3538 4871
rect 4042 4973 4076 5007
rect 4042 4903 4076 4937
rect 4042 4835 4076 4869
rect 4126 4973 4160 5007
rect 4126 4903 4160 4937
rect 4126 4835 4160 4869
rect 4210 4903 4244 4937
rect 4210 4835 4244 4869
rect 4294 4973 4328 5007
rect 4294 4903 4328 4937
rect 4294 4835 4328 4869
rect 4378 4903 4412 4937
rect 4378 4835 4412 4869
rect 4462 4973 4496 5007
rect 4462 4903 4496 4937
rect 4462 4835 4496 4869
rect 4546 4903 4580 4937
rect 4546 4835 4580 4869
rect 4630 4973 4664 5007
rect 4630 4903 4664 4937
rect 4630 4835 4664 4869
rect 4714 4903 4748 4937
rect 4714 4835 4748 4869
rect 4798 4973 4832 5007
rect 4798 4903 4832 4937
rect 4798 4835 4832 4869
rect 4882 4903 4916 4937
rect 4882 4835 4916 4869
rect 4966 4973 5000 5007
rect 4966 4903 5000 4937
rect 4966 4835 5000 4869
rect 5050 4903 5084 4937
rect 5050 4835 5084 4869
rect 5134 4973 5168 5007
rect 5134 4903 5168 4937
rect 5134 4835 5168 4869
rect 5218 4903 5252 4937
rect 5218 4835 5252 4869
rect 5302 4973 5336 5007
rect 5302 4903 5336 4937
rect 5302 4835 5336 4869
rect 5386 4903 5420 4937
rect 5386 4835 5420 4869
rect 17258 4975 17292 5009
rect 17258 4905 17292 4939
rect 17258 4837 17292 4871
rect 17342 4975 17376 5009
rect 17342 4905 17376 4939
rect 17342 4837 17376 4871
rect 17426 4905 17460 4939
rect 17426 4837 17460 4871
rect 17510 4975 17544 5009
rect 17510 4905 17544 4939
rect 17510 4837 17544 4871
rect 17594 4905 17628 4939
rect 17594 4837 17628 4871
rect 17678 4975 17712 5009
rect 17678 4905 17712 4939
rect 17678 4837 17712 4871
rect 17762 4905 17796 4939
rect 17762 4837 17796 4871
rect 17846 4975 17880 5009
rect 17846 4905 17880 4939
rect 17846 4837 17880 4871
rect 17930 4905 17964 4939
rect 17930 4837 17964 4871
rect 18014 4975 18048 5009
rect 18014 4905 18048 4939
rect 18014 4837 18048 4871
rect 18098 4905 18132 4939
rect 18098 4837 18132 4871
rect 18182 4975 18216 5009
rect 18182 4905 18216 4939
rect 18182 4837 18216 4871
rect 18266 4905 18300 4939
rect 18266 4837 18300 4871
rect 18350 4975 18384 5009
rect 18350 4905 18384 4939
rect 18350 4837 18384 4871
rect 18434 4905 18468 4939
rect 18434 4837 18468 4871
rect 18518 4975 18552 5009
rect 18518 4905 18552 4939
rect 18518 4837 18552 4871
rect 18602 4905 18636 4939
rect 18602 4837 18636 4871
rect 19140 4973 19174 5007
rect 19140 4903 19174 4937
rect 19140 4835 19174 4869
rect 19224 4973 19258 5007
rect 19224 4903 19258 4937
rect 19224 4835 19258 4869
rect 19308 4903 19342 4937
rect 19308 4835 19342 4869
rect 19392 4973 19426 5007
rect 19392 4903 19426 4937
rect 19392 4835 19426 4869
rect 19476 4903 19510 4937
rect 19476 4835 19510 4869
rect 19560 4973 19594 5007
rect 19560 4903 19594 4937
rect 19560 4835 19594 4869
rect 19644 4903 19678 4937
rect 19644 4835 19678 4869
rect 19728 4973 19762 5007
rect 19728 4903 19762 4937
rect 19728 4835 19762 4869
rect 19812 4903 19846 4937
rect 19812 4835 19846 4869
rect 19896 4973 19930 5007
rect 19896 4903 19930 4937
rect 19896 4835 19930 4869
rect 19980 4903 20014 4937
rect 19980 4835 20014 4869
rect 20064 4973 20098 5007
rect 20064 4903 20098 4937
rect 20064 4835 20098 4869
rect 20148 4903 20182 4937
rect 20148 4835 20182 4869
rect 20232 4973 20266 5007
rect 20232 4903 20266 4937
rect 20232 4835 20266 4869
rect 20316 4903 20350 4937
rect 20316 4835 20350 4869
rect 20400 4973 20434 5007
rect 20400 4903 20434 4937
rect 20400 4835 20434 4869
rect 20484 4903 20518 4937
rect 20484 4835 20518 4869
rect -3299 4605 -3265 4639
rect -3299 4537 -3265 4571
rect -3299 4469 -3265 4503
rect -3143 4605 -3109 4639
rect -2485 4605 -2451 4639
rect -3143 4537 -3109 4571
rect -2485 4537 -2451 4571
rect -3143 4469 -3109 4503
rect -2946 4437 -2912 4471
rect -2946 4369 -2912 4403
rect -2946 4301 -2912 4335
rect -2850 4437 -2816 4471
rect -2850 4369 -2816 4403
rect -2850 4301 -2816 4335
rect -2754 4437 -2720 4471
rect -2485 4469 -2451 4503
rect -2329 4605 -2295 4639
rect -2329 4537 -2295 4571
rect -2329 4469 -2295 4503
rect -1411 4605 -1377 4639
rect -1411 4537 -1377 4571
rect -1411 4469 -1377 4503
rect -1255 4605 -1221 4639
rect -597 4605 -563 4639
rect -1255 4537 -1221 4571
rect -597 4537 -563 4571
rect -1255 4469 -1221 4503
rect -2754 4369 -2720 4403
rect -2754 4301 -2720 4335
rect -1058 4437 -1024 4471
rect -1058 4369 -1024 4403
rect -1058 4301 -1024 4335
rect -962 4437 -928 4471
rect -962 4369 -928 4403
rect -962 4301 -928 4335
rect -866 4437 -832 4471
rect -597 4469 -563 4503
rect -441 4605 -407 4639
rect -441 4537 -407 4571
rect -441 4469 -407 4503
rect 477 4605 511 4639
rect 477 4537 511 4571
rect 477 4469 511 4503
rect 633 4605 667 4639
rect 1291 4605 1325 4639
rect 633 4537 667 4571
rect 1291 4537 1325 4571
rect 633 4469 667 4503
rect -866 4369 -832 4403
rect -866 4301 -832 4335
rect 830 4437 864 4471
rect 830 4369 864 4403
rect 830 4301 864 4335
rect 926 4437 960 4471
rect 926 4369 960 4403
rect 926 4301 960 4335
rect 1022 4437 1056 4471
rect 1291 4469 1325 4503
rect 1447 4605 1481 4639
rect 1447 4537 1481 4571
rect 1447 4469 1481 4503
rect 2365 4605 2399 4639
rect 2365 4537 2399 4571
rect 2365 4469 2399 4503
rect 2521 4605 2555 4639
rect 3179 4605 3213 4639
rect 2521 4537 2555 4571
rect 3179 4537 3213 4571
rect 2521 4469 2555 4503
rect 1022 4369 1056 4403
rect 1022 4301 1056 4335
rect 2718 4437 2752 4471
rect 2718 4369 2752 4403
rect 2718 4301 2752 4335
rect 2814 4437 2848 4471
rect 2814 4369 2848 4403
rect 2814 4301 2848 4335
rect 2910 4437 2944 4471
rect 3179 4469 3213 4503
rect 3335 4605 3369 4639
rect 3335 4537 3369 4571
rect 3335 4469 3369 4503
rect 4253 4605 4287 4639
rect 4253 4537 4287 4571
rect 4253 4469 4287 4503
rect 4409 4605 4443 4639
rect 5067 4605 5101 4639
rect 4409 4537 4443 4571
rect 5067 4537 5101 4571
rect 4409 4469 4443 4503
rect 2910 4369 2944 4403
rect 2910 4301 2944 4335
rect 4606 4437 4640 4471
rect 4606 4369 4640 4403
rect 4606 4301 4640 4335
rect 4702 4437 4736 4471
rect 4702 4369 4736 4403
rect 4702 4301 4736 4335
rect 4798 4437 4832 4471
rect 5067 4469 5101 4503
rect 5223 4605 5257 4639
rect 5223 4537 5257 4571
rect 5223 4469 5257 4503
rect 6141 4605 6175 4639
rect 6141 4537 6175 4571
rect 6141 4469 6175 4503
rect 6297 4605 6331 4639
rect 6955 4605 6989 4639
rect 6297 4537 6331 4571
rect 6955 4537 6989 4571
rect 6297 4469 6331 4503
rect 4798 4369 4832 4403
rect 4798 4301 4832 4335
rect 6494 4437 6528 4471
rect 6494 4369 6528 4403
rect 6494 4301 6528 4335
rect 6590 4437 6624 4471
rect 6590 4369 6624 4403
rect 6590 4301 6624 4335
rect 6686 4437 6720 4471
rect 6955 4469 6989 4503
rect 7111 4605 7145 4639
rect 7111 4537 7145 4571
rect 7111 4469 7145 4503
rect 8029 4605 8063 4639
rect 8029 4537 8063 4571
rect 8029 4469 8063 4503
rect 8185 4605 8219 4639
rect 8843 4605 8877 4639
rect 8185 4537 8219 4571
rect 8843 4537 8877 4571
rect 8185 4469 8219 4503
rect 6686 4369 6720 4403
rect 6686 4301 6720 4335
rect 8382 4437 8416 4471
rect 8382 4369 8416 4403
rect 8382 4301 8416 4335
rect 8478 4437 8512 4471
rect 8478 4369 8512 4403
rect 8478 4301 8512 4335
rect 8574 4437 8608 4471
rect 8843 4469 8877 4503
rect 8999 4605 9033 4639
rect 8999 4537 9033 4571
rect 8999 4469 9033 4503
rect 9917 4605 9951 4639
rect 9917 4537 9951 4571
rect 9917 4469 9951 4503
rect 10073 4605 10107 4639
rect 10731 4605 10765 4639
rect 10073 4537 10107 4571
rect 10731 4537 10765 4571
rect 10073 4469 10107 4503
rect 8574 4369 8608 4403
rect 8574 4301 8608 4335
rect 10270 4437 10304 4471
rect 10270 4369 10304 4403
rect 10270 4301 10304 4335
rect 10366 4437 10400 4471
rect 10366 4369 10400 4403
rect 10366 4301 10400 4335
rect 10462 4437 10496 4471
rect 10731 4469 10765 4503
rect 10887 4605 10921 4639
rect 10887 4537 10921 4571
rect 10887 4469 10921 4503
rect 11799 4605 11833 4639
rect 11799 4537 11833 4571
rect 11799 4469 11833 4503
rect 11955 4605 11989 4639
rect 12613 4605 12647 4639
rect 11955 4537 11989 4571
rect 12613 4537 12647 4571
rect 11955 4469 11989 4503
rect 10462 4369 10496 4403
rect 10462 4301 10496 4335
rect 12152 4437 12186 4471
rect 12152 4369 12186 4403
rect 12152 4301 12186 4335
rect 12248 4437 12282 4471
rect 12248 4369 12282 4403
rect 12248 4301 12282 4335
rect 12344 4437 12378 4471
rect 12613 4469 12647 4503
rect 12769 4605 12803 4639
rect 12769 4537 12803 4571
rect 12769 4469 12803 4503
rect 13687 4605 13721 4639
rect 13687 4537 13721 4571
rect 13687 4469 13721 4503
rect 13843 4605 13877 4639
rect 14501 4605 14535 4639
rect 13843 4537 13877 4571
rect 14501 4537 14535 4571
rect 13843 4469 13877 4503
rect 12344 4369 12378 4403
rect 12344 4301 12378 4335
rect 14040 4437 14074 4471
rect 14040 4369 14074 4403
rect 14040 4301 14074 4335
rect 14136 4437 14170 4471
rect 14136 4369 14170 4403
rect 14136 4301 14170 4335
rect 14232 4437 14266 4471
rect 14501 4469 14535 4503
rect 14657 4605 14691 4639
rect 14657 4537 14691 4571
rect 14657 4469 14691 4503
rect 15575 4605 15609 4639
rect 15575 4537 15609 4571
rect 15575 4469 15609 4503
rect 15731 4605 15765 4639
rect 16389 4605 16423 4639
rect 15731 4537 15765 4571
rect 16389 4537 16423 4571
rect 15731 4469 15765 4503
rect 14232 4369 14266 4403
rect 14232 4301 14266 4335
rect 15928 4437 15962 4471
rect 15928 4369 15962 4403
rect 15928 4301 15962 4335
rect 16024 4437 16058 4471
rect 16024 4369 16058 4403
rect 16024 4301 16058 4335
rect 16120 4437 16154 4471
rect 16389 4469 16423 4503
rect 16545 4605 16579 4639
rect 16545 4537 16579 4571
rect 16545 4469 16579 4503
rect 17463 4605 17497 4639
rect 17463 4537 17497 4571
rect 17463 4469 17497 4503
rect 17619 4605 17653 4639
rect 18277 4605 18311 4639
rect 17619 4537 17653 4571
rect 18277 4537 18311 4571
rect 17619 4469 17653 4503
rect 16120 4369 16154 4403
rect 16120 4301 16154 4335
rect 17816 4437 17850 4471
rect 17816 4369 17850 4403
rect 17816 4301 17850 4335
rect 17912 4437 17946 4471
rect 17912 4369 17946 4403
rect 17912 4301 17946 4335
rect 18008 4437 18042 4471
rect 18277 4469 18311 4503
rect 18433 4605 18467 4639
rect 18433 4537 18467 4571
rect 18433 4469 18467 4503
rect 19351 4605 19385 4639
rect 19351 4537 19385 4571
rect 19351 4469 19385 4503
rect 19507 4605 19541 4639
rect 20165 4605 20199 4639
rect 19507 4537 19541 4571
rect 20165 4537 20199 4571
rect 19507 4469 19541 4503
rect 18008 4369 18042 4403
rect 18008 4301 18042 4335
rect 19704 4437 19738 4471
rect 19704 4369 19738 4403
rect 19704 4301 19738 4335
rect 19800 4437 19834 4471
rect 19800 4369 19834 4403
rect 19800 4301 19834 4335
rect 19896 4437 19930 4471
rect 20165 4469 20199 4503
rect 20321 4605 20355 4639
rect 20321 4537 20355 4571
rect 20321 4469 20355 4503
rect 21239 4605 21273 4639
rect 21239 4537 21273 4571
rect 21239 4469 21273 4503
rect 21395 4605 21429 4639
rect 22053 4605 22087 4639
rect 21395 4537 21429 4571
rect 22053 4537 22087 4571
rect 21395 4469 21429 4503
rect 19896 4369 19930 4403
rect 19896 4301 19930 4335
rect 21592 4437 21626 4471
rect 21592 4369 21626 4403
rect 21592 4301 21626 4335
rect 21688 4437 21722 4471
rect 21688 4369 21722 4403
rect 21688 4301 21722 4335
rect 21784 4437 21818 4471
rect 22053 4469 22087 4503
rect 22209 4605 22243 4639
rect 22209 4537 22243 4571
rect 22209 4469 22243 4503
rect 23127 4605 23161 4639
rect 23127 4537 23161 4571
rect 23127 4469 23161 4503
rect 23283 4605 23317 4639
rect 23941 4605 23975 4639
rect 23283 4537 23317 4571
rect 23941 4537 23975 4571
rect 23283 4469 23317 4503
rect 21784 4369 21818 4403
rect 21784 4301 21818 4335
rect 23480 4437 23514 4471
rect 23480 4369 23514 4403
rect 23480 4301 23514 4335
rect 23576 4437 23610 4471
rect 23576 4369 23610 4403
rect 23576 4301 23610 4335
rect 23672 4437 23706 4471
rect 23941 4469 23975 4503
rect 24097 4605 24131 4639
rect 24097 4537 24131 4571
rect 24097 4469 24131 4503
rect 25015 4605 25049 4639
rect 25015 4537 25049 4571
rect 25015 4469 25049 4503
rect 25171 4605 25205 4639
rect 25829 4605 25863 4639
rect 25171 4537 25205 4571
rect 25829 4537 25863 4571
rect 25171 4469 25205 4503
rect 23672 4369 23706 4403
rect 23672 4301 23706 4335
rect 25368 4437 25402 4471
rect 25368 4369 25402 4403
rect 25368 4301 25402 4335
rect 25464 4437 25498 4471
rect 25464 4369 25498 4403
rect 25464 4301 25498 4335
rect 25560 4437 25594 4471
rect 25829 4469 25863 4503
rect 25985 4605 26019 4639
rect 25985 4537 26019 4571
rect 25985 4469 26019 4503
rect 25560 4369 25594 4403
rect 25560 4301 25594 4335
rect -3436 3551 -3402 3585
rect -3436 3483 -3402 3517
rect -3436 3415 -3402 3449
rect -3352 3551 -3318 3585
rect -3352 3483 -3318 3517
rect -3352 3415 -3318 3449
rect -3164 3541 -3130 3575
rect -3164 3473 -3130 3507
rect -3164 3405 -3130 3439
rect -3076 3541 -3042 3575
rect -2518 3541 -2484 3575
rect -3076 3473 -3042 3507
rect -3076 3405 -3042 3439
rect -2518 3473 -2484 3507
rect -2948 3381 -2914 3415
rect -2948 3313 -2914 3347
rect -2948 3245 -2914 3279
rect -2852 3381 -2818 3415
rect -2852 3313 -2818 3347
rect -2852 3245 -2818 3279
rect -2756 3381 -2722 3415
rect -2518 3405 -2484 3439
rect -2430 3541 -2396 3575
rect -2430 3473 -2396 3507
rect -2430 3405 -2396 3439
rect -2240 3559 -2206 3593
rect -2240 3491 -2206 3525
rect -2240 3423 -2206 3457
rect -2156 3559 -2122 3593
rect -2156 3491 -2122 3525
rect -2156 3423 -2122 3457
rect -1935 3549 -1901 3583
rect -1935 3481 -1901 3515
rect -1849 3549 -1815 3583
rect -1849 3481 -1815 3515
rect -1763 3549 -1729 3583
rect -1763 3468 -1729 3502
rect -1548 3551 -1514 3585
rect -1548 3483 -1514 3517
rect -2756 3313 -2722 3347
rect -1548 3415 -1514 3449
rect -1464 3551 -1430 3585
rect -1464 3483 -1430 3517
rect -1464 3415 -1430 3449
rect -1276 3541 -1242 3575
rect -1276 3473 -1242 3507
rect -1276 3405 -1242 3439
rect -1188 3541 -1154 3575
rect -630 3541 -596 3575
rect -1188 3473 -1154 3507
rect -1188 3405 -1154 3439
rect -630 3473 -596 3507
rect -1060 3381 -1026 3415
rect -2756 3245 -2722 3279
rect -1060 3313 -1026 3347
rect -1060 3245 -1026 3279
rect -964 3381 -930 3415
rect -964 3313 -930 3347
rect -964 3245 -930 3279
rect -868 3381 -834 3415
rect -630 3405 -596 3439
rect -542 3541 -508 3575
rect -542 3473 -508 3507
rect -542 3405 -508 3439
rect -352 3559 -318 3593
rect -352 3491 -318 3525
rect -352 3423 -318 3457
rect -268 3559 -234 3593
rect -268 3491 -234 3525
rect -268 3423 -234 3457
rect -47 3549 -13 3583
rect -47 3481 -13 3515
rect 39 3549 73 3583
rect 39 3481 73 3515
rect 125 3549 159 3583
rect 125 3468 159 3502
rect 340 3551 374 3585
rect 340 3483 374 3517
rect -868 3313 -834 3347
rect 340 3415 374 3449
rect 424 3551 458 3585
rect 424 3483 458 3517
rect 424 3415 458 3449
rect 612 3541 646 3575
rect 612 3473 646 3507
rect 612 3405 646 3439
rect 700 3541 734 3575
rect 1258 3541 1292 3575
rect 700 3473 734 3507
rect 700 3405 734 3439
rect 1258 3473 1292 3507
rect 828 3381 862 3415
rect -868 3245 -834 3279
rect 828 3313 862 3347
rect 828 3245 862 3279
rect 924 3381 958 3415
rect 924 3313 958 3347
rect 924 3245 958 3279
rect 1020 3381 1054 3415
rect 1258 3405 1292 3439
rect 1346 3541 1380 3575
rect 1346 3473 1380 3507
rect 1346 3405 1380 3439
rect 1536 3559 1570 3593
rect 1536 3491 1570 3525
rect 1536 3423 1570 3457
rect 1620 3559 1654 3593
rect 1620 3491 1654 3525
rect 1620 3423 1654 3457
rect 1841 3549 1875 3583
rect 1841 3481 1875 3515
rect 1927 3549 1961 3583
rect 1927 3481 1961 3515
rect 2013 3549 2047 3583
rect 2013 3468 2047 3502
rect 2228 3551 2262 3585
rect 2228 3483 2262 3517
rect 1020 3313 1054 3347
rect 2228 3415 2262 3449
rect 2312 3551 2346 3585
rect 2312 3483 2346 3517
rect 2312 3415 2346 3449
rect 2500 3541 2534 3575
rect 2500 3473 2534 3507
rect 2500 3405 2534 3439
rect 2588 3541 2622 3575
rect 3146 3541 3180 3575
rect 2588 3473 2622 3507
rect 2588 3405 2622 3439
rect 3146 3473 3180 3507
rect 2716 3381 2750 3415
rect 1020 3245 1054 3279
rect 2716 3313 2750 3347
rect 2716 3245 2750 3279
rect 2812 3381 2846 3415
rect 2812 3313 2846 3347
rect 2812 3245 2846 3279
rect 2908 3381 2942 3415
rect 3146 3405 3180 3439
rect 3234 3541 3268 3575
rect 3234 3473 3268 3507
rect 3234 3405 3268 3439
rect 3424 3559 3458 3593
rect 3424 3491 3458 3525
rect 3424 3423 3458 3457
rect 3508 3559 3542 3593
rect 3508 3491 3542 3525
rect 3508 3423 3542 3457
rect 3729 3549 3763 3583
rect 3729 3481 3763 3515
rect 3815 3549 3849 3583
rect 3815 3481 3849 3515
rect 3901 3549 3935 3583
rect 3901 3468 3935 3502
rect 4116 3551 4150 3585
rect 4116 3483 4150 3517
rect 2908 3313 2942 3347
rect 4116 3415 4150 3449
rect 4200 3551 4234 3585
rect 4200 3483 4234 3517
rect 4200 3415 4234 3449
rect 4388 3541 4422 3575
rect 4388 3473 4422 3507
rect 4388 3405 4422 3439
rect 4476 3541 4510 3575
rect 5034 3541 5068 3575
rect 4476 3473 4510 3507
rect 4476 3405 4510 3439
rect 5034 3473 5068 3507
rect 4604 3381 4638 3415
rect 2908 3245 2942 3279
rect 4604 3313 4638 3347
rect 4604 3245 4638 3279
rect 4700 3381 4734 3415
rect 4700 3313 4734 3347
rect 4700 3245 4734 3279
rect 4796 3381 4830 3415
rect 5034 3405 5068 3439
rect 5122 3541 5156 3575
rect 5122 3473 5156 3507
rect 5122 3405 5156 3439
rect 5312 3559 5346 3593
rect 5312 3491 5346 3525
rect 5312 3423 5346 3457
rect 5396 3559 5430 3593
rect 5396 3491 5430 3525
rect 5396 3423 5430 3457
rect 5617 3549 5651 3583
rect 5617 3481 5651 3515
rect 5703 3549 5737 3583
rect 5703 3481 5737 3515
rect 5789 3549 5823 3583
rect 5789 3468 5823 3502
rect 6004 3551 6038 3585
rect 6004 3483 6038 3517
rect 4796 3313 4830 3347
rect 6004 3415 6038 3449
rect 6088 3551 6122 3585
rect 6088 3483 6122 3517
rect 6088 3415 6122 3449
rect 6276 3541 6310 3575
rect 6276 3473 6310 3507
rect 6276 3405 6310 3439
rect 6364 3541 6398 3575
rect 6922 3541 6956 3575
rect 6364 3473 6398 3507
rect 6364 3405 6398 3439
rect 6922 3473 6956 3507
rect 6492 3381 6526 3415
rect 4796 3245 4830 3279
rect 6492 3313 6526 3347
rect 6492 3245 6526 3279
rect 6588 3381 6622 3415
rect 6588 3313 6622 3347
rect 6588 3245 6622 3279
rect 6684 3381 6718 3415
rect 6922 3405 6956 3439
rect 7010 3541 7044 3575
rect 7010 3473 7044 3507
rect 7010 3405 7044 3439
rect 7200 3559 7234 3593
rect 7200 3491 7234 3525
rect 7200 3423 7234 3457
rect 7284 3559 7318 3593
rect 7284 3491 7318 3525
rect 7284 3423 7318 3457
rect 7505 3549 7539 3583
rect 7505 3481 7539 3515
rect 7591 3549 7625 3583
rect 7591 3481 7625 3515
rect 7677 3549 7711 3583
rect 7677 3468 7711 3502
rect 7892 3551 7926 3585
rect 7892 3483 7926 3517
rect 6684 3313 6718 3347
rect 7892 3415 7926 3449
rect 7976 3551 8010 3585
rect 7976 3483 8010 3517
rect 7976 3415 8010 3449
rect 8164 3541 8198 3575
rect 8164 3473 8198 3507
rect 8164 3405 8198 3439
rect 8252 3541 8286 3575
rect 8810 3541 8844 3575
rect 8252 3473 8286 3507
rect 8252 3405 8286 3439
rect 8810 3473 8844 3507
rect 8380 3381 8414 3415
rect 6684 3245 6718 3279
rect 8380 3313 8414 3347
rect 8380 3245 8414 3279
rect 8476 3381 8510 3415
rect 8476 3313 8510 3347
rect 8476 3245 8510 3279
rect 8572 3381 8606 3415
rect 8810 3405 8844 3439
rect 8898 3541 8932 3575
rect 8898 3473 8932 3507
rect 8898 3405 8932 3439
rect 9088 3559 9122 3593
rect 9088 3491 9122 3525
rect 9088 3423 9122 3457
rect 9172 3559 9206 3593
rect 9172 3491 9206 3525
rect 9172 3423 9206 3457
rect 9393 3549 9427 3583
rect 9393 3481 9427 3515
rect 9479 3549 9513 3583
rect 9479 3481 9513 3515
rect 9565 3549 9599 3583
rect 9565 3468 9599 3502
rect 9780 3551 9814 3585
rect 9780 3483 9814 3517
rect 8572 3313 8606 3347
rect 9780 3415 9814 3449
rect 9864 3551 9898 3585
rect 9864 3483 9898 3517
rect 9864 3415 9898 3449
rect 10052 3541 10086 3575
rect 10052 3473 10086 3507
rect 10052 3405 10086 3439
rect 10140 3541 10174 3575
rect 10698 3541 10732 3575
rect 10140 3473 10174 3507
rect 10140 3405 10174 3439
rect 10698 3473 10732 3507
rect 10268 3381 10302 3415
rect 8572 3245 8606 3279
rect 10268 3313 10302 3347
rect 10268 3245 10302 3279
rect 10364 3381 10398 3415
rect 10364 3313 10398 3347
rect 10364 3245 10398 3279
rect 10460 3381 10494 3415
rect 10698 3405 10732 3439
rect 10786 3541 10820 3575
rect 10786 3473 10820 3507
rect 10786 3405 10820 3439
rect 10976 3559 11010 3593
rect 10976 3491 11010 3525
rect 10976 3423 11010 3457
rect 11060 3559 11094 3593
rect 11060 3491 11094 3525
rect 11060 3423 11094 3457
rect 11281 3549 11315 3583
rect 11281 3481 11315 3515
rect 11367 3549 11401 3583
rect 11367 3481 11401 3515
rect 11453 3549 11487 3583
rect 11453 3468 11487 3502
rect 11662 3551 11696 3585
rect 11662 3483 11696 3517
rect 10460 3313 10494 3347
rect 11662 3415 11696 3449
rect 11746 3551 11780 3585
rect 11746 3483 11780 3517
rect 11746 3415 11780 3449
rect 11934 3541 11968 3575
rect 11934 3473 11968 3507
rect 11934 3405 11968 3439
rect 12022 3541 12056 3575
rect 12580 3541 12614 3575
rect 12022 3473 12056 3507
rect 12022 3405 12056 3439
rect 12580 3473 12614 3507
rect 12150 3381 12184 3415
rect 10460 3245 10494 3279
rect 12150 3313 12184 3347
rect 12150 3245 12184 3279
rect 12246 3381 12280 3415
rect 12246 3313 12280 3347
rect 12246 3245 12280 3279
rect 12342 3381 12376 3415
rect 12580 3405 12614 3439
rect 12668 3541 12702 3575
rect 12668 3473 12702 3507
rect 12668 3405 12702 3439
rect 12858 3559 12892 3593
rect 12858 3491 12892 3525
rect 12858 3423 12892 3457
rect 12942 3559 12976 3593
rect 12942 3491 12976 3525
rect 12942 3423 12976 3457
rect 13163 3549 13197 3583
rect 13163 3481 13197 3515
rect 13249 3549 13283 3583
rect 13249 3481 13283 3515
rect 13335 3549 13369 3583
rect 13335 3468 13369 3502
rect 13550 3551 13584 3585
rect 13550 3483 13584 3517
rect 12342 3313 12376 3347
rect 13550 3415 13584 3449
rect 13634 3551 13668 3585
rect 13634 3483 13668 3517
rect 13634 3415 13668 3449
rect 13822 3541 13856 3575
rect 13822 3473 13856 3507
rect 13822 3405 13856 3439
rect 13910 3541 13944 3575
rect 14468 3541 14502 3575
rect 13910 3473 13944 3507
rect 13910 3405 13944 3439
rect 14468 3473 14502 3507
rect 14038 3381 14072 3415
rect 12342 3245 12376 3279
rect 14038 3313 14072 3347
rect 14038 3245 14072 3279
rect 14134 3381 14168 3415
rect 14134 3313 14168 3347
rect 14134 3245 14168 3279
rect 14230 3381 14264 3415
rect 14468 3405 14502 3439
rect 14556 3541 14590 3575
rect 14556 3473 14590 3507
rect 14556 3405 14590 3439
rect 14746 3559 14780 3593
rect 14746 3491 14780 3525
rect 14746 3423 14780 3457
rect 14830 3559 14864 3593
rect 14830 3491 14864 3525
rect 14830 3423 14864 3457
rect 15051 3549 15085 3583
rect 15051 3481 15085 3515
rect 15137 3549 15171 3583
rect 15137 3481 15171 3515
rect 15223 3549 15257 3583
rect 15223 3468 15257 3502
rect 15438 3551 15472 3585
rect 15438 3483 15472 3517
rect 14230 3313 14264 3347
rect 15438 3415 15472 3449
rect 15522 3551 15556 3585
rect 15522 3483 15556 3517
rect 15522 3415 15556 3449
rect 15710 3541 15744 3575
rect 15710 3473 15744 3507
rect 15710 3405 15744 3439
rect 15798 3541 15832 3575
rect 16356 3541 16390 3575
rect 15798 3473 15832 3507
rect 15798 3405 15832 3439
rect 16356 3473 16390 3507
rect 15926 3381 15960 3415
rect 14230 3245 14264 3279
rect 15926 3313 15960 3347
rect 15926 3245 15960 3279
rect 16022 3381 16056 3415
rect 16022 3313 16056 3347
rect 16022 3245 16056 3279
rect 16118 3381 16152 3415
rect 16356 3405 16390 3439
rect 16444 3541 16478 3575
rect 16444 3473 16478 3507
rect 16444 3405 16478 3439
rect 16634 3559 16668 3593
rect 16634 3491 16668 3525
rect 16634 3423 16668 3457
rect 16718 3559 16752 3593
rect 16718 3491 16752 3525
rect 16718 3423 16752 3457
rect 16939 3549 16973 3583
rect 16939 3481 16973 3515
rect 17025 3549 17059 3583
rect 17025 3481 17059 3515
rect 17111 3549 17145 3583
rect 17111 3468 17145 3502
rect 17326 3551 17360 3585
rect 17326 3483 17360 3517
rect 16118 3313 16152 3347
rect 17326 3415 17360 3449
rect 17410 3551 17444 3585
rect 17410 3483 17444 3517
rect 17410 3415 17444 3449
rect 17598 3541 17632 3575
rect 17598 3473 17632 3507
rect 17598 3405 17632 3439
rect 17686 3541 17720 3575
rect 18244 3541 18278 3575
rect 17686 3473 17720 3507
rect 17686 3405 17720 3439
rect 18244 3473 18278 3507
rect 17814 3381 17848 3415
rect 16118 3245 16152 3279
rect 17814 3313 17848 3347
rect 17814 3245 17848 3279
rect 17910 3381 17944 3415
rect 17910 3313 17944 3347
rect 17910 3245 17944 3279
rect 18006 3381 18040 3415
rect 18244 3405 18278 3439
rect 18332 3541 18366 3575
rect 18332 3473 18366 3507
rect 18332 3405 18366 3439
rect 18522 3559 18556 3593
rect 18522 3491 18556 3525
rect 18522 3423 18556 3457
rect 18606 3559 18640 3593
rect 18606 3491 18640 3525
rect 18606 3423 18640 3457
rect 18827 3549 18861 3583
rect 18827 3481 18861 3515
rect 18913 3549 18947 3583
rect 18913 3481 18947 3515
rect 18999 3549 19033 3583
rect 18999 3468 19033 3502
rect 19214 3551 19248 3585
rect 19214 3483 19248 3517
rect 18006 3313 18040 3347
rect 19214 3415 19248 3449
rect 19298 3551 19332 3585
rect 19298 3483 19332 3517
rect 19298 3415 19332 3449
rect 19486 3541 19520 3575
rect 19486 3473 19520 3507
rect 19486 3405 19520 3439
rect 19574 3541 19608 3575
rect 20132 3541 20166 3575
rect 19574 3473 19608 3507
rect 19574 3405 19608 3439
rect 20132 3473 20166 3507
rect 19702 3381 19736 3415
rect 18006 3245 18040 3279
rect 19702 3313 19736 3347
rect 19702 3245 19736 3279
rect 19798 3381 19832 3415
rect 19798 3313 19832 3347
rect 19798 3245 19832 3279
rect 19894 3381 19928 3415
rect 20132 3405 20166 3439
rect 20220 3541 20254 3575
rect 20220 3473 20254 3507
rect 20220 3405 20254 3439
rect 20410 3559 20444 3593
rect 20410 3491 20444 3525
rect 20410 3423 20444 3457
rect 20494 3559 20528 3593
rect 20494 3491 20528 3525
rect 20494 3423 20528 3457
rect 20715 3549 20749 3583
rect 20715 3481 20749 3515
rect 20801 3549 20835 3583
rect 20801 3481 20835 3515
rect 20887 3549 20921 3583
rect 20887 3468 20921 3502
rect 21102 3551 21136 3585
rect 21102 3483 21136 3517
rect 19894 3313 19928 3347
rect 21102 3415 21136 3449
rect 21186 3551 21220 3585
rect 21186 3483 21220 3517
rect 21186 3415 21220 3449
rect 21374 3541 21408 3575
rect 21374 3473 21408 3507
rect 21374 3405 21408 3439
rect 21462 3541 21496 3575
rect 22020 3541 22054 3575
rect 21462 3473 21496 3507
rect 21462 3405 21496 3439
rect 22020 3473 22054 3507
rect 21590 3381 21624 3415
rect 19894 3245 19928 3279
rect 21590 3313 21624 3347
rect 21590 3245 21624 3279
rect 21686 3381 21720 3415
rect 21686 3313 21720 3347
rect 21686 3245 21720 3279
rect 21782 3381 21816 3415
rect 22020 3405 22054 3439
rect 22108 3541 22142 3575
rect 22108 3473 22142 3507
rect 22108 3405 22142 3439
rect 22298 3559 22332 3593
rect 22298 3491 22332 3525
rect 22298 3423 22332 3457
rect 22382 3559 22416 3593
rect 22382 3491 22416 3525
rect 22382 3423 22416 3457
rect 22603 3549 22637 3583
rect 22603 3481 22637 3515
rect 22689 3549 22723 3583
rect 22689 3481 22723 3515
rect 22775 3549 22809 3583
rect 22775 3468 22809 3502
rect 22990 3551 23024 3585
rect 22990 3483 23024 3517
rect 21782 3313 21816 3347
rect 22990 3415 23024 3449
rect 23074 3551 23108 3585
rect 23074 3483 23108 3517
rect 23074 3415 23108 3449
rect 23262 3541 23296 3575
rect 23262 3473 23296 3507
rect 23262 3405 23296 3439
rect 23350 3541 23384 3575
rect 23908 3541 23942 3575
rect 23350 3473 23384 3507
rect 23350 3405 23384 3439
rect 23908 3473 23942 3507
rect 23478 3381 23512 3415
rect 21782 3245 21816 3279
rect 23478 3313 23512 3347
rect 23478 3245 23512 3279
rect 23574 3381 23608 3415
rect 23574 3313 23608 3347
rect 23574 3245 23608 3279
rect 23670 3381 23704 3415
rect 23908 3405 23942 3439
rect 23996 3541 24030 3575
rect 23996 3473 24030 3507
rect 23996 3405 24030 3439
rect 24186 3559 24220 3593
rect 24186 3491 24220 3525
rect 24186 3423 24220 3457
rect 24270 3559 24304 3593
rect 24270 3491 24304 3525
rect 24270 3423 24304 3457
rect 24491 3549 24525 3583
rect 24491 3481 24525 3515
rect 24577 3549 24611 3583
rect 24577 3481 24611 3515
rect 24663 3549 24697 3583
rect 24663 3468 24697 3502
rect 24878 3551 24912 3585
rect 24878 3483 24912 3517
rect 23670 3313 23704 3347
rect 24878 3415 24912 3449
rect 24962 3551 24996 3585
rect 24962 3483 24996 3517
rect 24962 3415 24996 3449
rect 25150 3541 25184 3575
rect 25150 3473 25184 3507
rect 25150 3405 25184 3439
rect 25238 3541 25272 3575
rect 25796 3541 25830 3575
rect 25238 3473 25272 3507
rect 25238 3405 25272 3439
rect 25796 3473 25830 3507
rect 25366 3381 25400 3415
rect 23670 3245 23704 3279
rect 25366 3313 25400 3347
rect 25366 3245 25400 3279
rect 25462 3381 25496 3415
rect 25462 3313 25496 3347
rect 25462 3245 25496 3279
rect 25558 3381 25592 3415
rect 25796 3405 25830 3439
rect 25884 3541 25918 3575
rect 25884 3473 25918 3507
rect 25884 3405 25918 3439
rect 26074 3559 26108 3593
rect 26074 3491 26108 3525
rect 26074 3423 26108 3457
rect 26158 3559 26192 3593
rect 26158 3491 26192 3525
rect 26158 3423 26192 3457
rect 26379 3549 26413 3583
rect 26379 3481 26413 3515
rect 26465 3549 26499 3583
rect 26465 3481 26499 3515
rect 26551 3549 26585 3583
rect 26551 3468 26585 3502
rect 25558 3313 25592 3347
rect 25558 3245 25592 3279
<< psubdiff >>
rect -2898 3814 -2738 3820
rect -2898 3780 -2841 3814
rect -2807 3780 -2738 3814
rect -2898 3772 -2738 3780
rect -1010 3814 -850 3820
rect -1010 3780 -953 3814
rect -919 3780 -850 3814
rect -1010 3772 -850 3780
rect 878 3814 1038 3820
rect 878 3780 935 3814
rect 969 3780 1038 3814
rect 878 3772 1038 3780
rect 2766 3814 2926 3820
rect 2766 3780 2823 3814
rect 2857 3780 2926 3814
rect 2766 3772 2926 3780
rect 4654 3814 4814 3820
rect 4654 3780 4711 3814
rect 4745 3780 4814 3814
rect 4654 3772 4814 3780
rect 6542 3814 6702 3820
rect 6542 3780 6599 3814
rect 6633 3780 6702 3814
rect 6542 3772 6702 3780
rect 8430 3814 8590 3820
rect 8430 3780 8487 3814
rect 8521 3780 8590 3814
rect 8430 3772 8590 3780
rect 10318 3814 10478 3820
rect 10318 3780 10375 3814
rect 10409 3780 10478 3814
rect 10318 3772 10478 3780
rect 12200 3814 12360 3820
rect 12200 3780 12257 3814
rect 12291 3780 12360 3814
rect 12200 3772 12360 3780
rect 14088 3814 14248 3820
rect 14088 3780 14145 3814
rect 14179 3780 14248 3814
rect 14088 3772 14248 3780
rect 15976 3814 16136 3820
rect 15976 3780 16033 3814
rect 16067 3780 16136 3814
rect 15976 3772 16136 3780
rect 17864 3814 18024 3820
rect 17864 3780 17921 3814
rect 17955 3780 18024 3814
rect 17864 3772 18024 3780
rect 19752 3814 19912 3820
rect 19752 3780 19809 3814
rect 19843 3780 19912 3814
rect 19752 3772 19912 3780
rect 21640 3814 21800 3820
rect 21640 3780 21697 3814
rect 21731 3780 21800 3814
rect 21640 3772 21800 3780
rect 23528 3814 23688 3820
rect 23528 3780 23585 3814
rect 23619 3780 23688 3814
rect 23528 3772 23688 3780
rect 25416 3814 25576 3820
rect 25416 3780 25473 3814
rect 25507 3780 25576 3814
rect 25416 3772 25576 3780
rect -2900 2758 -2740 2764
rect -2900 2724 -2843 2758
rect -2809 2724 -2740 2758
rect -2900 2716 -2740 2724
rect -1012 2758 -852 2764
rect -1012 2724 -955 2758
rect -921 2724 -852 2758
rect -1012 2716 -852 2724
rect 876 2758 1036 2764
rect 876 2724 933 2758
rect 967 2724 1036 2758
rect 876 2716 1036 2724
rect 2764 2758 2924 2764
rect 2764 2724 2821 2758
rect 2855 2724 2924 2758
rect 2764 2716 2924 2724
rect 4652 2758 4812 2764
rect 4652 2724 4709 2758
rect 4743 2724 4812 2758
rect 4652 2716 4812 2724
rect 6540 2758 6700 2764
rect 6540 2724 6597 2758
rect 6631 2724 6700 2758
rect 6540 2716 6700 2724
rect 8428 2758 8588 2764
rect 8428 2724 8485 2758
rect 8519 2724 8588 2758
rect 8428 2716 8588 2724
rect 10316 2758 10476 2764
rect 10316 2724 10373 2758
rect 10407 2724 10476 2758
rect 10316 2716 10476 2724
rect 12198 2758 12358 2764
rect 12198 2724 12255 2758
rect 12289 2724 12358 2758
rect 12198 2716 12358 2724
rect 14086 2758 14246 2764
rect 14086 2724 14143 2758
rect 14177 2724 14246 2758
rect 14086 2716 14246 2724
rect 15974 2758 16134 2764
rect 15974 2724 16031 2758
rect 16065 2724 16134 2758
rect 15974 2716 16134 2724
rect 17862 2758 18022 2764
rect 17862 2724 17919 2758
rect 17953 2724 18022 2758
rect 17862 2716 18022 2724
rect 19750 2758 19910 2764
rect 19750 2724 19807 2758
rect 19841 2724 19910 2758
rect 19750 2716 19910 2724
rect 21638 2758 21798 2764
rect 21638 2724 21695 2758
rect 21729 2724 21798 2758
rect 21638 2716 21798 2724
rect 23526 2758 23686 2764
rect 23526 2724 23583 2758
rect 23617 2724 23686 2758
rect 23526 2716 23686 2724
rect 25414 2758 25574 2764
rect 25414 2724 25471 2758
rect 25505 2724 25574 2758
rect 25414 2716 25574 2724
<< nsubdiff >>
rect -2780 4673 -2646 4690
rect -2780 4639 -2752 4673
rect -2718 4639 -2646 4673
rect -892 4673 -758 4690
rect -2780 4620 -2646 4639
rect -892 4639 -864 4673
rect -830 4639 -758 4673
rect 996 4673 1130 4690
rect -892 4620 -758 4639
rect 996 4639 1024 4673
rect 1058 4639 1130 4673
rect 2884 4673 3018 4690
rect 996 4620 1130 4639
rect 2884 4639 2912 4673
rect 2946 4639 3018 4673
rect 4772 4673 4906 4690
rect 2884 4620 3018 4639
rect 4772 4639 4800 4673
rect 4834 4639 4906 4673
rect 6660 4673 6794 4690
rect 4772 4620 4906 4639
rect 6660 4639 6688 4673
rect 6722 4639 6794 4673
rect 8548 4673 8682 4690
rect 6660 4620 6794 4639
rect 8548 4639 8576 4673
rect 8610 4639 8682 4673
rect 10436 4673 10570 4690
rect 8548 4620 8682 4639
rect 10436 4639 10464 4673
rect 10498 4639 10570 4673
rect 12318 4673 12452 4690
rect 10436 4620 10570 4639
rect 12318 4639 12346 4673
rect 12380 4639 12452 4673
rect 14206 4673 14340 4690
rect 12318 4620 12452 4639
rect 14206 4639 14234 4673
rect 14268 4639 14340 4673
rect 16094 4673 16228 4690
rect 14206 4620 14340 4639
rect 16094 4639 16122 4673
rect 16156 4639 16228 4673
rect 17982 4673 18116 4690
rect 16094 4620 16228 4639
rect 17982 4639 18010 4673
rect 18044 4639 18116 4673
rect 19870 4673 20004 4690
rect 17982 4620 18116 4639
rect 19870 4639 19898 4673
rect 19932 4639 20004 4673
rect 21758 4673 21892 4690
rect 19870 4620 20004 4639
rect 21758 4639 21786 4673
rect 21820 4639 21892 4673
rect 23646 4673 23780 4690
rect 21758 4620 21892 4639
rect 23646 4639 23674 4673
rect 23708 4639 23780 4673
rect 25534 4673 25668 4690
rect 23646 4620 23780 4639
rect 25534 4639 25562 4673
rect 25596 4639 25668 4673
rect 25534 4620 25668 4639
rect -2782 3617 -2648 3634
rect -2782 3583 -2754 3617
rect -2720 3583 -2648 3617
rect -2782 3564 -2648 3583
rect -894 3617 -760 3634
rect -894 3583 -866 3617
rect -832 3583 -760 3617
rect -894 3564 -760 3583
rect 994 3617 1128 3634
rect 994 3583 1022 3617
rect 1056 3583 1128 3617
rect 994 3564 1128 3583
rect 2882 3617 3016 3634
rect 2882 3583 2910 3617
rect 2944 3583 3016 3617
rect 2882 3564 3016 3583
rect 4770 3617 4904 3634
rect 4770 3583 4798 3617
rect 4832 3583 4904 3617
rect 4770 3564 4904 3583
rect 6658 3617 6792 3634
rect 6658 3583 6686 3617
rect 6720 3583 6792 3617
rect 6658 3564 6792 3583
rect 8546 3617 8680 3634
rect 8546 3583 8574 3617
rect 8608 3583 8680 3617
rect 8546 3564 8680 3583
rect 10434 3617 10568 3634
rect 10434 3583 10462 3617
rect 10496 3583 10568 3617
rect 10434 3564 10568 3583
rect 12316 3617 12450 3634
rect 12316 3583 12344 3617
rect 12378 3583 12450 3617
rect 12316 3564 12450 3583
rect 14204 3617 14338 3634
rect 14204 3583 14232 3617
rect 14266 3583 14338 3617
rect 14204 3564 14338 3583
rect 16092 3617 16226 3634
rect 16092 3583 16120 3617
rect 16154 3583 16226 3617
rect 16092 3564 16226 3583
rect 17980 3617 18114 3634
rect 17980 3583 18008 3617
rect 18042 3583 18114 3617
rect 17980 3564 18114 3583
rect 19868 3617 20002 3634
rect 19868 3583 19896 3617
rect 19930 3583 20002 3617
rect 19868 3564 20002 3583
rect 21756 3617 21890 3634
rect 21756 3583 21784 3617
rect 21818 3583 21890 3617
rect 21756 3564 21890 3583
rect 23644 3617 23778 3634
rect 23644 3583 23672 3617
rect 23706 3583 23778 3617
rect 23644 3564 23778 3583
rect 25532 3617 25666 3634
rect 25532 3583 25560 3617
rect 25594 3583 25666 3617
rect 25532 3564 25666 3583
<< psubdiffcont >>
rect -2841 3780 -2807 3814
rect -953 3780 -919 3814
rect 935 3780 969 3814
rect 2823 3780 2857 3814
rect 4711 3780 4745 3814
rect 6599 3780 6633 3814
rect 8487 3780 8521 3814
rect 10375 3780 10409 3814
rect 12257 3780 12291 3814
rect 14145 3780 14179 3814
rect 16033 3780 16067 3814
rect 17921 3780 17955 3814
rect 19809 3780 19843 3814
rect 21697 3780 21731 3814
rect 23585 3780 23619 3814
rect 25473 3780 25507 3814
rect -2843 2724 -2809 2758
rect -955 2724 -921 2758
rect 933 2724 967 2758
rect 2821 2724 2855 2758
rect 4709 2724 4743 2758
rect 6597 2724 6631 2758
rect 8485 2724 8519 2758
rect 10373 2724 10407 2758
rect 12255 2724 12289 2758
rect 14143 2724 14177 2758
rect 16031 2724 16065 2758
rect 17919 2724 17953 2758
rect 19807 2724 19841 2758
rect 21695 2724 21729 2758
rect 23583 2724 23617 2758
rect 25471 2724 25505 2758
<< nsubdiffcont >>
rect -2752 4639 -2718 4673
rect -864 4639 -830 4673
rect 1024 4639 1058 4673
rect 2912 4639 2946 4673
rect 4800 4639 4834 4673
rect 6688 4639 6722 4673
rect 8576 4639 8610 4673
rect 10464 4639 10498 4673
rect 12346 4639 12380 4673
rect 14234 4639 14268 4673
rect 16122 4639 16156 4673
rect 18010 4639 18044 4673
rect 19898 4639 19932 4673
rect 21786 4639 21820 4673
rect 23674 4639 23708 4673
rect 25562 4639 25596 4673
rect -2754 3583 -2720 3617
rect -866 3583 -832 3617
rect 1022 3583 1056 3617
rect 2910 3583 2944 3617
rect 4798 3583 4832 3617
rect 6686 3583 6720 3617
rect 8574 3583 8608 3617
rect 10462 3583 10496 3617
rect 12344 3583 12378 3617
rect 14232 3583 14266 3617
rect 16120 3583 16154 3617
rect 18008 3583 18042 3617
rect 19896 3583 19930 3617
rect 21784 3583 21818 3617
rect 23672 3583 23706 3617
rect 25560 3583 25594 3617
<< poly >>
rect 2204 5275 2234 5301
rect 2288 5275 2318 5301
rect 2372 5275 2402 5301
rect 2456 5275 2486 5301
rect 2540 5275 2570 5301
rect 2624 5275 2654 5301
rect 2708 5275 2738 5301
rect 2792 5275 2822 5301
rect 2876 5275 2906 5301
rect 2960 5275 2990 5301
rect 3044 5275 3074 5301
rect 3128 5275 3158 5301
rect 3212 5275 3242 5301
rect 3296 5275 3326 5301
rect 3380 5275 3410 5301
rect 3464 5275 3494 5301
rect 4086 5273 4116 5299
rect 4170 5273 4200 5299
rect 4254 5273 4284 5299
rect 4338 5273 4368 5299
rect 4422 5273 4452 5299
rect 4506 5273 4536 5299
rect 4590 5273 4620 5299
rect 4674 5273 4704 5299
rect 4758 5273 4788 5299
rect 4842 5273 4872 5299
rect 4926 5273 4956 5299
rect 5010 5273 5040 5299
rect 5094 5273 5124 5299
rect 5178 5273 5208 5299
rect 5262 5273 5292 5299
rect 5346 5273 5376 5299
rect 17302 5275 17332 5301
rect 17386 5275 17416 5301
rect 17470 5275 17500 5301
rect 17554 5275 17584 5301
rect 17638 5275 17668 5301
rect 17722 5275 17752 5301
rect 17806 5275 17836 5301
rect 17890 5275 17920 5301
rect 17974 5275 18004 5301
rect 18058 5275 18088 5301
rect 18142 5275 18172 5301
rect 18226 5275 18256 5301
rect 18310 5275 18340 5301
rect 18394 5275 18424 5301
rect 18478 5275 18508 5301
rect 18562 5275 18592 5301
rect 2204 5123 2234 5145
rect 2288 5123 2318 5145
rect 2372 5123 2402 5145
rect 2456 5123 2486 5145
rect 2540 5123 2570 5145
rect 2624 5123 2654 5145
rect 2708 5123 2738 5145
rect 2792 5123 2822 5145
rect 2876 5123 2906 5145
rect 2960 5123 2990 5145
rect 3044 5123 3074 5145
rect 3128 5123 3158 5145
rect 3212 5123 3242 5145
rect 3296 5123 3326 5145
rect 3380 5123 3410 5145
rect 3464 5123 3494 5145
rect 19184 5273 19214 5299
rect 19268 5273 19298 5299
rect 19352 5273 19382 5299
rect 19436 5273 19466 5299
rect 19520 5273 19550 5299
rect 19604 5273 19634 5299
rect 19688 5273 19718 5299
rect 19772 5273 19802 5299
rect 19856 5273 19886 5299
rect 19940 5273 19970 5299
rect 20024 5273 20054 5299
rect 20108 5273 20138 5299
rect 20192 5273 20222 5299
rect 20276 5273 20306 5299
rect 20360 5273 20390 5299
rect 20444 5273 20474 5299
rect 2138 5107 3494 5123
rect 4086 5121 4116 5143
rect 4170 5121 4200 5143
rect 4254 5121 4284 5143
rect 4338 5121 4368 5143
rect 4422 5121 4452 5143
rect 4506 5121 4536 5143
rect 4590 5121 4620 5143
rect 4674 5121 4704 5143
rect 4758 5121 4788 5143
rect 4842 5121 4872 5143
rect 4926 5121 4956 5143
rect 5010 5121 5040 5143
rect 5094 5121 5124 5143
rect 5178 5121 5208 5143
rect 5262 5121 5292 5143
rect 5346 5121 5376 5143
rect 17302 5123 17332 5145
rect 17386 5123 17416 5145
rect 17470 5123 17500 5145
rect 17554 5123 17584 5145
rect 17638 5123 17668 5145
rect 17722 5123 17752 5145
rect 17806 5123 17836 5145
rect 17890 5123 17920 5145
rect 17974 5123 18004 5145
rect 18058 5123 18088 5145
rect 18142 5123 18172 5145
rect 18226 5123 18256 5145
rect 18310 5123 18340 5145
rect 18394 5123 18424 5145
rect 18478 5123 18508 5145
rect 18562 5123 18592 5145
rect 2138 5073 2154 5107
rect 2188 5073 2328 5107
rect 2362 5073 2496 5107
rect 2530 5073 2665 5107
rect 2699 5073 2832 5107
rect 2866 5073 3000 5107
rect 3034 5073 3167 5107
rect 3201 5073 3494 5107
rect 2138 5057 3494 5073
rect 2204 5025 2234 5057
rect 2288 5025 2318 5057
rect 2372 5025 2402 5057
rect 2456 5025 2486 5057
rect 2540 5025 2570 5057
rect 2624 5025 2654 5057
rect 2708 5025 2738 5057
rect 2792 5025 2822 5057
rect 2876 5025 2906 5057
rect 2960 5025 2990 5057
rect 3044 5025 3074 5057
rect 3128 5025 3158 5057
rect 3212 5025 3242 5057
rect 3296 5025 3326 5057
rect 3380 5025 3410 5057
rect 3464 5025 3494 5057
rect 4020 5105 5376 5121
rect 4020 5071 4036 5105
rect 4070 5071 4210 5105
rect 4244 5071 4378 5105
rect 4412 5071 4547 5105
rect 4581 5071 4714 5105
rect 4748 5071 4882 5105
rect 4916 5071 5049 5105
rect 5083 5071 5376 5105
rect 4020 5055 5376 5071
rect 17236 5107 18592 5123
rect 19184 5121 19214 5143
rect 19268 5121 19298 5143
rect 19352 5121 19382 5143
rect 19436 5121 19466 5143
rect 19520 5121 19550 5143
rect 19604 5121 19634 5143
rect 19688 5121 19718 5143
rect 19772 5121 19802 5143
rect 19856 5121 19886 5143
rect 19940 5121 19970 5143
rect 20024 5121 20054 5143
rect 20108 5121 20138 5143
rect 20192 5121 20222 5143
rect 20276 5121 20306 5143
rect 20360 5121 20390 5143
rect 20444 5121 20474 5143
rect 17236 5073 17252 5107
rect 17286 5073 17426 5107
rect 17460 5073 17594 5107
rect 17628 5073 17763 5107
rect 17797 5073 17930 5107
rect 17964 5073 18098 5107
rect 18132 5073 18265 5107
rect 18299 5073 18592 5107
rect 17236 5057 18592 5073
rect 4086 5023 4116 5055
rect 4170 5023 4200 5055
rect 4254 5023 4284 5055
rect 4338 5023 4368 5055
rect 4422 5023 4452 5055
rect 4506 5023 4536 5055
rect 4590 5023 4620 5055
rect 4674 5023 4704 5055
rect 4758 5023 4788 5055
rect 4842 5023 4872 5055
rect 4926 5023 4956 5055
rect 5010 5023 5040 5055
rect 5094 5023 5124 5055
rect 5178 5023 5208 5055
rect 5262 5023 5292 5055
rect 5346 5023 5376 5055
rect 17302 5025 17332 5057
rect 17386 5025 17416 5057
rect 17470 5025 17500 5057
rect 17554 5025 17584 5057
rect 17638 5025 17668 5057
rect 17722 5025 17752 5057
rect 17806 5025 17836 5057
rect 17890 5025 17920 5057
rect 17974 5025 18004 5057
rect 18058 5025 18088 5057
rect 18142 5025 18172 5057
rect 18226 5025 18256 5057
rect 18310 5025 18340 5057
rect 18394 5025 18424 5057
rect 18478 5025 18508 5057
rect 18562 5025 18592 5057
rect 19118 5105 20474 5121
rect 19118 5071 19134 5105
rect 19168 5071 19308 5105
rect 19342 5071 19476 5105
rect 19510 5071 19645 5105
rect 19679 5071 19812 5105
rect 19846 5071 19980 5105
rect 20014 5071 20147 5105
rect 20181 5071 20474 5105
rect 19118 5055 20474 5071
rect 2204 4799 2234 4825
rect 2288 4799 2318 4825
rect 2372 4799 2402 4825
rect 2456 4799 2486 4825
rect 2540 4799 2570 4825
rect 2624 4799 2654 4825
rect 2708 4799 2738 4825
rect 2792 4799 2822 4825
rect 2876 4799 2906 4825
rect 2960 4799 2990 4825
rect 3044 4799 3074 4825
rect 3128 4799 3158 4825
rect 3212 4799 3242 4825
rect 3296 4799 3326 4825
rect 3380 4799 3410 4825
rect 3464 4799 3494 4825
rect 19184 5023 19214 5055
rect 19268 5023 19298 5055
rect 19352 5023 19382 5055
rect 19436 5023 19466 5055
rect 19520 5023 19550 5055
rect 19604 5023 19634 5055
rect 19688 5023 19718 5055
rect 19772 5023 19802 5055
rect 19856 5023 19886 5055
rect 19940 5023 19970 5055
rect 20024 5023 20054 5055
rect 20108 5023 20138 5055
rect 20192 5023 20222 5055
rect 20276 5023 20306 5055
rect 20360 5023 20390 5055
rect 20444 5023 20474 5055
rect 4086 4797 4116 4823
rect 4170 4797 4200 4823
rect 4254 4797 4284 4823
rect 4338 4797 4368 4823
rect 4422 4797 4452 4823
rect 4506 4797 4536 4823
rect 4590 4797 4620 4823
rect 4674 4797 4704 4823
rect 4758 4797 4788 4823
rect 4842 4797 4872 4823
rect 4926 4797 4956 4823
rect 5010 4797 5040 4823
rect 5094 4797 5124 4823
rect 5178 4797 5208 4823
rect 5262 4797 5292 4823
rect 5346 4797 5376 4823
rect 17302 4799 17332 4825
rect 17386 4799 17416 4825
rect 17470 4799 17500 4825
rect 17554 4799 17584 4825
rect 17638 4799 17668 4825
rect 17722 4799 17752 4825
rect 17806 4799 17836 4825
rect 17890 4799 17920 4825
rect 17974 4799 18004 4825
rect 18058 4799 18088 4825
rect 18142 4799 18172 4825
rect 18226 4799 18256 4825
rect 18310 4799 18340 4825
rect 18394 4799 18424 4825
rect 18478 4799 18508 4825
rect 18562 4799 18592 4825
rect 19184 4797 19214 4823
rect 19268 4797 19298 4823
rect 19352 4797 19382 4823
rect 19436 4797 19466 4823
rect 19520 4797 19550 4823
rect 19604 4797 19634 4823
rect 19688 4797 19718 4823
rect 19772 4797 19802 4823
rect 19856 4797 19886 4823
rect 19940 4797 19970 4823
rect 20024 4797 20054 4823
rect 20108 4797 20138 4823
rect 20192 4797 20222 4823
rect 20276 4797 20306 4823
rect 20360 4797 20390 4823
rect 20444 4797 20474 4823
rect -3255 4651 -3225 4677
rect -3183 4651 -3153 4677
rect -2441 4651 -2411 4677
rect -2369 4651 -2339 4677
rect -1367 4651 -1337 4677
rect -1295 4651 -1265 4677
rect -2818 4567 -2752 4583
rect -2818 4533 -2802 4567
rect -2768 4533 -2752 4567
rect -2818 4517 -2752 4533
rect -2896 4486 -2866 4512
rect -2800 4486 -2770 4517
rect -3255 4419 -3225 4451
rect -3312 4403 -3225 4419
rect -3312 4369 -3297 4403
rect -3263 4369 -3225 4403
rect -3183 4419 -3153 4451
rect -3183 4403 -3079 4419
rect -3183 4389 -3129 4403
rect -3312 4353 -3225 4369
rect -3255 4331 -3225 4353
rect -3171 4369 -3129 4389
rect -3095 4369 -3079 4403
rect -3171 4353 -3079 4369
rect -3171 4331 -3141 4353
rect -553 4651 -523 4677
rect -481 4651 -451 4677
rect 521 4651 551 4677
rect 593 4651 623 4677
rect -930 4567 -864 4583
rect -930 4533 -914 4567
rect -880 4533 -864 4567
rect -930 4517 -864 4533
rect -1008 4486 -978 4512
rect -912 4486 -882 4517
rect -2441 4419 -2411 4451
rect -2498 4403 -2411 4419
rect -2498 4369 -2483 4403
rect -2449 4369 -2411 4403
rect -2369 4419 -2339 4451
rect -1367 4419 -1337 4451
rect -2369 4403 -2265 4419
rect -2369 4389 -2315 4403
rect -2498 4353 -2411 4369
rect -2441 4331 -2411 4353
rect -2357 4369 -2315 4389
rect -2281 4369 -2265 4403
rect -2357 4353 -2265 4369
rect -1424 4403 -1337 4419
rect -1424 4369 -1409 4403
rect -1375 4369 -1337 4403
rect -1295 4419 -1265 4451
rect -1295 4403 -1191 4419
rect -1295 4389 -1241 4403
rect -1424 4353 -1337 4369
rect -2357 4331 -2327 4353
rect -1367 4331 -1337 4353
rect -1283 4369 -1241 4389
rect -1207 4369 -1191 4403
rect -1283 4353 -1191 4369
rect -1283 4331 -1253 4353
rect -2896 4255 -2866 4286
rect -2800 4260 -2770 4286
rect -2914 4239 -2848 4255
rect -2914 4205 -2898 4239
rect -2864 4218 -2848 4239
rect -2864 4205 -2736 4218
rect -3255 4175 -3225 4201
rect -3171 4175 -3141 4201
rect -2914 4186 -2736 4205
rect 1335 4651 1365 4677
rect 1407 4651 1437 4677
rect 2409 4651 2439 4677
rect 2481 4651 2511 4677
rect 958 4567 1024 4583
rect 958 4533 974 4567
rect 1008 4533 1024 4567
rect 958 4517 1024 4533
rect 880 4486 910 4512
rect 976 4486 1006 4517
rect -553 4419 -523 4451
rect -610 4403 -523 4419
rect -610 4369 -595 4403
rect -561 4369 -523 4403
rect -481 4419 -451 4451
rect 521 4419 551 4451
rect -481 4403 -377 4419
rect -481 4389 -427 4403
rect -610 4353 -523 4369
rect -553 4331 -523 4353
rect -469 4369 -427 4389
rect -393 4369 -377 4403
rect -469 4353 -377 4369
rect 464 4403 551 4419
rect 464 4369 479 4403
rect 513 4369 551 4403
rect 593 4419 623 4451
rect 593 4403 697 4419
rect 593 4389 647 4403
rect 464 4353 551 4369
rect -469 4331 -439 4353
rect 521 4331 551 4353
rect 605 4369 647 4389
rect 681 4369 697 4403
rect 605 4353 697 4369
rect 605 4331 635 4353
rect -1008 4255 -978 4286
rect -912 4260 -882 4286
rect -1026 4239 -960 4255
rect -1026 4205 -1010 4239
rect -976 4218 -960 4239
rect -976 4205 -848 4218
rect -2802 4158 -2736 4186
rect -2441 4175 -2411 4201
rect -2357 4175 -2327 4201
rect -1367 4175 -1337 4201
rect -1283 4175 -1253 4201
rect -1026 4186 -848 4205
rect 3223 4651 3253 4677
rect 3295 4651 3325 4677
rect 4297 4651 4327 4677
rect 4369 4651 4399 4677
rect 2846 4567 2912 4583
rect 2846 4533 2862 4567
rect 2896 4533 2912 4567
rect 2846 4517 2912 4533
rect 2768 4486 2798 4512
rect 2864 4486 2894 4517
rect 1335 4419 1365 4451
rect 1278 4403 1365 4419
rect 1278 4369 1293 4403
rect 1327 4369 1365 4403
rect 1407 4419 1437 4451
rect 2409 4419 2439 4451
rect 1407 4403 1511 4419
rect 1407 4389 1461 4403
rect 1278 4353 1365 4369
rect 1335 4331 1365 4353
rect 1419 4369 1461 4389
rect 1495 4369 1511 4403
rect 1419 4353 1511 4369
rect 2352 4403 2439 4419
rect 2352 4369 2367 4403
rect 2401 4369 2439 4403
rect 2481 4419 2511 4451
rect 2481 4403 2585 4419
rect 2481 4389 2535 4403
rect 2352 4353 2439 4369
rect 1419 4331 1449 4353
rect 2409 4331 2439 4353
rect 2493 4369 2535 4389
rect 2569 4369 2585 4403
rect 2493 4353 2585 4369
rect 2493 4331 2523 4353
rect 880 4255 910 4286
rect 976 4260 1006 4286
rect 862 4239 928 4255
rect 862 4205 878 4239
rect 912 4218 928 4239
rect 912 4205 1040 4218
rect -2802 4124 -2786 4158
rect -2752 4124 -2736 4158
rect -2880 4086 -2850 4112
rect -2802 4108 -2736 4124
rect -914 4158 -848 4186
rect -553 4175 -523 4201
rect -469 4175 -439 4201
rect 521 4175 551 4201
rect 605 4175 635 4201
rect 862 4186 1040 4205
rect 5111 4651 5141 4677
rect 5183 4651 5213 4677
rect 6185 4651 6215 4677
rect 6257 4651 6287 4677
rect 4734 4567 4800 4583
rect 4734 4533 4750 4567
rect 4784 4533 4800 4567
rect 4734 4517 4800 4533
rect 4656 4486 4686 4512
rect 4752 4486 4782 4517
rect 3223 4419 3253 4451
rect 3166 4403 3253 4419
rect 3166 4369 3181 4403
rect 3215 4369 3253 4403
rect 3295 4419 3325 4451
rect 4297 4419 4327 4451
rect 3295 4403 3399 4419
rect 3295 4389 3349 4403
rect 3166 4353 3253 4369
rect 3223 4331 3253 4353
rect 3307 4369 3349 4389
rect 3383 4369 3399 4403
rect 3307 4353 3399 4369
rect 4240 4403 4327 4419
rect 4240 4369 4255 4403
rect 4289 4369 4327 4403
rect 4369 4419 4399 4451
rect 4369 4403 4473 4419
rect 4369 4389 4423 4403
rect 4240 4353 4327 4369
rect 3307 4331 3337 4353
rect 4297 4331 4327 4353
rect 4381 4369 4423 4389
rect 4457 4369 4473 4403
rect 4381 4353 4473 4369
rect 4381 4331 4411 4353
rect 2768 4255 2798 4286
rect 2864 4260 2894 4286
rect 2750 4239 2816 4255
rect 2750 4205 2766 4239
rect 2800 4218 2816 4239
rect 2800 4205 2928 4218
rect -914 4124 -898 4158
rect -864 4124 -848 4158
rect -2784 4086 -2754 4108
rect -992 4086 -962 4112
rect -914 4108 -848 4124
rect 974 4158 1040 4186
rect 1335 4175 1365 4201
rect 1419 4175 1449 4201
rect 2409 4175 2439 4201
rect 2493 4175 2523 4201
rect 2750 4186 2928 4205
rect 6999 4651 7029 4677
rect 7071 4651 7101 4677
rect 8073 4651 8103 4677
rect 8145 4651 8175 4677
rect 6622 4567 6688 4583
rect 6622 4533 6638 4567
rect 6672 4533 6688 4567
rect 6622 4517 6688 4533
rect 6544 4486 6574 4512
rect 6640 4486 6670 4517
rect 5111 4419 5141 4451
rect 5054 4403 5141 4419
rect 5054 4369 5069 4403
rect 5103 4369 5141 4403
rect 5183 4419 5213 4451
rect 6185 4419 6215 4451
rect 5183 4403 5287 4419
rect 5183 4389 5237 4403
rect 5054 4353 5141 4369
rect 5111 4331 5141 4353
rect 5195 4369 5237 4389
rect 5271 4369 5287 4403
rect 5195 4353 5287 4369
rect 6128 4403 6215 4419
rect 6128 4369 6143 4403
rect 6177 4369 6215 4403
rect 6257 4419 6287 4451
rect 6257 4403 6361 4419
rect 6257 4389 6311 4403
rect 6128 4353 6215 4369
rect 5195 4331 5225 4353
rect 6185 4331 6215 4353
rect 6269 4369 6311 4389
rect 6345 4369 6361 4403
rect 6269 4353 6361 4369
rect 6269 4331 6299 4353
rect 4656 4255 4686 4286
rect 4752 4260 4782 4286
rect 4638 4239 4704 4255
rect 4638 4205 4654 4239
rect 4688 4218 4704 4239
rect 4688 4205 4816 4218
rect 974 4124 990 4158
rect 1024 4124 1040 4158
rect -896 4086 -866 4108
rect 896 4086 926 4112
rect 974 4108 1040 4124
rect 2862 4158 2928 4186
rect 3223 4175 3253 4201
rect 3307 4175 3337 4201
rect 4297 4175 4327 4201
rect 4381 4175 4411 4201
rect 4638 4186 4816 4205
rect 8887 4651 8917 4677
rect 8959 4651 8989 4677
rect 9961 4651 9991 4677
rect 10033 4651 10063 4677
rect 8510 4567 8576 4583
rect 8510 4533 8526 4567
rect 8560 4533 8576 4567
rect 8510 4517 8576 4533
rect 8432 4486 8462 4512
rect 8528 4486 8558 4517
rect 6999 4419 7029 4451
rect 6942 4403 7029 4419
rect 6942 4369 6957 4403
rect 6991 4369 7029 4403
rect 7071 4419 7101 4451
rect 8073 4419 8103 4451
rect 7071 4403 7175 4419
rect 7071 4389 7125 4403
rect 6942 4353 7029 4369
rect 6999 4331 7029 4353
rect 7083 4369 7125 4389
rect 7159 4369 7175 4403
rect 7083 4353 7175 4369
rect 8016 4403 8103 4419
rect 8016 4369 8031 4403
rect 8065 4369 8103 4403
rect 8145 4419 8175 4451
rect 8145 4403 8249 4419
rect 8145 4389 8199 4403
rect 8016 4353 8103 4369
rect 7083 4331 7113 4353
rect 8073 4331 8103 4353
rect 8157 4369 8199 4389
rect 8233 4369 8249 4403
rect 8157 4353 8249 4369
rect 8157 4331 8187 4353
rect 6544 4255 6574 4286
rect 6640 4260 6670 4286
rect 6526 4239 6592 4255
rect 6526 4205 6542 4239
rect 6576 4218 6592 4239
rect 6576 4205 6704 4218
rect 2862 4124 2878 4158
rect 2912 4124 2928 4158
rect 992 4086 1022 4108
rect 2784 4086 2814 4112
rect 2862 4108 2928 4124
rect 4750 4158 4816 4186
rect 5111 4175 5141 4201
rect 5195 4175 5225 4201
rect 6185 4175 6215 4201
rect 6269 4175 6299 4201
rect 6526 4186 6704 4205
rect 10775 4651 10805 4677
rect 10847 4651 10877 4677
rect 11843 4651 11873 4677
rect 11915 4651 11945 4677
rect 10398 4567 10464 4583
rect 10398 4533 10414 4567
rect 10448 4533 10464 4567
rect 10398 4517 10464 4533
rect 10320 4486 10350 4512
rect 10416 4486 10446 4517
rect 8887 4419 8917 4451
rect 8830 4403 8917 4419
rect 8830 4369 8845 4403
rect 8879 4369 8917 4403
rect 8959 4419 8989 4451
rect 9961 4419 9991 4451
rect 8959 4403 9063 4419
rect 8959 4389 9013 4403
rect 8830 4353 8917 4369
rect 8887 4331 8917 4353
rect 8971 4369 9013 4389
rect 9047 4369 9063 4403
rect 8971 4353 9063 4369
rect 9904 4403 9991 4419
rect 9904 4369 9919 4403
rect 9953 4369 9991 4403
rect 10033 4419 10063 4451
rect 10033 4403 10137 4419
rect 10033 4389 10087 4403
rect 9904 4353 9991 4369
rect 8971 4331 9001 4353
rect 9961 4331 9991 4353
rect 10045 4369 10087 4389
rect 10121 4369 10137 4403
rect 10045 4353 10137 4369
rect 10045 4331 10075 4353
rect 8432 4255 8462 4286
rect 8528 4260 8558 4286
rect 8414 4239 8480 4255
rect 8414 4205 8430 4239
rect 8464 4218 8480 4239
rect 8464 4205 8592 4218
rect 4750 4124 4766 4158
rect 4800 4124 4816 4158
rect 2880 4086 2910 4108
rect 4672 4086 4702 4112
rect 4750 4108 4816 4124
rect 6638 4158 6704 4186
rect 6999 4175 7029 4201
rect 7083 4175 7113 4201
rect 8073 4175 8103 4201
rect 8157 4175 8187 4201
rect 8414 4186 8592 4205
rect 12657 4651 12687 4677
rect 12729 4651 12759 4677
rect 13731 4651 13761 4677
rect 13803 4651 13833 4677
rect 12280 4567 12346 4583
rect 12280 4533 12296 4567
rect 12330 4533 12346 4567
rect 12280 4517 12346 4533
rect 12202 4486 12232 4512
rect 12298 4486 12328 4517
rect 10775 4419 10805 4451
rect 10718 4403 10805 4419
rect 10718 4369 10733 4403
rect 10767 4369 10805 4403
rect 10847 4419 10877 4451
rect 11843 4419 11873 4451
rect 10847 4403 10951 4419
rect 10847 4389 10901 4403
rect 10718 4353 10805 4369
rect 10775 4331 10805 4353
rect 10859 4369 10901 4389
rect 10935 4369 10951 4403
rect 10859 4353 10951 4369
rect 11786 4403 11873 4419
rect 11786 4369 11801 4403
rect 11835 4369 11873 4403
rect 11915 4419 11945 4451
rect 11915 4403 12019 4419
rect 11915 4389 11969 4403
rect 11786 4353 11873 4369
rect 10859 4331 10889 4353
rect 11843 4331 11873 4353
rect 11927 4369 11969 4389
rect 12003 4369 12019 4403
rect 11927 4353 12019 4369
rect 11927 4331 11957 4353
rect 10320 4255 10350 4286
rect 10416 4260 10446 4286
rect 10302 4239 10368 4255
rect 10302 4205 10318 4239
rect 10352 4218 10368 4239
rect 10352 4205 10480 4218
rect 6638 4124 6654 4158
rect 6688 4124 6704 4158
rect 4768 4086 4798 4108
rect 6560 4086 6590 4112
rect 6638 4108 6704 4124
rect 8526 4158 8592 4186
rect 8887 4175 8917 4201
rect 8971 4175 9001 4201
rect 9961 4175 9991 4201
rect 10045 4175 10075 4201
rect 10302 4186 10480 4205
rect 14545 4651 14575 4677
rect 14617 4651 14647 4677
rect 15619 4651 15649 4677
rect 15691 4651 15721 4677
rect 14168 4567 14234 4583
rect 14168 4533 14184 4567
rect 14218 4533 14234 4567
rect 14168 4517 14234 4533
rect 14090 4486 14120 4512
rect 14186 4486 14216 4517
rect 12657 4419 12687 4451
rect 12600 4403 12687 4419
rect 12600 4369 12615 4403
rect 12649 4369 12687 4403
rect 12729 4419 12759 4451
rect 13731 4419 13761 4451
rect 12729 4403 12833 4419
rect 12729 4389 12783 4403
rect 12600 4353 12687 4369
rect 12657 4331 12687 4353
rect 12741 4369 12783 4389
rect 12817 4369 12833 4403
rect 12741 4353 12833 4369
rect 13674 4403 13761 4419
rect 13674 4369 13689 4403
rect 13723 4369 13761 4403
rect 13803 4419 13833 4451
rect 13803 4403 13907 4419
rect 13803 4389 13857 4403
rect 13674 4353 13761 4369
rect 12741 4331 12771 4353
rect 13731 4331 13761 4353
rect 13815 4369 13857 4389
rect 13891 4369 13907 4403
rect 13815 4353 13907 4369
rect 13815 4331 13845 4353
rect 12202 4255 12232 4286
rect 12298 4260 12328 4286
rect 12184 4239 12250 4255
rect 12184 4205 12200 4239
rect 12234 4218 12250 4239
rect 12234 4205 12362 4218
rect 8526 4124 8542 4158
rect 8576 4124 8592 4158
rect 6656 4086 6686 4108
rect 8448 4086 8478 4112
rect 8526 4108 8592 4124
rect 10414 4158 10480 4186
rect 10775 4175 10805 4201
rect 10859 4175 10889 4201
rect 11843 4175 11873 4201
rect 11927 4175 11957 4201
rect 12184 4186 12362 4205
rect 16433 4651 16463 4677
rect 16505 4651 16535 4677
rect 17507 4651 17537 4677
rect 17579 4651 17609 4677
rect 16056 4567 16122 4583
rect 16056 4533 16072 4567
rect 16106 4533 16122 4567
rect 16056 4517 16122 4533
rect 15978 4486 16008 4512
rect 16074 4486 16104 4517
rect 14545 4419 14575 4451
rect 14488 4403 14575 4419
rect 14488 4369 14503 4403
rect 14537 4369 14575 4403
rect 14617 4419 14647 4451
rect 15619 4419 15649 4451
rect 14617 4403 14721 4419
rect 14617 4389 14671 4403
rect 14488 4353 14575 4369
rect 14545 4331 14575 4353
rect 14629 4369 14671 4389
rect 14705 4369 14721 4403
rect 14629 4353 14721 4369
rect 15562 4403 15649 4419
rect 15562 4369 15577 4403
rect 15611 4369 15649 4403
rect 15691 4419 15721 4451
rect 15691 4403 15795 4419
rect 15691 4389 15745 4403
rect 15562 4353 15649 4369
rect 14629 4331 14659 4353
rect 15619 4331 15649 4353
rect 15703 4369 15745 4389
rect 15779 4369 15795 4403
rect 15703 4353 15795 4369
rect 15703 4331 15733 4353
rect 14090 4255 14120 4286
rect 14186 4260 14216 4286
rect 14072 4239 14138 4255
rect 14072 4205 14088 4239
rect 14122 4218 14138 4239
rect 14122 4205 14250 4218
rect 10414 4124 10430 4158
rect 10464 4124 10480 4158
rect 8544 4086 8574 4108
rect 10336 4086 10366 4112
rect 10414 4108 10480 4124
rect 12296 4158 12362 4186
rect 12657 4175 12687 4201
rect 12741 4175 12771 4201
rect 13731 4175 13761 4201
rect 13815 4175 13845 4201
rect 14072 4186 14250 4205
rect 18321 4651 18351 4677
rect 18393 4651 18423 4677
rect 19395 4651 19425 4677
rect 19467 4651 19497 4677
rect 17944 4567 18010 4583
rect 17944 4533 17960 4567
rect 17994 4533 18010 4567
rect 17944 4517 18010 4533
rect 17866 4486 17896 4512
rect 17962 4486 17992 4517
rect 16433 4419 16463 4451
rect 16376 4403 16463 4419
rect 16376 4369 16391 4403
rect 16425 4369 16463 4403
rect 16505 4419 16535 4451
rect 17507 4419 17537 4451
rect 16505 4403 16609 4419
rect 16505 4389 16559 4403
rect 16376 4353 16463 4369
rect 16433 4331 16463 4353
rect 16517 4369 16559 4389
rect 16593 4369 16609 4403
rect 16517 4353 16609 4369
rect 17450 4403 17537 4419
rect 17450 4369 17465 4403
rect 17499 4369 17537 4403
rect 17579 4419 17609 4451
rect 17579 4403 17683 4419
rect 17579 4389 17633 4403
rect 17450 4353 17537 4369
rect 16517 4331 16547 4353
rect 17507 4331 17537 4353
rect 17591 4369 17633 4389
rect 17667 4369 17683 4403
rect 17591 4353 17683 4369
rect 17591 4331 17621 4353
rect 15978 4255 16008 4286
rect 16074 4260 16104 4286
rect 15960 4239 16026 4255
rect 15960 4205 15976 4239
rect 16010 4218 16026 4239
rect 16010 4205 16138 4218
rect 12296 4124 12312 4158
rect 12346 4124 12362 4158
rect 10432 4086 10462 4108
rect 12218 4086 12248 4112
rect 12296 4108 12362 4124
rect 14184 4158 14250 4186
rect 14545 4175 14575 4201
rect 14629 4175 14659 4201
rect 15619 4175 15649 4201
rect 15703 4175 15733 4201
rect 15960 4186 16138 4205
rect 20209 4651 20239 4677
rect 20281 4651 20311 4677
rect 21283 4651 21313 4677
rect 21355 4651 21385 4677
rect 19832 4567 19898 4583
rect 19832 4533 19848 4567
rect 19882 4533 19898 4567
rect 19832 4517 19898 4533
rect 19754 4486 19784 4512
rect 19850 4486 19880 4517
rect 18321 4419 18351 4451
rect 18264 4403 18351 4419
rect 18264 4369 18279 4403
rect 18313 4369 18351 4403
rect 18393 4419 18423 4451
rect 19395 4419 19425 4451
rect 18393 4403 18497 4419
rect 18393 4389 18447 4403
rect 18264 4353 18351 4369
rect 18321 4331 18351 4353
rect 18405 4369 18447 4389
rect 18481 4369 18497 4403
rect 18405 4353 18497 4369
rect 19338 4403 19425 4419
rect 19338 4369 19353 4403
rect 19387 4369 19425 4403
rect 19467 4419 19497 4451
rect 19467 4403 19571 4419
rect 19467 4389 19521 4403
rect 19338 4353 19425 4369
rect 18405 4331 18435 4353
rect 19395 4331 19425 4353
rect 19479 4369 19521 4389
rect 19555 4369 19571 4403
rect 19479 4353 19571 4369
rect 19479 4331 19509 4353
rect 17866 4255 17896 4286
rect 17962 4260 17992 4286
rect 17848 4239 17914 4255
rect 17848 4205 17864 4239
rect 17898 4218 17914 4239
rect 17898 4205 18026 4218
rect 14184 4124 14200 4158
rect 14234 4124 14250 4158
rect 12314 4086 12344 4108
rect 14106 4086 14136 4112
rect 14184 4108 14250 4124
rect 16072 4158 16138 4186
rect 16433 4175 16463 4201
rect 16517 4175 16547 4201
rect 17507 4175 17537 4201
rect 17591 4175 17621 4201
rect 17848 4186 18026 4205
rect 22097 4651 22127 4677
rect 22169 4651 22199 4677
rect 23171 4651 23201 4677
rect 23243 4651 23273 4677
rect 21720 4567 21786 4583
rect 21720 4533 21736 4567
rect 21770 4533 21786 4567
rect 21720 4517 21786 4533
rect 21642 4486 21672 4512
rect 21738 4486 21768 4517
rect 20209 4419 20239 4451
rect 20152 4403 20239 4419
rect 20152 4369 20167 4403
rect 20201 4369 20239 4403
rect 20281 4419 20311 4451
rect 21283 4419 21313 4451
rect 20281 4403 20385 4419
rect 20281 4389 20335 4403
rect 20152 4353 20239 4369
rect 20209 4331 20239 4353
rect 20293 4369 20335 4389
rect 20369 4369 20385 4403
rect 20293 4353 20385 4369
rect 21226 4403 21313 4419
rect 21226 4369 21241 4403
rect 21275 4369 21313 4403
rect 21355 4419 21385 4451
rect 21355 4403 21459 4419
rect 21355 4389 21409 4403
rect 21226 4353 21313 4369
rect 20293 4331 20323 4353
rect 21283 4331 21313 4353
rect 21367 4369 21409 4389
rect 21443 4369 21459 4403
rect 21367 4353 21459 4369
rect 21367 4331 21397 4353
rect 19754 4255 19784 4286
rect 19850 4260 19880 4286
rect 19736 4239 19802 4255
rect 19736 4205 19752 4239
rect 19786 4218 19802 4239
rect 19786 4205 19914 4218
rect 16072 4124 16088 4158
rect 16122 4124 16138 4158
rect 14202 4086 14232 4108
rect 15994 4086 16024 4112
rect 16072 4108 16138 4124
rect 17960 4158 18026 4186
rect 18321 4175 18351 4201
rect 18405 4175 18435 4201
rect 19395 4175 19425 4201
rect 19479 4175 19509 4201
rect 19736 4186 19914 4205
rect 23985 4651 24015 4677
rect 24057 4651 24087 4677
rect 25059 4651 25089 4677
rect 25131 4651 25161 4677
rect 23608 4567 23674 4583
rect 23608 4533 23624 4567
rect 23658 4533 23674 4567
rect 23608 4517 23674 4533
rect 23530 4486 23560 4512
rect 23626 4486 23656 4517
rect 22097 4419 22127 4451
rect 22040 4403 22127 4419
rect 22040 4369 22055 4403
rect 22089 4369 22127 4403
rect 22169 4419 22199 4451
rect 23171 4419 23201 4451
rect 22169 4403 22273 4419
rect 22169 4389 22223 4403
rect 22040 4353 22127 4369
rect 22097 4331 22127 4353
rect 22181 4369 22223 4389
rect 22257 4369 22273 4403
rect 22181 4353 22273 4369
rect 23114 4403 23201 4419
rect 23114 4369 23129 4403
rect 23163 4369 23201 4403
rect 23243 4419 23273 4451
rect 23243 4403 23347 4419
rect 23243 4389 23297 4403
rect 23114 4353 23201 4369
rect 22181 4331 22211 4353
rect 23171 4331 23201 4353
rect 23255 4369 23297 4389
rect 23331 4369 23347 4403
rect 23255 4353 23347 4369
rect 23255 4331 23285 4353
rect 21642 4255 21672 4286
rect 21738 4260 21768 4286
rect 21624 4239 21690 4255
rect 21624 4205 21640 4239
rect 21674 4218 21690 4239
rect 21674 4205 21802 4218
rect 17960 4124 17976 4158
rect 18010 4124 18026 4158
rect 16090 4086 16120 4108
rect 17882 4086 17912 4112
rect 17960 4108 18026 4124
rect 19848 4158 19914 4186
rect 20209 4175 20239 4201
rect 20293 4175 20323 4201
rect 21283 4175 21313 4201
rect 21367 4175 21397 4201
rect 21624 4186 21802 4205
rect 25873 4651 25903 4677
rect 25945 4651 25975 4677
rect 25496 4567 25562 4583
rect 25496 4533 25512 4567
rect 25546 4533 25562 4567
rect 25496 4517 25562 4533
rect 25418 4486 25448 4512
rect 25514 4486 25544 4517
rect 23985 4419 24015 4451
rect 23928 4403 24015 4419
rect 23928 4369 23943 4403
rect 23977 4369 24015 4403
rect 24057 4419 24087 4451
rect 25059 4419 25089 4451
rect 24057 4403 24161 4419
rect 24057 4389 24111 4403
rect 23928 4353 24015 4369
rect 23985 4331 24015 4353
rect 24069 4369 24111 4389
rect 24145 4369 24161 4403
rect 24069 4353 24161 4369
rect 25002 4403 25089 4419
rect 25002 4369 25017 4403
rect 25051 4369 25089 4403
rect 25131 4419 25161 4451
rect 25131 4403 25235 4419
rect 25131 4389 25185 4403
rect 25002 4353 25089 4369
rect 24069 4331 24099 4353
rect 25059 4331 25089 4353
rect 25143 4369 25185 4389
rect 25219 4369 25235 4403
rect 25143 4353 25235 4369
rect 25143 4331 25173 4353
rect 23530 4255 23560 4286
rect 23626 4260 23656 4286
rect 23512 4239 23578 4255
rect 23512 4205 23528 4239
rect 23562 4218 23578 4239
rect 23562 4205 23690 4218
rect 19848 4124 19864 4158
rect 19898 4124 19914 4158
rect 17978 4086 18008 4108
rect 19770 4086 19800 4112
rect 19848 4108 19914 4124
rect 21736 4158 21802 4186
rect 22097 4175 22127 4201
rect 22181 4175 22211 4201
rect 23171 4175 23201 4201
rect 23255 4175 23285 4201
rect 23512 4186 23690 4205
rect 25873 4419 25903 4451
rect 25816 4403 25903 4419
rect 25816 4369 25831 4403
rect 25865 4369 25903 4403
rect 25945 4419 25975 4451
rect 25945 4403 26049 4419
rect 25945 4389 25999 4403
rect 25816 4353 25903 4369
rect 25873 4331 25903 4353
rect 25957 4369 25999 4389
rect 26033 4369 26049 4403
rect 25957 4353 26049 4369
rect 25957 4331 25987 4353
rect 25418 4255 25448 4286
rect 25514 4260 25544 4286
rect 25400 4239 25466 4255
rect 25400 4205 25416 4239
rect 25450 4218 25466 4239
rect 25450 4205 25578 4218
rect 21736 4124 21752 4158
rect 21786 4124 21802 4158
rect 19866 4086 19896 4108
rect 21658 4086 21688 4112
rect 21736 4108 21802 4124
rect 23624 4158 23690 4186
rect 23985 4175 24015 4201
rect 24069 4175 24099 4201
rect 25059 4175 25089 4201
rect 25143 4175 25173 4201
rect 25400 4186 25578 4205
rect 23624 4124 23640 4158
rect 23674 4124 23690 4158
rect 21754 4086 21784 4108
rect 23546 4086 23576 4112
rect 23624 4108 23690 4124
rect 25512 4158 25578 4186
rect 25873 4175 25903 4201
rect 25957 4175 25987 4201
rect 25512 4124 25528 4158
rect 25562 4124 25578 4158
rect 23642 4086 23672 4108
rect 25434 4086 25464 4112
rect 25512 4108 25578 4124
rect 25530 4086 25560 4108
rect -2880 3934 -2850 3956
rect -2898 3918 -2832 3934
rect -2898 3884 -2882 3918
rect -2848 3884 -2832 3918
rect -2784 3930 -2754 3956
rect -992 3934 -962 3956
rect -2784 3900 -2650 3930
rect -2898 3868 -2832 3884
rect -2680 3732 -2650 3900
rect -1010 3918 -944 3934
rect -1010 3884 -994 3918
rect -960 3884 -944 3918
rect -896 3930 -866 3956
rect 896 3934 926 3956
rect -896 3900 -762 3930
rect -1010 3868 -944 3884
rect -792 3732 -762 3900
rect 878 3918 944 3934
rect 878 3884 894 3918
rect 928 3884 944 3918
rect 992 3930 1022 3956
rect 2784 3934 2814 3956
rect 992 3900 1126 3930
rect 878 3868 944 3884
rect 1096 3732 1126 3900
rect 2766 3918 2832 3934
rect 2766 3884 2782 3918
rect 2816 3884 2832 3918
rect 2880 3930 2910 3956
rect 4672 3934 4702 3956
rect 2880 3900 3014 3930
rect 2766 3868 2832 3884
rect 2984 3732 3014 3900
rect 4654 3918 4720 3934
rect 4654 3884 4670 3918
rect 4704 3884 4720 3918
rect 4768 3930 4798 3956
rect 6560 3934 6590 3956
rect 4768 3900 4902 3930
rect 4654 3868 4720 3884
rect 4872 3732 4902 3900
rect 6542 3918 6608 3934
rect 6542 3884 6558 3918
rect 6592 3884 6608 3918
rect 6656 3930 6686 3956
rect 8448 3934 8478 3956
rect 6656 3900 6790 3930
rect 6542 3868 6608 3884
rect 6760 3732 6790 3900
rect 8430 3918 8496 3934
rect 8430 3884 8446 3918
rect 8480 3884 8496 3918
rect 8544 3930 8574 3956
rect 10336 3934 10366 3956
rect 8544 3900 8678 3930
rect 8430 3868 8496 3884
rect 8648 3732 8678 3900
rect 10318 3918 10384 3934
rect 10318 3884 10334 3918
rect 10368 3884 10384 3918
rect 10432 3930 10462 3956
rect 12218 3934 12248 3956
rect 10432 3900 10566 3930
rect 10318 3868 10384 3884
rect 10536 3732 10566 3900
rect 12200 3918 12266 3934
rect 12200 3884 12216 3918
rect 12250 3884 12266 3918
rect 12314 3930 12344 3956
rect 14106 3934 14136 3956
rect 12314 3900 12448 3930
rect 12200 3868 12266 3884
rect 12418 3732 12448 3900
rect 14088 3918 14154 3934
rect 14088 3884 14104 3918
rect 14138 3884 14154 3918
rect 14202 3930 14232 3956
rect 15994 3934 16024 3956
rect 14202 3900 14336 3930
rect 14088 3868 14154 3884
rect 14306 3732 14336 3900
rect 15976 3918 16042 3934
rect 15976 3884 15992 3918
rect 16026 3884 16042 3918
rect 16090 3930 16120 3956
rect 17882 3934 17912 3956
rect 16090 3900 16224 3930
rect 15976 3868 16042 3884
rect 16194 3732 16224 3900
rect 17864 3918 17930 3934
rect 17864 3884 17880 3918
rect 17914 3884 17930 3918
rect 17978 3930 18008 3956
rect 19770 3934 19800 3956
rect 17978 3900 18112 3930
rect 17864 3868 17930 3884
rect 18082 3732 18112 3900
rect 19752 3918 19818 3934
rect 19752 3884 19768 3918
rect 19802 3884 19818 3918
rect 19866 3930 19896 3956
rect 21658 3934 21688 3956
rect 19866 3900 20000 3930
rect 19752 3868 19818 3884
rect 19970 3732 20000 3900
rect 21640 3918 21706 3934
rect 21640 3884 21656 3918
rect 21690 3884 21706 3918
rect 21754 3930 21784 3956
rect 23546 3934 23576 3956
rect 21754 3900 21888 3930
rect 21640 3868 21706 3884
rect 21858 3732 21888 3900
rect 23528 3918 23594 3934
rect 23528 3884 23544 3918
rect 23578 3884 23594 3918
rect 23642 3930 23672 3956
rect 25434 3934 25464 3956
rect 23642 3900 23776 3930
rect 23528 3868 23594 3884
rect 23746 3732 23776 3900
rect 25416 3918 25482 3934
rect 25416 3884 25432 3918
rect 25466 3884 25482 3918
rect 25530 3930 25560 3956
rect 25530 3900 25664 3930
rect 25416 3868 25482 3884
rect 25634 3732 25664 3900
rect -2954 3702 -2472 3732
rect -3136 3671 -3070 3687
rect -3136 3637 -3120 3671
rect -3086 3637 -3070 3671
rect -3392 3597 -3362 3623
rect -3136 3621 -3070 3637
rect -3118 3590 -3088 3621
rect -3392 3365 -3362 3397
rect -2954 3544 -2924 3702
rect -2504 3687 -2472 3702
rect -1066 3702 -584 3732
rect -2504 3671 -2424 3687
rect -2504 3637 -2474 3671
rect -2440 3637 -2424 3671
rect -2504 3621 -2424 3637
rect -1248 3671 -1182 3687
rect -1248 3637 -1232 3671
rect -1198 3637 -1182 3671
rect -2504 3620 -2442 3621
rect -2472 3590 -2442 3620
rect -2196 3605 -2166 3631
rect -2954 3514 -2868 3544
rect -2898 3430 -2868 3514
rect -2820 3511 -2754 3527
rect -2820 3477 -2804 3511
rect -2770 3477 -2754 3511
rect -2820 3461 -2754 3477
rect -2802 3430 -2772 3461
rect -3448 3349 -3362 3365
rect -3118 3359 -3088 3390
rect -3448 3315 -3432 3349
rect -3398 3315 -3362 3349
rect -3448 3299 -3362 3315
rect -3392 3277 -3362 3299
rect -3136 3343 -3070 3359
rect -3136 3309 -3120 3343
rect -3086 3309 -3070 3343
rect -3136 3293 -3070 3309
rect -1891 3603 -1861 3629
rect -1803 3603 -1773 3629
rect -1504 3597 -1474 3623
rect -1248 3621 -1182 3637
rect -1891 3430 -1861 3445
rect -1897 3406 -1861 3430
rect -2472 3359 -2442 3390
rect -2196 3373 -2166 3405
rect -2490 3343 -2424 3359
rect -2490 3309 -2474 3343
rect -2440 3309 -2424 3343
rect -2490 3293 -2424 3309
rect -2252 3357 -2166 3373
rect -1897 3371 -1867 3406
rect -1803 3384 -1773 3445
rect -1230 3590 -1200 3621
rect -2252 3323 -2236 3357
rect -2202 3323 -2166 3357
rect -2252 3307 -2166 3323
rect -2196 3285 -2166 3307
rect -1943 3355 -1867 3371
rect -1943 3321 -1933 3355
rect -1899 3321 -1867 3355
rect -1943 3305 -1867 3321
rect -1825 3368 -1771 3384
rect -1825 3334 -1815 3368
rect -1781 3334 -1771 3368
rect -1504 3365 -1474 3397
rect -1066 3544 -1036 3702
rect -616 3687 -584 3702
rect 822 3702 1304 3732
rect -616 3671 -536 3687
rect -616 3637 -586 3671
rect -552 3637 -536 3671
rect -616 3621 -536 3637
rect 640 3671 706 3687
rect 640 3637 656 3671
rect 690 3637 706 3671
rect -616 3620 -554 3621
rect -584 3590 -554 3620
rect -308 3605 -278 3631
rect -1066 3514 -980 3544
rect -1010 3430 -980 3514
rect -932 3511 -866 3527
rect -932 3477 -916 3511
rect -882 3477 -866 3511
rect -932 3461 -866 3477
rect -914 3430 -884 3461
rect -1825 3318 -1771 3334
rect -1560 3349 -1474 3365
rect -1230 3359 -1200 3390
rect -1897 3296 -1867 3305
rect -2898 3199 -2868 3230
rect -2802 3204 -2772 3230
rect -2916 3183 -2850 3199
rect -2916 3149 -2900 3183
rect -2866 3162 -2850 3183
rect -2866 3149 -2738 3162
rect -1897 3272 -1861 3296
rect -1891 3257 -1861 3272
rect -1803 3257 -1773 3318
rect -1560 3315 -1544 3349
rect -1510 3315 -1474 3349
rect -1560 3299 -1474 3315
rect -1504 3277 -1474 3299
rect -1248 3343 -1182 3359
rect -1248 3309 -1232 3343
rect -1198 3309 -1182 3343
rect -1248 3293 -1182 3309
rect -3392 3121 -3362 3147
rect -2916 3130 -2738 3149
rect -2804 3102 -2738 3130
rect -2196 3129 -2166 3155
rect -1891 3127 -1861 3153
rect -1803 3127 -1773 3153
rect -3 3603 27 3629
rect 85 3603 115 3629
rect 384 3597 414 3623
rect 640 3621 706 3637
rect -3 3430 27 3445
rect -9 3406 27 3430
rect -584 3359 -554 3390
rect -308 3373 -278 3405
rect -602 3343 -536 3359
rect -602 3309 -586 3343
rect -552 3309 -536 3343
rect -602 3293 -536 3309
rect -364 3357 -278 3373
rect -9 3371 21 3406
rect 85 3384 115 3445
rect 658 3590 688 3621
rect -364 3323 -348 3357
rect -314 3323 -278 3357
rect -364 3307 -278 3323
rect -308 3285 -278 3307
rect -55 3355 21 3371
rect -55 3321 -45 3355
rect -11 3321 21 3355
rect -55 3305 21 3321
rect 63 3368 117 3384
rect 63 3334 73 3368
rect 107 3334 117 3368
rect 384 3365 414 3397
rect 822 3544 852 3702
rect 1272 3687 1304 3702
rect 2710 3702 3192 3732
rect 1272 3671 1352 3687
rect 1272 3637 1302 3671
rect 1336 3637 1352 3671
rect 1272 3621 1352 3637
rect 2528 3671 2594 3687
rect 2528 3637 2544 3671
rect 2578 3637 2594 3671
rect 1272 3620 1334 3621
rect 1304 3590 1334 3620
rect 1580 3605 1610 3631
rect 822 3514 908 3544
rect 878 3430 908 3514
rect 956 3511 1022 3527
rect 956 3477 972 3511
rect 1006 3477 1022 3511
rect 956 3461 1022 3477
rect 974 3430 1004 3461
rect 63 3318 117 3334
rect 328 3349 414 3365
rect 658 3359 688 3390
rect -9 3296 21 3305
rect -1010 3199 -980 3230
rect -914 3204 -884 3230
rect -1028 3183 -962 3199
rect -1028 3149 -1012 3183
rect -978 3162 -962 3183
rect -978 3149 -850 3162
rect -9 3272 27 3296
rect -3 3257 27 3272
rect 85 3257 115 3318
rect 328 3315 344 3349
rect 378 3315 414 3349
rect 328 3299 414 3315
rect 384 3277 414 3299
rect 640 3343 706 3359
rect 640 3309 656 3343
rect 690 3309 706 3343
rect 640 3293 706 3309
rect -1504 3121 -1474 3147
rect -1028 3130 -850 3149
rect -2804 3068 -2788 3102
rect -2754 3068 -2738 3102
rect -2882 3030 -2852 3056
rect -2804 3052 -2738 3068
rect -916 3102 -850 3130
rect -308 3129 -278 3155
rect -3 3127 27 3153
rect 85 3127 115 3153
rect 1885 3603 1915 3629
rect 1973 3603 2003 3629
rect 2272 3597 2302 3623
rect 2528 3621 2594 3637
rect 1885 3430 1915 3445
rect 1879 3406 1915 3430
rect 1304 3359 1334 3390
rect 1580 3373 1610 3405
rect 1286 3343 1352 3359
rect 1286 3309 1302 3343
rect 1336 3309 1352 3343
rect 1286 3293 1352 3309
rect 1524 3357 1610 3373
rect 1879 3371 1909 3406
rect 1973 3384 2003 3445
rect 2546 3590 2576 3621
rect 1524 3323 1540 3357
rect 1574 3323 1610 3357
rect 1524 3307 1610 3323
rect 1580 3285 1610 3307
rect 1833 3355 1909 3371
rect 1833 3321 1843 3355
rect 1877 3321 1909 3355
rect 1833 3305 1909 3321
rect 1951 3368 2005 3384
rect 1951 3334 1961 3368
rect 1995 3334 2005 3368
rect 2272 3365 2302 3397
rect 2710 3544 2740 3702
rect 3160 3687 3192 3702
rect 4598 3702 5080 3732
rect 3160 3671 3240 3687
rect 3160 3637 3190 3671
rect 3224 3637 3240 3671
rect 3160 3621 3240 3637
rect 4416 3671 4482 3687
rect 4416 3637 4432 3671
rect 4466 3637 4482 3671
rect 3160 3620 3222 3621
rect 3192 3590 3222 3620
rect 3468 3605 3498 3631
rect 2710 3514 2796 3544
rect 2766 3430 2796 3514
rect 2844 3511 2910 3527
rect 2844 3477 2860 3511
rect 2894 3477 2910 3511
rect 2844 3461 2910 3477
rect 2862 3430 2892 3461
rect 1951 3318 2005 3334
rect 2216 3349 2302 3365
rect 2546 3359 2576 3390
rect 1879 3296 1909 3305
rect 878 3199 908 3230
rect 974 3204 1004 3230
rect 860 3183 926 3199
rect 860 3149 876 3183
rect 910 3162 926 3183
rect 910 3149 1038 3162
rect 1879 3272 1915 3296
rect 1885 3257 1915 3272
rect 1973 3257 2003 3318
rect 2216 3315 2232 3349
rect 2266 3315 2302 3349
rect 2216 3299 2302 3315
rect 2272 3277 2302 3299
rect 2528 3343 2594 3359
rect 2528 3309 2544 3343
rect 2578 3309 2594 3343
rect 2528 3293 2594 3309
rect 384 3121 414 3147
rect 860 3130 1038 3149
rect -916 3068 -900 3102
rect -866 3068 -850 3102
rect -2786 3030 -2756 3052
rect -994 3030 -964 3056
rect -916 3052 -850 3068
rect 972 3102 1038 3130
rect 1580 3129 1610 3155
rect 1885 3127 1915 3153
rect 1973 3127 2003 3153
rect 3773 3603 3803 3629
rect 3861 3603 3891 3629
rect 4160 3597 4190 3623
rect 4416 3621 4482 3637
rect 3773 3430 3803 3445
rect 3767 3406 3803 3430
rect 3192 3359 3222 3390
rect 3468 3373 3498 3405
rect 3174 3343 3240 3359
rect 3174 3309 3190 3343
rect 3224 3309 3240 3343
rect 3174 3293 3240 3309
rect 3412 3357 3498 3373
rect 3767 3371 3797 3406
rect 3861 3384 3891 3445
rect 4434 3590 4464 3621
rect 3412 3323 3428 3357
rect 3462 3323 3498 3357
rect 3412 3307 3498 3323
rect 3468 3285 3498 3307
rect 3721 3355 3797 3371
rect 3721 3321 3731 3355
rect 3765 3321 3797 3355
rect 3721 3305 3797 3321
rect 3839 3368 3893 3384
rect 3839 3334 3849 3368
rect 3883 3334 3893 3368
rect 4160 3365 4190 3397
rect 4598 3544 4628 3702
rect 5048 3687 5080 3702
rect 6486 3702 6968 3732
rect 5048 3671 5128 3687
rect 5048 3637 5078 3671
rect 5112 3637 5128 3671
rect 5048 3621 5128 3637
rect 6304 3671 6370 3687
rect 6304 3637 6320 3671
rect 6354 3637 6370 3671
rect 5048 3620 5110 3621
rect 5080 3590 5110 3620
rect 5356 3605 5386 3631
rect 4598 3514 4684 3544
rect 4654 3430 4684 3514
rect 4732 3511 4798 3527
rect 4732 3477 4748 3511
rect 4782 3477 4798 3511
rect 4732 3461 4798 3477
rect 4750 3430 4780 3461
rect 3839 3318 3893 3334
rect 4104 3349 4190 3365
rect 4434 3359 4464 3390
rect 3767 3296 3797 3305
rect 2766 3199 2796 3230
rect 2862 3204 2892 3230
rect 2748 3183 2814 3199
rect 2748 3149 2764 3183
rect 2798 3162 2814 3183
rect 2798 3149 2926 3162
rect 3767 3272 3803 3296
rect 3773 3257 3803 3272
rect 3861 3257 3891 3318
rect 4104 3315 4120 3349
rect 4154 3315 4190 3349
rect 4104 3299 4190 3315
rect 4160 3277 4190 3299
rect 4416 3343 4482 3359
rect 4416 3309 4432 3343
rect 4466 3309 4482 3343
rect 4416 3293 4482 3309
rect 2272 3121 2302 3147
rect 2748 3130 2926 3149
rect 972 3068 988 3102
rect 1022 3068 1038 3102
rect -898 3030 -868 3052
rect 894 3030 924 3056
rect 972 3052 1038 3068
rect 2860 3102 2926 3130
rect 3468 3129 3498 3155
rect 3773 3127 3803 3153
rect 3861 3127 3891 3153
rect 5661 3603 5691 3629
rect 5749 3603 5779 3629
rect 6048 3597 6078 3623
rect 6304 3621 6370 3637
rect 5661 3430 5691 3445
rect 5655 3406 5691 3430
rect 5080 3359 5110 3390
rect 5356 3373 5386 3405
rect 5062 3343 5128 3359
rect 5062 3309 5078 3343
rect 5112 3309 5128 3343
rect 5062 3293 5128 3309
rect 5300 3357 5386 3373
rect 5655 3371 5685 3406
rect 5749 3384 5779 3445
rect 6322 3590 6352 3621
rect 5300 3323 5316 3357
rect 5350 3323 5386 3357
rect 5300 3307 5386 3323
rect 5356 3285 5386 3307
rect 5609 3355 5685 3371
rect 5609 3321 5619 3355
rect 5653 3321 5685 3355
rect 5609 3305 5685 3321
rect 5727 3368 5781 3384
rect 5727 3334 5737 3368
rect 5771 3334 5781 3368
rect 6048 3365 6078 3397
rect 6486 3544 6516 3702
rect 6936 3687 6968 3702
rect 8374 3702 8856 3732
rect 6936 3671 7016 3687
rect 6936 3637 6966 3671
rect 7000 3637 7016 3671
rect 6936 3621 7016 3637
rect 8192 3671 8258 3687
rect 8192 3637 8208 3671
rect 8242 3637 8258 3671
rect 6936 3620 6998 3621
rect 6968 3590 6998 3620
rect 7244 3605 7274 3631
rect 6486 3514 6572 3544
rect 6542 3430 6572 3514
rect 6620 3511 6686 3527
rect 6620 3477 6636 3511
rect 6670 3477 6686 3511
rect 6620 3461 6686 3477
rect 6638 3430 6668 3461
rect 5727 3318 5781 3334
rect 5992 3349 6078 3365
rect 6322 3359 6352 3390
rect 5655 3296 5685 3305
rect 4654 3199 4684 3230
rect 4750 3204 4780 3230
rect 4636 3183 4702 3199
rect 4636 3149 4652 3183
rect 4686 3162 4702 3183
rect 4686 3149 4814 3162
rect 5655 3272 5691 3296
rect 5661 3257 5691 3272
rect 5749 3257 5779 3318
rect 5992 3315 6008 3349
rect 6042 3315 6078 3349
rect 5992 3299 6078 3315
rect 6048 3277 6078 3299
rect 6304 3343 6370 3359
rect 6304 3309 6320 3343
rect 6354 3309 6370 3343
rect 6304 3293 6370 3309
rect 4160 3121 4190 3147
rect 4636 3130 4814 3149
rect 2860 3068 2876 3102
rect 2910 3068 2926 3102
rect 990 3030 1020 3052
rect 2782 3030 2812 3056
rect 2860 3052 2926 3068
rect 4748 3102 4814 3130
rect 5356 3129 5386 3155
rect 5661 3127 5691 3153
rect 5749 3127 5779 3153
rect 7549 3603 7579 3629
rect 7637 3603 7667 3629
rect 7936 3597 7966 3623
rect 8192 3621 8258 3637
rect 7549 3430 7579 3445
rect 7543 3406 7579 3430
rect 6968 3359 6998 3390
rect 7244 3373 7274 3405
rect 6950 3343 7016 3359
rect 6950 3309 6966 3343
rect 7000 3309 7016 3343
rect 6950 3293 7016 3309
rect 7188 3357 7274 3373
rect 7543 3371 7573 3406
rect 7637 3384 7667 3445
rect 8210 3590 8240 3621
rect 7188 3323 7204 3357
rect 7238 3323 7274 3357
rect 7188 3307 7274 3323
rect 7244 3285 7274 3307
rect 7497 3355 7573 3371
rect 7497 3321 7507 3355
rect 7541 3321 7573 3355
rect 7497 3305 7573 3321
rect 7615 3368 7669 3384
rect 7615 3334 7625 3368
rect 7659 3334 7669 3368
rect 7936 3365 7966 3397
rect 8374 3544 8404 3702
rect 8824 3687 8856 3702
rect 10262 3702 10744 3732
rect 8824 3671 8904 3687
rect 8824 3637 8854 3671
rect 8888 3637 8904 3671
rect 8824 3621 8904 3637
rect 10080 3671 10146 3687
rect 10080 3637 10096 3671
rect 10130 3637 10146 3671
rect 8824 3620 8886 3621
rect 8856 3590 8886 3620
rect 9132 3605 9162 3631
rect 8374 3514 8460 3544
rect 8430 3430 8460 3514
rect 8508 3511 8574 3527
rect 8508 3477 8524 3511
rect 8558 3477 8574 3511
rect 8508 3461 8574 3477
rect 8526 3430 8556 3461
rect 7615 3318 7669 3334
rect 7880 3349 7966 3365
rect 8210 3359 8240 3390
rect 7543 3296 7573 3305
rect 6542 3199 6572 3230
rect 6638 3204 6668 3230
rect 6524 3183 6590 3199
rect 6524 3149 6540 3183
rect 6574 3162 6590 3183
rect 6574 3149 6702 3162
rect 7543 3272 7579 3296
rect 7549 3257 7579 3272
rect 7637 3257 7667 3318
rect 7880 3315 7896 3349
rect 7930 3315 7966 3349
rect 7880 3299 7966 3315
rect 7936 3277 7966 3299
rect 8192 3343 8258 3359
rect 8192 3309 8208 3343
rect 8242 3309 8258 3343
rect 8192 3293 8258 3309
rect 6048 3121 6078 3147
rect 6524 3130 6702 3149
rect 4748 3068 4764 3102
rect 4798 3068 4814 3102
rect 2878 3030 2908 3052
rect 4670 3030 4700 3056
rect 4748 3052 4814 3068
rect 6636 3102 6702 3130
rect 7244 3129 7274 3155
rect 7549 3127 7579 3153
rect 7637 3127 7667 3153
rect 9437 3603 9467 3629
rect 9525 3603 9555 3629
rect 9824 3597 9854 3623
rect 10080 3621 10146 3637
rect 9437 3430 9467 3445
rect 9431 3406 9467 3430
rect 8856 3359 8886 3390
rect 9132 3373 9162 3405
rect 8838 3343 8904 3359
rect 8838 3309 8854 3343
rect 8888 3309 8904 3343
rect 8838 3293 8904 3309
rect 9076 3357 9162 3373
rect 9431 3371 9461 3406
rect 9525 3384 9555 3445
rect 10098 3590 10128 3621
rect 9076 3323 9092 3357
rect 9126 3323 9162 3357
rect 9076 3307 9162 3323
rect 9132 3285 9162 3307
rect 9385 3355 9461 3371
rect 9385 3321 9395 3355
rect 9429 3321 9461 3355
rect 9385 3305 9461 3321
rect 9503 3368 9557 3384
rect 9503 3334 9513 3368
rect 9547 3334 9557 3368
rect 9824 3365 9854 3397
rect 10262 3544 10292 3702
rect 10712 3687 10744 3702
rect 12144 3702 12626 3732
rect 10712 3671 10792 3687
rect 10712 3637 10742 3671
rect 10776 3637 10792 3671
rect 10712 3621 10792 3637
rect 11962 3671 12028 3687
rect 11962 3637 11978 3671
rect 12012 3637 12028 3671
rect 10712 3620 10774 3621
rect 10744 3590 10774 3620
rect 11020 3605 11050 3631
rect 10262 3514 10348 3544
rect 10318 3430 10348 3514
rect 10396 3511 10462 3527
rect 10396 3477 10412 3511
rect 10446 3477 10462 3511
rect 10396 3461 10462 3477
rect 10414 3430 10444 3461
rect 9503 3318 9557 3334
rect 9768 3349 9854 3365
rect 10098 3359 10128 3390
rect 9431 3296 9461 3305
rect 8430 3199 8460 3230
rect 8526 3204 8556 3230
rect 8412 3183 8478 3199
rect 8412 3149 8428 3183
rect 8462 3162 8478 3183
rect 8462 3149 8590 3162
rect 9431 3272 9467 3296
rect 9437 3257 9467 3272
rect 9525 3257 9555 3318
rect 9768 3315 9784 3349
rect 9818 3315 9854 3349
rect 9768 3299 9854 3315
rect 9824 3277 9854 3299
rect 10080 3343 10146 3359
rect 10080 3309 10096 3343
rect 10130 3309 10146 3343
rect 10080 3293 10146 3309
rect 7936 3121 7966 3147
rect 8412 3130 8590 3149
rect 6636 3068 6652 3102
rect 6686 3068 6702 3102
rect 4766 3030 4796 3052
rect 6558 3030 6588 3056
rect 6636 3052 6702 3068
rect 8524 3102 8590 3130
rect 9132 3129 9162 3155
rect 9437 3127 9467 3153
rect 9525 3127 9555 3153
rect 11325 3603 11355 3629
rect 11413 3603 11443 3629
rect 11706 3597 11736 3623
rect 11962 3621 12028 3637
rect 11325 3430 11355 3445
rect 11319 3406 11355 3430
rect 10744 3359 10774 3390
rect 11020 3373 11050 3405
rect 10726 3343 10792 3359
rect 10726 3309 10742 3343
rect 10776 3309 10792 3343
rect 10726 3293 10792 3309
rect 10964 3357 11050 3373
rect 11319 3371 11349 3406
rect 11413 3384 11443 3445
rect 11980 3590 12010 3621
rect 10964 3323 10980 3357
rect 11014 3323 11050 3357
rect 10964 3307 11050 3323
rect 11020 3285 11050 3307
rect 11273 3355 11349 3371
rect 11273 3321 11283 3355
rect 11317 3321 11349 3355
rect 11273 3305 11349 3321
rect 11391 3368 11445 3384
rect 11391 3334 11401 3368
rect 11435 3334 11445 3368
rect 11706 3365 11736 3397
rect 12144 3544 12174 3702
rect 12594 3687 12626 3702
rect 14032 3702 14514 3732
rect 12594 3671 12674 3687
rect 12594 3637 12624 3671
rect 12658 3637 12674 3671
rect 12594 3621 12674 3637
rect 13850 3671 13916 3687
rect 13850 3637 13866 3671
rect 13900 3637 13916 3671
rect 12594 3620 12656 3621
rect 12626 3590 12656 3620
rect 12902 3605 12932 3631
rect 12144 3514 12230 3544
rect 12200 3430 12230 3514
rect 12278 3511 12344 3527
rect 12278 3477 12294 3511
rect 12328 3477 12344 3511
rect 12278 3461 12344 3477
rect 12296 3430 12326 3461
rect 11391 3318 11445 3334
rect 11650 3349 11736 3365
rect 11980 3359 12010 3390
rect 11319 3296 11349 3305
rect 10318 3199 10348 3230
rect 10414 3204 10444 3230
rect 10300 3183 10366 3199
rect 10300 3149 10316 3183
rect 10350 3162 10366 3183
rect 10350 3149 10478 3162
rect 11319 3272 11355 3296
rect 11325 3257 11355 3272
rect 11413 3257 11443 3318
rect 11650 3315 11666 3349
rect 11700 3315 11736 3349
rect 11650 3299 11736 3315
rect 11706 3277 11736 3299
rect 11962 3343 12028 3359
rect 11962 3309 11978 3343
rect 12012 3309 12028 3343
rect 11962 3293 12028 3309
rect 9824 3121 9854 3147
rect 10300 3130 10478 3149
rect 8524 3068 8540 3102
rect 8574 3068 8590 3102
rect 6654 3030 6684 3052
rect 8446 3030 8476 3056
rect 8524 3052 8590 3068
rect 10412 3102 10478 3130
rect 11020 3129 11050 3155
rect 11325 3127 11355 3153
rect 11413 3127 11443 3153
rect 13207 3603 13237 3629
rect 13295 3603 13325 3629
rect 13594 3597 13624 3623
rect 13850 3621 13916 3637
rect 13207 3430 13237 3445
rect 13201 3406 13237 3430
rect 12626 3359 12656 3390
rect 12902 3373 12932 3405
rect 12608 3343 12674 3359
rect 12608 3309 12624 3343
rect 12658 3309 12674 3343
rect 12608 3293 12674 3309
rect 12846 3357 12932 3373
rect 13201 3371 13231 3406
rect 13295 3384 13325 3445
rect 13868 3590 13898 3621
rect 12846 3323 12862 3357
rect 12896 3323 12932 3357
rect 12846 3307 12932 3323
rect 12902 3285 12932 3307
rect 13155 3355 13231 3371
rect 13155 3321 13165 3355
rect 13199 3321 13231 3355
rect 13155 3305 13231 3321
rect 13273 3368 13327 3384
rect 13273 3334 13283 3368
rect 13317 3334 13327 3368
rect 13594 3365 13624 3397
rect 14032 3544 14062 3702
rect 14482 3687 14514 3702
rect 15920 3702 16402 3732
rect 14482 3671 14562 3687
rect 14482 3637 14512 3671
rect 14546 3637 14562 3671
rect 14482 3621 14562 3637
rect 15738 3671 15804 3687
rect 15738 3637 15754 3671
rect 15788 3637 15804 3671
rect 14482 3620 14544 3621
rect 14514 3590 14544 3620
rect 14790 3605 14820 3631
rect 14032 3514 14118 3544
rect 14088 3430 14118 3514
rect 14166 3511 14232 3527
rect 14166 3477 14182 3511
rect 14216 3477 14232 3511
rect 14166 3461 14232 3477
rect 14184 3430 14214 3461
rect 13273 3318 13327 3334
rect 13538 3349 13624 3365
rect 13868 3359 13898 3390
rect 13201 3296 13231 3305
rect 12200 3199 12230 3230
rect 12296 3204 12326 3230
rect 12182 3183 12248 3199
rect 12182 3149 12198 3183
rect 12232 3162 12248 3183
rect 12232 3149 12360 3162
rect 13201 3272 13237 3296
rect 13207 3257 13237 3272
rect 13295 3257 13325 3318
rect 13538 3315 13554 3349
rect 13588 3315 13624 3349
rect 13538 3299 13624 3315
rect 13594 3277 13624 3299
rect 13850 3343 13916 3359
rect 13850 3309 13866 3343
rect 13900 3309 13916 3343
rect 13850 3293 13916 3309
rect 11706 3121 11736 3147
rect 12182 3130 12360 3149
rect 10412 3068 10428 3102
rect 10462 3068 10478 3102
rect 8542 3030 8572 3052
rect 10334 3030 10364 3056
rect 10412 3052 10478 3068
rect 12294 3102 12360 3130
rect 12902 3129 12932 3155
rect 13207 3127 13237 3153
rect 13295 3127 13325 3153
rect 15095 3603 15125 3629
rect 15183 3603 15213 3629
rect 15482 3597 15512 3623
rect 15738 3621 15804 3637
rect 15095 3430 15125 3445
rect 15089 3406 15125 3430
rect 14514 3359 14544 3390
rect 14790 3373 14820 3405
rect 14496 3343 14562 3359
rect 14496 3309 14512 3343
rect 14546 3309 14562 3343
rect 14496 3293 14562 3309
rect 14734 3357 14820 3373
rect 15089 3371 15119 3406
rect 15183 3384 15213 3445
rect 15756 3590 15786 3621
rect 14734 3323 14750 3357
rect 14784 3323 14820 3357
rect 14734 3307 14820 3323
rect 14790 3285 14820 3307
rect 15043 3355 15119 3371
rect 15043 3321 15053 3355
rect 15087 3321 15119 3355
rect 15043 3305 15119 3321
rect 15161 3368 15215 3384
rect 15161 3334 15171 3368
rect 15205 3334 15215 3368
rect 15482 3365 15512 3397
rect 15920 3544 15950 3702
rect 16370 3687 16402 3702
rect 17808 3702 18290 3732
rect 16370 3671 16450 3687
rect 16370 3637 16400 3671
rect 16434 3637 16450 3671
rect 16370 3621 16450 3637
rect 17626 3671 17692 3687
rect 17626 3637 17642 3671
rect 17676 3637 17692 3671
rect 16370 3620 16432 3621
rect 16402 3590 16432 3620
rect 16678 3605 16708 3631
rect 15920 3514 16006 3544
rect 15976 3430 16006 3514
rect 16054 3511 16120 3527
rect 16054 3477 16070 3511
rect 16104 3477 16120 3511
rect 16054 3461 16120 3477
rect 16072 3430 16102 3461
rect 15161 3318 15215 3334
rect 15426 3349 15512 3365
rect 15756 3359 15786 3390
rect 15089 3296 15119 3305
rect 14088 3199 14118 3230
rect 14184 3204 14214 3230
rect 14070 3183 14136 3199
rect 14070 3149 14086 3183
rect 14120 3162 14136 3183
rect 14120 3149 14248 3162
rect 15089 3272 15125 3296
rect 15095 3257 15125 3272
rect 15183 3257 15213 3318
rect 15426 3315 15442 3349
rect 15476 3315 15512 3349
rect 15426 3299 15512 3315
rect 15482 3277 15512 3299
rect 15738 3343 15804 3359
rect 15738 3309 15754 3343
rect 15788 3309 15804 3343
rect 15738 3293 15804 3309
rect 13594 3121 13624 3147
rect 14070 3130 14248 3149
rect 12294 3068 12310 3102
rect 12344 3068 12360 3102
rect 10430 3030 10460 3052
rect 12216 3030 12246 3056
rect 12294 3052 12360 3068
rect 14182 3102 14248 3130
rect 14790 3129 14820 3155
rect 15095 3127 15125 3153
rect 15183 3127 15213 3153
rect 16983 3603 17013 3629
rect 17071 3603 17101 3629
rect 17370 3597 17400 3623
rect 17626 3621 17692 3637
rect 16983 3430 17013 3445
rect 16977 3406 17013 3430
rect 16402 3359 16432 3390
rect 16678 3373 16708 3405
rect 16384 3343 16450 3359
rect 16384 3309 16400 3343
rect 16434 3309 16450 3343
rect 16384 3293 16450 3309
rect 16622 3357 16708 3373
rect 16977 3371 17007 3406
rect 17071 3384 17101 3445
rect 17644 3590 17674 3621
rect 16622 3323 16638 3357
rect 16672 3323 16708 3357
rect 16622 3307 16708 3323
rect 16678 3285 16708 3307
rect 16931 3355 17007 3371
rect 16931 3321 16941 3355
rect 16975 3321 17007 3355
rect 16931 3305 17007 3321
rect 17049 3368 17103 3384
rect 17049 3334 17059 3368
rect 17093 3334 17103 3368
rect 17370 3365 17400 3397
rect 17808 3544 17838 3702
rect 18258 3687 18290 3702
rect 19696 3702 20178 3732
rect 18258 3671 18338 3687
rect 18258 3637 18288 3671
rect 18322 3637 18338 3671
rect 18258 3621 18338 3637
rect 19514 3671 19580 3687
rect 19514 3637 19530 3671
rect 19564 3637 19580 3671
rect 18258 3620 18320 3621
rect 18290 3590 18320 3620
rect 18566 3605 18596 3631
rect 17808 3514 17894 3544
rect 17864 3430 17894 3514
rect 17942 3511 18008 3527
rect 17942 3477 17958 3511
rect 17992 3477 18008 3511
rect 17942 3461 18008 3477
rect 17960 3430 17990 3461
rect 17049 3318 17103 3334
rect 17314 3349 17400 3365
rect 17644 3359 17674 3390
rect 16977 3296 17007 3305
rect 15976 3199 16006 3230
rect 16072 3204 16102 3230
rect 15958 3183 16024 3199
rect 15958 3149 15974 3183
rect 16008 3162 16024 3183
rect 16008 3149 16136 3162
rect 16977 3272 17013 3296
rect 16983 3257 17013 3272
rect 17071 3257 17101 3318
rect 17314 3315 17330 3349
rect 17364 3315 17400 3349
rect 17314 3299 17400 3315
rect 17370 3277 17400 3299
rect 17626 3343 17692 3359
rect 17626 3309 17642 3343
rect 17676 3309 17692 3343
rect 17626 3293 17692 3309
rect 15482 3121 15512 3147
rect 15958 3130 16136 3149
rect 14182 3068 14198 3102
rect 14232 3068 14248 3102
rect 12312 3030 12342 3052
rect 14104 3030 14134 3056
rect 14182 3052 14248 3068
rect 16070 3102 16136 3130
rect 16678 3129 16708 3155
rect 16983 3127 17013 3153
rect 17071 3127 17101 3153
rect 18871 3603 18901 3629
rect 18959 3603 18989 3629
rect 19258 3597 19288 3623
rect 19514 3621 19580 3637
rect 18871 3430 18901 3445
rect 18865 3406 18901 3430
rect 18290 3359 18320 3390
rect 18566 3373 18596 3405
rect 18272 3343 18338 3359
rect 18272 3309 18288 3343
rect 18322 3309 18338 3343
rect 18272 3293 18338 3309
rect 18510 3357 18596 3373
rect 18865 3371 18895 3406
rect 18959 3384 18989 3445
rect 19532 3590 19562 3621
rect 18510 3323 18526 3357
rect 18560 3323 18596 3357
rect 18510 3307 18596 3323
rect 18566 3285 18596 3307
rect 18819 3355 18895 3371
rect 18819 3321 18829 3355
rect 18863 3321 18895 3355
rect 18819 3305 18895 3321
rect 18937 3368 18991 3384
rect 18937 3334 18947 3368
rect 18981 3334 18991 3368
rect 19258 3365 19288 3397
rect 19696 3544 19726 3702
rect 20146 3687 20178 3702
rect 21584 3702 22066 3732
rect 20146 3671 20226 3687
rect 20146 3637 20176 3671
rect 20210 3637 20226 3671
rect 20146 3621 20226 3637
rect 21402 3671 21468 3687
rect 21402 3637 21418 3671
rect 21452 3637 21468 3671
rect 20146 3620 20208 3621
rect 20178 3590 20208 3620
rect 20454 3605 20484 3631
rect 19696 3514 19782 3544
rect 19752 3430 19782 3514
rect 19830 3511 19896 3527
rect 19830 3477 19846 3511
rect 19880 3477 19896 3511
rect 19830 3461 19896 3477
rect 19848 3430 19878 3461
rect 18937 3318 18991 3334
rect 19202 3349 19288 3365
rect 19532 3359 19562 3390
rect 18865 3296 18895 3305
rect 17864 3199 17894 3230
rect 17960 3204 17990 3230
rect 17846 3183 17912 3199
rect 17846 3149 17862 3183
rect 17896 3162 17912 3183
rect 17896 3149 18024 3162
rect 18865 3272 18901 3296
rect 18871 3257 18901 3272
rect 18959 3257 18989 3318
rect 19202 3315 19218 3349
rect 19252 3315 19288 3349
rect 19202 3299 19288 3315
rect 19258 3277 19288 3299
rect 19514 3343 19580 3359
rect 19514 3309 19530 3343
rect 19564 3309 19580 3343
rect 19514 3293 19580 3309
rect 17370 3121 17400 3147
rect 17846 3130 18024 3149
rect 16070 3068 16086 3102
rect 16120 3068 16136 3102
rect 14200 3030 14230 3052
rect 15992 3030 16022 3056
rect 16070 3052 16136 3068
rect 17958 3102 18024 3130
rect 18566 3129 18596 3155
rect 18871 3127 18901 3153
rect 18959 3127 18989 3153
rect 20759 3603 20789 3629
rect 20847 3603 20877 3629
rect 21146 3597 21176 3623
rect 21402 3621 21468 3637
rect 20759 3430 20789 3445
rect 20753 3406 20789 3430
rect 20178 3359 20208 3390
rect 20454 3373 20484 3405
rect 20160 3343 20226 3359
rect 20160 3309 20176 3343
rect 20210 3309 20226 3343
rect 20160 3293 20226 3309
rect 20398 3357 20484 3373
rect 20753 3371 20783 3406
rect 20847 3384 20877 3445
rect 21420 3590 21450 3621
rect 20398 3323 20414 3357
rect 20448 3323 20484 3357
rect 20398 3307 20484 3323
rect 20454 3285 20484 3307
rect 20707 3355 20783 3371
rect 20707 3321 20717 3355
rect 20751 3321 20783 3355
rect 20707 3305 20783 3321
rect 20825 3368 20879 3384
rect 20825 3334 20835 3368
rect 20869 3334 20879 3368
rect 21146 3365 21176 3397
rect 21584 3544 21614 3702
rect 22034 3687 22066 3702
rect 23472 3702 23954 3732
rect 22034 3671 22114 3687
rect 22034 3637 22064 3671
rect 22098 3637 22114 3671
rect 22034 3621 22114 3637
rect 23290 3671 23356 3687
rect 23290 3637 23306 3671
rect 23340 3637 23356 3671
rect 22034 3620 22096 3621
rect 22066 3590 22096 3620
rect 22342 3605 22372 3631
rect 21584 3514 21670 3544
rect 21640 3430 21670 3514
rect 21718 3511 21784 3527
rect 21718 3477 21734 3511
rect 21768 3477 21784 3511
rect 21718 3461 21784 3477
rect 21736 3430 21766 3461
rect 20825 3318 20879 3334
rect 21090 3349 21176 3365
rect 21420 3359 21450 3390
rect 20753 3296 20783 3305
rect 19752 3199 19782 3230
rect 19848 3204 19878 3230
rect 19734 3183 19800 3199
rect 19734 3149 19750 3183
rect 19784 3162 19800 3183
rect 19784 3149 19912 3162
rect 20753 3272 20789 3296
rect 20759 3257 20789 3272
rect 20847 3257 20877 3318
rect 21090 3315 21106 3349
rect 21140 3315 21176 3349
rect 21090 3299 21176 3315
rect 21146 3277 21176 3299
rect 21402 3343 21468 3359
rect 21402 3309 21418 3343
rect 21452 3309 21468 3343
rect 21402 3293 21468 3309
rect 19258 3121 19288 3147
rect 19734 3130 19912 3149
rect 17958 3068 17974 3102
rect 18008 3068 18024 3102
rect 16088 3030 16118 3052
rect 17880 3030 17910 3056
rect 17958 3052 18024 3068
rect 19846 3102 19912 3130
rect 20454 3129 20484 3155
rect 20759 3127 20789 3153
rect 20847 3127 20877 3153
rect 22647 3603 22677 3629
rect 22735 3603 22765 3629
rect 23034 3597 23064 3623
rect 23290 3621 23356 3637
rect 22647 3430 22677 3445
rect 22641 3406 22677 3430
rect 22066 3359 22096 3390
rect 22342 3373 22372 3405
rect 22048 3343 22114 3359
rect 22048 3309 22064 3343
rect 22098 3309 22114 3343
rect 22048 3293 22114 3309
rect 22286 3357 22372 3373
rect 22641 3371 22671 3406
rect 22735 3384 22765 3445
rect 23308 3590 23338 3621
rect 22286 3323 22302 3357
rect 22336 3323 22372 3357
rect 22286 3307 22372 3323
rect 22342 3285 22372 3307
rect 22595 3355 22671 3371
rect 22595 3321 22605 3355
rect 22639 3321 22671 3355
rect 22595 3305 22671 3321
rect 22713 3368 22767 3384
rect 22713 3334 22723 3368
rect 22757 3334 22767 3368
rect 23034 3365 23064 3397
rect 23472 3544 23502 3702
rect 23922 3687 23954 3702
rect 25360 3702 25842 3732
rect 23922 3671 24002 3687
rect 23922 3637 23952 3671
rect 23986 3637 24002 3671
rect 23922 3621 24002 3637
rect 25178 3671 25244 3687
rect 25178 3637 25194 3671
rect 25228 3637 25244 3671
rect 23922 3620 23984 3621
rect 23954 3590 23984 3620
rect 24230 3605 24260 3631
rect 23472 3514 23558 3544
rect 23528 3430 23558 3514
rect 23606 3511 23672 3527
rect 23606 3477 23622 3511
rect 23656 3477 23672 3511
rect 23606 3461 23672 3477
rect 23624 3430 23654 3461
rect 22713 3318 22767 3334
rect 22978 3349 23064 3365
rect 23308 3359 23338 3390
rect 22641 3296 22671 3305
rect 21640 3199 21670 3230
rect 21736 3204 21766 3230
rect 21622 3183 21688 3199
rect 21622 3149 21638 3183
rect 21672 3162 21688 3183
rect 21672 3149 21800 3162
rect 22641 3272 22677 3296
rect 22647 3257 22677 3272
rect 22735 3257 22765 3318
rect 22978 3315 22994 3349
rect 23028 3315 23064 3349
rect 22978 3299 23064 3315
rect 23034 3277 23064 3299
rect 23290 3343 23356 3359
rect 23290 3309 23306 3343
rect 23340 3309 23356 3343
rect 23290 3293 23356 3309
rect 21146 3121 21176 3147
rect 21622 3130 21800 3149
rect 19846 3068 19862 3102
rect 19896 3068 19912 3102
rect 17976 3030 18006 3052
rect 19768 3030 19798 3056
rect 19846 3052 19912 3068
rect 21734 3102 21800 3130
rect 22342 3129 22372 3155
rect 22647 3127 22677 3153
rect 22735 3127 22765 3153
rect 24535 3603 24565 3629
rect 24623 3603 24653 3629
rect 24922 3597 24952 3623
rect 25178 3621 25244 3637
rect 24535 3430 24565 3445
rect 24529 3406 24565 3430
rect 23954 3359 23984 3390
rect 24230 3373 24260 3405
rect 23936 3343 24002 3359
rect 23936 3309 23952 3343
rect 23986 3309 24002 3343
rect 23936 3293 24002 3309
rect 24174 3357 24260 3373
rect 24529 3371 24559 3406
rect 24623 3384 24653 3445
rect 25196 3590 25226 3621
rect 24174 3323 24190 3357
rect 24224 3323 24260 3357
rect 24174 3307 24260 3323
rect 24230 3285 24260 3307
rect 24483 3355 24559 3371
rect 24483 3321 24493 3355
rect 24527 3321 24559 3355
rect 24483 3305 24559 3321
rect 24601 3368 24655 3384
rect 24601 3334 24611 3368
rect 24645 3334 24655 3368
rect 24922 3365 24952 3397
rect 25360 3544 25390 3702
rect 25810 3687 25842 3702
rect 25810 3671 25890 3687
rect 25810 3637 25840 3671
rect 25874 3637 25890 3671
rect 25810 3621 25890 3637
rect 25810 3620 25872 3621
rect 25842 3590 25872 3620
rect 26118 3605 26148 3631
rect 25360 3514 25446 3544
rect 25416 3430 25446 3514
rect 25494 3511 25560 3527
rect 25494 3477 25510 3511
rect 25544 3477 25560 3511
rect 25494 3461 25560 3477
rect 25512 3430 25542 3461
rect 24601 3318 24655 3334
rect 24866 3349 24952 3365
rect 25196 3359 25226 3390
rect 24529 3296 24559 3305
rect 23528 3199 23558 3230
rect 23624 3204 23654 3230
rect 23510 3183 23576 3199
rect 23510 3149 23526 3183
rect 23560 3162 23576 3183
rect 23560 3149 23688 3162
rect 24529 3272 24565 3296
rect 24535 3257 24565 3272
rect 24623 3257 24653 3318
rect 24866 3315 24882 3349
rect 24916 3315 24952 3349
rect 24866 3299 24952 3315
rect 24922 3277 24952 3299
rect 25178 3343 25244 3359
rect 25178 3309 25194 3343
rect 25228 3309 25244 3343
rect 25178 3293 25244 3309
rect 23034 3121 23064 3147
rect 23510 3130 23688 3149
rect 21734 3068 21750 3102
rect 21784 3068 21800 3102
rect 19864 3030 19894 3052
rect 21656 3030 21686 3056
rect 21734 3052 21800 3068
rect 23622 3102 23688 3130
rect 24230 3129 24260 3155
rect 24535 3127 24565 3153
rect 24623 3127 24653 3153
rect 26423 3603 26453 3629
rect 26511 3603 26541 3629
rect 26423 3430 26453 3445
rect 26417 3406 26453 3430
rect 25842 3359 25872 3390
rect 26118 3373 26148 3405
rect 25824 3343 25890 3359
rect 25824 3309 25840 3343
rect 25874 3309 25890 3343
rect 25824 3293 25890 3309
rect 26062 3357 26148 3373
rect 26417 3371 26447 3406
rect 26511 3384 26541 3445
rect 26062 3323 26078 3357
rect 26112 3323 26148 3357
rect 26062 3307 26148 3323
rect 26118 3285 26148 3307
rect 26371 3355 26447 3371
rect 26371 3321 26381 3355
rect 26415 3321 26447 3355
rect 26371 3305 26447 3321
rect 26489 3368 26543 3384
rect 26489 3334 26499 3368
rect 26533 3334 26543 3368
rect 26489 3318 26543 3334
rect 26417 3296 26447 3305
rect 25416 3199 25446 3230
rect 25512 3204 25542 3230
rect 25398 3183 25464 3199
rect 25398 3149 25414 3183
rect 25448 3162 25464 3183
rect 25448 3149 25576 3162
rect 26417 3272 26453 3296
rect 26423 3257 26453 3272
rect 26511 3257 26541 3318
rect 24922 3121 24952 3147
rect 25398 3130 25576 3149
rect 23622 3068 23638 3102
rect 23672 3068 23688 3102
rect 21752 3030 21782 3052
rect 23544 3030 23574 3056
rect 23622 3052 23688 3068
rect 25510 3102 25576 3130
rect 26118 3129 26148 3155
rect 26423 3127 26453 3153
rect 26511 3127 26541 3153
rect 25510 3068 25526 3102
rect 25560 3068 25576 3102
rect 23640 3030 23670 3052
rect 25432 3030 25462 3056
rect 25510 3052 25576 3068
rect 25528 3030 25558 3052
rect -2882 2878 -2852 2900
rect -2900 2862 -2834 2878
rect -2786 2874 -2756 2900
rect -994 2878 -964 2900
rect -2900 2828 -2884 2862
rect -2850 2828 -2834 2862
rect -2900 2812 -2834 2828
rect -1012 2862 -946 2878
rect -898 2874 -868 2900
rect 894 2878 924 2900
rect -1012 2828 -996 2862
rect -962 2828 -946 2862
rect -1012 2812 -946 2828
rect 876 2862 942 2878
rect 990 2874 1020 2900
rect 2782 2878 2812 2900
rect 876 2828 892 2862
rect 926 2828 942 2862
rect 876 2812 942 2828
rect 2764 2862 2830 2878
rect 2878 2874 2908 2900
rect 4670 2878 4700 2900
rect 2764 2828 2780 2862
rect 2814 2828 2830 2862
rect 2764 2812 2830 2828
rect 4652 2862 4718 2878
rect 4766 2874 4796 2900
rect 6558 2878 6588 2900
rect 4652 2828 4668 2862
rect 4702 2828 4718 2862
rect 4652 2812 4718 2828
rect 6540 2862 6606 2878
rect 6654 2874 6684 2900
rect 8446 2878 8476 2900
rect 6540 2828 6556 2862
rect 6590 2828 6606 2862
rect 6540 2812 6606 2828
rect 8428 2862 8494 2878
rect 8542 2874 8572 2900
rect 10334 2878 10364 2900
rect 8428 2828 8444 2862
rect 8478 2828 8494 2862
rect 8428 2812 8494 2828
rect 10316 2862 10382 2878
rect 10430 2874 10460 2900
rect 12216 2878 12246 2900
rect 10316 2828 10332 2862
rect 10366 2828 10382 2862
rect 10316 2812 10382 2828
rect 12198 2862 12264 2878
rect 12312 2874 12342 2900
rect 14104 2878 14134 2900
rect 12198 2828 12214 2862
rect 12248 2828 12264 2862
rect 12198 2812 12264 2828
rect 14086 2862 14152 2878
rect 14200 2874 14230 2900
rect 15992 2878 16022 2900
rect 14086 2828 14102 2862
rect 14136 2828 14152 2862
rect 14086 2812 14152 2828
rect 15974 2862 16040 2878
rect 16088 2874 16118 2900
rect 17880 2878 17910 2900
rect 15974 2828 15990 2862
rect 16024 2828 16040 2862
rect 15974 2812 16040 2828
rect 17862 2862 17928 2878
rect 17976 2874 18006 2900
rect 19768 2878 19798 2900
rect 17862 2828 17878 2862
rect 17912 2828 17928 2862
rect 17862 2812 17928 2828
rect 19750 2862 19816 2878
rect 19864 2874 19894 2900
rect 21656 2878 21686 2900
rect 19750 2828 19766 2862
rect 19800 2828 19816 2862
rect 19750 2812 19816 2828
rect 21638 2862 21704 2878
rect 21752 2874 21782 2900
rect 23544 2878 23574 2900
rect 21638 2828 21654 2862
rect 21688 2828 21704 2862
rect 21638 2812 21704 2828
rect 23526 2862 23592 2878
rect 23640 2874 23670 2900
rect 25432 2878 25462 2900
rect 23526 2828 23542 2862
rect 23576 2828 23592 2862
rect 23526 2812 23592 2828
rect 25414 2862 25480 2878
rect 25528 2874 25558 2900
rect 25414 2828 25430 2862
rect 25464 2828 25480 2862
rect 25414 2812 25480 2828
<< polycont >>
rect 2154 5073 2188 5107
rect 2328 5073 2362 5107
rect 2496 5073 2530 5107
rect 2665 5073 2699 5107
rect 2832 5073 2866 5107
rect 3000 5073 3034 5107
rect 3167 5073 3201 5107
rect 4036 5071 4070 5105
rect 4210 5071 4244 5105
rect 4378 5071 4412 5105
rect 4547 5071 4581 5105
rect 4714 5071 4748 5105
rect 4882 5071 4916 5105
rect 5049 5071 5083 5105
rect 17252 5073 17286 5107
rect 17426 5073 17460 5107
rect 17594 5073 17628 5107
rect 17763 5073 17797 5107
rect 17930 5073 17964 5107
rect 18098 5073 18132 5107
rect 18265 5073 18299 5107
rect 19134 5071 19168 5105
rect 19308 5071 19342 5105
rect 19476 5071 19510 5105
rect 19645 5071 19679 5105
rect 19812 5071 19846 5105
rect 19980 5071 20014 5105
rect 20147 5071 20181 5105
rect -2802 4533 -2768 4567
rect -3297 4369 -3263 4403
rect -3129 4369 -3095 4403
rect -914 4533 -880 4567
rect -2483 4369 -2449 4403
rect -2315 4369 -2281 4403
rect -1409 4369 -1375 4403
rect -1241 4369 -1207 4403
rect -2898 4205 -2864 4239
rect 974 4533 1008 4567
rect -595 4369 -561 4403
rect -427 4369 -393 4403
rect 479 4369 513 4403
rect 647 4369 681 4403
rect -1010 4205 -976 4239
rect 2862 4533 2896 4567
rect 1293 4369 1327 4403
rect 1461 4369 1495 4403
rect 2367 4369 2401 4403
rect 2535 4369 2569 4403
rect 878 4205 912 4239
rect -2786 4124 -2752 4158
rect 4750 4533 4784 4567
rect 3181 4369 3215 4403
rect 3349 4369 3383 4403
rect 4255 4369 4289 4403
rect 4423 4369 4457 4403
rect 2766 4205 2800 4239
rect -898 4124 -864 4158
rect 6638 4533 6672 4567
rect 5069 4369 5103 4403
rect 5237 4369 5271 4403
rect 6143 4369 6177 4403
rect 6311 4369 6345 4403
rect 4654 4205 4688 4239
rect 990 4124 1024 4158
rect 8526 4533 8560 4567
rect 6957 4369 6991 4403
rect 7125 4369 7159 4403
rect 8031 4369 8065 4403
rect 8199 4369 8233 4403
rect 6542 4205 6576 4239
rect 2878 4124 2912 4158
rect 10414 4533 10448 4567
rect 8845 4369 8879 4403
rect 9013 4369 9047 4403
rect 9919 4369 9953 4403
rect 10087 4369 10121 4403
rect 8430 4205 8464 4239
rect 4766 4124 4800 4158
rect 12296 4533 12330 4567
rect 10733 4369 10767 4403
rect 10901 4369 10935 4403
rect 11801 4369 11835 4403
rect 11969 4369 12003 4403
rect 10318 4205 10352 4239
rect 6654 4124 6688 4158
rect 14184 4533 14218 4567
rect 12615 4369 12649 4403
rect 12783 4369 12817 4403
rect 13689 4369 13723 4403
rect 13857 4369 13891 4403
rect 12200 4205 12234 4239
rect 8542 4124 8576 4158
rect 16072 4533 16106 4567
rect 14503 4369 14537 4403
rect 14671 4369 14705 4403
rect 15577 4369 15611 4403
rect 15745 4369 15779 4403
rect 14088 4205 14122 4239
rect 10430 4124 10464 4158
rect 17960 4533 17994 4567
rect 16391 4369 16425 4403
rect 16559 4369 16593 4403
rect 17465 4369 17499 4403
rect 17633 4369 17667 4403
rect 15976 4205 16010 4239
rect 12312 4124 12346 4158
rect 19848 4533 19882 4567
rect 18279 4369 18313 4403
rect 18447 4369 18481 4403
rect 19353 4369 19387 4403
rect 19521 4369 19555 4403
rect 17864 4205 17898 4239
rect 14200 4124 14234 4158
rect 21736 4533 21770 4567
rect 20167 4369 20201 4403
rect 20335 4369 20369 4403
rect 21241 4369 21275 4403
rect 21409 4369 21443 4403
rect 19752 4205 19786 4239
rect 16088 4124 16122 4158
rect 23624 4533 23658 4567
rect 22055 4369 22089 4403
rect 22223 4369 22257 4403
rect 23129 4369 23163 4403
rect 23297 4369 23331 4403
rect 21640 4205 21674 4239
rect 17976 4124 18010 4158
rect 25512 4533 25546 4567
rect 23943 4369 23977 4403
rect 24111 4369 24145 4403
rect 25017 4369 25051 4403
rect 25185 4369 25219 4403
rect 23528 4205 23562 4239
rect 19864 4124 19898 4158
rect 25831 4369 25865 4403
rect 25999 4369 26033 4403
rect 25416 4205 25450 4239
rect 21752 4124 21786 4158
rect 23640 4124 23674 4158
rect 25528 4124 25562 4158
rect -2882 3884 -2848 3918
rect -994 3884 -960 3918
rect 894 3884 928 3918
rect 2782 3884 2816 3918
rect 4670 3884 4704 3918
rect 6558 3884 6592 3918
rect 8446 3884 8480 3918
rect 10334 3884 10368 3918
rect 12216 3884 12250 3918
rect 14104 3884 14138 3918
rect 15992 3884 16026 3918
rect 17880 3884 17914 3918
rect 19768 3884 19802 3918
rect 21656 3884 21690 3918
rect 23544 3884 23578 3918
rect 25432 3884 25466 3918
rect -3120 3637 -3086 3671
rect -2474 3637 -2440 3671
rect -1232 3637 -1198 3671
rect -2804 3477 -2770 3511
rect -3432 3315 -3398 3349
rect -3120 3309 -3086 3343
rect -2474 3309 -2440 3343
rect -2236 3323 -2202 3357
rect -1933 3321 -1899 3355
rect -1815 3334 -1781 3368
rect -586 3637 -552 3671
rect 656 3637 690 3671
rect -916 3477 -882 3511
rect -2900 3149 -2866 3183
rect -1544 3315 -1510 3349
rect -1232 3309 -1198 3343
rect -586 3309 -552 3343
rect -348 3323 -314 3357
rect -45 3321 -11 3355
rect 73 3334 107 3368
rect 1302 3637 1336 3671
rect 2544 3637 2578 3671
rect 972 3477 1006 3511
rect -1012 3149 -978 3183
rect 344 3315 378 3349
rect 656 3309 690 3343
rect -2788 3068 -2754 3102
rect 1302 3309 1336 3343
rect 1540 3323 1574 3357
rect 1843 3321 1877 3355
rect 1961 3334 1995 3368
rect 3190 3637 3224 3671
rect 4432 3637 4466 3671
rect 2860 3477 2894 3511
rect 876 3149 910 3183
rect 2232 3315 2266 3349
rect 2544 3309 2578 3343
rect -900 3068 -866 3102
rect 3190 3309 3224 3343
rect 3428 3323 3462 3357
rect 3731 3321 3765 3355
rect 3849 3334 3883 3368
rect 5078 3637 5112 3671
rect 6320 3637 6354 3671
rect 4748 3477 4782 3511
rect 2764 3149 2798 3183
rect 4120 3315 4154 3349
rect 4432 3309 4466 3343
rect 988 3068 1022 3102
rect 5078 3309 5112 3343
rect 5316 3323 5350 3357
rect 5619 3321 5653 3355
rect 5737 3334 5771 3368
rect 6966 3637 7000 3671
rect 8208 3637 8242 3671
rect 6636 3477 6670 3511
rect 4652 3149 4686 3183
rect 6008 3315 6042 3349
rect 6320 3309 6354 3343
rect 2876 3068 2910 3102
rect 6966 3309 7000 3343
rect 7204 3323 7238 3357
rect 7507 3321 7541 3355
rect 7625 3334 7659 3368
rect 8854 3637 8888 3671
rect 10096 3637 10130 3671
rect 8524 3477 8558 3511
rect 6540 3149 6574 3183
rect 7896 3315 7930 3349
rect 8208 3309 8242 3343
rect 4764 3068 4798 3102
rect 8854 3309 8888 3343
rect 9092 3323 9126 3357
rect 9395 3321 9429 3355
rect 9513 3334 9547 3368
rect 10742 3637 10776 3671
rect 11978 3637 12012 3671
rect 10412 3477 10446 3511
rect 8428 3149 8462 3183
rect 9784 3315 9818 3349
rect 10096 3309 10130 3343
rect 6652 3068 6686 3102
rect 10742 3309 10776 3343
rect 10980 3323 11014 3357
rect 11283 3321 11317 3355
rect 11401 3334 11435 3368
rect 12624 3637 12658 3671
rect 13866 3637 13900 3671
rect 12294 3477 12328 3511
rect 10316 3149 10350 3183
rect 11666 3315 11700 3349
rect 11978 3309 12012 3343
rect 8540 3068 8574 3102
rect 12624 3309 12658 3343
rect 12862 3323 12896 3357
rect 13165 3321 13199 3355
rect 13283 3334 13317 3368
rect 14512 3637 14546 3671
rect 15754 3637 15788 3671
rect 14182 3477 14216 3511
rect 12198 3149 12232 3183
rect 13554 3315 13588 3349
rect 13866 3309 13900 3343
rect 10428 3068 10462 3102
rect 14512 3309 14546 3343
rect 14750 3323 14784 3357
rect 15053 3321 15087 3355
rect 15171 3334 15205 3368
rect 16400 3637 16434 3671
rect 17642 3637 17676 3671
rect 16070 3477 16104 3511
rect 14086 3149 14120 3183
rect 15442 3315 15476 3349
rect 15754 3309 15788 3343
rect 12310 3068 12344 3102
rect 16400 3309 16434 3343
rect 16638 3323 16672 3357
rect 16941 3321 16975 3355
rect 17059 3334 17093 3368
rect 18288 3637 18322 3671
rect 19530 3637 19564 3671
rect 17958 3477 17992 3511
rect 15974 3149 16008 3183
rect 17330 3315 17364 3349
rect 17642 3309 17676 3343
rect 14198 3068 14232 3102
rect 18288 3309 18322 3343
rect 18526 3323 18560 3357
rect 18829 3321 18863 3355
rect 18947 3334 18981 3368
rect 20176 3637 20210 3671
rect 21418 3637 21452 3671
rect 19846 3477 19880 3511
rect 17862 3149 17896 3183
rect 19218 3315 19252 3349
rect 19530 3309 19564 3343
rect 16086 3068 16120 3102
rect 20176 3309 20210 3343
rect 20414 3323 20448 3357
rect 20717 3321 20751 3355
rect 20835 3334 20869 3368
rect 22064 3637 22098 3671
rect 23306 3637 23340 3671
rect 21734 3477 21768 3511
rect 19750 3149 19784 3183
rect 21106 3315 21140 3349
rect 21418 3309 21452 3343
rect 17974 3068 18008 3102
rect 22064 3309 22098 3343
rect 22302 3323 22336 3357
rect 22605 3321 22639 3355
rect 22723 3334 22757 3368
rect 23952 3637 23986 3671
rect 25194 3637 25228 3671
rect 23622 3477 23656 3511
rect 21638 3149 21672 3183
rect 22994 3315 23028 3349
rect 23306 3309 23340 3343
rect 19862 3068 19896 3102
rect 23952 3309 23986 3343
rect 24190 3323 24224 3357
rect 24493 3321 24527 3355
rect 24611 3334 24645 3368
rect 25840 3637 25874 3671
rect 25510 3477 25544 3511
rect 23526 3149 23560 3183
rect 24882 3315 24916 3349
rect 25194 3309 25228 3343
rect 21750 3068 21784 3102
rect 25840 3309 25874 3343
rect 26078 3323 26112 3357
rect 26381 3321 26415 3355
rect 26499 3334 26533 3368
rect 25414 3149 25448 3183
rect 23638 3068 23672 3102
rect 25526 3068 25560 3102
rect -2884 2828 -2850 2862
rect -996 2828 -962 2862
rect 892 2828 926 2862
rect 2780 2828 2814 2862
rect 4668 2828 4702 2862
rect 6556 2828 6590 2862
rect 8444 2828 8478 2862
rect 10332 2828 10366 2862
rect 12214 2828 12248 2862
rect 14102 2828 14136 2862
rect 15990 2828 16024 2862
rect 17878 2828 17912 2862
rect 19766 2828 19800 2862
rect 21654 2828 21688 2862
rect 23542 2828 23576 2862
rect 25430 2828 25464 2862
<< locali >>
rect 2112 5305 2141 5339
rect 2175 5305 2233 5339
rect 2267 5305 2325 5339
rect 2359 5305 2417 5339
rect 2451 5305 2509 5339
rect 2543 5305 2601 5339
rect 2635 5305 2693 5339
rect 2727 5305 2785 5339
rect 2819 5305 2877 5339
rect 2911 5305 2969 5339
rect 3003 5305 3061 5339
rect 3095 5305 3153 5339
rect 3187 5305 3245 5339
rect 3279 5305 3337 5339
rect 3371 5305 3429 5339
rect 3463 5305 3521 5339
rect 3555 5305 3584 5339
rect 2148 5263 2194 5305
rect 2148 5229 2160 5263
rect 2148 5195 2194 5229
rect 2148 5161 2160 5195
rect 2148 5145 2194 5161
rect 2228 5263 2294 5271
rect 2228 5229 2244 5263
rect 2278 5229 2294 5263
rect 2228 5195 2294 5229
rect 2328 5263 2362 5305
rect 2328 5213 2362 5229
rect 2396 5263 2462 5271
rect 2396 5229 2412 5263
rect 2446 5229 2462 5263
rect 2228 5161 2244 5195
rect 2278 5179 2294 5195
rect 2396 5195 2462 5229
rect 2496 5263 2530 5305
rect 2496 5213 2530 5229
rect 2564 5263 2630 5271
rect 2564 5229 2580 5263
rect 2614 5229 2630 5263
rect 2396 5179 2412 5195
rect 2278 5161 2412 5179
rect 2446 5179 2462 5195
rect 2564 5195 2630 5229
rect 2664 5263 2698 5305
rect 2664 5213 2698 5229
rect 2732 5263 2798 5271
rect 2732 5229 2748 5263
rect 2782 5229 2798 5263
rect 2564 5179 2580 5195
rect 2446 5161 2580 5179
rect 2614 5179 2630 5195
rect 2732 5195 2798 5229
rect 2832 5263 2866 5305
rect 2832 5213 2866 5229
rect 2900 5263 2966 5271
rect 2900 5229 2916 5263
rect 2950 5229 2966 5263
rect 2732 5179 2748 5195
rect 2614 5161 2748 5179
rect 2782 5179 2798 5195
rect 2900 5195 2966 5229
rect 3000 5263 3034 5305
rect 3000 5213 3034 5229
rect 3068 5263 3134 5271
rect 3068 5229 3084 5263
rect 3118 5229 3134 5263
rect 2900 5179 2916 5195
rect 2782 5161 2916 5179
rect 2950 5179 2966 5195
rect 3068 5195 3134 5229
rect 3168 5263 3202 5305
rect 3168 5213 3202 5229
rect 3236 5263 3302 5271
rect 3236 5229 3252 5263
rect 3286 5229 3302 5263
rect 3068 5179 3084 5195
rect 2950 5161 3084 5179
rect 3118 5179 3134 5195
rect 3236 5195 3302 5229
rect 3336 5263 3370 5305
rect 3336 5213 3370 5229
rect 3404 5263 3470 5271
rect 3404 5229 3420 5263
rect 3454 5229 3470 5263
rect 3236 5179 3252 5195
rect 3118 5161 3252 5179
rect 3286 5179 3302 5195
rect 3404 5195 3470 5229
rect 3404 5179 3420 5195
rect 3286 5161 3420 5179
rect 3454 5161 3470 5195
rect 2228 5141 3470 5161
rect 3504 5263 3546 5305
rect 3994 5303 4023 5337
rect 4057 5303 4115 5337
rect 4149 5303 4207 5337
rect 4241 5303 4299 5337
rect 4333 5303 4391 5337
rect 4425 5303 4483 5337
rect 4517 5303 4575 5337
rect 4609 5303 4667 5337
rect 4701 5303 4759 5337
rect 4793 5303 4851 5337
rect 4885 5303 4943 5337
rect 4977 5303 5035 5337
rect 5069 5303 5127 5337
rect 5161 5303 5219 5337
rect 5253 5303 5311 5337
rect 5345 5303 5403 5337
rect 5437 5303 5466 5337
rect 17210 5305 17239 5339
rect 17273 5305 17331 5339
rect 17365 5305 17423 5339
rect 17457 5305 17515 5339
rect 17549 5305 17607 5339
rect 17641 5305 17699 5339
rect 17733 5305 17791 5339
rect 17825 5305 17883 5339
rect 17917 5305 17975 5339
rect 18009 5305 18067 5339
rect 18101 5305 18159 5339
rect 18193 5305 18251 5339
rect 18285 5305 18343 5339
rect 18377 5305 18435 5339
rect 18469 5305 18527 5339
rect 18561 5305 18619 5339
rect 18653 5305 18682 5339
rect 3538 5229 3546 5263
rect 3504 5195 3546 5229
rect 3538 5161 3546 5195
rect 3504 5145 3546 5161
rect 4030 5261 4076 5303
rect 4030 5227 4042 5261
rect 4030 5193 4076 5227
rect 4030 5159 4042 5193
rect 4030 5143 4076 5159
rect 4110 5261 4176 5269
rect 4110 5227 4126 5261
rect 4160 5227 4176 5261
rect 4110 5193 4176 5227
rect 4210 5261 4244 5303
rect 4210 5211 4244 5227
rect 4278 5261 4344 5269
rect 4278 5227 4294 5261
rect 4328 5227 4344 5261
rect 4110 5159 4126 5193
rect 4160 5177 4176 5193
rect 4278 5193 4344 5227
rect 4378 5261 4412 5303
rect 4378 5211 4412 5227
rect 4446 5261 4512 5269
rect 4446 5227 4462 5261
rect 4496 5227 4512 5261
rect 4278 5177 4294 5193
rect 4160 5159 4294 5177
rect 4328 5177 4344 5193
rect 4446 5193 4512 5227
rect 4546 5261 4580 5303
rect 4546 5211 4580 5227
rect 4614 5261 4680 5269
rect 4614 5227 4630 5261
rect 4664 5227 4680 5261
rect 4446 5177 4462 5193
rect 4328 5159 4462 5177
rect 4496 5177 4512 5193
rect 4614 5193 4680 5227
rect 4714 5261 4748 5303
rect 4714 5211 4748 5227
rect 4782 5261 4848 5269
rect 4782 5227 4798 5261
rect 4832 5227 4848 5261
rect 4614 5177 4630 5193
rect 4496 5159 4630 5177
rect 4664 5177 4680 5193
rect 4782 5193 4848 5227
rect 4882 5261 4916 5303
rect 4882 5211 4916 5227
rect 4950 5261 5016 5269
rect 4950 5227 4966 5261
rect 5000 5227 5016 5261
rect 4782 5177 4798 5193
rect 4664 5159 4798 5177
rect 4832 5177 4848 5193
rect 4950 5193 5016 5227
rect 5050 5261 5084 5303
rect 5050 5211 5084 5227
rect 5118 5261 5184 5269
rect 5118 5227 5134 5261
rect 5168 5227 5184 5261
rect 4950 5177 4966 5193
rect 4832 5159 4966 5177
rect 5000 5177 5016 5193
rect 5118 5193 5184 5227
rect 5218 5261 5252 5303
rect 5218 5211 5252 5227
rect 5286 5261 5352 5269
rect 5286 5227 5302 5261
rect 5336 5227 5352 5261
rect 5118 5177 5134 5193
rect 5000 5159 5134 5177
rect 5168 5177 5184 5193
rect 5286 5193 5352 5227
rect 5286 5177 5302 5193
rect 5168 5159 5302 5177
rect 5336 5159 5352 5193
rect 2129 5073 2154 5107
rect 2188 5102 2328 5107
rect 2188 5073 2268 5102
rect 2129 5068 2268 5073
rect 2302 5073 2328 5102
rect 2362 5102 2496 5107
rect 2530 5102 2665 5107
rect 2362 5073 2381 5102
rect 2302 5068 2381 5073
rect 2415 5068 2494 5102
rect 2530 5073 2607 5102
rect 2528 5068 2607 5073
rect 2641 5073 2665 5102
rect 2699 5102 2832 5107
rect 2866 5102 3000 5107
rect 2699 5073 2720 5102
rect 2641 5068 2720 5073
rect 2754 5073 2832 5102
rect 2754 5068 2833 5073
rect 2867 5068 2946 5102
rect 2980 5073 3000 5102
rect 3034 5102 3167 5107
rect 3034 5073 3062 5102
rect 2980 5068 3062 5073
rect 3096 5068 3166 5102
rect 3201 5073 3217 5107
rect 3200 5068 3217 5073
rect 2129 5059 3217 5068
rect 2152 5009 2194 5025
rect 3404 5023 3470 5141
rect 4110 5139 5352 5159
rect 5386 5261 5428 5303
rect 5420 5227 5428 5261
rect 5386 5193 5428 5227
rect 5420 5159 5428 5193
rect 5386 5143 5428 5159
rect 17246 5263 17292 5305
rect 17246 5229 17258 5263
rect 17246 5195 17292 5229
rect 17246 5161 17258 5195
rect 17246 5145 17292 5161
rect 17326 5263 17392 5271
rect 17326 5229 17342 5263
rect 17376 5229 17392 5263
rect 17326 5195 17392 5229
rect 17426 5263 17460 5305
rect 17426 5213 17460 5229
rect 17494 5263 17560 5271
rect 17494 5229 17510 5263
rect 17544 5229 17560 5263
rect 17326 5161 17342 5195
rect 17376 5179 17392 5195
rect 17494 5195 17560 5229
rect 17594 5263 17628 5305
rect 17594 5213 17628 5229
rect 17662 5263 17728 5271
rect 17662 5229 17678 5263
rect 17712 5229 17728 5263
rect 17494 5179 17510 5195
rect 17376 5161 17510 5179
rect 17544 5179 17560 5195
rect 17662 5195 17728 5229
rect 17762 5263 17796 5305
rect 17762 5213 17796 5229
rect 17830 5263 17896 5271
rect 17830 5229 17846 5263
rect 17880 5229 17896 5263
rect 17662 5179 17678 5195
rect 17544 5161 17678 5179
rect 17712 5179 17728 5195
rect 17830 5195 17896 5229
rect 17930 5263 17964 5305
rect 17930 5213 17964 5229
rect 17998 5263 18064 5271
rect 17998 5229 18014 5263
rect 18048 5229 18064 5263
rect 17830 5179 17846 5195
rect 17712 5161 17846 5179
rect 17880 5179 17896 5195
rect 17998 5195 18064 5229
rect 18098 5263 18132 5305
rect 18098 5213 18132 5229
rect 18166 5263 18232 5271
rect 18166 5229 18182 5263
rect 18216 5229 18232 5263
rect 17998 5179 18014 5195
rect 17880 5161 18014 5179
rect 18048 5179 18064 5195
rect 18166 5195 18232 5229
rect 18266 5263 18300 5305
rect 18266 5213 18300 5229
rect 18334 5263 18400 5271
rect 18334 5229 18350 5263
rect 18384 5229 18400 5263
rect 18166 5179 18182 5195
rect 18048 5161 18182 5179
rect 18216 5179 18232 5195
rect 18334 5195 18400 5229
rect 18434 5263 18468 5305
rect 18434 5213 18468 5229
rect 18502 5263 18568 5271
rect 18502 5229 18518 5263
rect 18552 5229 18568 5263
rect 18334 5179 18350 5195
rect 18216 5161 18350 5179
rect 18384 5179 18400 5195
rect 18502 5195 18568 5229
rect 18502 5179 18518 5195
rect 18384 5161 18518 5179
rect 18552 5161 18568 5195
rect 17326 5141 18568 5161
rect 18602 5263 18644 5305
rect 19092 5303 19121 5337
rect 19155 5303 19213 5337
rect 19247 5303 19305 5337
rect 19339 5303 19397 5337
rect 19431 5303 19489 5337
rect 19523 5303 19581 5337
rect 19615 5303 19673 5337
rect 19707 5303 19765 5337
rect 19799 5303 19857 5337
rect 19891 5303 19949 5337
rect 19983 5303 20041 5337
rect 20075 5303 20133 5337
rect 20167 5303 20225 5337
rect 20259 5303 20317 5337
rect 20351 5303 20409 5337
rect 20443 5303 20501 5337
rect 20535 5303 20564 5337
rect 18636 5229 18644 5263
rect 18602 5195 18644 5229
rect 18636 5161 18644 5195
rect 18602 5145 18644 5161
rect 19128 5261 19174 5303
rect 19128 5227 19140 5261
rect 19128 5193 19174 5227
rect 19128 5159 19140 5193
rect 19128 5143 19174 5159
rect 19208 5261 19274 5269
rect 19208 5227 19224 5261
rect 19258 5227 19274 5261
rect 19208 5193 19274 5227
rect 19308 5261 19342 5303
rect 19308 5211 19342 5227
rect 19376 5261 19442 5269
rect 19376 5227 19392 5261
rect 19426 5227 19442 5261
rect 19208 5159 19224 5193
rect 19258 5177 19274 5193
rect 19376 5193 19442 5227
rect 19476 5261 19510 5303
rect 19476 5211 19510 5227
rect 19544 5261 19610 5269
rect 19544 5227 19560 5261
rect 19594 5227 19610 5261
rect 19376 5177 19392 5193
rect 19258 5159 19392 5177
rect 19426 5177 19442 5193
rect 19544 5193 19610 5227
rect 19644 5261 19678 5303
rect 19644 5211 19678 5227
rect 19712 5261 19778 5269
rect 19712 5227 19728 5261
rect 19762 5227 19778 5261
rect 19544 5177 19560 5193
rect 19426 5159 19560 5177
rect 19594 5177 19610 5193
rect 19712 5193 19778 5227
rect 19812 5261 19846 5303
rect 19812 5211 19846 5227
rect 19880 5261 19946 5269
rect 19880 5227 19896 5261
rect 19930 5227 19946 5261
rect 19712 5177 19728 5193
rect 19594 5159 19728 5177
rect 19762 5177 19778 5193
rect 19880 5193 19946 5227
rect 19980 5261 20014 5303
rect 19980 5211 20014 5227
rect 20048 5261 20114 5269
rect 20048 5227 20064 5261
rect 20098 5227 20114 5261
rect 19880 5177 19896 5193
rect 19762 5159 19896 5177
rect 19930 5177 19946 5193
rect 20048 5193 20114 5227
rect 20148 5261 20182 5303
rect 20148 5211 20182 5227
rect 20216 5261 20282 5269
rect 20216 5227 20232 5261
rect 20266 5227 20282 5261
rect 20048 5177 20064 5193
rect 19930 5159 20064 5177
rect 20098 5177 20114 5193
rect 20216 5193 20282 5227
rect 20316 5261 20350 5303
rect 20316 5211 20350 5227
rect 20384 5261 20450 5269
rect 20384 5227 20400 5261
rect 20434 5227 20450 5261
rect 20216 5177 20232 5193
rect 20098 5159 20232 5177
rect 20266 5177 20282 5193
rect 20384 5193 20450 5227
rect 20384 5177 20400 5193
rect 20266 5159 20400 5177
rect 20434 5159 20450 5193
rect 4011 5102 4036 5105
rect 4070 5102 4210 5105
rect 4011 5068 4022 5102
rect 4070 5071 4141 5102
rect 4056 5068 4141 5071
rect 4175 5071 4210 5102
rect 4244 5102 4378 5105
rect 4412 5102 4547 5105
rect 4244 5071 4260 5102
rect 4175 5068 4260 5071
rect 4294 5071 4378 5102
rect 4294 5068 4379 5071
rect 4413 5068 4498 5102
rect 4532 5071 4547 5102
rect 4581 5102 4714 5105
rect 4748 5102 4882 5105
rect 4581 5071 4617 5102
rect 4532 5068 4617 5071
rect 4651 5071 4714 5102
rect 4770 5071 4882 5102
rect 4916 5071 5049 5105
rect 5083 5071 5099 5105
rect 4651 5068 4736 5071
rect 4770 5068 5099 5071
rect 4011 5057 5099 5068
rect 2152 4975 2160 5009
rect 2152 4939 2194 4975
rect 2152 4905 2160 4939
rect 2152 4871 2194 4905
rect 2152 4837 2160 4871
rect 2152 4795 2194 4837
rect 2228 5009 3470 5023
rect 2228 4975 2244 5009
rect 2278 5007 2412 5009
rect 2279 5005 2412 5007
rect 2279 4989 2411 5005
rect 2228 4973 2245 4975
rect 2279 4973 2294 4989
rect 2228 4939 2294 4973
rect 2396 4971 2411 4989
rect 2446 5003 2580 5009
rect 2614 5005 2748 5009
rect 2446 4989 2575 5003
rect 2446 4975 2462 4989
rect 2445 4971 2462 4975
rect 2228 4905 2244 4939
rect 2278 4905 2294 4939
rect 2228 4871 2294 4905
rect 2228 4837 2244 4871
rect 2278 4837 2294 4871
rect 2228 4829 2294 4837
rect 2328 4939 2362 4955
rect 2328 4871 2362 4905
rect 2328 4795 2362 4837
rect 2396 4939 2462 4971
rect 2564 4969 2575 4989
rect 2614 4989 2746 5005
rect 2614 4975 2630 4989
rect 2609 4969 2630 4975
rect 2396 4905 2412 4939
rect 2446 4905 2462 4939
rect 2396 4871 2462 4905
rect 2396 4837 2412 4871
rect 2446 4837 2462 4871
rect 2396 4829 2462 4837
rect 2496 4939 2530 4955
rect 2496 4871 2530 4905
rect 2496 4795 2530 4837
rect 2564 4939 2630 4969
rect 2732 4971 2746 4989
rect 2782 5001 2916 5009
rect 2782 4989 2915 5001
rect 2782 4975 2798 4989
rect 2780 4971 2798 4975
rect 2564 4905 2580 4939
rect 2614 4905 2630 4939
rect 2564 4871 2630 4905
rect 2564 4837 2580 4871
rect 2614 4837 2630 4871
rect 2564 4829 2630 4837
rect 2664 4939 2698 4955
rect 2664 4871 2698 4905
rect 2664 4795 2698 4837
rect 2732 4939 2798 4971
rect 2900 4967 2915 4989
rect 2950 4989 3084 5009
rect 3118 5006 3252 5009
rect 2950 4975 2966 4989
rect 2949 4967 2966 4975
rect 2732 4905 2748 4939
rect 2782 4905 2798 4939
rect 2732 4871 2798 4905
rect 2732 4837 2748 4871
rect 2782 4837 2798 4871
rect 2732 4829 2798 4837
rect 2832 4939 2866 4955
rect 2832 4871 2866 4905
rect 2832 4795 2866 4837
rect 2900 4939 2966 4967
rect 3068 4966 3084 4989
rect 3118 4989 3250 5006
rect 3118 4966 3134 4989
rect 2900 4905 2916 4939
rect 2950 4905 2966 4939
rect 2900 4871 2966 4905
rect 2900 4837 2916 4871
rect 2950 4837 2966 4871
rect 2900 4829 2966 4837
rect 3000 4939 3034 4955
rect 3000 4871 3034 4905
rect 3000 4795 3034 4837
rect 3068 4939 3134 4966
rect 3236 4972 3250 4989
rect 3286 4989 3420 5009
rect 3286 4975 3302 4989
rect 3284 4972 3302 4975
rect 3068 4905 3084 4939
rect 3118 4905 3134 4939
rect 3068 4871 3134 4905
rect 3068 4837 3084 4871
rect 3118 4837 3134 4871
rect 3068 4829 3134 4837
rect 3168 4939 3202 4955
rect 3168 4871 3202 4905
rect 3168 4795 3202 4837
rect 3236 4939 3302 4972
rect 3404 4974 3420 4989
rect 3454 4974 3470 5009
rect 3236 4905 3252 4939
rect 3286 4905 3302 4939
rect 3236 4871 3302 4905
rect 3236 4837 3252 4871
rect 3286 4837 3302 4871
rect 3236 4829 3302 4837
rect 3336 4939 3370 4955
rect 3336 4871 3370 4905
rect 3336 4795 3370 4837
rect 3404 4939 3470 4974
rect 4034 5007 4076 5023
rect 5286 5021 5352 5139
rect 17227 5073 17252 5107
rect 17286 5073 17426 5107
rect 17460 5102 17594 5107
rect 17227 5068 17434 5073
rect 17468 5068 17531 5102
rect 17565 5073 17594 5102
rect 17628 5102 17763 5107
rect 17565 5068 17628 5073
rect 17662 5068 17725 5102
rect 17759 5073 17763 5102
rect 17797 5102 17930 5107
rect 17964 5102 18098 5107
rect 18132 5102 18265 5107
rect 17797 5073 17822 5102
rect 17759 5068 17822 5073
rect 17856 5068 17919 5102
rect 17964 5073 18016 5102
rect 17953 5068 18016 5073
rect 18050 5073 18098 5102
rect 18050 5068 18113 5073
rect 18147 5068 18264 5102
rect 18299 5073 18315 5107
rect 18298 5068 18315 5073
rect 17227 5059 18315 5068
rect 4034 4973 4042 5007
rect 3404 4905 3420 4939
rect 3454 4905 3470 4939
rect 3404 4871 3470 4905
rect 3404 4837 3420 4871
rect 3454 4837 3470 4871
rect 3404 4829 3470 4837
rect 3504 4939 3546 4955
rect 3538 4905 3546 4939
rect 3504 4871 3546 4905
rect 3538 4837 3546 4871
rect 3504 4795 3546 4837
rect 4034 4937 4076 4973
rect 4034 4903 4042 4937
rect 4034 4869 4076 4903
rect 4034 4835 4042 4869
rect 2112 4761 2141 4795
rect 2175 4761 2233 4795
rect 2267 4761 2325 4795
rect 2359 4761 2417 4795
rect 2451 4761 2509 4795
rect 2543 4761 2601 4795
rect 2635 4761 2693 4795
rect 2727 4761 2785 4795
rect 2819 4761 2877 4795
rect 2911 4761 2969 4795
rect 3003 4761 3061 4795
rect 3095 4761 3153 4795
rect 3187 4761 3245 4795
rect 3279 4761 3337 4795
rect 3371 4761 3429 4795
rect 3463 4761 3521 4795
rect 3555 4761 3584 4795
rect 4034 4793 4076 4835
rect 4110 5009 5352 5021
rect 4110 5007 4630 5009
rect 4664 5007 5352 5009
rect 4110 4973 4126 5007
rect 4160 5005 4294 5007
rect 4168 4987 4294 5005
rect 4110 4971 4134 4973
rect 4168 4971 4176 4987
rect 4110 4937 4176 4971
rect 4278 4971 4294 4987
rect 4328 4999 4462 5007
rect 4328 4987 4461 4999
rect 4328 4971 4344 4987
rect 4110 4903 4126 4937
rect 4160 4903 4176 4937
rect 4110 4869 4176 4903
rect 4110 4835 4126 4869
rect 4160 4835 4176 4869
rect 4110 4827 4176 4835
rect 4210 4937 4244 4953
rect 4210 4869 4244 4903
rect 4210 4793 4244 4835
rect 4278 4937 4344 4971
rect 4446 4965 4461 4987
rect 4496 4987 4630 5007
rect 4496 4973 4512 4987
rect 4495 4965 4512 4973
rect 4278 4903 4294 4937
rect 4328 4903 4344 4937
rect 4278 4869 4344 4903
rect 4278 4835 4294 4869
rect 4328 4835 4344 4869
rect 4278 4827 4344 4835
rect 4378 4937 4412 4953
rect 4378 4869 4412 4903
rect 4378 4793 4412 4835
rect 4446 4937 4512 4965
rect 4614 4973 4630 4987
rect 4664 4996 4798 5007
rect 4832 5002 4966 5007
rect 4664 4987 4794 4996
rect 4664 4973 4680 4987
rect 4446 4903 4462 4937
rect 4496 4903 4512 4937
rect 4446 4869 4512 4903
rect 4446 4835 4462 4869
rect 4496 4835 4512 4869
rect 4446 4827 4512 4835
rect 4546 4937 4580 4953
rect 4546 4869 4580 4903
rect 4546 4793 4580 4835
rect 4614 4937 4680 4973
rect 4782 4962 4794 4987
rect 4832 4987 4964 5002
rect 4832 4973 4848 4987
rect 4828 4962 4848 4973
rect 4614 4903 4630 4937
rect 4664 4903 4680 4937
rect 4614 4869 4680 4903
rect 4614 4835 4630 4869
rect 4664 4835 4680 4869
rect 4614 4827 4680 4835
rect 4714 4937 4748 4953
rect 4714 4869 4748 4903
rect 4714 4793 4748 4835
rect 4782 4937 4848 4962
rect 4950 4968 4964 4987
rect 5000 4987 5134 5007
rect 5168 5006 5302 5007
rect 5000 4973 5016 4987
rect 4998 4968 5016 4973
rect 4782 4903 4798 4937
rect 4832 4903 4848 4937
rect 4782 4869 4848 4903
rect 4782 4835 4798 4869
rect 4832 4835 4848 4869
rect 4782 4827 4848 4835
rect 4882 4937 4916 4953
rect 4882 4869 4916 4903
rect 4882 4793 4916 4835
rect 4950 4937 5016 4968
rect 5118 4970 5134 4987
rect 5168 4987 5293 5006
rect 5168 4970 5184 4987
rect 4950 4903 4966 4937
rect 5000 4903 5016 4937
rect 4950 4869 5016 4903
rect 4950 4835 4966 4869
rect 5000 4835 5016 4869
rect 4950 4827 5016 4835
rect 5050 4937 5084 4953
rect 5050 4869 5084 4903
rect 5050 4793 5084 4835
rect 5118 4937 5184 4970
rect 5286 4972 5293 4987
rect 5336 4973 5352 5007
rect 5327 4972 5352 4973
rect 5118 4903 5134 4937
rect 5168 4903 5184 4937
rect 5118 4869 5184 4903
rect 5118 4835 5134 4869
rect 5168 4835 5184 4869
rect 5118 4827 5184 4835
rect 5218 4937 5252 4953
rect 5218 4869 5252 4903
rect 5218 4793 5252 4835
rect 5286 4937 5352 4972
rect 17250 5009 17292 5025
rect 18502 5023 18568 5141
rect 19208 5139 20450 5159
rect 20484 5261 20526 5303
rect 20518 5227 20526 5261
rect 20484 5193 20526 5227
rect 20518 5159 20526 5193
rect 20484 5143 20526 5159
rect 19109 5102 19134 5105
rect 19168 5102 19308 5105
rect 19342 5102 19476 5105
rect 19510 5102 19645 5105
rect 19679 5102 19812 5105
rect 19109 5068 19120 5102
rect 19168 5071 19228 5102
rect 19154 5068 19228 5071
rect 19262 5071 19308 5102
rect 19262 5068 19336 5071
rect 19370 5068 19444 5102
rect 19510 5071 19552 5102
rect 19478 5068 19552 5071
rect 19586 5071 19645 5102
rect 19586 5068 19660 5071
rect 19694 5068 19768 5102
rect 19802 5071 19812 5102
rect 19846 5102 19980 5105
rect 19846 5071 19876 5102
rect 19802 5068 19876 5071
rect 19910 5071 19980 5102
rect 20014 5071 20147 5105
rect 20181 5071 20197 5105
rect 19910 5068 20197 5071
rect 19109 5057 20197 5068
rect 17250 4975 17258 5009
rect 5286 4903 5302 4937
rect 5336 4903 5352 4937
rect 5286 4869 5352 4903
rect 5286 4835 5302 4869
rect 5336 4835 5352 4869
rect 5286 4827 5352 4835
rect 5386 4937 5428 4953
rect 5420 4903 5428 4937
rect 5386 4869 5428 4903
rect 5420 4835 5428 4869
rect 5386 4793 5428 4835
rect 17250 4939 17292 4975
rect 17250 4905 17258 4939
rect 17250 4871 17292 4905
rect 17250 4837 17258 4871
rect 17250 4795 17292 4837
rect 17326 5009 18568 5023
rect 17326 4975 17342 5009
rect 17376 5001 17510 5009
rect 17377 4996 17510 5001
rect 17377 4989 17506 4996
rect 17326 4967 17343 4975
rect 17377 4967 17392 4989
rect 17326 4939 17392 4967
rect 17494 4962 17506 4989
rect 17544 4989 17678 5009
rect 17712 5005 17846 5009
rect 17712 5000 17844 5005
rect 17544 4975 17560 4989
rect 17540 4962 17560 4975
rect 17326 4905 17342 4939
rect 17376 4905 17392 4939
rect 17326 4871 17392 4905
rect 17326 4837 17342 4871
rect 17376 4837 17392 4871
rect 17326 4829 17392 4837
rect 17426 4939 17460 4955
rect 17426 4871 17460 4905
rect 17426 4795 17460 4837
rect 17494 4939 17560 4962
rect 17662 4975 17678 4989
rect 17713 4989 17844 5000
rect 17662 4966 17679 4975
rect 17713 4966 17728 4989
rect 17494 4905 17510 4939
rect 17544 4905 17560 4939
rect 17494 4871 17560 4905
rect 17494 4837 17510 4871
rect 17544 4837 17560 4871
rect 17494 4829 17560 4837
rect 17594 4939 17628 4955
rect 17594 4871 17628 4905
rect 17594 4795 17628 4837
rect 17662 4939 17728 4966
rect 17830 4971 17844 4989
rect 17880 4992 18014 5009
rect 17880 4989 18011 4992
rect 17880 4975 17896 4989
rect 17878 4971 17896 4975
rect 17662 4905 17678 4939
rect 17712 4905 17728 4939
rect 17662 4871 17728 4905
rect 17662 4837 17678 4871
rect 17712 4837 17728 4871
rect 17662 4829 17728 4837
rect 17762 4939 17796 4955
rect 17762 4871 17796 4905
rect 17762 4795 17796 4837
rect 17830 4939 17896 4971
rect 17998 4958 18011 4989
rect 18048 4990 18182 5009
rect 18216 4999 18350 5009
rect 18048 4989 18179 4990
rect 18048 4975 18064 4989
rect 18045 4958 18064 4975
rect 17830 4905 17846 4939
rect 17880 4905 17896 4939
rect 17830 4871 17896 4905
rect 17830 4837 17846 4871
rect 17880 4837 17896 4871
rect 17830 4829 17896 4837
rect 17930 4939 17964 4955
rect 17930 4871 17964 4905
rect 17930 4795 17964 4837
rect 17998 4939 18064 4958
rect 18166 4956 18179 4989
rect 18216 4989 18349 4999
rect 18216 4975 18232 4989
rect 18213 4956 18232 4975
rect 17998 4905 18014 4939
rect 18048 4905 18064 4939
rect 17998 4871 18064 4905
rect 17998 4837 18014 4871
rect 18048 4837 18064 4871
rect 17998 4829 18064 4837
rect 18098 4939 18132 4955
rect 18098 4871 18132 4905
rect 18098 4795 18132 4837
rect 18166 4939 18232 4956
rect 18334 4965 18349 4989
rect 18384 4989 18518 5009
rect 18384 4975 18400 4989
rect 18383 4965 18400 4975
rect 18166 4905 18182 4939
rect 18216 4905 18232 4939
rect 18166 4871 18232 4905
rect 18166 4837 18182 4871
rect 18216 4837 18232 4871
rect 18166 4829 18232 4837
rect 18266 4939 18300 4955
rect 18266 4871 18300 4905
rect 18266 4795 18300 4837
rect 18334 4939 18400 4965
rect 18502 4975 18518 4989
rect 18552 4975 18568 5009
rect 18334 4905 18350 4939
rect 18384 4905 18400 4939
rect 18334 4871 18400 4905
rect 18334 4837 18350 4871
rect 18384 4837 18400 4871
rect 18334 4829 18400 4837
rect 18434 4939 18468 4955
rect 18434 4871 18468 4905
rect 18434 4795 18468 4837
rect 18502 4939 18568 4975
rect 19132 5007 19174 5023
rect 20384 5021 20450 5139
rect 19132 4973 19140 5007
rect 18502 4905 18518 4939
rect 18552 4905 18568 4939
rect 18502 4871 18568 4905
rect 18502 4837 18518 4871
rect 18552 4837 18568 4871
rect 18502 4829 18568 4837
rect 18602 4939 18644 4955
rect 18636 4905 18644 4939
rect 18602 4871 18644 4905
rect 18636 4837 18644 4871
rect 18602 4795 18644 4837
rect 19132 4937 19174 4973
rect 19132 4903 19140 4937
rect 19132 4869 19174 4903
rect 19132 4835 19140 4869
rect 3994 4759 4023 4793
rect 4057 4759 4115 4793
rect 4149 4759 4207 4793
rect 4241 4759 4299 4793
rect 4333 4759 4391 4793
rect 4425 4759 4483 4793
rect 4517 4759 4575 4793
rect 4609 4759 4667 4793
rect 4701 4759 4759 4793
rect 4793 4759 4851 4793
rect 4885 4759 4943 4793
rect 4977 4759 5035 4793
rect 5069 4759 5127 4793
rect 5161 4759 5219 4793
rect 5253 4759 5311 4793
rect 5345 4759 5403 4793
rect 5437 4759 5466 4793
rect 17210 4761 17239 4795
rect 17273 4761 17331 4795
rect 17365 4761 17423 4795
rect 17457 4761 17515 4795
rect 17549 4761 17607 4795
rect 17641 4761 17699 4795
rect 17733 4761 17791 4795
rect 17825 4761 17883 4795
rect 17917 4761 17975 4795
rect 18009 4761 18067 4795
rect 18101 4761 18159 4795
rect 18193 4761 18251 4795
rect 18285 4761 18343 4795
rect 18377 4761 18435 4795
rect 18469 4761 18527 4795
rect 18561 4761 18619 4795
rect 18653 4761 18682 4795
rect 19132 4793 19174 4835
rect 19208 5009 20450 5021
rect 19208 5007 19728 5009
rect 19762 5007 20450 5009
rect 19208 5000 19224 5007
rect 19208 4966 19222 5000
rect 19258 4987 19392 5007
rect 19426 5006 19560 5007
rect 19426 5001 19557 5006
rect 19258 4973 19274 4987
rect 19256 4966 19274 4973
rect 19208 4937 19274 4966
rect 19376 4973 19392 4987
rect 19429 4987 19557 5001
rect 19376 4967 19395 4973
rect 19429 4967 19442 4987
rect 19208 4903 19224 4937
rect 19258 4903 19274 4937
rect 19208 4869 19274 4903
rect 19208 4835 19224 4869
rect 19258 4835 19274 4869
rect 19208 4827 19274 4835
rect 19308 4937 19342 4953
rect 19308 4869 19342 4903
rect 19308 4793 19342 4835
rect 19376 4937 19442 4967
rect 19544 4972 19557 4987
rect 19594 4987 19728 5007
rect 19594 4973 19610 4987
rect 19591 4972 19610 4973
rect 19376 4903 19392 4937
rect 19426 4903 19442 4937
rect 19376 4869 19442 4903
rect 19376 4835 19392 4869
rect 19426 4835 19442 4869
rect 19376 4827 19442 4835
rect 19476 4937 19510 4953
rect 19476 4869 19510 4903
rect 19476 4793 19510 4835
rect 19544 4937 19610 4972
rect 19712 4973 19728 4987
rect 19762 4987 19896 5007
rect 19930 4995 20064 5007
rect 19762 4973 19778 4987
rect 19544 4903 19560 4937
rect 19594 4903 19610 4937
rect 19544 4869 19610 4903
rect 19544 4835 19560 4869
rect 19594 4835 19610 4869
rect 19544 4827 19610 4835
rect 19644 4937 19678 4953
rect 19644 4869 19678 4903
rect 19644 4793 19678 4835
rect 19712 4937 19778 4973
rect 19880 4973 19896 4987
rect 19931 4987 20062 4995
rect 19880 4961 19897 4973
rect 19931 4961 19946 4987
rect 19712 4903 19728 4937
rect 19762 4903 19778 4937
rect 19712 4869 19778 4903
rect 19712 4835 19728 4869
rect 19762 4835 19778 4869
rect 19712 4827 19778 4835
rect 19812 4937 19846 4953
rect 19812 4869 19846 4903
rect 19812 4793 19846 4835
rect 19880 4937 19946 4961
rect 20048 4961 20062 4987
rect 20098 4987 20232 5007
rect 20266 4997 20400 5007
rect 20098 4973 20114 4987
rect 20096 4961 20114 4973
rect 19880 4903 19896 4937
rect 19930 4903 19946 4937
rect 19880 4869 19946 4903
rect 19880 4835 19896 4869
rect 19930 4835 19946 4869
rect 19880 4827 19946 4835
rect 19980 4937 20014 4953
rect 19980 4869 20014 4903
rect 19980 4793 20014 4835
rect 20048 4937 20114 4961
rect 20216 4959 20232 4987
rect 20266 4987 20395 4997
rect 20266 4959 20282 4987
rect 20048 4903 20064 4937
rect 20098 4903 20114 4937
rect 20048 4869 20114 4903
rect 20048 4835 20064 4869
rect 20098 4835 20114 4869
rect 20048 4827 20114 4835
rect 20148 4937 20182 4953
rect 20148 4869 20182 4903
rect 20148 4793 20182 4835
rect 20216 4937 20282 4959
rect 20384 4963 20395 4987
rect 20434 4973 20450 5007
rect 20429 4963 20450 4973
rect 20216 4903 20232 4937
rect 20266 4903 20282 4937
rect 20216 4869 20282 4903
rect 20216 4835 20232 4869
rect 20266 4835 20282 4869
rect 20216 4827 20282 4835
rect 20316 4937 20350 4953
rect 20316 4869 20350 4903
rect 20316 4793 20350 4835
rect 20384 4937 20450 4963
rect 20384 4903 20400 4937
rect 20434 4903 20450 4937
rect 20384 4869 20450 4903
rect 20384 4835 20400 4869
rect 20434 4835 20450 4869
rect 20384 4827 20450 4835
rect 20484 4937 20526 4953
rect 20518 4903 20526 4937
rect 20484 4869 20526 4903
rect 20518 4835 20526 4869
rect 20484 4793 20526 4835
rect 19092 4759 19121 4793
rect 19155 4759 19213 4793
rect 19247 4759 19305 4793
rect 19339 4759 19397 4793
rect 19431 4759 19489 4793
rect 19523 4759 19581 4793
rect 19615 4759 19673 4793
rect 19707 4759 19765 4793
rect 19799 4759 19857 4793
rect 19891 4759 19949 4793
rect 19983 4759 20041 4793
rect 20075 4759 20133 4793
rect 20167 4759 20225 4793
rect 20259 4759 20317 4793
rect 20351 4759 20409 4793
rect 20443 4759 20501 4793
rect 20535 4759 20564 4793
rect -3376 4715 -3314 4716
rect -2910 4715 -2520 4716
rect -1488 4715 -1426 4716
rect -1022 4715 -632 4716
rect 400 4715 462 4716
rect 866 4715 1256 4716
rect 2288 4715 2350 4716
rect 2754 4715 3144 4716
rect 4176 4715 4238 4716
rect 4642 4715 5032 4716
rect 6064 4715 6126 4716
rect 6530 4715 6920 4716
rect 7952 4715 8014 4716
rect 8418 4715 8808 4716
rect 9840 4715 9902 4716
rect 10306 4715 10696 4716
rect 11722 4715 11784 4716
rect 12188 4715 12578 4716
rect 13610 4715 13672 4716
rect 14076 4715 14466 4716
rect 15498 4715 15560 4716
rect 15964 4715 16354 4716
rect 17386 4715 17448 4716
rect 17852 4715 18242 4716
rect 19274 4715 19336 4716
rect 19740 4715 20130 4716
rect 21162 4715 21224 4716
rect 21628 4715 22018 4716
rect 23050 4715 23112 4716
rect 23516 4715 23906 4716
rect 24938 4715 25000 4716
rect 25404 4715 25794 4716
rect -3376 4682 -3305 4715
rect -3334 4681 -3305 4682
rect -3271 4681 -3213 4715
rect -3179 4681 -3121 4715
rect -3087 4681 -2491 4715
rect -2457 4681 -2399 4715
rect -2365 4681 -2307 4715
rect -2273 4681 -2244 4715
rect -1488 4682 -1417 4715
rect -1446 4681 -1417 4682
rect -1383 4681 -1325 4715
rect -1291 4681 -1233 4715
rect -1199 4681 -603 4715
rect -569 4681 -511 4715
rect -477 4681 -419 4715
rect -385 4681 -356 4715
rect 400 4682 471 4715
rect 442 4681 471 4682
rect 505 4681 563 4715
rect 597 4681 655 4715
rect 689 4681 1285 4715
rect 1319 4681 1377 4715
rect 1411 4681 1469 4715
rect 1503 4681 1532 4715
rect 2288 4682 2359 4715
rect 2330 4681 2359 4682
rect 2393 4681 2451 4715
rect 2485 4681 2543 4715
rect 2577 4681 3173 4715
rect 3207 4681 3265 4715
rect 3299 4681 3357 4715
rect 3391 4681 3420 4715
rect 4176 4682 4247 4715
rect 4218 4681 4247 4682
rect 4281 4681 4339 4715
rect 4373 4681 4431 4715
rect 4465 4681 5061 4715
rect 5095 4681 5153 4715
rect 5187 4681 5245 4715
rect 5279 4681 5308 4715
rect 6064 4682 6135 4715
rect 6106 4681 6135 4682
rect 6169 4681 6227 4715
rect 6261 4681 6319 4715
rect 6353 4681 6949 4715
rect 6983 4681 7041 4715
rect 7075 4681 7133 4715
rect 7167 4681 7196 4715
rect 7952 4682 8023 4715
rect 7994 4681 8023 4682
rect 8057 4681 8115 4715
rect 8149 4681 8207 4715
rect 8241 4681 8837 4715
rect 8871 4681 8929 4715
rect 8963 4681 9021 4715
rect 9055 4681 9084 4715
rect 9840 4682 9911 4715
rect 9882 4681 9911 4682
rect 9945 4681 10003 4715
rect 10037 4681 10095 4715
rect 10129 4681 10725 4715
rect 10759 4681 10817 4715
rect 10851 4681 10909 4715
rect 10943 4681 10972 4715
rect 11722 4682 11793 4715
rect 11764 4681 11793 4682
rect 11827 4681 11885 4715
rect 11919 4681 11977 4715
rect 12011 4681 12607 4715
rect 12641 4681 12699 4715
rect 12733 4681 12791 4715
rect 12825 4681 12854 4715
rect 13610 4682 13681 4715
rect 13652 4681 13681 4682
rect 13715 4681 13773 4715
rect 13807 4681 13865 4715
rect 13899 4681 14495 4715
rect 14529 4681 14587 4715
rect 14621 4681 14679 4715
rect 14713 4681 14742 4715
rect 15498 4682 15569 4715
rect 15540 4681 15569 4682
rect 15603 4681 15661 4715
rect 15695 4681 15753 4715
rect 15787 4681 16383 4715
rect 16417 4681 16475 4715
rect 16509 4681 16567 4715
rect 16601 4681 16630 4715
rect 17386 4682 17457 4715
rect 17428 4681 17457 4682
rect 17491 4681 17549 4715
rect 17583 4681 17641 4715
rect 17675 4681 18271 4715
rect 18305 4681 18363 4715
rect 18397 4681 18455 4715
rect 18489 4681 18518 4715
rect 19274 4682 19345 4715
rect 19316 4681 19345 4682
rect 19379 4681 19437 4715
rect 19471 4681 19529 4715
rect 19563 4681 20159 4715
rect 20193 4681 20251 4715
rect 20285 4681 20343 4715
rect 20377 4681 20406 4715
rect 21162 4682 21233 4715
rect 21204 4681 21233 4682
rect 21267 4681 21325 4715
rect 21359 4681 21417 4715
rect 21451 4681 22047 4715
rect 22081 4681 22139 4715
rect 22173 4681 22231 4715
rect 22265 4681 22294 4715
rect 23050 4682 23121 4715
rect 23092 4681 23121 4682
rect 23155 4681 23213 4715
rect 23247 4681 23305 4715
rect 23339 4681 23935 4715
rect 23969 4681 24027 4715
rect 24061 4681 24119 4715
rect 24153 4681 24182 4715
rect 24938 4682 25009 4715
rect 24980 4681 25009 4682
rect 25043 4681 25101 4715
rect 25135 4681 25193 4715
rect 25227 4681 25823 4715
rect 25857 4681 25915 4715
rect 25949 4681 26007 4715
rect 26041 4681 26070 4715
rect -3315 4639 -3249 4644
rect -3315 4605 -3299 4639
rect -3265 4605 -3249 4639
rect -3315 4571 -3249 4605
rect -3315 4537 -3299 4571
rect -3265 4537 -3249 4571
rect -3315 4503 -3249 4537
rect -3315 4469 -3299 4503
rect -3265 4487 -3249 4503
rect -3143 4639 -3077 4681
rect -3109 4605 -3077 4639
rect -2910 4675 -2628 4681
rect -2910 4641 -2871 4675
rect -2837 4673 -2628 4675
rect -2837 4641 -2752 4673
rect -2910 4639 -2752 4641
rect -2718 4639 -2628 4673
rect -2910 4606 -2628 4639
rect -2501 4639 -2435 4644
rect -3143 4571 -3077 4605
rect -3109 4537 -3077 4571
rect -2501 4605 -2485 4639
rect -2451 4605 -2435 4639
rect -2501 4571 -2435 4605
rect -3143 4503 -3077 4537
rect -3265 4469 -3179 4487
rect -3315 4453 -3179 4469
rect -3109 4469 -3077 4503
rect -3143 4453 -3077 4469
rect -3018 4567 -2752 4568
rect -3018 4533 -2802 4567
rect -2768 4533 -2752 4567
rect -3018 4532 -2752 4533
rect -3317 4412 -3247 4419
rect -3317 4378 -3299 4412
rect -3265 4403 -3247 4412
rect -3317 4369 -3297 4378
rect -3263 4369 -3247 4403
rect -3213 4333 -3179 4453
rect -3145 4408 -3075 4419
rect -3145 4403 -3126 4408
rect -3145 4369 -3129 4403
rect -3092 4374 -3075 4408
rect -3095 4369 -3075 4374
rect -3313 4317 -3265 4333
rect -3313 4283 -3299 4317
rect -3313 4249 -3265 4283
rect -3313 4215 -3299 4249
rect -3313 4171 -3265 4215
rect -3231 4317 -3165 4333
rect -3231 4292 -3215 4317
rect -3231 4258 -3217 4292
rect -3181 4283 -3165 4317
rect -3183 4258 -3165 4283
rect -3231 4249 -3165 4258
rect -3231 4215 -3215 4249
rect -3181 4215 -3165 4249
rect -3231 4205 -3165 4215
rect -3131 4317 -3077 4333
rect -3097 4283 -3077 4317
rect -3131 4249 -3077 4283
rect -3097 4215 -3077 4249
rect -3131 4171 -3077 4215
rect -3334 4137 -3305 4171
rect -3271 4137 -3213 4171
rect -3179 4137 -3121 4171
rect -3087 4137 -3058 4171
rect -3334 3926 -3300 4137
rect -3103 3834 -3069 4137
rect -3018 3918 -2984 4532
rect -2818 4530 -2752 4532
rect -2501 4537 -2485 4571
rect -2451 4537 -2435 4571
rect -2501 4503 -2435 4537
rect -2946 4471 -2912 4490
rect -2946 4403 -2912 4405
rect -2946 4367 -2912 4369
rect -2946 4282 -2912 4301
rect -2850 4471 -2816 4490
rect -2850 4403 -2816 4405
rect -2850 4367 -2816 4369
rect -2850 4282 -2816 4301
rect -2754 4471 -2720 4490
rect -2501 4469 -2485 4503
rect -2451 4487 -2435 4503
rect -2329 4639 -2263 4681
rect -2295 4605 -2263 4639
rect -2329 4571 -2263 4605
rect -2295 4537 -2263 4571
rect -2329 4503 -2263 4537
rect -2451 4469 -2365 4487
rect -2501 4453 -2365 4469
rect -2295 4469 -2263 4503
rect -2329 4453 -2263 4469
rect -1427 4639 -1361 4644
rect -1427 4605 -1411 4639
rect -1377 4605 -1361 4639
rect -1427 4571 -1361 4605
rect -1427 4537 -1411 4571
rect -1377 4537 -1361 4571
rect -1427 4503 -1361 4537
rect -1427 4469 -1411 4503
rect -1377 4487 -1361 4503
rect -1255 4639 -1189 4681
rect -1221 4605 -1189 4639
rect -1022 4675 -740 4681
rect -1022 4641 -983 4675
rect -949 4673 -740 4675
rect -949 4641 -864 4673
rect -1022 4639 -864 4641
rect -830 4639 -740 4673
rect -1022 4606 -740 4639
rect -613 4639 -547 4644
rect -1255 4571 -1189 4605
rect -1221 4537 -1189 4571
rect -613 4605 -597 4639
rect -563 4605 -547 4639
rect -613 4571 -547 4605
rect -1255 4503 -1189 4537
rect -1377 4469 -1291 4487
rect -1427 4453 -1291 4469
rect -1221 4469 -1189 4503
rect -1255 4453 -1189 4469
rect -1130 4567 -864 4568
rect -1130 4533 -914 4567
rect -880 4533 -864 4567
rect -1130 4532 -864 4533
rect -2754 4403 -2720 4405
rect -2503 4410 -2433 4419
rect -2503 4376 -2487 4410
rect -2453 4403 -2433 4410
rect -2503 4369 -2483 4376
rect -2449 4369 -2433 4403
rect -2754 4367 -2720 4369
rect -2399 4333 -2365 4453
rect -2331 4410 -2261 4419
rect -2331 4403 -2313 4410
rect -2331 4369 -2315 4403
rect -2279 4376 -2261 4410
rect -2281 4369 -2261 4376
rect -1429 4412 -1359 4419
rect -1429 4378 -1411 4412
rect -1377 4403 -1359 4412
rect -1429 4369 -1409 4378
rect -1375 4369 -1359 4403
rect -1325 4333 -1291 4453
rect -1257 4408 -1187 4419
rect -1257 4403 -1238 4408
rect -1257 4369 -1241 4403
rect -1204 4374 -1187 4408
rect -1207 4369 -1187 4374
rect -2754 4282 -2720 4301
rect -2499 4317 -2451 4333
rect -2499 4283 -2485 4317
rect -2499 4249 -2451 4283
rect -2914 4205 -2898 4239
rect -2864 4205 -2848 4239
rect -2499 4215 -2485 4249
rect -2499 4171 -2451 4215
rect -2417 4317 -2351 4333
rect -2417 4283 -2401 4317
rect -2367 4287 -2351 4317
rect -2417 4253 -2399 4283
rect -2365 4253 -2351 4287
rect -2417 4249 -2351 4253
rect -2417 4215 -2401 4249
rect -2367 4215 -2351 4249
rect -2417 4205 -2351 4215
rect -2317 4317 -2263 4333
rect -2283 4283 -2263 4317
rect -2317 4249 -2263 4283
rect -2283 4215 -2263 4249
rect -2317 4171 -2263 4215
rect -1425 4317 -1377 4333
rect -1425 4283 -1411 4317
rect -1425 4249 -1377 4283
rect -1425 4215 -1411 4249
rect -1425 4171 -1377 4215
rect -1343 4317 -1277 4333
rect -1343 4292 -1327 4317
rect -1343 4258 -1329 4292
rect -1293 4283 -1277 4317
rect -1295 4258 -1277 4283
rect -1343 4249 -1277 4258
rect -1343 4215 -1327 4249
rect -1293 4215 -1277 4249
rect -1343 4205 -1277 4215
rect -1243 4317 -1189 4333
rect -1209 4283 -1189 4317
rect -1243 4249 -1189 4283
rect -1209 4215 -1189 4249
rect -1243 4171 -1189 4215
rect -2802 4124 -2786 4158
rect -2752 4124 -2736 4158
rect -2520 4137 -2491 4171
rect -2457 4137 -2399 4171
rect -2365 4137 -2307 4171
rect -2273 4137 -2244 4171
rect -1446 4137 -1417 4171
rect -1383 4137 -1325 4171
rect -1291 4137 -1233 4171
rect -1199 4137 -1170 4171
rect -2930 4074 -2896 4090
rect -2930 4004 -2896 4038
rect -2930 3952 -2896 3968
rect -2834 4074 -2800 4090
rect -2834 4004 -2800 4038
rect -2834 3952 -2800 3968
rect -2738 4074 -2704 4090
rect -2738 4004 -2704 4038
rect -2704 3968 -2356 3992
rect -2738 3952 -2356 3968
rect -3018 3884 -2882 3918
rect -2848 3884 -2832 3918
rect -3103 3814 -2708 3834
rect -3103 3809 -2841 3814
rect -3103 3800 -2962 3809
rect -2978 3775 -2962 3800
rect -2928 3780 -2841 3809
rect -2807 3790 -2708 3814
rect -2536 3792 -2490 3794
rect -2536 3790 -2532 3792
rect -2807 3780 -2532 3790
rect -2928 3775 -2532 3780
rect -2978 3758 -2532 3775
rect -2498 3758 -2490 3792
rect -2978 3756 -2490 3758
rect -2536 3750 -2490 3756
rect -3437 3661 -3403 3668
rect -3512 3627 -3483 3661
rect -3449 3627 -3391 3661
rect -3357 3627 -3299 3661
rect -3265 3627 -3236 3661
rect -3136 3637 -3120 3671
rect -3086 3637 -3070 3671
rect -2912 3658 -2798 3660
rect -3444 3585 -3402 3627
rect -2912 3619 -2630 3658
rect -2490 3637 -2474 3671
rect -2440 3637 -2424 3671
rect -2912 3594 -2873 3619
rect -3444 3551 -3436 3585
rect -3444 3517 -3402 3551
rect -3444 3483 -3436 3517
rect -3444 3449 -3402 3483
rect -3444 3415 -3436 3449
rect -3444 3399 -3402 3415
rect -3368 3585 -3302 3593
rect -3368 3551 -3352 3585
rect -3318 3551 -3302 3585
rect -3368 3517 -3302 3551
rect -3368 3483 -3352 3517
rect -3318 3483 -3302 3517
rect -3368 3449 -3302 3483
rect -3368 3415 -3352 3449
rect -3318 3415 -3302 3449
rect -3368 3397 -3302 3415
rect -3448 3360 -3382 3363
rect -3448 3326 -3434 3360
rect -3400 3349 -3382 3360
rect -3448 3315 -3432 3326
rect -3398 3315 -3382 3349
rect -3448 3265 -3402 3281
rect -3348 3277 -3302 3397
rect -3164 3575 -3130 3594
rect -3078 3585 -2873 3594
rect -2839 3617 -2630 3619
rect -2839 3585 -2754 3617
rect -3078 3583 -2754 3585
rect -2720 3594 -2630 3617
rect -2390 3594 -2356 3952
rect -1446 3926 -1412 4137
rect -1215 3834 -1181 4137
rect -1130 3918 -1096 4532
rect -930 4530 -864 4532
rect -613 4537 -597 4571
rect -563 4537 -547 4571
rect -613 4503 -547 4537
rect -1058 4471 -1024 4490
rect -1058 4403 -1024 4405
rect -1058 4367 -1024 4369
rect -1058 4282 -1024 4301
rect -962 4471 -928 4490
rect -962 4403 -928 4405
rect -962 4367 -928 4369
rect -962 4282 -928 4301
rect -866 4471 -832 4490
rect -613 4469 -597 4503
rect -563 4487 -547 4503
rect -441 4639 -375 4681
rect -407 4605 -375 4639
rect -441 4571 -375 4605
rect -407 4537 -375 4571
rect -441 4503 -375 4537
rect -563 4469 -477 4487
rect -613 4453 -477 4469
rect -407 4469 -375 4503
rect -441 4453 -375 4469
rect 461 4639 527 4644
rect 461 4605 477 4639
rect 511 4605 527 4639
rect 461 4571 527 4605
rect 461 4537 477 4571
rect 511 4537 527 4571
rect 461 4503 527 4537
rect 461 4469 477 4503
rect 511 4487 527 4503
rect 633 4639 699 4681
rect 667 4605 699 4639
rect 866 4675 1148 4681
rect 866 4641 905 4675
rect 939 4673 1148 4675
rect 939 4641 1024 4673
rect 866 4639 1024 4641
rect 1058 4639 1148 4673
rect 866 4606 1148 4639
rect 1275 4639 1341 4644
rect 633 4571 699 4605
rect 667 4537 699 4571
rect 1275 4605 1291 4639
rect 1325 4605 1341 4639
rect 1275 4571 1341 4605
rect 633 4503 699 4537
rect 511 4469 597 4487
rect 461 4453 597 4469
rect 667 4469 699 4503
rect 633 4453 699 4469
rect 758 4567 1024 4568
rect 758 4533 974 4567
rect 1008 4533 1024 4567
rect 758 4532 1024 4533
rect -866 4403 -832 4405
rect -615 4410 -545 4419
rect -615 4376 -599 4410
rect -565 4403 -545 4410
rect -615 4369 -595 4376
rect -561 4369 -545 4403
rect -866 4367 -832 4369
rect -511 4333 -477 4453
rect -443 4410 -373 4419
rect -443 4403 -425 4410
rect -443 4369 -427 4403
rect -391 4376 -373 4410
rect -393 4369 -373 4376
rect 459 4412 529 4419
rect 459 4378 477 4412
rect 511 4403 529 4412
rect 459 4369 479 4378
rect 513 4369 529 4403
rect 563 4333 597 4453
rect 631 4408 701 4419
rect 631 4403 650 4408
rect 631 4369 647 4403
rect 684 4374 701 4408
rect 681 4369 701 4374
rect -866 4282 -832 4301
rect -611 4317 -563 4333
rect -611 4283 -597 4317
rect -611 4249 -563 4283
rect -1026 4205 -1010 4239
rect -976 4205 -960 4239
rect -611 4215 -597 4249
rect -611 4171 -563 4215
rect -529 4317 -463 4333
rect -529 4283 -513 4317
rect -479 4287 -463 4317
rect -529 4253 -511 4283
rect -477 4253 -463 4287
rect -529 4249 -463 4253
rect -529 4215 -513 4249
rect -479 4215 -463 4249
rect -529 4205 -463 4215
rect -429 4317 -375 4333
rect -395 4283 -375 4317
rect -429 4249 -375 4283
rect -395 4215 -375 4249
rect -429 4171 -375 4215
rect 463 4317 511 4333
rect 463 4283 477 4317
rect 463 4249 511 4283
rect 463 4215 477 4249
rect 463 4171 511 4215
rect 545 4317 611 4333
rect 545 4292 561 4317
rect 545 4258 559 4292
rect 595 4283 611 4317
rect 593 4258 611 4283
rect 545 4249 611 4258
rect 545 4215 561 4249
rect 595 4215 611 4249
rect 545 4205 611 4215
rect 645 4317 699 4333
rect 679 4283 699 4317
rect 645 4249 699 4283
rect 679 4215 699 4249
rect 645 4171 699 4215
rect -914 4124 -898 4158
rect -864 4124 -848 4158
rect -632 4137 -603 4171
rect -569 4137 -511 4171
rect -477 4137 -419 4171
rect -385 4137 -356 4171
rect 442 4137 471 4171
rect 505 4137 563 4171
rect 597 4137 655 4171
rect 689 4137 718 4171
rect -1042 4074 -1008 4090
rect -1042 4004 -1008 4038
rect -1042 3952 -1008 3968
rect -946 4074 -912 4090
rect -946 4004 -912 4038
rect -946 3952 -912 3968
rect -850 4074 -816 4090
rect -850 4004 -816 4038
rect -816 3968 -468 3992
rect -850 3952 -468 3968
rect -1130 3884 -994 3918
rect -960 3884 -944 3918
rect -1215 3814 -820 3834
rect -1215 3809 -953 3814
rect -1215 3800 -1074 3809
rect -1090 3775 -1074 3800
rect -1040 3780 -953 3809
rect -919 3790 -820 3814
rect -648 3792 -602 3794
rect -648 3790 -644 3792
rect -919 3780 -644 3790
rect -1040 3775 -644 3780
rect -1090 3758 -644 3775
rect -610 3758 -602 3792
rect -1090 3756 -602 3758
rect -648 3750 -602 3756
rect -2316 3635 -2287 3669
rect -2253 3635 -2195 3669
rect -2161 3635 -2103 3669
rect -2069 3635 -2040 3669
rect -2720 3583 -2484 3594
rect -3078 3575 -2484 3583
rect -3078 3550 -3076 3575
rect -3164 3507 -3130 3509
rect -3164 3471 -3130 3473
rect -3164 3386 -3130 3405
rect -3042 3550 -2518 3575
rect -2432 3575 -2356 3594
rect -2432 3554 -2430 3575
rect -3076 3507 -3042 3509
rect -2820 3477 -2804 3511
rect -2770 3477 -2754 3511
rect -2518 3507 -2484 3509
rect -3076 3471 -3042 3473
rect -2518 3471 -2484 3473
rect -3076 3386 -3042 3405
rect -2948 3415 -2914 3434
rect -2948 3347 -2914 3349
rect -3136 3309 -3120 3343
rect -3086 3309 -3070 3343
rect -2948 3311 -2914 3313
rect -3448 3231 -3436 3265
rect -3448 3197 -3402 3231
rect -3448 3163 -3436 3197
rect -3448 3117 -3402 3163
rect -3368 3265 -3302 3277
rect -3368 3231 -3352 3265
rect -3318 3231 -3302 3265
rect -3368 3218 -3302 3231
rect -2948 3226 -2914 3245
rect -2852 3415 -2818 3434
rect -2852 3347 -2818 3349
rect -2852 3311 -2818 3313
rect -2852 3226 -2818 3245
rect -2756 3415 -2722 3434
rect -2518 3386 -2484 3405
rect -2396 3554 -2356 3575
rect -2248 3593 -2206 3635
rect -1970 3633 -1941 3667
rect -1907 3633 -1849 3667
rect -1815 3633 -1757 3667
rect -1723 3633 -1694 3667
rect -1549 3661 -1515 3668
rect -2248 3559 -2240 3593
rect -2430 3507 -2396 3509
rect -2430 3471 -2396 3473
rect -2248 3525 -2206 3559
rect -2248 3491 -2240 3525
rect -2248 3457 -2206 3491
rect -2248 3423 -2240 3457
rect -2248 3407 -2206 3423
rect -2172 3593 -2106 3601
rect -2172 3559 -2156 3593
rect -2122 3559 -2106 3593
rect -2172 3525 -2106 3559
rect -2172 3491 -2156 3525
rect -2122 3491 -2106 3525
rect -2172 3457 -2106 3491
rect -2172 3423 -2156 3457
rect -2122 3423 -2106 3457
rect -2172 3405 -2106 3423
rect -1937 3583 -1901 3599
rect -1937 3549 -1935 3583
rect -1937 3515 -1901 3549
rect -1937 3481 -1935 3515
rect -1865 3583 -1799 3633
rect -1624 3627 -1595 3661
rect -1561 3627 -1503 3661
rect -1469 3627 -1411 3661
rect -1377 3627 -1348 3661
rect -1248 3637 -1232 3671
rect -1198 3637 -1182 3671
rect -1024 3658 -910 3660
rect -1865 3549 -1849 3583
rect -1815 3549 -1799 3583
rect -1865 3515 -1799 3549
rect -1865 3481 -1849 3515
rect -1815 3481 -1799 3515
rect -1765 3583 -1711 3599
rect -1765 3549 -1763 3583
rect -1729 3549 -1711 3583
rect -1765 3502 -1711 3549
rect -1937 3447 -1901 3481
rect -1765 3468 -1763 3502
rect -1729 3468 -1711 3502
rect -1937 3413 -1802 3447
rect -1765 3418 -1711 3468
rect -2430 3386 -2396 3405
rect -2756 3347 -2722 3349
rect -2344 3371 -2200 3372
rect -2344 3357 -2186 3371
rect -2756 3311 -2722 3313
rect -2490 3344 -2424 3346
rect -2344 3344 -2236 3357
rect -2490 3343 -2236 3344
rect -2490 3309 -2474 3343
rect -2440 3330 -2236 3343
rect -2440 3310 -2304 3330
rect -2252 3323 -2236 3330
rect -2202 3323 -2186 3357
rect -2440 3309 -2424 3310
rect -2252 3273 -2206 3289
rect -2152 3285 -2106 3405
rect -1836 3384 -1802 3413
rect -1949 3355 -1881 3377
rect -1949 3354 -1933 3355
rect -1949 3320 -1935 3354
rect -1899 3321 -1881 3355
rect -1901 3320 -1881 3321
rect -1949 3303 -1881 3320
rect -1836 3368 -1781 3384
rect -1836 3334 -1815 3368
rect -1836 3318 -1781 3334
rect -1747 3368 -1711 3418
rect -1556 3585 -1514 3627
rect -1024 3619 -742 3658
rect -602 3637 -586 3671
rect -552 3637 -536 3671
rect -1024 3594 -985 3619
rect -1556 3551 -1548 3585
rect -1556 3517 -1514 3551
rect -1556 3483 -1548 3517
rect -1556 3449 -1514 3483
rect -1556 3415 -1548 3449
rect -1556 3399 -1514 3415
rect -1480 3585 -1414 3593
rect -1480 3551 -1464 3585
rect -1430 3551 -1414 3585
rect -1480 3517 -1414 3551
rect -1480 3483 -1464 3517
rect -1430 3483 -1414 3517
rect -1480 3449 -1414 3483
rect -1480 3415 -1464 3449
rect -1430 3415 -1414 3449
rect -1480 3397 -1414 3415
rect -1747 3366 -1706 3368
rect -1747 3332 -1742 3366
rect -1708 3332 -1706 3366
rect -1747 3330 -1706 3332
rect -1560 3360 -1494 3363
rect -2722 3245 -2476 3262
rect -2756 3228 -2476 3245
rect -2756 3226 -2722 3228
rect -3368 3197 -3026 3218
rect -3368 3163 -3352 3197
rect -3318 3186 -3026 3197
rect -3318 3183 -2850 3186
rect -3318 3182 -2900 3183
rect -3318 3163 -3296 3182
rect -3368 3158 -3296 3163
rect -3368 3151 -3302 3158
rect -3062 3150 -2900 3182
rect -2916 3149 -2900 3150
rect -2866 3149 -2850 3183
rect -2524 3140 -2476 3228
rect -3512 3083 -3483 3117
rect -3449 3083 -3391 3117
rect -3357 3083 -3299 3117
rect -3265 3083 -3236 3117
rect -3154 3112 -3108 3122
rect -3154 3078 -3148 3112
rect -3114 3092 -3108 3112
rect -2524 3106 -2516 3140
rect -2482 3106 -2476 3140
rect -2252 3239 -2240 3273
rect -2252 3205 -2206 3239
rect -2252 3171 -2240 3205
rect -2252 3125 -2206 3171
rect -2172 3273 -2106 3285
rect -2172 3222 -2156 3273
rect -2122 3222 -2106 3273
rect -1836 3267 -1802 3318
rect -2172 3205 -2106 3222
rect -2172 3171 -2156 3205
rect -2122 3171 -2106 3205
rect -2172 3159 -2106 3171
rect -1935 3233 -1802 3267
rect -1747 3258 -1711 3330
rect -1560 3326 -1546 3360
rect -1512 3349 -1494 3360
rect -1560 3315 -1544 3326
rect -1510 3315 -1494 3349
rect -1935 3212 -1901 3233
rect -1763 3229 -1711 3258
rect -1935 3157 -1901 3178
rect -1865 3165 -1849 3199
rect -1815 3165 -1799 3199
rect -3114 3078 -3104 3092
rect -3154 3008 -3104 3078
rect -2804 3068 -2788 3102
rect -2754 3068 -2738 3102
rect -2524 3094 -2476 3106
rect -2316 3091 -2287 3125
rect -2253 3091 -2195 3125
rect -2161 3091 -2103 3125
rect -2069 3091 -2040 3125
rect -1865 3123 -1799 3165
rect -1729 3195 -1711 3229
rect -1763 3157 -1711 3195
rect -1560 3265 -1514 3281
rect -1460 3277 -1414 3397
rect -1276 3575 -1242 3594
rect -1190 3585 -985 3594
rect -951 3617 -742 3619
rect -951 3585 -866 3617
rect -1190 3583 -866 3585
rect -832 3594 -742 3617
rect -502 3594 -468 3952
rect 442 3926 476 4137
rect 673 3834 707 4137
rect 758 3918 792 4532
rect 958 4530 1024 4532
rect 1275 4537 1291 4571
rect 1325 4537 1341 4571
rect 1275 4503 1341 4537
rect 830 4471 864 4490
rect 830 4403 864 4405
rect 830 4367 864 4369
rect 830 4282 864 4301
rect 926 4471 960 4490
rect 926 4403 960 4405
rect 926 4367 960 4369
rect 926 4282 960 4301
rect 1022 4471 1056 4490
rect 1275 4469 1291 4503
rect 1325 4487 1341 4503
rect 1447 4639 1513 4681
rect 1481 4605 1513 4639
rect 1447 4571 1513 4605
rect 1481 4537 1513 4571
rect 1447 4503 1513 4537
rect 1325 4469 1411 4487
rect 1275 4453 1411 4469
rect 1481 4469 1513 4503
rect 1447 4453 1513 4469
rect 2349 4639 2415 4644
rect 2349 4605 2365 4639
rect 2399 4605 2415 4639
rect 2349 4571 2415 4605
rect 2349 4537 2365 4571
rect 2399 4537 2415 4571
rect 2349 4503 2415 4537
rect 2349 4469 2365 4503
rect 2399 4487 2415 4503
rect 2521 4639 2587 4681
rect 2555 4605 2587 4639
rect 2754 4675 3036 4681
rect 2754 4641 2793 4675
rect 2827 4673 3036 4675
rect 2827 4641 2912 4673
rect 2754 4639 2912 4641
rect 2946 4639 3036 4673
rect 2754 4606 3036 4639
rect 3163 4639 3229 4644
rect 2521 4571 2587 4605
rect 2555 4537 2587 4571
rect 3163 4605 3179 4639
rect 3213 4605 3229 4639
rect 3163 4571 3229 4605
rect 2521 4503 2587 4537
rect 2399 4469 2485 4487
rect 2349 4453 2485 4469
rect 2555 4469 2587 4503
rect 2521 4453 2587 4469
rect 2646 4567 2912 4568
rect 2646 4533 2862 4567
rect 2896 4533 2912 4567
rect 2646 4532 2912 4533
rect 1022 4403 1056 4405
rect 1273 4410 1343 4419
rect 1273 4376 1289 4410
rect 1323 4403 1343 4410
rect 1273 4369 1293 4376
rect 1327 4369 1343 4403
rect 1022 4367 1056 4369
rect 1377 4333 1411 4453
rect 1445 4410 1515 4419
rect 1445 4403 1463 4410
rect 1445 4369 1461 4403
rect 1497 4376 1515 4410
rect 1495 4369 1515 4376
rect 2347 4412 2417 4419
rect 2347 4378 2365 4412
rect 2399 4403 2417 4412
rect 2347 4369 2367 4378
rect 2401 4369 2417 4403
rect 2451 4333 2485 4453
rect 2519 4408 2589 4419
rect 2519 4403 2538 4408
rect 2519 4369 2535 4403
rect 2572 4374 2589 4408
rect 2569 4369 2589 4374
rect 1022 4282 1056 4301
rect 1277 4317 1325 4333
rect 1277 4283 1291 4317
rect 1277 4249 1325 4283
rect 862 4205 878 4239
rect 912 4205 928 4239
rect 1277 4215 1291 4249
rect 1277 4171 1325 4215
rect 1359 4317 1425 4333
rect 1359 4283 1375 4317
rect 1409 4287 1425 4317
rect 1359 4253 1377 4283
rect 1411 4253 1425 4287
rect 1359 4249 1425 4253
rect 1359 4215 1375 4249
rect 1409 4215 1425 4249
rect 1359 4205 1425 4215
rect 1459 4317 1513 4333
rect 1493 4283 1513 4317
rect 1459 4249 1513 4283
rect 1493 4215 1513 4249
rect 1459 4171 1513 4215
rect 2351 4317 2399 4333
rect 2351 4283 2365 4317
rect 2351 4249 2399 4283
rect 2351 4215 2365 4249
rect 2351 4171 2399 4215
rect 2433 4317 2499 4333
rect 2433 4292 2449 4317
rect 2433 4258 2447 4292
rect 2483 4283 2499 4317
rect 2481 4258 2499 4283
rect 2433 4249 2499 4258
rect 2433 4215 2449 4249
rect 2483 4215 2499 4249
rect 2433 4205 2499 4215
rect 2533 4317 2587 4333
rect 2567 4283 2587 4317
rect 2533 4249 2587 4283
rect 2567 4215 2587 4249
rect 2533 4171 2587 4215
rect 974 4124 990 4158
rect 1024 4124 1040 4158
rect 1256 4137 1285 4171
rect 1319 4137 1377 4171
rect 1411 4137 1469 4171
rect 1503 4137 1532 4171
rect 2330 4137 2359 4171
rect 2393 4137 2451 4171
rect 2485 4137 2543 4171
rect 2577 4137 2606 4171
rect 846 4074 880 4090
rect 846 4004 880 4038
rect 846 3952 880 3968
rect 942 4074 976 4090
rect 942 4004 976 4038
rect 942 3952 976 3968
rect 1038 4074 1072 4090
rect 1038 4004 1072 4038
rect 1072 3968 1420 3992
rect 1038 3952 1420 3968
rect 758 3884 894 3918
rect 928 3884 944 3918
rect 673 3814 1068 3834
rect 673 3809 935 3814
rect 673 3800 814 3809
rect 798 3775 814 3800
rect 848 3780 935 3809
rect 969 3790 1068 3814
rect 1240 3792 1286 3794
rect 1240 3790 1244 3792
rect 969 3780 1244 3790
rect 848 3775 1244 3780
rect 798 3758 1244 3775
rect 1278 3758 1286 3792
rect 798 3756 1286 3758
rect 1240 3750 1286 3756
rect -428 3635 -399 3669
rect -365 3635 -307 3669
rect -273 3635 -215 3669
rect -181 3635 -152 3669
rect -832 3583 -596 3594
rect -1190 3575 -596 3583
rect -1190 3550 -1188 3575
rect -1276 3507 -1242 3509
rect -1276 3471 -1242 3473
rect -1276 3386 -1242 3405
rect -1154 3550 -630 3575
rect -544 3575 -468 3594
rect -544 3554 -542 3575
rect -1188 3507 -1154 3509
rect -932 3477 -916 3511
rect -882 3477 -866 3511
rect -630 3507 -596 3509
rect -1188 3471 -1154 3473
rect -630 3471 -596 3473
rect -1188 3386 -1154 3405
rect -1060 3415 -1026 3434
rect -1060 3347 -1026 3349
rect -1248 3309 -1232 3343
rect -1198 3309 -1182 3343
rect -1060 3311 -1026 3313
rect -1560 3231 -1548 3265
rect -1560 3197 -1514 3231
rect -1560 3163 -1548 3197
rect -1970 3089 -1941 3123
rect -1907 3089 -1849 3123
rect -1815 3089 -1757 3123
rect -1723 3089 -1694 3123
rect -1560 3117 -1514 3163
rect -1480 3265 -1414 3277
rect -1480 3231 -1464 3265
rect -1430 3231 -1414 3265
rect -1480 3218 -1414 3231
rect -1060 3226 -1026 3245
rect -964 3415 -930 3434
rect -964 3347 -930 3349
rect -964 3311 -930 3313
rect -964 3226 -930 3245
rect -868 3415 -834 3434
rect -630 3386 -596 3405
rect -508 3554 -468 3575
rect -360 3593 -318 3635
rect -82 3633 -53 3667
rect -19 3633 39 3667
rect 73 3633 131 3667
rect 165 3633 194 3667
rect 339 3661 373 3668
rect -360 3559 -352 3593
rect -542 3507 -508 3509
rect -542 3471 -508 3473
rect -360 3525 -318 3559
rect -360 3491 -352 3525
rect -360 3457 -318 3491
rect -360 3423 -352 3457
rect -360 3407 -318 3423
rect -284 3593 -218 3601
rect -284 3559 -268 3593
rect -234 3559 -218 3593
rect -284 3525 -218 3559
rect -284 3491 -268 3525
rect -234 3491 -218 3525
rect -284 3457 -218 3491
rect -284 3423 -268 3457
rect -234 3423 -218 3457
rect -284 3405 -218 3423
rect -49 3583 -13 3599
rect -49 3549 -47 3583
rect -49 3515 -13 3549
rect -49 3481 -47 3515
rect 23 3583 89 3633
rect 264 3627 293 3661
rect 327 3627 385 3661
rect 419 3627 477 3661
rect 511 3627 540 3661
rect 640 3637 656 3671
rect 690 3637 706 3671
rect 864 3658 978 3660
rect 23 3549 39 3583
rect 73 3549 89 3583
rect 23 3515 89 3549
rect 23 3481 39 3515
rect 73 3481 89 3515
rect 123 3583 177 3599
rect 123 3549 125 3583
rect 159 3549 177 3583
rect 123 3502 177 3549
rect -49 3447 -13 3481
rect 123 3468 125 3502
rect 159 3468 177 3502
rect -49 3413 86 3447
rect 123 3418 177 3468
rect -542 3386 -508 3405
rect -868 3347 -834 3349
rect -456 3371 -312 3372
rect -456 3357 -298 3371
rect -868 3311 -834 3313
rect -602 3344 -536 3346
rect -456 3344 -348 3357
rect -602 3343 -348 3344
rect -602 3309 -586 3343
rect -552 3330 -348 3343
rect -552 3310 -416 3330
rect -364 3323 -348 3330
rect -314 3323 -298 3357
rect -552 3309 -536 3310
rect -364 3273 -318 3289
rect -264 3285 -218 3405
rect 52 3384 86 3413
rect -61 3355 7 3377
rect -61 3354 -45 3355
rect -61 3320 -47 3354
rect -11 3321 7 3355
rect -13 3320 7 3321
rect -61 3303 7 3320
rect 52 3368 107 3384
rect 52 3334 73 3368
rect 52 3318 107 3334
rect 141 3368 177 3418
rect 332 3585 374 3627
rect 864 3619 1146 3658
rect 1286 3637 1302 3671
rect 1336 3637 1352 3671
rect 864 3594 903 3619
rect 332 3551 340 3585
rect 332 3517 374 3551
rect 332 3483 340 3517
rect 332 3449 374 3483
rect 332 3415 340 3449
rect 332 3399 374 3415
rect 408 3585 474 3593
rect 408 3551 424 3585
rect 458 3551 474 3585
rect 408 3517 474 3551
rect 408 3483 424 3517
rect 458 3483 474 3517
rect 408 3449 474 3483
rect 408 3415 424 3449
rect 458 3415 474 3449
rect 408 3397 474 3415
rect 141 3366 182 3368
rect 141 3332 146 3366
rect 180 3332 182 3366
rect 141 3330 182 3332
rect 328 3360 394 3363
rect -834 3245 -588 3262
rect -868 3228 -588 3245
rect -868 3226 -834 3228
rect -1480 3197 -1138 3218
rect -1480 3163 -1464 3197
rect -1430 3186 -1138 3197
rect -1430 3183 -962 3186
rect -1430 3182 -1012 3183
rect -1430 3163 -1408 3182
rect -1480 3158 -1408 3163
rect -1480 3151 -1414 3158
rect -1174 3150 -1012 3182
rect -1028 3149 -1012 3150
rect -978 3149 -962 3183
rect -636 3140 -588 3228
rect -1624 3083 -1595 3117
rect -1561 3083 -1503 3117
rect -1469 3083 -1411 3117
rect -1377 3083 -1348 3117
rect -1266 3112 -1220 3122
rect -1266 3078 -1260 3112
rect -1226 3092 -1220 3112
rect -636 3106 -628 3140
rect -594 3106 -588 3140
rect -364 3239 -352 3273
rect -364 3205 -318 3239
rect -364 3171 -352 3205
rect -364 3125 -318 3171
rect -284 3273 -218 3285
rect -284 3222 -268 3273
rect -234 3222 -218 3273
rect 52 3267 86 3318
rect -284 3205 -218 3222
rect -284 3171 -268 3205
rect -234 3171 -218 3205
rect -284 3159 -218 3171
rect -47 3233 86 3267
rect 141 3258 177 3330
rect 328 3326 342 3360
rect 376 3349 394 3360
rect 328 3315 344 3326
rect 378 3315 394 3349
rect -47 3212 -13 3233
rect 125 3229 177 3258
rect -47 3157 -13 3178
rect 23 3165 39 3199
rect 73 3165 89 3199
rect -1226 3078 -1216 3092
rect -3236 2972 -3104 3008
rect -2932 3018 -2898 3034
rect -2836 3018 -2802 3034
rect -2898 2982 -2897 2983
rect -3236 2924 -3200 2972
rect -2932 2948 -2897 2982
rect -2898 2946 -2897 2948
rect -2836 2948 -2802 2982
rect -3052 2924 -2932 2946
rect -3236 2912 -2932 2924
rect -2898 2912 -2896 2946
rect -3236 2910 -2896 2912
rect -3236 2888 -3016 2910
rect -2932 2896 -2898 2910
rect -2836 2896 -2802 2912
rect -2740 3018 -2706 3034
rect -1266 3008 -1216 3078
rect -916 3068 -900 3102
rect -866 3068 -850 3102
rect -636 3094 -588 3106
rect -428 3091 -399 3125
rect -365 3091 -307 3125
rect -273 3091 -215 3125
rect -181 3091 -152 3125
rect 23 3123 89 3165
rect 159 3195 177 3229
rect 125 3157 177 3195
rect 328 3265 374 3281
rect 428 3277 474 3397
rect 612 3575 646 3594
rect 698 3585 903 3594
rect 937 3617 1146 3619
rect 937 3585 1022 3617
rect 698 3583 1022 3585
rect 1056 3594 1146 3617
rect 1386 3594 1420 3952
rect 2330 3926 2364 4137
rect 2561 3834 2595 4137
rect 2646 3918 2680 4532
rect 2846 4530 2912 4532
rect 3163 4537 3179 4571
rect 3213 4537 3229 4571
rect 3163 4503 3229 4537
rect 2718 4471 2752 4490
rect 2718 4403 2752 4405
rect 2718 4367 2752 4369
rect 2718 4282 2752 4301
rect 2814 4471 2848 4490
rect 2814 4403 2848 4405
rect 2814 4367 2848 4369
rect 2814 4282 2848 4301
rect 2910 4471 2944 4490
rect 3163 4469 3179 4503
rect 3213 4487 3229 4503
rect 3335 4639 3401 4681
rect 3369 4605 3401 4639
rect 3335 4571 3401 4605
rect 3369 4537 3401 4571
rect 3335 4503 3401 4537
rect 3213 4469 3299 4487
rect 3163 4453 3299 4469
rect 3369 4469 3401 4503
rect 3335 4453 3401 4469
rect 4237 4639 4303 4644
rect 4237 4605 4253 4639
rect 4287 4605 4303 4639
rect 4237 4571 4303 4605
rect 4237 4537 4253 4571
rect 4287 4537 4303 4571
rect 4237 4503 4303 4537
rect 4237 4469 4253 4503
rect 4287 4487 4303 4503
rect 4409 4639 4475 4681
rect 4443 4605 4475 4639
rect 4642 4675 4924 4681
rect 4642 4641 4681 4675
rect 4715 4673 4924 4675
rect 4715 4641 4800 4673
rect 4642 4639 4800 4641
rect 4834 4639 4924 4673
rect 4642 4606 4924 4639
rect 5051 4639 5117 4644
rect 4409 4571 4475 4605
rect 4443 4537 4475 4571
rect 5051 4605 5067 4639
rect 5101 4605 5117 4639
rect 5051 4571 5117 4605
rect 4409 4503 4475 4537
rect 4287 4469 4373 4487
rect 4237 4453 4373 4469
rect 4443 4469 4475 4503
rect 4409 4453 4475 4469
rect 4534 4567 4800 4568
rect 4534 4533 4750 4567
rect 4784 4533 4800 4567
rect 4534 4532 4800 4533
rect 2910 4403 2944 4405
rect 3161 4410 3231 4419
rect 3161 4376 3177 4410
rect 3211 4403 3231 4410
rect 3161 4369 3181 4376
rect 3215 4369 3231 4403
rect 2910 4367 2944 4369
rect 3265 4333 3299 4453
rect 3333 4410 3403 4419
rect 3333 4403 3351 4410
rect 3333 4369 3349 4403
rect 3385 4376 3403 4410
rect 3383 4369 3403 4376
rect 4235 4412 4305 4419
rect 4235 4378 4253 4412
rect 4287 4403 4305 4412
rect 4235 4369 4255 4378
rect 4289 4369 4305 4403
rect 4339 4333 4373 4453
rect 4407 4408 4477 4419
rect 4407 4403 4426 4408
rect 4407 4369 4423 4403
rect 4460 4374 4477 4408
rect 4457 4369 4477 4374
rect 2910 4282 2944 4301
rect 3165 4317 3213 4333
rect 3165 4283 3179 4317
rect 3165 4249 3213 4283
rect 2750 4205 2766 4239
rect 2800 4205 2816 4239
rect 3165 4215 3179 4249
rect 3165 4171 3213 4215
rect 3247 4317 3313 4333
rect 3247 4283 3263 4317
rect 3297 4287 3313 4317
rect 3247 4253 3265 4283
rect 3299 4253 3313 4287
rect 3247 4249 3313 4253
rect 3247 4215 3263 4249
rect 3297 4215 3313 4249
rect 3247 4205 3313 4215
rect 3347 4317 3401 4333
rect 3381 4283 3401 4317
rect 3347 4249 3401 4283
rect 3381 4215 3401 4249
rect 3347 4171 3401 4215
rect 4239 4317 4287 4333
rect 4239 4283 4253 4317
rect 4239 4249 4287 4283
rect 4239 4215 4253 4249
rect 4239 4171 4287 4215
rect 4321 4317 4387 4333
rect 4321 4292 4337 4317
rect 4321 4258 4335 4292
rect 4371 4283 4387 4317
rect 4369 4258 4387 4283
rect 4321 4249 4387 4258
rect 4321 4215 4337 4249
rect 4371 4215 4387 4249
rect 4321 4205 4387 4215
rect 4421 4317 4475 4333
rect 4455 4283 4475 4317
rect 4421 4249 4475 4283
rect 4455 4215 4475 4249
rect 4421 4171 4475 4215
rect 2862 4124 2878 4158
rect 2912 4124 2928 4158
rect 3144 4137 3173 4171
rect 3207 4137 3265 4171
rect 3299 4137 3357 4171
rect 3391 4137 3420 4171
rect 4218 4137 4247 4171
rect 4281 4137 4339 4171
rect 4373 4137 4431 4171
rect 4465 4137 4494 4171
rect 2734 4074 2768 4090
rect 2734 4004 2768 4038
rect 2734 3952 2768 3968
rect 2830 4074 2864 4090
rect 2830 4004 2864 4038
rect 2830 3952 2864 3968
rect 2926 4074 2960 4090
rect 2926 4004 2960 4038
rect 2960 3968 3308 3992
rect 2926 3952 3308 3968
rect 2646 3884 2782 3918
rect 2816 3884 2832 3918
rect 2561 3814 2956 3834
rect 2561 3809 2823 3814
rect 2561 3800 2702 3809
rect 2686 3775 2702 3800
rect 2736 3780 2823 3809
rect 2857 3790 2956 3814
rect 3128 3792 3174 3794
rect 3128 3790 3132 3792
rect 2857 3780 3132 3790
rect 2736 3775 3132 3780
rect 2686 3758 3132 3775
rect 3166 3758 3174 3792
rect 2686 3756 3174 3758
rect 3128 3750 3174 3756
rect 1460 3635 1489 3669
rect 1523 3635 1581 3669
rect 1615 3635 1673 3669
rect 1707 3635 1736 3669
rect 1056 3583 1292 3594
rect 698 3575 1292 3583
rect 698 3550 700 3575
rect 612 3507 646 3509
rect 612 3471 646 3473
rect 612 3386 646 3405
rect 734 3550 1258 3575
rect 1344 3575 1420 3594
rect 1344 3554 1346 3575
rect 700 3507 734 3509
rect 956 3477 972 3511
rect 1006 3477 1022 3511
rect 1258 3507 1292 3509
rect 700 3471 734 3473
rect 1258 3471 1292 3473
rect 700 3386 734 3405
rect 828 3415 862 3434
rect 828 3347 862 3349
rect 640 3309 656 3343
rect 690 3309 706 3343
rect 828 3311 862 3313
rect 328 3231 340 3265
rect 328 3197 374 3231
rect 328 3163 340 3197
rect -82 3089 -53 3123
rect -19 3089 39 3123
rect 73 3089 131 3123
rect 165 3089 194 3123
rect 328 3117 374 3163
rect 408 3265 474 3277
rect 408 3231 424 3265
rect 458 3231 474 3265
rect 408 3218 474 3231
rect 828 3226 862 3245
rect 924 3415 958 3434
rect 924 3347 958 3349
rect 924 3311 958 3313
rect 924 3226 958 3245
rect 1020 3415 1054 3434
rect 1258 3386 1292 3405
rect 1380 3554 1420 3575
rect 1528 3593 1570 3635
rect 1806 3633 1835 3667
rect 1869 3633 1927 3667
rect 1961 3633 2019 3667
rect 2053 3633 2082 3667
rect 2227 3661 2261 3668
rect 1528 3559 1536 3593
rect 1346 3507 1380 3509
rect 1346 3471 1380 3473
rect 1528 3525 1570 3559
rect 1528 3491 1536 3525
rect 1528 3457 1570 3491
rect 1528 3423 1536 3457
rect 1528 3407 1570 3423
rect 1604 3593 1670 3601
rect 1604 3559 1620 3593
rect 1654 3559 1670 3593
rect 1604 3525 1670 3559
rect 1604 3491 1620 3525
rect 1654 3491 1670 3525
rect 1604 3457 1670 3491
rect 1604 3423 1620 3457
rect 1654 3423 1670 3457
rect 1604 3405 1670 3423
rect 1839 3583 1875 3599
rect 1839 3549 1841 3583
rect 1839 3515 1875 3549
rect 1839 3481 1841 3515
rect 1911 3583 1977 3633
rect 2152 3627 2181 3661
rect 2215 3627 2273 3661
rect 2307 3627 2365 3661
rect 2399 3627 2428 3661
rect 2528 3637 2544 3671
rect 2578 3637 2594 3671
rect 2752 3658 2866 3660
rect 1911 3549 1927 3583
rect 1961 3549 1977 3583
rect 1911 3515 1977 3549
rect 1911 3481 1927 3515
rect 1961 3481 1977 3515
rect 2011 3583 2065 3599
rect 2011 3549 2013 3583
rect 2047 3549 2065 3583
rect 2011 3502 2065 3549
rect 1839 3447 1875 3481
rect 2011 3468 2013 3502
rect 2047 3468 2065 3502
rect 1839 3413 1974 3447
rect 2011 3418 2065 3468
rect 1346 3386 1380 3405
rect 1020 3347 1054 3349
rect 1432 3371 1576 3372
rect 1432 3357 1590 3371
rect 1020 3311 1054 3313
rect 1286 3344 1352 3346
rect 1432 3344 1540 3357
rect 1286 3343 1540 3344
rect 1286 3309 1302 3343
rect 1336 3330 1540 3343
rect 1336 3310 1472 3330
rect 1524 3323 1540 3330
rect 1574 3323 1590 3357
rect 1336 3309 1352 3310
rect 1524 3273 1570 3289
rect 1624 3285 1670 3405
rect 1940 3384 1974 3413
rect 1827 3355 1895 3377
rect 1827 3354 1843 3355
rect 1827 3320 1841 3354
rect 1877 3321 1895 3355
rect 1875 3320 1895 3321
rect 1827 3303 1895 3320
rect 1940 3368 1995 3384
rect 1940 3334 1961 3368
rect 1940 3318 1995 3334
rect 2029 3368 2065 3418
rect 2220 3585 2262 3627
rect 2752 3619 3034 3658
rect 3174 3637 3190 3671
rect 3224 3637 3240 3671
rect 2752 3594 2791 3619
rect 2220 3551 2228 3585
rect 2220 3517 2262 3551
rect 2220 3483 2228 3517
rect 2220 3449 2262 3483
rect 2220 3415 2228 3449
rect 2220 3399 2262 3415
rect 2296 3585 2362 3593
rect 2296 3551 2312 3585
rect 2346 3551 2362 3585
rect 2296 3517 2362 3551
rect 2296 3483 2312 3517
rect 2346 3483 2362 3517
rect 2296 3449 2362 3483
rect 2296 3415 2312 3449
rect 2346 3415 2362 3449
rect 2296 3397 2362 3415
rect 2029 3366 2070 3368
rect 2029 3332 2034 3366
rect 2068 3332 2070 3366
rect 2029 3330 2070 3332
rect 2216 3360 2282 3363
rect 1054 3245 1300 3262
rect 1020 3228 1300 3245
rect 1020 3226 1054 3228
rect 408 3197 750 3218
rect 408 3163 424 3197
rect 458 3186 750 3197
rect 458 3183 926 3186
rect 458 3182 876 3183
rect 458 3163 480 3182
rect 408 3158 480 3163
rect 408 3151 474 3158
rect 714 3150 876 3182
rect 860 3149 876 3150
rect 910 3149 926 3183
rect 1252 3140 1300 3228
rect 264 3083 293 3117
rect 327 3083 385 3117
rect 419 3083 477 3117
rect 511 3083 540 3117
rect 622 3112 668 3122
rect 622 3078 628 3112
rect 662 3092 668 3112
rect 1252 3106 1260 3140
rect 1294 3106 1300 3140
rect 1524 3239 1536 3273
rect 1524 3205 1570 3239
rect 1524 3171 1536 3205
rect 1524 3125 1570 3171
rect 1604 3273 1670 3285
rect 1604 3222 1620 3273
rect 1654 3222 1670 3273
rect 1940 3267 1974 3318
rect 1604 3205 1670 3222
rect 1604 3171 1620 3205
rect 1654 3171 1670 3205
rect 1604 3159 1670 3171
rect 1841 3233 1974 3267
rect 2029 3258 2065 3330
rect 2216 3326 2230 3360
rect 2264 3349 2282 3360
rect 2216 3315 2232 3326
rect 2266 3315 2282 3349
rect 1841 3212 1875 3233
rect 2013 3229 2065 3258
rect 1841 3157 1875 3178
rect 1911 3165 1927 3199
rect 1961 3165 1977 3199
rect 662 3078 672 3092
rect -2740 2948 -2706 2982
rect -2740 2896 -2706 2912
rect -1348 2972 -1216 3008
rect -1044 3018 -1010 3034
rect -948 3018 -914 3034
rect -1010 2982 -1009 2983
rect -1348 2924 -1312 2972
rect -1044 2948 -1009 2982
rect -1010 2946 -1009 2948
rect -948 2948 -914 2982
rect -1164 2924 -1044 2946
rect -1348 2912 -1044 2924
rect -1010 2912 -1008 2946
rect -1348 2910 -1008 2912
rect -1348 2888 -1128 2910
rect -1044 2896 -1010 2910
rect -948 2896 -914 2912
rect -852 3018 -818 3034
rect 622 3008 672 3078
rect 972 3068 988 3102
rect 1022 3068 1038 3102
rect 1252 3094 1300 3106
rect 1460 3091 1489 3125
rect 1523 3091 1581 3125
rect 1615 3091 1673 3125
rect 1707 3091 1736 3125
rect 1911 3123 1977 3165
rect 2047 3195 2065 3229
rect 2013 3157 2065 3195
rect 2216 3265 2262 3281
rect 2316 3277 2362 3397
rect 2500 3575 2534 3594
rect 2586 3585 2791 3594
rect 2825 3617 3034 3619
rect 2825 3585 2910 3617
rect 2586 3583 2910 3585
rect 2944 3594 3034 3617
rect 3274 3594 3308 3952
rect 4218 3926 4252 4137
rect 4449 3834 4483 4137
rect 4534 3918 4568 4532
rect 4734 4530 4800 4532
rect 5051 4537 5067 4571
rect 5101 4537 5117 4571
rect 5051 4503 5117 4537
rect 4606 4471 4640 4490
rect 4606 4403 4640 4405
rect 4606 4367 4640 4369
rect 4606 4282 4640 4301
rect 4702 4471 4736 4490
rect 4702 4403 4736 4405
rect 4702 4367 4736 4369
rect 4702 4282 4736 4301
rect 4798 4471 4832 4490
rect 5051 4469 5067 4503
rect 5101 4487 5117 4503
rect 5223 4639 5289 4681
rect 5257 4605 5289 4639
rect 5223 4571 5289 4605
rect 5257 4537 5289 4571
rect 5223 4503 5289 4537
rect 5101 4469 5187 4487
rect 5051 4453 5187 4469
rect 5257 4469 5289 4503
rect 5223 4453 5289 4469
rect 6125 4639 6191 4644
rect 6125 4605 6141 4639
rect 6175 4605 6191 4639
rect 6125 4571 6191 4605
rect 6125 4537 6141 4571
rect 6175 4537 6191 4571
rect 6125 4503 6191 4537
rect 6125 4469 6141 4503
rect 6175 4487 6191 4503
rect 6297 4639 6363 4681
rect 6331 4605 6363 4639
rect 6530 4675 6812 4681
rect 6530 4641 6569 4675
rect 6603 4673 6812 4675
rect 6603 4641 6688 4673
rect 6530 4639 6688 4641
rect 6722 4639 6812 4673
rect 6530 4606 6812 4639
rect 6939 4639 7005 4644
rect 6297 4571 6363 4605
rect 6331 4537 6363 4571
rect 6939 4605 6955 4639
rect 6989 4605 7005 4639
rect 6939 4571 7005 4605
rect 6297 4503 6363 4537
rect 6175 4469 6261 4487
rect 6125 4453 6261 4469
rect 6331 4469 6363 4503
rect 6297 4453 6363 4469
rect 6422 4567 6688 4568
rect 6422 4533 6638 4567
rect 6672 4533 6688 4567
rect 6422 4532 6688 4533
rect 4798 4403 4832 4405
rect 5049 4410 5119 4419
rect 5049 4376 5065 4410
rect 5099 4403 5119 4410
rect 5049 4369 5069 4376
rect 5103 4369 5119 4403
rect 4798 4367 4832 4369
rect 5153 4333 5187 4453
rect 5221 4410 5291 4419
rect 5221 4403 5239 4410
rect 5221 4369 5237 4403
rect 5273 4376 5291 4410
rect 5271 4369 5291 4376
rect 6123 4412 6193 4419
rect 6123 4378 6141 4412
rect 6175 4403 6193 4412
rect 6123 4369 6143 4378
rect 6177 4369 6193 4403
rect 6227 4333 6261 4453
rect 6295 4408 6365 4419
rect 6295 4403 6314 4408
rect 6295 4369 6311 4403
rect 6348 4374 6365 4408
rect 6345 4369 6365 4374
rect 4798 4282 4832 4301
rect 5053 4317 5101 4333
rect 5053 4283 5067 4317
rect 5053 4249 5101 4283
rect 4638 4205 4654 4239
rect 4688 4205 4704 4239
rect 5053 4215 5067 4249
rect 5053 4171 5101 4215
rect 5135 4317 5201 4333
rect 5135 4283 5151 4317
rect 5185 4287 5201 4317
rect 5135 4253 5153 4283
rect 5187 4253 5201 4287
rect 5135 4249 5201 4253
rect 5135 4215 5151 4249
rect 5185 4215 5201 4249
rect 5135 4205 5201 4215
rect 5235 4317 5289 4333
rect 5269 4283 5289 4317
rect 5235 4249 5289 4283
rect 5269 4215 5289 4249
rect 5235 4171 5289 4215
rect 6127 4317 6175 4333
rect 6127 4283 6141 4317
rect 6127 4249 6175 4283
rect 6127 4215 6141 4249
rect 6127 4171 6175 4215
rect 6209 4317 6275 4333
rect 6209 4292 6225 4317
rect 6209 4258 6223 4292
rect 6259 4283 6275 4317
rect 6257 4258 6275 4283
rect 6209 4249 6275 4258
rect 6209 4215 6225 4249
rect 6259 4215 6275 4249
rect 6209 4205 6275 4215
rect 6309 4317 6363 4333
rect 6343 4283 6363 4317
rect 6309 4249 6363 4283
rect 6343 4215 6363 4249
rect 6309 4171 6363 4215
rect 4750 4124 4766 4158
rect 4800 4124 4816 4158
rect 5032 4137 5061 4171
rect 5095 4137 5153 4171
rect 5187 4137 5245 4171
rect 5279 4137 5308 4171
rect 6106 4137 6135 4171
rect 6169 4137 6227 4171
rect 6261 4137 6319 4171
rect 6353 4137 6382 4171
rect 4622 4074 4656 4090
rect 4622 4004 4656 4038
rect 4622 3952 4656 3968
rect 4718 4074 4752 4090
rect 4718 4004 4752 4038
rect 4718 3952 4752 3968
rect 4814 4074 4848 4090
rect 4814 4004 4848 4038
rect 4848 3968 5196 3992
rect 4814 3952 5196 3968
rect 4534 3884 4670 3918
rect 4704 3884 4720 3918
rect 4449 3814 4844 3834
rect 4449 3809 4711 3814
rect 4449 3800 4590 3809
rect 4574 3775 4590 3800
rect 4624 3780 4711 3809
rect 4745 3790 4844 3814
rect 5016 3792 5062 3794
rect 5016 3790 5020 3792
rect 4745 3780 5020 3790
rect 4624 3775 5020 3780
rect 4574 3758 5020 3775
rect 5054 3758 5062 3792
rect 4574 3756 5062 3758
rect 5016 3750 5062 3756
rect 3348 3635 3377 3669
rect 3411 3635 3469 3669
rect 3503 3635 3561 3669
rect 3595 3635 3624 3669
rect 2944 3583 3180 3594
rect 2586 3575 3180 3583
rect 2586 3550 2588 3575
rect 2500 3507 2534 3509
rect 2500 3471 2534 3473
rect 2500 3386 2534 3405
rect 2622 3550 3146 3575
rect 3232 3575 3308 3594
rect 3232 3554 3234 3575
rect 2588 3507 2622 3509
rect 2844 3477 2860 3511
rect 2894 3477 2910 3511
rect 3146 3507 3180 3509
rect 2588 3471 2622 3473
rect 3146 3471 3180 3473
rect 2588 3386 2622 3405
rect 2716 3415 2750 3434
rect 2716 3347 2750 3349
rect 2528 3309 2544 3343
rect 2578 3309 2594 3343
rect 2716 3311 2750 3313
rect 2216 3231 2228 3265
rect 2216 3197 2262 3231
rect 2216 3163 2228 3197
rect 1806 3089 1835 3123
rect 1869 3089 1927 3123
rect 1961 3089 2019 3123
rect 2053 3089 2082 3123
rect 2216 3117 2262 3163
rect 2296 3265 2362 3277
rect 2296 3231 2312 3265
rect 2346 3231 2362 3265
rect 2296 3218 2362 3231
rect 2716 3226 2750 3245
rect 2812 3415 2846 3434
rect 2812 3347 2846 3349
rect 2812 3311 2846 3313
rect 2812 3226 2846 3245
rect 2908 3415 2942 3434
rect 3146 3386 3180 3405
rect 3268 3554 3308 3575
rect 3416 3593 3458 3635
rect 3694 3633 3723 3667
rect 3757 3633 3815 3667
rect 3849 3633 3907 3667
rect 3941 3633 3970 3667
rect 4115 3661 4149 3668
rect 3416 3559 3424 3593
rect 3234 3507 3268 3509
rect 3234 3471 3268 3473
rect 3416 3525 3458 3559
rect 3416 3491 3424 3525
rect 3416 3457 3458 3491
rect 3416 3423 3424 3457
rect 3416 3407 3458 3423
rect 3492 3593 3558 3601
rect 3492 3559 3508 3593
rect 3542 3559 3558 3593
rect 3492 3525 3558 3559
rect 3492 3491 3508 3525
rect 3542 3491 3558 3525
rect 3492 3457 3558 3491
rect 3492 3423 3508 3457
rect 3542 3423 3558 3457
rect 3492 3405 3558 3423
rect 3727 3583 3763 3599
rect 3727 3549 3729 3583
rect 3727 3515 3763 3549
rect 3727 3481 3729 3515
rect 3799 3583 3865 3633
rect 4040 3627 4069 3661
rect 4103 3627 4161 3661
rect 4195 3627 4253 3661
rect 4287 3627 4316 3661
rect 4416 3637 4432 3671
rect 4466 3637 4482 3671
rect 4640 3658 4754 3660
rect 3799 3549 3815 3583
rect 3849 3549 3865 3583
rect 3799 3515 3865 3549
rect 3799 3481 3815 3515
rect 3849 3481 3865 3515
rect 3899 3583 3953 3599
rect 3899 3549 3901 3583
rect 3935 3549 3953 3583
rect 3899 3502 3953 3549
rect 3727 3447 3763 3481
rect 3899 3468 3901 3502
rect 3935 3468 3953 3502
rect 3727 3413 3862 3447
rect 3899 3418 3953 3468
rect 3234 3386 3268 3405
rect 2908 3347 2942 3349
rect 3320 3371 3464 3372
rect 3320 3357 3478 3371
rect 2908 3311 2942 3313
rect 3174 3344 3240 3346
rect 3320 3344 3428 3357
rect 3174 3343 3428 3344
rect 3174 3309 3190 3343
rect 3224 3330 3428 3343
rect 3224 3310 3360 3330
rect 3412 3323 3428 3330
rect 3462 3323 3478 3357
rect 3224 3309 3240 3310
rect 3412 3273 3458 3289
rect 3512 3285 3558 3405
rect 3828 3384 3862 3413
rect 3715 3355 3783 3377
rect 3715 3354 3731 3355
rect 3715 3320 3729 3354
rect 3765 3321 3783 3355
rect 3763 3320 3783 3321
rect 3715 3303 3783 3320
rect 3828 3368 3883 3384
rect 3828 3334 3849 3368
rect 3828 3318 3883 3334
rect 3917 3368 3953 3418
rect 4108 3585 4150 3627
rect 4640 3619 4922 3658
rect 5062 3637 5078 3671
rect 5112 3637 5128 3671
rect 4640 3594 4679 3619
rect 4108 3551 4116 3585
rect 4108 3517 4150 3551
rect 4108 3483 4116 3517
rect 4108 3449 4150 3483
rect 4108 3415 4116 3449
rect 4108 3399 4150 3415
rect 4184 3585 4250 3593
rect 4184 3551 4200 3585
rect 4234 3551 4250 3585
rect 4184 3517 4250 3551
rect 4184 3483 4200 3517
rect 4234 3483 4250 3517
rect 4184 3449 4250 3483
rect 4184 3415 4200 3449
rect 4234 3415 4250 3449
rect 4184 3397 4250 3415
rect 3917 3366 3958 3368
rect 3917 3332 3922 3366
rect 3956 3332 3958 3366
rect 3917 3330 3958 3332
rect 4104 3360 4170 3363
rect 2942 3245 3188 3262
rect 2908 3228 3188 3245
rect 2908 3226 2942 3228
rect 2296 3197 2638 3218
rect 2296 3163 2312 3197
rect 2346 3186 2638 3197
rect 2346 3183 2814 3186
rect 2346 3182 2764 3183
rect 2346 3163 2368 3182
rect 2296 3158 2368 3163
rect 2296 3151 2362 3158
rect 2602 3150 2764 3182
rect 2748 3149 2764 3150
rect 2798 3149 2814 3183
rect 3140 3140 3188 3228
rect 2152 3083 2181 3117
rect 2215 3083 2273 3117
rect 2307 3083 2365 3117
rect 2399 3083 2428 3117
rect 2510 3112 2556 3122
rect 2510 3078 2516 3112
rect 2550 3092 2556 3112
rect 3140 3106 3148 3140
rect 3182 3106 3188 3140
rect 3412 3239 3424 3273
rect 3412 3205 3458 3239
rect 3412 3171 3424 3205
rect 3412 3125 3458 3171
rect 3492 3273 3558 3285
rect 3492 3222 3508 3273
rect 3542 3222 3558 3273
rect 3828 3267 3862 3318
rect 3492 3205 3558 3222
rect 3492 3171 3508 3205
rect 3542 3171 3558 3205
rect 3492 3159 3558 3171
rect 3729 3233 3862 3267
rect 3917 3258 3953 3330
rect 4104 3326 4118 3360
rect 4152 3349 4170 3360
rect 4104 3315 4120 3326
rect 4154 3315 4170 3349
rect 3729 3212 3763 3233
rect 3901 3229 3953 3258
rect 3729 3157 3763 3178
rect 3799 3165 3815 3199
rect 3849 3165 3865 3199
rect 2550 3078 2560 3092
rect -852 2948 -818 2982
rect -852 2896 -818 2912
rect 540 2972 672 3008
rect 844 3018 878 3034
rect 940 3018 974 3034
rect 878 2982 879 2983
rect 540 2924 576 2972
rect 844 2948 879 2982
rect 878 2946 879 2948
rect 940 2948 974 2982
rect 724 2924 844 2946
rect 540 2912 844 2924
rect 878 2912 880 2946
rect 540 2910 880 2912
rect 540 2888 760 2910
rect 844 2896 878 2910
rect 940 2896 974 2912
rect 1036 3018 1070 3034
rect 2510 3008 2560 3078
rect 2860 3068 2876 3102
rect 2910 3068 2926 3102
rect 3140 3094 3188 3106
rect 3348 3091 3377 3125
rect 3411 3091 3469 3125
rect 3503 3091 3561 3125
rect 3595 3091 3624 3125
rect 3799 3123 3865 3165
rect 3935 3195 3953 3229
rect 3901 3157 3953 3195
rect 4104 3265 4150 3281
rect 4204 3277 4250 3397
rect 4388 3575 4422 3594
rect 4474 3585 4679 3594
rect 4713 3617 4922 3619
rect 4713 3585 4798 3617
rect 4474 3583 4798 3585
rect 4832 3594 4922 3617
rect 5162 3594 5196 3952
rect 6106 3926 6140 4137
rect 6337 3834 6371 4137
rect 6422 3918 6456 4532
rect 6622 4530 6688 4532
rect 6939 4537 6955 4571
rect 6989 4537 7005 4571
rect 6939 4503 7005 4537
rect 6494 4471 6528 4490
rect 6494 4403 6528 4405
rect 6494 4367 6528 4369
rect 6494 4282 6528 4301
rect 6590 4471 6624 4490
rect 6590 4403 6624 4405
rect 6590 4367 6624 4369
rect 6590 4282 6624 4301
rect 6686 4471 6720 4490
rect 6939 4469 6955 4503
rect 6989 4487 7005 4503
rect 7111 4639 7177 4681
rect 7145 4605 7177 4639
rect 7111 4571 7177 4605
rect 7145 4537 7177 4571
rect 7111 4503 7177 4537
rect 6989 4469 7075 4487
rect 6939 4453 7075 4469
rect 7145 4469 7177 4503
rect 7111 4453 7177 4469
rect 8013 4639 8079 4644
rect 8013 4605 8029 4639
rect 8063 4605 8079 4639
rect 8013 4571 8079 4605
rect 8013 4537 8029 4571
rect 8063 4537 8079 4571
rect 8013 4503 8079 4537
rect 8013 4469 8029 4503
rect 8063 4487 8079 4503
rect 8185 4639 8251 4681
rect 8219 4605 8251 4639
rect 8418 4675 8700 4681
rect 8418 4641 8457 4675
rect 8491 4673 8700 4675
rect 8491 4641 8576 4673
rect 8418 4639 8576 4641
rect 8610 4639 8700 4673
rect 8418 4606 8700 4639
rect 8827 4639 8893 4644
rect 8185 4571 8251 4605
rect 8219 4537 8251 4571
rect 8827 4605 8843 4639
rect 8877 4605 8893 4639
rect 8827 4571 8893 4605
rect 8185 4503 8251 4537
rect 8063 4469 8149 4487
rect 8013 4453 8149 4469
rect 8219 4469 8251 4503
rect 8185 4453 8251 4469
rect 8310 4567 8576 4568
rect 8310 4533 8526 4567
rect 8560 4533 8576 4567
rect 8310 4532 8576 4533
rect 6686 4403 6720 4405
rect 6937 4410 7007 4419
rect 6937 4376 6953 4410
rect 6987 4403 7007 4410
rect 6937 4369 6957 4376
rect 6991 4369 7007 4403
rect 6686 4367 6720 4369
rect 7041 4333 7075 4453
rect 7109 4410 7179 4419
rect 7109 4403 7127 4410
rect 7109 4369 7125 4403
rect 7161 4376 7179 4410
rect 7159 4369 7179 4376
rect 8011 4412 8081 4419
rect 8011 4378 8029 4412
rect 8063 4403 8081 4412
rect 8011 4369 8031 4378
rect 8065 4369 8081 4403
rect 8115 4333 8149 4453
rect 8183 4408 8253 4419
rect 8183 4403 8202 4408
rect 8183 4369 8199 4403
rect 8236 4374 8253 4408
rect 8233 4369 8253 4374
rect 6686 4282 6720 4301
rect 6941 4317 6989 4333
rect 6941 4283 6955 4317
rect 6941 4249 6989 4283
rect 6526 4205 6542 4239
rect 6576 4205 6592 4239
rect 6941 4215 6955 4249
rect 6941 4171 6989 4215
rect 7023 4317 7089 4333
rect 7023 4283 7039 4317
rect 7073 4287 7089 4317
rect 7023 4253 7041 4283
rect 7075 4253 7089 4287
rect 7023 4249 7089 4253
rect 7023 4215 7039 4249
rect 7073 4215 7089 4249
rect 7023 4205 7089 4215
rect 7123 4317 7177 4333
rect 7157 4283 7177 4317
rect 7123 4249 7177 4283
rect 7157 4215 7177 4249
rect 7123 4171 7177 4215
rect 8015 4317 8063 4333
rect 8015 4283 8029 4317
rect 8015 4249 8063 4283
rect 8015 4215 8029 4249
rect 8015 4171 8063 4215
rect 8097 4317 8163 4333
rect 8097 4292 8113 4317
rect 8097 4258 8111 4292
rect 8147 4283 8163 4317
rect 8145 4258 8163 4283
rect 8097 4249 8163 4258
rect 8097 4215 8113 4249
rect 8147 4215 8163 4249
rect 8097 4205 8163 4215
rect 8197 4317 8251 4333
rect 8231 4283 8251 4317
rect 8197 4249 8251 4283
rect 8231 4215 8251 4249
rect 8197 4171 8251 4215
rect 6638 4124 6654 4158
rect 6688 4124 6704 4158
rect 6920 4137 6949 4171
rect 6983 4137 7041 4171
rect 7075 4137 7133 4171
rect 7167 4137 7196 4171
rect 7994 4137 8023 4171
rect 8057 4137 8115 4171
rect 8149 4137 8207 4171
rect 8241 4137 8270 4171
rect 6510 4074 6544 4090
rect 6510 4004 6544 4038
rect 6510 3952 6544 3968
rect 6606 4074 6640 4090
rect 6606 4004 6640 4038
rect 6606 3952 6640 3968
rect 6702 4074 6736 4090
rect 6702 4004 6736 4038
rect 6736 3968 7084 3992
rect 6702 3952 7084 3968
rect 6422 3884 6558 3918
rect 6592 3884 6608 3918
rect 6337 3814 6732 3834
rect 6337 3809 6599 3814
rect 6337 3800 6478 3809
rect 6462 3775 6478 3800
rect 6512 3780 6599 3809
rect 6633 3790 6732 3814
rect 6904 3792 6950 3794
rect 6904 3790 6908 3792
rect 6633 3780 6908 3790
rect 6512 3775 6908 3780
rect 6462 3758 6908 3775
rect 6942 3758 6950 3792
rect 6462 3756 6950 3758
rect 6904 3750 6950 3756
rect 5236 3635 5265 3669
rect 5299 3635 5357 3669
rect 5391 3635 5449 3669
rect 5483 3635 5512 3669
rect 4832 3583 5068 3594
rect 4474 3575 5068 3583
rect 4474 3550 4476 3575
rect 4388 3507 4422 3509
rect 4388 3471 4422 3473
rect 4388 3386 4422 3405
rect 4510 3550 5034 3575
rect 5120 3575 5196 3594
rect 5120 3554 5122 3575
rect 4476 3507 4510 3509
rect 4732 3477 4748 3511
rect 4782 3477 4798 3511
rect 5034 3507 5068 3509
rect 4476 3471 4510 3473
rect 5034 3471 5068 3473
rect 4476 3386 4510 3405
rect 4604 3415 4638 3434
rect 4604 3347 4638 3349
rect 4416 3309 4432 3343
rect 4466 3309 4482 3343
rect 4604 3311 4638 3313
rect 4104 3231 4116 3265
rect 4104 3197 4150 3231
rect 4104 3163 4116 3197
rect 3694 3089 3723 3123
rect 3757 3089 3815 3123
rect 3849 3089 3907 3123
rect 3941 3089 3970 3123
rect 4104 3117 4150 3163
rect 4184 3265 4250 3277
rect 4184 3231 4200 3265
rect 4234 3231 4250 3265
rect 4184 3218 4250 3231
rect 4604 3226 4638 3245
rect 4700 3415 4734 3434
rect 4700 3347 4734 3349
rect 4700 3311 4734 3313
rect 4700 3226 4734 3245
rect 4796 3415 4830 3434
rect 5034 3386 5068 3405
rect 5156 3554 5196 3575
rect 5304 3593 5346 3635
rect 5582 3633 5611 3667
rect 5645 3633 5703 3667
rect 5737 3633 5795 3667
rect 5829 3633 5858 3667
rect 6003 3661 6037 3668
rect 5304 3559 5312 3593
rect 5122 3507 5156 3509
rect 5122 3471 5156 3473
rect 5304 3525 5346 3559
rect 5304 3491 5312 3525
rect 5304 3457 5346 3491
rect 5304 3423 5312 3457
rect 5304 3407 5346 3423
rect 5380 3593 5446 3601
rect 5380 3559 5396 3593
rect 5430 3559 5446 3593
rect 5380 3525 5446 3559
rect 5380 3491 5396 3525
rect 5430 3491 5446 3525
rect 5380 3457 5446 3491
rect 5380 3423 5396 3457
rect 5430 3423 5446 3457
rect 5380 3405 5446 3423
rect 5615 3583 5651 3599
rect 5615 3549 5617 3583
rect 5615 3515 5651 3549
rect 5615 3481 5617 3515
rect 5687 3583 5753 3633
rect 5928 3627 5957 3661
rect 5991 3627 6049 3661
rect 6083 3627 6141 3661
rect 6175 3627 6204 3661
rect 6304 3637 6320 3671
rect 6354 3637 6370 3671
rect 6528 3658 6642 3660
rect 5687 3549 5703 3583
rect 5737 3549 5753 3583
rect 5687 3515 5753 3549
rect 5687 3481 5703 3515
rect 5737 3481 5753 3515
rect 5787 3583 5841 3599
rect 5787 3549 5789 3583
rect 5823 3549 5841 3583
rect 5787 3502 5841 3549
rect 5615 3447 5651 3481
rect 5787 3468 5789 3502
rect 5823 3468 5841 3502
rect 5615 3413 5750 3447
rect 5787 3418 5841 3468
rect 5122 3386 5156 3405
rect 4796 3347 4830 3349
rect 5208 3371 5352 3372
rect 5208 3357 5366 3371
rect 4796 3311 4830 3313
rect 5062 3344 5128 3346
rect 5208 3344 5316 3357
rect 5062 3343 5316 3344
rect 5062 3309 5078 3343
rect 5112 3330 5316 3343
rect 5112 3310 5248 3330
rect 5300 3323 5316 3330
rect 5350 3323 5366 3357
rect 5112 3309 5128 3310
rect 5300 3273 5346 3289
rect 5400 3285 5446 3405
rect 5716 3384 5750 3413
rect 5603 3355 5671 3377
rect 5603 3354 5619 3355
rect 5603 3320 5617 3354
rect 5653 3321 5671 3355
rect 5651 3320 5671 3321
rect 5603 3303 5671 3320
rect 5716 3368 5771 3384
rect 5716 3334 5737 3368
rect 5716 3318 5771 3334
rect 5805 3368 5841 3418
rect 5996 3585 6038 3627
rect 6528 3619 6810 3658
rect 6950 3637 6966 3671
rect 7000 3637 7016 3671
rect 6528 3594 6567 3619
rect 5996 3551 6004 3585
rect 5996 3517 6038 3551
rect 5996 3483 6004 3517
rect 5996 3449 6038 3483
rect 5996 3415 6004 3449
rect 5996 3399 6038 3415
rect 6072 3585 6138 3593
rect 6072 3551 6088 3585
rect 6122 3551 6138 3585
rect 6072 3517 6138 3551
rect 6072 3483 6088 3517
rect 6122 3483 6138 3517
rect 6072 3449 6138 3483
rect 6072 3415 6088 3449
rect 6122 3415 6138 3449
rect 6072 3397 6138 3415
rect 5805 3366 5846 3368
rect 5805 3332 5810 3366
rect 5844 3332 5846 3366
rect 5805 3330 5846 3332
rect 5992 3360 6058 3363
rect 4830 3245 5076 3262
rect 4796 3228 5076 3245
rect 4796 3226 4830 3228
rect 4184 3197 4526 3218
rect 4184 3163 4200 3197
rect 4234 3186 4526 3197
rect 4234 3183 4702 3186
rect 4234 3182 4652 3183
rect 4234 3163 4256 3182
rect 4184 3158 4256 3163
rect 4184 3151 4250 3158
rect 4490 3150 4652 3182
rect 4636 3149 4652 3150
rect 4686 3149 4702 3183
rect 5028 3140 5076 3228
rect 4040 3083 4069 3117
rect 4103 3083 4161 3117
rect 4195 3083 4253 3117
rect 4287 3083 4316 3117
rect 4398 3112 4444 3122
rect 4398 3078 4404 3112
rect 4438 3092 4444 3112
rect 5028 3106 5036 3140
rect 5070 3106 5076 3140
rect 5300 3239 5312 3273
rect 5300 3205 5346 3239
rect 5300 3171 5312 3205
rect 5300 3125 5346 3171
rect 5380 3273 5446 3285
rect 5380 3222 5396 3273
rect 5430 3222 5446 3273
rect 5716 3267 5750 3318
rect 5380 3205 5446 3222
rect 5380 3171 5396 3205
rect 5430 3171 5446 3205
rect 5380 3159 5446 3171
rect 5617 3233 5750 3267
rect 5805 3258 5841 3330
rect 5992 3326 6006 3360
rect 6040 3349 6058 3360
rect 5992 3315 6008 3326
rect 6042 3315 6058 3349
rect 5617 3212 5651 3233
rect 5789 3229 5841 3258
rect 5617 3157 5651 3178
rect 5687 3165 5703 3199
rect 5737 3165 5753 3199
rect 4438 3078 4448 3092
rect 1036 2948 1070 2982
rect 1036 2896 1070 2912
rect 2428 2972 2560 3008
rect 2732 3018 2766 3034
rect 2828 3018 2862 3034
rect 2766 2982 2767 2983
rect 2428 2924 2464 2972
rect 2732 2948 2767 2982
rect 2766 2946 2767 2948
rect 2828 2948 2862 2982
rect 2612 2924 2732 2946
rect 2428 2912 2732 2924
rect 2766 2912 2768 2946
rect 2428 2910 2768 2912
rect 2428 2888 2648 2910
rect 2732 2896 2766 2910
rect 2828 2896 2862 2912
rect 2924 3018 2958 3034
rect 4398 3008 4448 3078
rect 4748 3068 4764 3102
rect 4798 3068 4814 3102
rect 5028 3094 5076 3106
rect 5236 3091 5265 3125
rect 5299 3091 5357 3125
rect 5391 3091 5449 3125
rect 5483 3091 5512 3125
rect 5687 3123 5753 3165
rect 5823 3195 5841 3229
rect 5789 3157 5841 3195
rect 5992 3265 6038 3281
rect 6092 3277 6138 3397
rect 6276 3575 6310 3594
rect 6362 3585 6567 3594
rect 6601 3617 6810 3619
rect 6601 3585 6686 3617
rect 6362 3583 6686 3585
rect 6720 3594 6810 3617
rect 7050 3594 7084 3952
rect 7994 3926 8028 4137
rect 8225 3834 8259 4137
rect 8310 3918 8344 4532
rect 8510 4530 8576 4532
rect 8827 4537 8843 4571
rect 8877 4537 8893 4571
rect 8827 4503 8893 4537
rect 8382 4471 8416 4490
rect 8382 4403 8416 4405
rect 8382 4367 8416 4369
rect 8382 4282 8416 4301
rect 8478 4471 8512 4490
rect 8478 4403 8512 4405
rect 8478 4367 8512 4369
rect 8478 4282 8512 4301
rect 8574 4471 8608 4490
rect 8827 4469 8843 4503
rect 8877 4487 8893 4503
rect 8999 4639 9065 4681
rect 9033 4605 9065 4639
rect 8999 4571 9065 4605
rect 9033 4537 9065 4571
rect 8999 4503 9065 4537
rect 8877 4469 8963 4487
rect 8827 4453 8963 4469
rect 9033 4469 9065 4503
rect 8999 4453 9065 4469
rect 9901 4639 9967 4644
rect 9901 4605 9917 4639
rect 9951 4605 9967 4639
rect 9901 4571 9967 4605
rect 9901 4537 9917 4571
rect 9951 4537 9967 4571
rect 9901 4503 9967 4537
rect 9901 4469 9917 4503
rect 9951 4487 9967 4503
rect 10073 4639 10139 4681
rect 10107 4605 10139 4639
rect 10306 4675 10588 4681
rect 10306 4641 10345 4675
rect 10379 4673 10588 4675
rect 10379 4641 10464 4673
rect 10306 4639 10464 4641
rect 10498 4639 10588 4673
rect 10306 4606 10588 4639
rect 10715 4639 10781 4644
rect 10073 4571 10139 4605
rect 10107 4537 10139 4571
rect 10715 4605 10731 4639
rect 10765 4605 10781 4639
rect 10715 4571 10781 4605
rect 10073 4503 10139 4537
rect 9951 4469 10037 4487
rect 9901 4453 10037 4469
rect 10107 4469 10139 4503
rect 10073 4453 10139 4469
rect 10198 4567 10464 4568
rect 10198 4533 10414 4567
rect 10448 4533 10464 4567
rect 10198 4532 10464 4533
rect 8574 4403 8608 4405
rect 8825 4410 8895 4419
rect 8825 4376 8841 4410
rect 8875 4403 8895 4410
rect 8825 4369 8845 4376
rect 8879 4369 8895 4403
rect 8574 4367 8608 4369
rect 8929 4333 8963 4453
rect 8997 4410 9067 4419
rect 8997 4403 9015 4410
rect 8997 4369 9013 4403
rect 9049 4376 9067 4410
rect 9047 4369 9067 4376
rect 9899 4412 9969 4419
rect 9899 4378 9917 4412
rect 9951 4403 9969 4412
rect 9899 4369 9919 4378
rect 9953 4369 9969 4403
rect 10003 4333 10037 4453
rect 10071 4408 10141 4419
rect 10071 4403 10090 4408
rect 10071 4369 10087 4403
rect 10124 4374 10141 4408
rect 10121 4369 10141 4374
rect 8574 4282 8608 4301
rect 8829 4317 8877 4333
rect 8829 4283 8843 4317
rect 8829 4249 8877 4283
rect 8414 4205 8430 4239
rect 8464 4205 8480 4239
rect 8829 4215 8843 4249
rect 8829 4171 8877 4215
rect 8911 4317 8977 4333
rect 8911 4283 8927 4317
rect 8961 4287 8977 4317
rect 8911 4253 8929 4283
rect 8963 4253 8977 4287
rect 8911 4249 8977 4253
rect 8911 4215 8927 4249
rect 8961 4215 8977 4249
rect 8911 4205 8977 4215
rect 9011 4317 9065 4333
rect 9045 4283 9065 4317
rect 9011 4249 9065 4283
rect 9045 4215 9065 4249
rect 9011 4171 9065 4215
rect 9903 4317 9951 4333
rect 9903 4283 9917 4317
rect 9903 4249 9951 4283
rect 9903 4215 9917 4249
rect 9903 4171 9951 4215
rect 9985 4317 10051 4333
rect 9985 4292 10001 4317
rect 9985 4258 9999 4292
rect 10035 4283 10051 4317
rect 10033 4258 10051 4283
rect 9985 4249 10051 4258
rect 9985 4215 10001 4249
rect 10035 4215 10051 4249
rect 9985 4205 10051 4215
rect 10085 4317 10139 4333
rect 10119 4283 10139 4317
rect 10085 4249 10139 4283
rect 10119 4215 10139 4249
rect 10085 4171 10139 4215
rect 8526 4124 8542 4158
rect 8576 4124 8592 4158
rect 8808 4137 8837 4171
rect 8871 4137 8929 4171
rect 8963 4137 9021 4171
rect 9055 4137 9084 4171
rect 9882 4137 9911 4171
rect 9945 4137 10003 4171
rect 10037 4137 10095 4171
rect 10129 4137 10158 4171
rect 8398 4074 8432 4090
rect 8398 4004 8432 4038
rect 8398 3952 8432 3968
rect 8494 4074 8528 4090
rect 8494 4004 8528 4038
rect 8494 3952 8528 3968
rect 8590 4074 8624 4090
rect 8590 4004 8624 4038
rect 8624 3968 8972 3992
rect 8590 3952 8972 3968
rect 8310 3884 8446 3918
rect 8480 3884 8496 3918
rect 8225 3814 8620 3834
rect 8225 3809 8487 3814
rect 8225 3800 8366 3809
rect 8350 3775 8366 3800
rect 8400 3780 8487 3809
rect 8521 3790 8620 3814
rect 8792 3792 8838 3794
rect 8792 3790 8796 3792
rect 8521 3780 8796 3790
rect 8400 3775 8796 3780
rect 8350 3758 8796 3775
rect 8830 3758 8838 3792
rect 8350 3756 8838 3758
rect 8792 3750 8838 3756
rect 7124 3635 7153 3669
rect 7187 3635 7245 3669
rect 7279 3635 7337 3669
rect 7371 3635 7400 3669
rect 6720 3583 6956 3594
rect 6362 3575 6956 3583
rect 6362 3550 6364 3575
rect 6276 3507 6310 3509
rect 6276 3471 6310 3473
rect 6276 3386 6310 3405
rect 6398 3550 6922 3575
rect 7008 3575 7084 3594
rect 7008 3554 7010 3575
rect 6364 3507 6398 3509
rect 6620 3477 6636 3511
rect 6670 3477 6686 3511
rect 6922 3507 6956 3509
rect 6364 3471 6398 3473
rect 6922 3471 6956 3473
rect 6364 3386 6398 3405
rect 6492 3415 6526 3434
rect 6492 3347 6526 3349
rect 6304 3309 6320 3343
rect 6354 3309 6370 3343
rect 6492 3311 6526 3313
rect 5992 3231 6004 3265
rect 5992 3197 6038 3231
rect 5992 3163 6004 3197
rect 5582 3089 5611 3123
rect 5645 3089 5703 3123
rect 5737 3089 5795 3123
rect 5829 3089 5858 3123
rect 5992 3117 6038 3163
rect 6072 3265 6138 3277
rect 6072 3231 6088 3265
rect 6122 3231 6138 3265
rect 6072 3218 6138 3231
rect 6492 3226 6526 3245
rect 6588 3415 6622 3434
rect 6588 3347 6622 3349
rect 6588 3311 6622 3313
rect 6588 3226 6622 3245
rect 6684 3415 6718 3434
rect 6922 3386 6956 3405
rect 7044 3554 7084 3575
rect 7192 3593 7234 3635
rect 7470 3633 7499 3667
rect 7533 3633 7591 3667
rect 7625 3633 7683 3667
rect 7717 3633 7746 3667
rect 7891 3661 7925 3668
rect 7192 3559 7200 3593
rect 7010 3507 7044 3509
rect 7010 3471 7044 3473
rect 7192 3525 7234 3559
rect 7192 3491 7200 3525
rect 7192 3457 7234 3491
rect 7192 3423 7200 3457
rect 7192 3407 7234 3423
rect 7268 3593 7334 3601
rect 7268 3559 7284 3593
rect 7318 3559 7334 3593
rect 7268 3525 7334 3559
rect 7268 3491 7284 3525
rect 7318 3491 7334 3525
rect 7268 3457 7334 3491
rect 7268 3423 7284 3457
rect 7318 3423 7334 3457
rect 7268 3405 7334 3423
rect 7503 3583 7539 3599
rect 7503 3549 7505 3583
rect 7503 3515 7539 3549
rect 7503 3481 7505 3515
rect 7575 3583 7641 3633
rect 7816 3627 7845 3661
rect 7879 3627 7937 3661
rect 7971 3627 8029 3661
rect 8063 3627 8092 3661
rect 8192 3637 8208 3671
rect 8242 3637 8258 3671
rect 8416 3658 8530 3660
rect 7575 3549 7591 3583
rect 7625 3549 7641 3583
rect 7575 3515 7641 3549
rect 7575 3481 7591 3515
rect 7625 3481 7641 3515
rect 7675 3583 7729 3599
rect 7675 3549 7677 3583
rect 7711 3549 7729 3583
rect 7675 3502 7729 3549
rect 7503 3447 7539 3481
rect 7675 3468 7677 3502
rect 7711 3468 7729 3502
rect 7503 3413 7638 3447
rect 7675 3418 7729 3468
rect 7010 3386 7044 3405
rect 6684 3347 6718 3349
rect 7096 3371 7240 3372
rect 7096 3357 7254 3371
rect 6684 3311 6718 3313
rect 6950 3344 7016 3346
rect 7096 3344 7204 3357
rect 6950 3343 7204 3344
rect 6950 3309 6966 3343
rect 7000 3330 7204 3343
rect 7000 3310 7136 3330
rect 7188 3323 7204 3330
rect 7238 3323 7254 3357
rect 7000 3309 7016 3310
rect 7188 3273 7234 3289
rect 7288 3285 7334 3405
rect 7604 3384 7638 3413
rect 7491 3355 7559 3377
rect 7491 3354 7507 3355
rect 7491 3320 7505 3354
rect 7541 3321 7559 3355
rect 7539 3320 7559 3321
rect 7491 3303 7559 3320
rect 7604 3368 7659 3384
rect 7604 3334 7625 3368
rect 7604 3318 7659 3334
rect 7693 3368 7729 3418
rect 7884 3585 7926 3627
rect 8416 3619 8698 3658
rect 8838 3637 8854 3671
rect 8888 3637 8904 3671
rect 8416 3594 8455 3619
rect 7884 3551 7892 3585
rect 7884 3517 7926 3551
rect 7884 3483 7892 3517
rect 7884 3449 7926 3483
rect 7884 3415 7892 3449
rect 7884 3399 7926 3415
rect 7960 3585 8026 3593
rect 7960 3551 7976 3585
rect 8010 3551 8026 3585
rect 7960 3517 8026 3551
rect 7960 3483 7976 3517
rect 8010 3483 8026 3517
rect 7960 3449 8026 3483
rect 7960 3415 7976 3449
rect 8010 3415 8026 3449
rect 7960 3397 8026 3415
rect 7693 3366 7734 3368
rect 7693 3332 7698 3366
rect 7732 3332 7734 3366
rect 7693 3330 7734 3332
rect 7880 3360 7946 3363
rect 6718 3245 6964 3262
rect 6684 3228 6964 3245
rect 6684 3226 6718 3228
rect 6072 3197 6414 3218
rect 6072 3163 6088 3197
rect 6122 3186 6414 3197
rect 6122 3183 6590 3186
rect 6122 3182 6540 3183
rect 6122 3163 6144 3182
rect 6072 3158 6144 3163
rect 6072 3151 6138 3158
rect 6378 3150 6540 3182
rect 6524 3149 6540 3150
rect 6574 3149 6590 3183
rect 6916 3140 6964 3228
rect 5928 3083 5957 3117
rect 5991 3083 6049 3117
rect 6083 3083 6141 3117
rect 6175 3083 6204 3117
rect 6286 3112 6332 3122
rect 6286 3078 6292 3112
rect 6326 3092 6332 3112
rect 6916 3106 6924 3140
rect 6958 3106 6964 3140
rect 7188 3239 7200 3273
rect 7188 3205 7234 3239
rect 7188 3171 7200 3205
rect 7188 3125 7234 3171
rect 7268 3273 7334 3285
rect 7268 3222 7284 3273
rect 7318 3222 7334 3273
rect 7604 3267 7638 3318
rect 7268 3205 7334 3222
rect 7268 3171 7284 3205
rect 7318 3171 7334 3205
rect 7268 3159 7334 3171
rect 7505 3233 7638 3267
rect 7693 3258 7729 3330
rect 7880 3326 7894 3360
rect 7928 3349 7946 3360
rect 7880 3315 7896 3326
rect 7930 3315 7946 3349
rect 7505 3212 7539 3233
rect 7677 3229 7729 3258
rect 7505 3157 7539 3178
rect 7575 3165 7591 3199
rect 7625 3165 7641 3199
rect 6326 3078 6336 3092
rect 2924 2948 2958 2982
rect 2924 2896 2958 2912
rect 4316 2972 4448 3008
rect 4620 3018 4654 3034
rect 4716 3018 4750 3034
rect 4654 2982 4655 2983
rect 4316 2924 4352 2972
rect 4620 2948 4655 2982
rect 4654 2946 4655 2948
rect 4716 2948 4750 2982
rect 4500 2924 4620 2946
rect 4316 2912 4620 2924
rect 4654 2912 4656 2946
rect 4316 2910 4656 2912
rect 4316 2888 4536 2910
rect 4620 2896 4654 2910
rect 4716 2896 4750 2912
rect 4812 3018 4846 3034
rect 6286 3008 6336 3078
rect 6636 3068 6652 3102
rect 6686 3068 6702 3102
rect 6916 3094 6964 3106
rect 7124 3091 7153 3125
rect 7187 3091 7245 3125
rect 7279 3091 7337 3125
rect 7371 3091 7400 3125
rect 7575 3123 7641 3165
rect 7711 3195 7729 3229
rect 7677 3157 7729 3195
rect 7880 3265 7926 3281
rect 7980 3277 8026 3397
rect 8164 3575 8198 3594
rect 8250 3585 8455 3594
rect 8489 3617 8698 3619
rect 8489 3585 8574 3617
rect 8250 3583 8574 3585
rect 8608 3594 8698 3617
rect 8938 3594 8972 3952
rect 9882 3926 9916 4137
rect 10113 3834 10147 4137
rect 10198 3918 10232 4532
rect 10398 4530 10464 4532
rect 10715 4537 10731 4571
rect 10765 4537 10781 4571
rect 10715 4503 10781 4537
rect 10270 4471 10304 4490
rect 10270 4403 10304 4405
rect 10270 4367 10304 4369
rect 10270 4282 10304 4301
rect 10366 4471 10400 4490
rect 10366 4403 10400 4405
rect 10366 4367 10400 4369
rect 10366 4282 10400 4301
rect 10462 4471 10496 4490
rect 10715 4469 10731 4503
rect 10765 4487 10781 4503
rect 10887 4639 10953 4681
rect 10921 4605 10953 4639
rect 10887 4571 10953 4605
rect 10921 4537 10953 4571
rect 10887 4503 10953 4537
rect 10765 4469 10851 4487
rect 10715 4453 10851 4469
rect 10921 4469 10953 4503
rect 10887 4453 10953 4469
rect 11783 4639 11849 4644
rect 11783 4605 11799 4639
rect 11833 4605 11849 4639
rect 11783 4571 11849 4605
rect 11783 4537 11799 4571
rect 11833 4537 11849 4571
rect 11783 4503 11849 4537
rect 11783 4469 11799 4503
rect 11833 4487 11849 4503
rect 11955 4639 12021 4681
rect 11989 4605 12021 4639
rect 12188 4675 12470 4681
rect 12188 4641 12227 4675
rect 12261 4673 12470 4675
rect 12261 4641 12346 4673
rect 12188 4639 12346 4641
rect 12380 4639 12470 4673
rect 12188 4606 12470 4639
rect 12597 4639 12663 4644
rect 11955 4571 12021 4605
rect 11989 4537 12021 4571
rect 12597 4605 12613 4639
rect 12647 4605 12663 4639
rect 12597 4571 12663 4605
rect 11955 4503 12021 4537
rect 11833 4469 11919 4487
rect 11783 4453 11919 4469
rect 11989 4469 12021 4503
rect 11955 4453 12021 4469
rect 12080 4567 12346 4568
rect 12080 4533 12296 4567
rect 12330 4533 12346 4567
rect 12080 4532 12346 4533
rect 10462 4403 10496 4405
rect 10713 4410 10783 4419
rect 10713 4376 10729 4410
rect 10763 4403 10783 4410
rect 10713 4369 10733 4376
rect 10767 4369 10783 4403
rect 10462 4367 10496 4369
rect 10817 4333 10851 4453
rect 10885 4410 10955 4419
rect 10885 4403 10903 4410
rect 10885 4369 10901 4403
rect 10937 4376 10955 4410
rect 10935 4369 10955 4376
rect 11781 4412 11851 4419
rect 11781 4378 11799 4412
rect 11833 4403 11851 4412
rect 11781 4369 11801 4378
rect 11835 4369 11851 4403
rect 11885 4333 11919 4453
rect 11953 4408 12023 4419
rect 11953 4403 11972 4408
rect 11953 4369 11969 4403
rect 12006 4374 12023 4408
rect 12003 4369 12023 4374
rect 10462 4282 10496 4301
rect 10717 4317 10765 4333
rect 10717 4283 10731 4317
rect 10717 4249 10765 4283
rect 10302 4205 10318 4239
rect 10352 4205 10368 4239
rect 10717 4215 10731 4249
rect 10717 4171 10765 4215
rect 10799 4317 10865 4333
rect 10799 4283 10815 4317
rect 10849 4287 10865 4317
rect 10799 4253 10817 4283
rect 10851 4253 10865 4287
rect 10799 4249 10865 4253
rect 10799 4215 10815 4249
rect 10849 4215 10865 4249
rect 10799 4205 10865 4215
rect 10899 4317 10953 4333
rect 10933 4283 10953 4317
rect 10899 4249 10953 4283
rect 10933 4215 10953 4249
rect 10899 4171 10953 4215
rect 11785 4317 11833 4333
rect 11785 4283 11799 4317
rect 11785 4249 11833 4283
rect 11785 4215 11799 4249
rect 11785 4171 11833 4215
rect 11867 4317 11933 4333
rect 11867 4292 11883 4317
rect 11867 4258 11881 4292
rect 11917 4283 11933 4317
rect 11915 4258 11933 4283
rect 11867 4249 11933 4258
rect 11867 4215 11883 4249
rect 11917 4215 11933 4249
rect 11867 4205 11933 4215
rect 11967 4317 12021 4333
rect 12001 4283 12021 4317
rect 11967 4249 12021 4283
rect 12001 4215 12021 4249
rect 11967 4171 12021 4215
rect 10414 4124 10430 4158
rect 10464 4124 10480 4158
rect 10696 4137 10725 4171
rect 10759 4137 10817 4171
rect 10851 4137 10909 4171
rect 10943 4137 10972 4171
rect 11764 4137 11793 4171
rect 11827 4137 11885 4171
rect 11919 4137 11977 4171
rect 12011 4137 12040 4171
rect 10286 4074 10320 4090
rect 10286 4004 10320 4038
rect 10286 3952 10320 3968
rect 10382 4074 10416 4090
rect 10382 4004 10416 4038
rect 10382 3952 10416 3968
rect 10478 4074 10512 4090
rect 10478 4004 10512 4038
rect 10512 3968 10860 3992
rect 10478 3952 10860 3968
rect 10198 3884 10334 3918
rect 10368 3884 10384 3918
rect 10113 3814 10508 3834
rect 10113 3809 10375 3814
rect 10113 3800 10254 3809
rect 10238 3775 10254 3800
rect 10288 3780 10375 3809
rect 10409 3790 10508 3814
rect 10680 3792 10726 3794
rect 10680 3790 10684 3792
rect 10409 3780 10684 3790
rect 10288 3775 10684 3780
rect 10238 3758 10684 3775
rect 10718 3758 10726 3792
rect 10238 3756 10726 3758
rect 10680 3750 10726 3756
rect 9012 3635 9041 3669
rect 9075 3635 9133 3669
rect 9167 3635 9225 3669
rect 9259 3635 9288 3669
rect 8608 3583 8844 3594
rect 8250 3575 8844 3583
rect 8250 3550 8252 3575
rect 8164 3507 8198 3509
rect 8164 3471 8198 3473
rect 8164 3386 8198 3405
rect 8286 3550 8810 3575
rect 8896 3575 8972 3594
rect 8896 3554 8898 3575
rect 8252 3507 8286 3509
rect 8508 3477 8524 3511
rect 8558 3477 8574 3511
rect 8810 3507 8844 3509
rect 8252 3471 8286 3473
rect 8810 3471 8844 3473
rect 8252 3386 8286 3405
rect 8380 3415 8414 3434
rect 8380 3347 8414 3349
rect 8192 3309 8208 3343
rect 8242 3309 8258 3343
rect 8380 3311 8414 3313
rect 7880 3231 7892 3265
rect 7880 3197 7926 3231
rect 7880 3163 7892 3197
rect 7470 3089 7499 3123
rect 7533 3089 7591 3123
rect 7625 3089 7683 3123
rect 7717 3089 7746 3123
rect 7880 3117 7926 3163
rect 7960 3265 8026 3277
rect 7960 3231 7976 3265
rect 8010 3231 8026 3265
rect 7960 3218 8026 3231
rect 8380 3226 8414 3245
rect 8476 3415 8510 3434
rect 8476 3347 8510 3349
rect 8476 3311 8510 3313
rect 8476 3226 8510 3245
rect 8572 3415 8606 3434
rect 8810 3386 8844 3405
rect 8932 3554 8972 3575
rect 9080 3593 9122 3635
rect 9358 3633 9387 3667
rect 9421 3633 9479 3667
rect 9513 3633 9571 3667
rect 9605 3633 9634 3667
rect 9779 3661 9813 3668
rect 9080 3559 9088 3593
rect 8898 3507 8932 3509
rect 8898 3471 8932 3473
rect 9080 3525 9122 3559
rect 9080 3491 9088 3525
rect 9080 3457 9122 3491
rect 9080 3423 9088 3457
rect 9080 3407 9122 3423
rect 9156 3593 9222 3601
rect 9156 3559 9172 3593
rect 9206 3559 9222 3593
rect 9156 3525 9222 3559
rect 9156 3491 9172 3525
rect 9206 3491 9222 3525
rect 9156 3457 9222 3491
rect 9156 3423 9172 3457
rect 9206 3423 9222 3457
rect 9156 3405 9222 3423
rect 9391 3583 9427 3599
rect 9391 3549 9393 3583
rect 9391 3515 9427 3549
rect 9391 3481 9393 3515
rect 9463 3583 9529 3633
rect 9704 3627 9733 3661
rect 9767 3627 9825 3661
rect 9859 3627 9917 3661
rect 9951 3627 9980 3661
rect 10080 3637 10096 3671
rect 10130 3637 10146 3671
rect 10304 3658 10418 3660
rect 9463 3549 9479 3583
rect 9513 3549 9529 3583
rect 9463 3515 9529 3549
rect 9463 3481 9479 3515
rect 9513 3481 9529 3515
rect 9563 3583 9617 3599
rect 9563 3549 9565 3583
rect 9599 3549 9617 3583
rect 9563 3502 9617 3549
rect 9391 3447 9427 3481
rect 9563 3468 9565 3502
rect 9599 3468 9617 3502
rect 9391 3413 9526 3447
rect 9563 3418 9617 3468
rect 8898 3386 8932 3405
rect 8572 3347 8606 3349
rect 8984 3371 9128 3372
rect 8984 3357 9142 3371
rect 8572 3311 8606 3313
rect 8838 3344 8904 3346
rect 8984 3344 9092 3357
rect 8838 3343 9092 3344
rect 8838 3309 8854 3343
rect 8888 3330 9092 3343
rect 8888 3310 9024 3330
rect 9076 3323 9092 3330
rect 9126 3323 9142 3357
rect 8888 3309 8904 3310
rect 9076 3273 9122 3289
rect 9176 3285 9222 3405
rect 9492 3384 9526 3413
rect 9379 3355 9447 3377
rect 9379 3354 9395 3355
rect 9379 3320 9393 3354
rect 9429 3321 9447 3355
rect 9427 3320 9447 3321
rect 9379 3303 9447 3320
rect 9492 3368 9547 3384
rect 9492 3334 9513 3368
rect 9492 3318 9547 3334
rect 9581 3368 9617 3418
rect 9772 3585 9814 3627
rect 10304 3619 10586 3658
rect 10726 3637 10742 3671
rect 10776 3637 10792 3671
rect 10304 3594 10343 3619
rect 9772 3551 9780 3585
rect 9772 3517 9814 3551
rect 9772 3483 9780 3517
rect 9772 3449 9814 3483
rect 9772 3415 9780 3449
rect 9772 3399 9814 3415
rect 9848 3585 9914 3593
rect 9848 3551 9864 3585
rect 9898 3551 9914 3585
rect 9848 3517 9914 3551
rect 9848 3483 9864 3517
rect 9898 3483 9914 3517
rect 9848 3449 9914 3483
rect 9848 3415 9864 3449
rect 9898 3415 9914 3449
rect 9848 3397 9914 3415
rect 9581 3366 9622 3368
rect 9581 3332 9586 3366
rect 9620 3332 9622 3366
rect 9581 3330 9622 3332
rect 9768 3360 9834 3363
rect 8606 3245 8852 3262
rect 8572 3228 8852 3245
rect 8572 3226 8606 3228
rect 7960 3197 8302 3218
rect 7960 3163 7976 3197
rect 8010 3186 8302 3197
rect 8010 3183 8478 3186
rect 8010 3182 8428 3183
rect 8010 3163 8032 3182
rect 7960 3158 8032 3163
rect 7960 3151 8026 3158
rect 8266 3150 8428 3182
rect 8412 3149 8428 3150
rect 8462 3149 8478 3183
rect 8804 3140 8852 3228
rect 7816 3083 7845 3117
rect 7879 3083 7937 3117
rect 7971 3083 8029 3117
rect 8063 3083 8092 3117
rect 8174 3112 8220 3122
rect 8174 3078 8180 3112
rect 8214 3092 8220 3112
rect 8804 3106 8812 3140
rect 8846 3106 8852 3140
rect 9076 3239 9088 3273
rect 9076 3205 9122 3239
rect 9076 3171 9088 3205
rect 9076 3125 9122 3171
rect 9156 3273 9222 3285
rect 9156 3222 9172 3273
rect 9206 3222 9222 3273
rect 9492 3267 9526 3318
rect 9156 3205 9222 3222
rect 9156 3171 9172 3205
rect 9206 3171 9222 3205
rect 9156 3159 9222 3171
rect 9393 3233 9526 3267
rect 9581 3258 9617 3330
rect 9768 3326 9782 3360
rect 9816 3349 9834 3360
rect 9768 3315 9784 3326
rect 9818 3315 9834 3349
rect 9393 3212 9427 3233
rect 9565 3229 9617 3258
rect 9393 3157 9427 3178
rect 9463 3165 9479 3199
rect 9513 3165 9529 3199
rect 8214 3078 8224 3092
rect 4812 2948 4846 2982
rect 4812 2896 4846 2912
rect 6204 2972 6336 3008
rect 6508 3018 6542 3034
rect 6604 3018 6638 3034
rect 6542 2982 6543 2983
rect 6204 2924 6240 2972
rect 6508 2948 6543 2982
rect 6542 2946 6543 2948
rect 6604 2948 6638 2982
rect 6388 2924 6508 2946
rect 6204 2912 6508 2924
rect 6542 2912 6544 2946
rect 6204 2910 6544 2912
rect 6204 2888 6424 2910
rect 6508 2896 6542 2910
rect 6604 2896 6638 2912
rect 6700 3018 6734 3034
rect 8174 3008 8224 3078
rect 8524 3068 8540 3102
rect 8574 3068 8590 3102
rect 8804 3094 8852 3106
rect 9012 3091 9041 3125
rect 9075 3091 9133 3125
rect 9167 3091 9225 3125
rect 9259 3091 9288 3125
rect 9463 3123 9529 3165
rect 9599 3195 9617 3229
rect 9565 3157 9617 3195
rect 9768 3265 9814 3281
rect 9868 3277 9914 3397
rect 10052 3575 10086 3594
rect 10138 3585 10343 3594
rect 10377 3617 10586 3619
rect 10377 3585 10462 3617
rect 10138 3583 10462 3585
rect 10496 3594 10586 3617
rect 10826 3594 10860 3952
rect 11764 3926 11798 4137
rect 11995 3834 12029 4137
rect 12080 3918 12114 4532
rect 12280 4530 12346 4532
rect 12597 4537 12613 4571
rect 12647 4537 12663 4571
rect 12597 4503 12663 4537
rect 12152 4471 12186 4490
rect 12152 4403 12186 4405
rect 12152 4367 12186 4369
rect 12152 4282 12186 4301
rect 12248 4471 12282 4490
rect 12248 4403 12282 4405
rect 12248 4367 12282 4369
rect 12248 4282 12282 4301
rect 12344 4471 12378 4490
rect 12597 4469 12613 4503
rect 12647 4487 12663 4503
rect 12769 4639 12835 4681
rect 12803 4605 12835 4639
rect 12769 4571 12835 4605
rect 12803 4537 12835 4571
rect 12769 4503 12835 4537
rect 12647 4469 12733 4487
rect 12597 4453 12733 4469
rect 12803 4469 12835 4503
rect 12769 4453 12835 4469
rect 13671 4639 13737 4644
rect 13671 4605 13687 4639
rect 13721 4605 13737 4639
rect 13671 4571 13737 4605
rect 13671 4537 13687 4571
rect 13721 4537 13737 4571
rect 13671 4503 13737 4537
rect 13671 4469 13687 4503
rect 13721 4487 13737 4503
rect 13843 4639 13909 4681
rect 13877 4605 13909 4639
rect 14076 4675 14358 4681
rect 14076 4641 14115 4675
rect 14149 4673 14358 4675
rect 14149 4641 14234 4673
rect 14076 4639 14234 4641
rect 14268 4639 14358 4673
rect 14076 4606 14358 4639
rect 14485 4639 14551 4644
rect 13843 4571 13909 4605
rect 13877 4537 13909 4571
rect 14485 4605 14501 4639
rect 14535 4605 14551 4639
rect 14485 4571 14551 4605
rect 13843 4503 13909 4537
rect 13721 4469 13807 4487
rect 13671 4453 13807 4469
rect 13877 4469 13909 4503
rect 13843 4453 13909 4469
rect 13968 4567 14234 4568
rect 13968 4533 14184 4567
rect 14218 4533 14234 4567
rect 13968 4532 14234 4533
rect 12344 4403 12378 4405
rect 12595 4410 12665 4419
rect 12595 4376 12611 4410
rect 12645 4403 12665 4410
rect 12595 4369 12615 4376
rect 12649 4369 12665 4403
rect 12344 4367 12378 4369
rect 12699 4333 12733 4453
rect 12767 4410 12837 4419
rect 12767 4403 12785 4410
rect 12767 4369 12783 4403
rect 12819 4376 12837 4410
rect 12817 4369 12837 4376
rect 13669 4412 13739 4419
rect 13669 4378 13687 4412
rect 13721 4403 13739 4412
rect 13669 4369 13689 4378
rect 13723 4369 13739 4403
rect 13773 4333 13807 4453
rect 13841 4408 13911 4419
rect 13841 4403 13860 4408
rect 13841 4369 13857 4403
rect 13894 4374 13911 4408
rect 13891 4369 13911 4374
rect 12344 4282 12378 4301
rect 12599 4317 12647 4333
rect 12599 4283 12613 4317
rect 12599 4249 12647 4283
rect 12184 4205 12200 4239
rect 12234 4205 12250 4239
rect 12599 4215 12613 4249
rect 12599 4171 12647 4215
rect 12681 4317 12747 4333
rect 12681 4283 12697 4317
rect 12731 4287 12747 4317
rect 12681 4253 12699 4283
rect 12733 4253 12747 4287
rect 12681 4249 12747 4253
rect 12681 4215 12697 4249
rect 12731 4215 12747 4249
rect 12681 4205 12747 4215
rect 12781 4317 12835 4333
rect 12815 4283 12835 4317
rect 12781 4249 12835 4283
rect 12815 4215 12835 4249
rect 12781 4171 12835 4215
rect 13673 4317 13721 4333
rect 13673 4283 13687 4317
rect 13673 4249 13721 4283
rect 13673 4215 13687 4249
rect 13673 4171 13721 4215
rect 13755 4317 13821 4333
rect 13755 4292 13771 4317
rect 13755 4258 13769 4292
rect 13805 4283 13821 4317
rect 13803 4258 13821 4283
rect 13755 4249 13821 4258
rect 13755 4215 13771 4249
rect 13805 4215 13821 4249
rect 13755 4205 13821 4215
rect 13855 4317 13909 4333
rect 13889 4283 13909 4317
rect 13855 4249 13909 4283
rect 13889 4215 13909 4249
rect 13855 4171 13909 4215
rect 12296 4124 12312 4158
rect 12346 4124 12362 4158
rect 12578 4137 12607 4171
rect 12641 4137 12699 4171
rect 12733 4137 12791 4171
rect 12825 4137 12854 4171
rect 13652 4137 13681 4171
rect 13715 4137 13773 4171
rect 13807 4137 13865 4171
rect 13899 4137 13928 4171
rect 12168 4074 12202 4090
rect 12168 4004 12202 4038
rect 12168 3952 12202 3968
rect 12264 4074 12298 4090
rect 12264 4004 12298 4038
rect 12264 3952 12298 3968
rect 12360 4074 12394 4090
rect 12360 4004 12394 4038
rect 12394 3968 12742 3992
rect 12360 3952 12742 3968
rect 12080 3884 12216 3918
rect 12250 3884 12266 3918
rect 11995 3814 12390 3834
rect 11995 3809 12257 3814
rect 11995 3800 12136 3809
rect 12120 3775 12136 3800
rect 12170 3780 12257 3809
rect 12291 3790 12390 3814
rect 12562 3792 12608 3794
rect 12562 3790 12566 3792
rect 12291 3780 12566 3790
rect 12170 3775 12566 3780
rect 12120 3758 12566 3775
rect 12600 3758 12608 3792
rect 12120 3756 12608 3758
rect 12562 3750 12608 3756
rect 10900 3635 10929 3669
rect 10963 3635 11021 3669
rect 11055 3635 11113 3669
rect 11147 3635 11176 3669
rect 10496 3583 10732 3594
rect 10138 3575 10732 3583
rect 10138 3550 10140 3575
rect 10052 3507 10086 3509
rect 10052 3471 10086 3473
rect 10052 3386 10086 3405
rect 10174 3550 10698 3575
rect 10784 3575 10860 3594
rect 10784 3554 10786 3575
rect 10140 3507 10174 3509
rect 10396 3477 10412 3511
rect 10446 3477 10462 3511
rect 10698 3507 10732 3509
rect 10140 3471 10174 3473
rect 10698 3471 10732 3473
rect 10140 3386 10174 3405
rect 10268 3415 10302 3434
rect 10268 3347 10302 3349
rect 10080 3309 10096 3343
rect 10130 3309 10146 3343
rect 10268 3311 10302 3313
rect 9768 3231 9780 3265
rect 9768 3197 9814 3231
rect 9768 3163 9780 3197
rect 9358 3089 9387 3123
rect 9421 3089 9479 3123
rect 9513 3089 9571 3123
rect 9605 3089 9634 3123
rect 9768 3117 9814 3163
rect 9848 3265 9914 3277
rect 9848 3231 9864 3265
rect 9898 3231 9914 3265
rect 9848 3218 9914 3231
rect 10268 3226 10302 3245
rect 10364 3415 10398 3434
rect 10364 3347 10398 3349
rect 10364 3311 10398 3313
rect 10364 3226 10398 3245
rect 10460 3415 10494 3434
rect 10698 3386 10732 3405
rect 10820 3554 10860 3575
rect 10968 3593 11010 3635
rect 11246 3633 11275 3667
rect 11309 3633 11367 3667
rect 11401 3633 11459 3667
rect 11493 3633 11522 3667
rect 11661 3661 11695 3668
rect 10968 3559 10976 3593
rect 10786 3507 10820 3509
rect 10786 3471 10820 3473
rect 10968 3525 11010 3559
rect 10968 3491 10976 3525
rect 10968 3457 11010 3491
rect 10968 3423 10976 3457
rect 10968 3407 11010 3423
rect 11044 3593 11110 3601
rect 11044 3559 11060 3593
rect 11094 3559 11110 3593
rect 11044 3525 11110 3559
rect 11044 3491 11060 3525
rect 11094 3491 11110 3525
rect 11044 3457 11110 3491
rect 11044 3423 11060 3457
rect 11094 3423 11110 3457
rect 11044 3405 11110 3423
rect 11279 3583 11315 3599
rect 11279 3549 11281 3583
rect 11279 3515 11315 3549
rect 11279 3481 11281 3515
rect 11351 3583 11417 3633
rect 11586 3627 11615 3661
rect 11649 3627 11707 3661
rect 11741 3627 11799 3661
rect 11833 3627 11862 3661
rect 11962 3637 11978 3671
rect 12012 3637 12028 3671
rect 12186 3658 12300 3660
rect 11351 3549 11367 3583
rect 11401 3549 11417 3583
rect 11351 3515 11417 3549
rect 11351 3481 11367 3515
rect 11401 3481 11417 3515
rect 11451 3583 11505 3599
rect 11451 3549 11453 3583
rect 11487 3549 11505 3583
rect 11451 3502 11505 3549
rect 11279 3447 11315 3481
rect 11451 3468 11453 3502
rect 11487 3468 11505 3502
rect 11279 3413 11414 3447
rect 11451 3418 11505 3468
rect 10786 3386 10820 3405
rect 10460 3347 10494 3349
rect 10872 3371 11016 3372
rect 10872 3357 11030 3371
rect 10460 3311 10494 3313
rect 10726 3344 10792 3346
rect 10872 3344 10980 3357
rect 10726 3343 10980 3344
rect 10726 3309 10742 3343
rect 10776 3330 10980 3343
rect 10776 3310 10912 3330
rect 10964 3323 10980 3330
rect 11014 3323 11030 3357
rect 10776 3309 10792 3310
rect 10964 3273 11010 3289
rect 11064 3285 11110 3405
rect 11380 3384 11414 3413
rect 11267 3355 11335 3377
rect 11267 3354 11283 3355
rect 11267 3320 11281 3354
rect 11317 3321 11335 3355
rect 11315 3320 11335 3321
rect 11267 3303 11335 3320
rect 11380 3368 11435 3384
rect 11380 3334 11401 3368
rect 11380 3318 11435 3334
rect 11469 3368 11505 3418
rect 11654 3585 11696 3627
rect 12186 3619 12468 3658
rect 12608 3637 12624 3671
rect 12658 3637 12674 3671
rect 12186 3594 12225 3619
rect 11654 3551 11662 3585
rect 11654 3517 11696 3551
rect 11654 3483 11662 3517
rect 11654 3449 11696 3483
rect 11654 3415 11662 3449
rect 11654 3399 11696 3415
rect 11730 3585 11796 3593
rect 11730 3551 11746 3585
rect 11780 3551 11796 3585
rect 11730 3517 11796 3551
rect 11730 3483 11746 3517
rect 11780 3483 11796 3517
rect 11730 3449 11796 3483
rect 11730 3415 11746 3449
rect 11780 3415 11796 3449
rect 11730 3397 11796 3415
rect 11469 3366 11510 3368
rect 11469 3332 11474 3366
rect 11508 3332 11510 3366
rect 11469 3330 11510 3332
rect 11650 3360 11716 3363
rect 10494 3245 10740 3262
rect 10460 3228 10740 3245
rect 10460 3226 10494 3228
rect 9848 3197 10190 3218
rect 9848 3163 9864 3197
rect 9898 3186 10190 3197
rect 9898 3183 10366 3186
rect 9898 3182 10316 3183
rect 9898 3163 9920 3182
rect 9848 3158 9920 3163
rect 9848 3151 9914 3158
rect 10154 3150 10316 3182
rect 10300 3149 10316 3150
rect 10350 3149 10366 3183
rect 10692 3140 10740 3228
rect 9704 3083 9733 3117
rect 9767 3083 9825 3117
rect 9859 3083 9917 3117
rect 9951 3083 9980 3117
rect 10062 3112 10108 3122
rect 10062 3078 10068 3112
rect 10102 3092 10108 3112
rect 10692 3106 10700 3140
rect 10734 3106 10740 3140
rect 10964 3239 10976 3273
rect 10964 3205 11010 3239
rect 10964 3171 10976 3205
rect 10964 3125 11010 3171
rect 11044 3273 11110 3285
rect 11044 3222 11060 3273
rect 11094 3222 11110 3273
rect 11380 3267 11414 3318
rect 11044 3205 11110 3222
rect 11044 3171 11060 3205
rect 11094 3171 11110 3205
rect 11044 3159 11110 3171
rect 11281 3233 11414 3267
rect 11469 3258 11505 3330
rect 11650 3326 11664 3360
rect 11698 3349 11716 3360
rect 11650 3315 11666 3326
rect 11700 3315 11716 3349
rect 11281 3212 11315 3233
rect 11453 3229 11505 3258
rect 11281 3157 11315 3178
rect 11351 3165 11367 3199
rect 11401 3165 11417 3199
rect 10102 3078 10112 3092
rect 6700 2948 6734 2982
rect 6700 2896 6734 2912
rect 8092 2972 8224 3008
rect 8396 3018 8430 3034
rect 8492 3018 8526 3034
rect 8430 2982 8431 2983
rect 8092 2924 8128 2972
rect 8396 2948 8431 2982
rect 8430 2946 8431 2948
rect 8492 2948 8526 2982
rect 8276 2924 8396 2946
rect 8092 2912 8396 2924
rect 8430 2912 8432 2946
rect 8092 2910 8432 2912
rect 8092 2888 8312 2910
rect 8396 2896 8430 2910
rect 8492 2896 8526 2912
rect 8588 3018 8622 3034
rect 10062 3008 10112 3078
rect 10412 3068 10428 3102
rect 10462 3068 10478 3102
rect 10692 3094 10740 3106
rect 10900 3091 10929 3125
rect 10963 3091 11021 3125
rect 11055 3091 11113 3125
rect 11147 3091 11176 3125
rect 11351 3123 11417 3165
rect 11487 3195 11505 3229
rect 11453 3157 11505 3195
rect 11650 3265 11696 3281
rect 11750 3277 11796 3397
rect 11934 3575 11968 3594
rect 12020 3585 12225 3594
rect 12259 3617 12468 3619
rect 12259 3585 12344 3617
rect 12020 3583 12344 3585
rect 12378 3594 12468 3617
rect 12708 3594 12742 3952
rect 13652 3926 13686 4137
rect 13883 3834 13917 4137
rect 13968 3918 14002 4532
rect 14168 4530 14234 4532
rect 14485 4537 14501 4571
rect 14535 4537 14551 4571
rect 14485 4503 14551 4537
rect 14040 4471 14074 4490
rect 14040 4403 14074 4405
rect 14040 4367 14074 4369
rect 14040 4282 14074 4301
rect 14136 4471 14170 4490
rect 14136 4403 14170 4405
rect 14136 4367 14170 4369
rect 14136 4282 14170 4301
rect 14232 4471 14266 4490
rect 14485 4469 14501 4503
rect 14535 4487 14551 4503
rect 14657 4639 14723 4681
rect 14691 4605 14723 4639
rect 14657 4571 14723 4605
rect 14691 4537 14723 4571
rect 14657 4503 14723 4537
rect 14535 4469 14621 4487
rect 14485 4453 14621 4469
rect 14691 4469 14723 4503
rect 14657 4453 14723 4469
rect 15559 4639 15625 4644
rect 15559 4605 15575 4639
rect 15609 4605 15625 4639
rect 15559 4571 15625 4605
rect 15559 4537 15575 4571
rect 15609 4537 15625 4571
rect 15559 4503 15625 4537
rect 15559 4469 15575 4503
rect 15609 4487 15625 4503
rect 15731 4639 15797 4681
rect 15765 4605 15797 4639
rect 15964 4675 16246 4681
rect 15964 4641 16003 4675
rect 16037 4673 16246 4675
rect 16037 4641 16122 4673
rect 15964 4639 16122 4641
rect 16156 4639 16246 4673
rect 15964 4606 16246 4639
rect 16373 4639 16439 4644
rect 15731 4571 15797 4605
rect 15765 4537 15797 4571
rect 16373 4605 16389 4639
rect 16423 4605 16439 4639
rect 16373 4571 16439 4605
rect 15731 4503 15797 4537
rect 15609 4469 15695 4487
rect 15559 4453 15695 4469
rect 15765 4469 15797 4503
rect 15731 4453 15797 4469
rect 15856 4567 16122 4568
rect 15856 4533 16072 4567
rect 16106 4533 16122 4567
rect 15856 4532 16122 4533
rect 14232 4403 14266 4405
rect 14483 4410 14553 4419
rect 14483 4376 14499 4410
rect 14533 4403 14553 4410
rect 14483 4369 14503 4376
rect 14537 4369 14553 4403
rect 14232 4367 14266 4369
rect 14587 4333 14621 4453
rect 14655 4410 14725 4419
rect 14655 4403 14673 4410
rect 14655 4369 14671 4403
rect 14707 4376 14725 4410
rect 14705 4369 14725 4376
rect 15557 4412 15627 4419
rect 15557 4378 15575 4412
rect 15609 4403 15627 4412
rect 15557 4369 15577 4378
rect 15611 4369 15627 4403
rect 15661 4333 15695 4453
rect 15729 4408 15799 4419
rect 15729 4403 15748 4408
rect 15729 4369 15745 4403
rect 15782 4374 15799 4408
rect 15779 4369 15799 4374
rect 14232 4282 14266 4301
rect 14487 4317 14535 4333
rect 14487 4283 14501 4317
rect 14487 4249 14535 4283
rect 14072 4205 14088 4239
rect 14122 4205 14138 4239
rect 14487 4215 14501 4249
rect 14487 4171 14535 4215
rect 14569 4317 14635 4333
rect 14569 4283 14585 4317
rect 14619 4287 14635 4317
rect 14569 4253 14587 4283
rect 14621 4253 14635 4287
rect 14569 4249 14635 4253
rect 14569 4215 14585 4249
rect 14619 4215 14635 4249
rect 14569 4205 14635 4215
rect 14669 4317 14723 4333
rect 14703 4283 14723 4317
rect 14669 4249 14723 4283
rect 14703 4215 14723 4249
rect 14669 4171 14723 4215
rect 15561 4317 15609 4333
rect 15561 4283 15575 4317
rect 15561 4249 15609 4283
rect 15561 4215 15575 4249
rect 15561 4171 15609 4215
rect 15643 4317 15709 4333
rect 15643 4292 15659 4317
rect 15643 4258 15657 4292
rect 15693 4283 15709 4317
rect 15691 4258 15709 4283
rect 15643 4249 15709 4258
rect 15643 4215 15659 4249
rect 15693 4215 15709 4249
rect 15643 4205 15709 4215
rect 15743 4317 15797 4333
rect 15777 4283 15797 4317
rect 15743 4249 15797 4283
rect 15777 4215 15797 4249
rect 15743 4171 15797 4215
rect 14184 4124 14200 4158
rect 14234 4124 14250 4158
rect 14466 4137 14495 4171
rect 14529 4137 14587 4171
rect 14621 4137 14679 4171
rect 14713 4137 14742 4171
rect 15540 4137 15569 4171
rect 15603 4137 15661 4171
rect 15695 4137 15753 4171
rect 15787 4137 15816 4171
rect 14056 4074 14090 4090
rect 14056 4004 14090 4038
rect 14056 3952 14090 3968
rect 14152 4074 14186 4090
rect 14152 4004 14186 4038
rect 14152 3952 14186 3968
rect 14248 4074 14282 4090
rect 14248 4004 14282 4038
rect 14282 3968 14630 3992
rect 14248 3952 14630 3968
rect 13968 3884 14104 3918
rect 14138 3884 14154 3918
rect 13883 3814 14278 3834
rect 13883 3809 14145 3814
rect 13883 3800 14024 3809
rect 14008 3775 14024 3800
rect 14058 3780 14145 3809
rect 14179 3790 14278 3814
rect 14450 3792 14496 3794
rect 14450 3790 14454 3792
rect 14179 3780 14454 3790
rect 14058 3775 14454 3780
rect 14008 3758 14454 3775
rect 14488 3758 14496 3792
rect 14008 3756 14496 3758
rect 14450 3750 14496 3756
rect 12782 3635 12811 3669
rect 12845 3635 12903 3669
rect 12937 3635 12995 3669
rect 13029 3635 13058 3669
rect 12378 3583 12614 3594
rect 12020 3575 12614 3583
rect 12020 3550 12022 3575
rect 11934 3507 11968 3509
rect 11934 3471 11968 3473
rect 11934 3386 11968 3405
rect 12056 3550 12580 3575
rect 12666 3575 12742 3594
rect 12666 3554 12668 3575
rect 12022 3507 12056 3509
rect 12278 3477 12294 3511
rect 12328 3477 12344 3511
rect 12580 3507 12614 3509
rect 12022 3471 12056 3473
rect 12580 3471 12614 3473
rect 12022 3386 12056 3405
rect 12150 3415 12184 3434
rect 12150 3347 12184 3349
rect 11962 3309 11978 3343
rect 12012 3309 12028 3343
rect 12150 3311 12184 3313
rect 11650 3231 11662 3265
rect 11650 3197 11696 3231
rect 11650 3163 11662 3197
rect 11246 3089 11275 3123
rect 11309 3089 11367 3123
rect 11401 3089 11459 3123
rect 11493 3089 11522 3123
rect 11650 3117 11696 3163
rect 11730 3265 11796 3277
rect 11730 3231 11746 3265
rect 11780 3231 11796 3265
rect 11730 3218 11796 3231
rect 12150 3226 12184 3245
rect 12246 3415 12280 3434
rect 12246 3347 12280 3349
rect 12246 3311 12280 3313
rect 12246 3226 12280 3245
rect 12342 3415 12376 3434
rect 12580 3386 12614 3405
rect 12702 3554 12742 3575
rect 12850 3593 12892 3635
rect 13128 3633 13157 3667
rect 13191 3633 13249 3667
rect 13283 3633 13341 3667
rect 13375 3633 13404 3667
rect 13549 3661 13583 3668
rect 12850 3559 12858 3593
rect 12668 3507 12702 3509
rect 12668 3471 12702 3473
rect 12850 3525 12892 3559
rect 12850 3491 12858 3525
rect 12850 3457 12892 3491
rect 12850 3423 12858 3457
rect 12850 3407 12892 3423
rect 12926 3593 12992 3601
rect 12926 3559 12942 3593
rect 12976 3559 12992 3593
rect 12926 3525 12992 3559
rect 12926 3491 12942 3525
rect 12976 3491 12992 3525
rect 12926 3457 12992 3491
rect 12926 3423 12942 3457
rect 12976 3423 12992 3457
rect 12926 3405 12992 3423
rect 13161 3583 13197 3599
rect 13161 3549 13163 3583
rect 13161 3515 13197 3549
rect 13161 3481 13163 3515
rect 13233 3583 13299 3633
rect 13474 3627 13503 3661
rect 13537 3627 13595 3661
rect 13629 3627 13687 3661
rect 13721 3627 13750 3661
rect 13850 3637 13866 3671
rect 13900 3637 13916 3671
rect 14074 3658 14188 3660
rect 13233 3549 13249 3583
rect 13283 3549 13299 3583
rect 13233 3515 13299 3549
rect 13233 3481 13249 3515
rect 13283 3481 13299 3515
rect 13333 3583 13387 3599
rect 13333 3549 13335 3583
rect 13369 3549 13387 3583
rect 13333 3502 13387 3549
rect 13161 3447 13197 3481
rect 13333 3468 13335 3502
rect 13369 3468 13387 3502
rect 13161 3413 13296 3447
rect 13333 3418 13387 3468
rect 12668 3386 12702 3405
rect 12342 3347 12376 3349
rect 12754 3371 12898 3372
rect 12754 3357 12912 3371
rect 12342 3311 12376 3313
rect 12608 3344 12674 3346
rect 12754 3344 12862 3357
rect 12608 3343 12862 3344
rect 12608 3309 12624 3343
rect 12658 3330 12862 3343
rect 12658 3310 12794 3330
rect 12846 3323 12862 3330
rect 12896 3323 12912 3357
rect 12658 3309 12674 3310
rect 12846 3273 12892 3289
rect 12946 3285 12992 3405
rect 13262 3384 13296 3413
rect 13149 3355 13217 3377
rect 13149 3354 13165 3355
rect 13149 3320 13163 3354
rect 13199 3321 13217 3355
rect 13197 3320 13217 3321
rect 13149 3303 13217 3320
rect 13262 3368 13317 3384
rect 13262 3334 13283 3368
rect 13262 3318 13317 3334
rect 13351 3368 13387 3418
rect 13542 3585 13584 3627
rect 14074 3619 14356 3658
rect 14496 3637 14512 3671
rect 14546 3637 14562 3671
rect 14074 3594 14113 3619
rect 13542 3551 13550 3585
rect 13542 3517 13584 3551
rect 13542 3483 13550 3517
rect 13542 3449 13584 3483
rect 13542 3415 13550 3449
rect 13542 3399 13584 3415
rect 13618 3585 13684 3593
rect 13618 3551 13634 3585
rect 13668 3551 13684 3585
rect 13618 3517 13684 3551
rect 13618 3483 13634 3517
rect 13668 3483 13684 3517
rect 13618 3449 13684 3483
rect 13618 3415 13634 3449
rect 13668 3415 13684 3449
rect 13618 3397 13684 3415
rect 13351 3366 13392 3368
rect 13351 3332 13356 3366
rect 13390 3332 13392 3366
rect 13351 3330 13392 3332
rect 13538 3360 13604 3363
rect 12376 3245 12622 3262
rect 12342 3228 12622 3245
rect 12342 3226 12376 3228
rect 11730 3197 12072 3218
rect 11730 3163 11746 3197
rect 11780 3186 12072 3197
rect 11780 3183 12248 3186
rect 11780 3182 12198 3183
rect 11780 3163 11802 3182
rect 11730 3158 11802 3163
rect 11730 3151 11796 3158
rect 12036 3150 12198 3182
rect 12182 3149 12198 3150
rect 12232 3149 12248 3183
rect 12574 3140 12622 3228
rect 11586 3083 11615 3117
rect 11649 3083 11707 3117
rect 11741 3083 11799 3117
rect 11833 3083 11862 3117
rect 11944 3112 11990 3122
rect 11944 3078 11950 3112
rect 11984 3092 11990 3112
rect 12574 3106 12582 3140
rect 12616 3106 12622 3140
rect 12846 3239 12858 3273
rect 12846 3205 12892 3239
rect 12846 3171 12858 3205
rect 12846 3125 12892 3171
rect 12926 3273 12992 3285
rect 12926 3222 12942 3273
rect 12976 3222 12992 3273
rect 13262 3267 13296 3318
rect 12926 3205 12992 3222
rect 12926 3171 12942 3205
rect 12976 3171 12992 3205
rect 12926 3159 12992 3171
rect 13163 3233 13296 3267
rect 13351 3258 13387 3330
rect 13538 3326 13552 3360
rect 13586 3349 13604 3360
rect 13538 3315 13554 3326
rect 13588 3315 13604 3349
rect 13163 3212 13197 3233
rect 13335 3229 13387 3258
rect 13163 3157 13197 3178
rect 13233 3165 13249 3199
rect 13283 3165 13299 3199
rect 11984 3078 11994 3092
rect 8588 2948 8622 2982
rect 8588 2896 8622 2912
rect 9980 2972 10112 3008
rect 10284 3018 10318 3034
rect 10380 3018 10414 3034
rect 10318 2982 10319 2983
rect 9980 2924 10016 2972
rect 10284 2948 10319 2982
rect 10318 2946 10319 2948
rect 10380 2948 10414 2982
rect 10164 2924 10284 2946
rect 9980 2912 10284 2924
rect 10318 2912 10320 2946
rect 9980 2910 10320 2912
rect 9980 2888 10200 2910
rect 10284 2896 10318 2910
rect 10380 2896 10414 2912
rect 10476 3018 10510 3034
rect 11944 3008 11994 3078
rect 12294 3068 12310 3102
rect 12344 3068 12360 3102
rect 12574 3094 12622 3106
rect 12782 3091 12811 3125
rect 12845 3091 12903 3125
rect 12937 3091 12995 3125
rect 13029 3091 13058 3125
rect 13233 3123 13299 3165
rect 13369 3195 13387 3229
rect 13335 3157 13387 3195
rect 13538 3265 13584 3281
rect 13638 3277 13684 3397
rect 13822 3575 13856 3594
rect 13908 3585 14113 3594
rect 14147 3617 14356 3619
rect 14147 3585 14232 3617
rect 13908 3583 14232 3585
rect 14266 3594 14356 3617
rect 14596 3594 14630 3952
rect 15540 3926 15574 4137
rect 15771 3834 15805 4137
rect 15856 3918 15890 4532
rect 16056 4530 16122 4532
rect 16373 4537 16389 4571
rect 16423 4537 16439 4571
rect 16373 4503 16439 4537
rect 15928 4471 15962 4490
rect 15928 4403 15962 4405
rect 15928 4367 15962 4369
rect 15928 4282 15962 4301
rect 16024 4471 16058 4490
rect 16024 4403 16058 4405
rect 16024 4367 16058 4369
rect 16024 4282 16058 4301
rect 16120 4471 16154 4490
rect 16373 4469 16389 4503
rect 16423 4487 16439 4503
rect 16545 4639 16611 4681
rect 16579 4605 16611 4639
rect 16545 4571 16611 4605
rect 16579 4537 16611 4571
rect 16545 4503 16611 4537
rect 16423 4469 16509 4487
rect 16373 4453 16509 4469
rect 16579 4469 16611 4503
rect 16545 4453 16611 4469
rect 17447 4639 17513 4644
rect 17447 4605 17463 4639
rect 17497 4605 17513 4639
rect 17447 4571 17513 4605
rect 17447 4537 17463 4571
rect 17497 4537 17513 4571
rect 17447 4503 17513 4537
rect 17447 4469 17463 4503
rect 17497 4487 17513 4503
rect 17619 4639 17685 4681
rect 17653 4605 17685 4639
rect 17852 4675 18134 4681
rect 17852 4641 17891 4675
rect 17925 4673 18134 4675
rect 17925 4641 18010 4673
rect 17852 4639 18010 4641
rect 18044 4639 18134 4673
rect 17852 4606 18134 4639
rect 18261 4639 18327 4644
rect 17619 4571 17685 4605
rect 17653 4537 17685 4571
rect 18261 4605 18277 4639
rect 18311 4605 18327 4639
rect 18261 4571 18327 4605
rect 17619 4503 17685 4537
rect 17497 4469 17583 4487
rect 17447 4453 17583 4469
rect 17653 4469 17685 4503
rect 17619 4453 17685 4469
rect 17744 4567 18010 4568
rect 17744 4533 17960 4567
rect 17994 4533 18010 4567
rect 17744 4532 18010 4533
rect 16120 4403 16154 4405
rect 16371 4410 16441 4419
rect 16371 4376 16387 4410
rect 16421 4403 16441 4410
rect 16371 4369 16391 4376
rect 16425 4369 16441 4403
rect 16120 4367 16154 4369
rect 16475 4333 16509 4453
rect 16543 4410 16613 4419
rect 16543 4403 16561 4410
rect 16543 4369 16559 4403
rect 16595 4376 16613 4410
rect 16593 4369 16613 4376
rect 17445 4412 17515 4419
rect 17445 4378 17463 4412
rect 17497 4403 17515 4412
rect 17445 4369 17465 4378
rect 17499 4369 17515 4403
rect 17549 4333 17583 4453
rect 17617 4408 17687 4419
rect 17617 4403 17636 4408
rect 17617 4369 17633 4403
rect 17670 4374 17687 4408
rect 17667 4369 17687 4374
rect 16120 4282 16154 4301
rect 16375 4317 16423 4333
rect 16375 4283 16389 4317
rect 16375 4249 16423 4283
rect 15960 4205 15976 4239
rect 16010 4205 16026 4239
rect 16375 4215 16389 4249
rect 16375 4171 16423 4215
rect 16457 4317 16523 4333
rect 16457 4283 16473 4317
rect 16507 4287 16523 4317
rect 16457 4253 16475 4283
rect 16509 4253 16523 4287
rect 16457 4249 16523 4253
rect 16457 4215 16473 4249
rect 16507 4215 16523 4249
rect 16457 4205 16523 4215
rect 16557 4317 16611 4333
rect 16591 4283 16611 4317
rect 16557 4249 16611 4283
rect 16591 4215 16611 4249
rect 16557 4171 16611 4215
rect 17449 4317 17497 4333
rect 17449 4283 17463 4317
rect 17449 4249 17497 4283
rect 17449 4215 17463 4249
rect 17449 4171 17497 4215
rect 17531 4317 17597 4333
rect 17531 4292 17547 4317
rect 17531 4258 17545 4292
rect 17581 4283 17597 4317
rect 17579 4258 17597 4283
rect 17531 4249 17597 4258
rect 17531 4215 17547 4249
rect 17581 4215 17597 4249
rect 17531 4205 17597 4215
rect 17631 4317 17685 4333
rect 17665 4283 17685 4317
rect 17631 4249 17685 4283
rect 17665 4215 17685 4249
rect 17631 4171 17685 4215
rect 16072 4124 16088 4158
rect 16122 4124 16138 4158
rect 16354 4137 16383 4171
rect 16417 4137 16475 4171
rect 16509 4137 16567 4171
rect 16601 4137 16630 4171
rect 17428 4137 17457 4171
rect 17491 4137 17549 4171
rect 17583 4137 17641 4171
rect 17675 4137 17704 4171
rect 15944 4074 15978 4090
rect 15944 4004 15978 4038
rect 15944 3952 15978 3968
rect 16040 4074 16074 4090
rect 16040 4004 16074 4038
rect 16040 3952 16074 3968
rect 16136 4074 16170 4090
rect 16136 4004 16170 4038
rect 16170 3968 16518 3992
rect 16136 3952 16518 3968
rect 15856 3884 15992 3918
rect 16026 3884 16042 3918
rect 15771 3814 16166 3834
rect 15771 3809 16033 3814
rect 15771 3800 15912 3809
rect 15896 3775 15912 3800
rect 15946 3780 16033 3809
rect 16067 3790 16166 3814
rect 16338 3792 16384 3794
rect 16338 3790 16342 3792
rect 16067 3780 16342 3790
rect 15946 3775 16342 3780
rect 15896 3758 16342 3775
rect 16376 3758 16384 3792
rect 15896 3756 16384 3758
rect 16338 3750 16384 3756
rect 14670 3635 14699 3669
rect 14733 3635 14791 3669
rect 14825 3635 14883 3669
rect 14917 3635 14946 3669
rect 14266 3583 14502 3594
rect 13908 3575 14502 3583
rect 13908 3550 13910 3575
rect 13822 3507 13856 3509
rect 13822 3471 13856 3473
rect 13822 3386 13856 3405
rect 13944 3550 14468 3575
rect 14554 3575 14630 3594
rect 14554 3554 14556 3575
rect 13910 3507 13944 3509
rect 14166 3477 14182 3511
rect 14216 3477 14232 3511
rect 14468 3507 14502 3509
rect 13910 3471 13944 3473
rect 14468 3471 14502 3473
rect 13910 3386 13944 3405
rect 14038 3415 14072 3434
rect 14038 3347 14072 3349
rect 13850 3309 13866 3343
rect 13900 3309 13916 3343
rect 14038 3311 14072 3313
rect 13538 3231 13550 3265
rect 13538 3197 13584 3231
rect 13538 3163 13550 3197
rect 13128 3089 13157 3123
rect 13191 3089 13249 3123
rect 13283 3089 13341 3123
rect 13375 3089 13404 3123
rect 13538 3117 13584 3163
rect 13618 3265 13684 3277
rect 13618 3231 13634 3265
rect 13668 3231 13684 3265
rect 13618 3218 13684 3231
rect 14038 3226 14072 3245
rect 14134 3415 14168 3434
rect 14134 3347 14168 3349
rect 14134 3311 14168 3313
rect 14134 3226 14168 3245
rect 14230 3415 14264 3434
rect 14468 3386 14502 3405
rect 14590 3554 14630 3575
rect 14738 3593 14780 3635
rect 15016 3633 15045 3667
rect 15079 3633 15137 3667
rect 15171 3633 15229 3667
rect 15263 3633 15292 3667
rect 15437 3661 15471 3668
rect 14738 3559 14746 3593
rect 14556 3507 14590 3509
rect 14556 3471 14590 3473
rect 14738 3525 14780 3559
rect 14738 3491 14746 3525
rect 14738 3457 14780 3491
rect 14738 3423 14746 3457
rect 14738 3407 14780 3423
rect 14814 3593 14880 3601
rect 14814 3559 14830 3593
rect 14864 3559 14880 3593
rect 14814 3525 14880 3559
rect 14814 3491 14830 3525
rect 14864 3491 14880 3525
rect 14814 3457 14880 3491
rect 14814 3423 14830 3457
rect 14864 3423 14880 3457
rect 14814 3405 14880 3423
rect 15049 3583 15085 3599
rect 15049 3549 15051 3583
rect 15049 3515 15085 3549
rect 15049 3481 15051 3515
rect 15121 3583 15187 3633
rect 15362 3627 15391 3661
rect 15425 3627 15483 3661
rect 15517 3627 15575 3661
rect 15609 3627 15638 3661
rect 15738 3637 15754 3671
rect 15788 3637 15804 3671
rect 15962 3658 16076 3660
rect 15121 3549 15137 3583
rect 15171 3549 15187 3583
rect 15121 3515 15187 3549
rect 15121 3481 15137 3515
rect 15171 3481 15187 3515
rect 15221 3583 15275 3599
rect 15221 3549 15223 3583
rect 15257 3549 15275 3583
rect 15221 3502 15275 3549
rect 15049 3447 15085 3481
rect 15221 3468 15223 3502
rect 15257 3468 15275 3502
rect 15049 3413 15184 3447
rect 15221 3418 15275 3468
rect 14556 3386 14590 3405
rect 14230 3347 14264 3349
rect 14642 3371 14786 3372
rect 14642 3357 14800 3371
rect 14230 3311 14264 3313
rect 14496 3344 14562 3346
rect 14642 3344 14750 3357
rect 14496 3343 14750 3344
rect 14496 3309 14512 3343
rect 14546 3330 14750 3343
rect 14546 3310 14682 3330
rect 14734 3323 14750 3330
rect 14784 3323 14800 3357
rect 14546 3309 14562 3310
rect 14734 3273 14780 3289
rect 14834 3285 14880 3405
rect 15150 3384 15184 3413
rect 15037 3355 15105 3377
rect 15037 3354 15053 3355
rect 15037 3320 15051 3354
rect 15087 3321 15105 3355
rect 15085 3320 15105 3321
rect 15037 3303 15105 3320
rect 15150 3368 15205 3384
rect 15150 3334 15171 3368
rect 15150 3318 15205 3334
rect 15239 3368 15275 3418
rect 15430 3585 15472 3627
rect 15962 3619 16244 3658
rect 16384 3637 16400 3671
rect 16434 3637 16450 3671
rect 15962 3594 16001 3619
rect 15430 3551 15438 3585
rect 15430 3517 15472 3551
rect 15430 3483 15438 3517
rect 15430 3449 15472 3483
rect 15430 3415 15438 3449
rect 15430 3399 15472 3415
rect 15506 3585 15572 3593
rect 15506 3551 15522 3585
rect 15556 3551 15572 3585
rect 15506 3517 15572 3551
rect 15506 3483 15522 3517
rect 15556 3483 15572 3517
rect 15506 3449 15572 3483
rect 15506 3415 15522 3449
rect 15556 3415 15572 3449
rect 15506 3397 15572 3415
rect 15239 3366 15280 3368
rect 15239 3332 15244 3366
rect 15278 3332 15280 3366
rect 15239 3330 15280 3332
rect 15426 3360 15492 3363
rect 14264 3245 14510 3262
rect 14230 3228 14510 3245
rect 14230 3226 14264 3228
rect 13618 3197 13960 3218
rect 13618 3163 13634 3197
rect 13668 3186 13960 3197
rect 13668 3183 14136 3186
rect 13668 3182 14086 3183
rect 13668 3163 13690 3182
rect 13618 3158 13690 3163
rect 13618 3151 13684 3158
rect 13924 3150 14086 3182
rect 14070 3149 14086 3150
rect 14120 3149 14136 3183
rect 14462 3140 14510 3228
rect 13474 3083 13503 3117
rect 13537 3083 13595 3117
rect 13629 3083 13687 3117
rect 13721 3083 13750 3117
rect 13832 3112 13878 3122
rect 13832 3078 13838 3112
rect 13872 3092 13878 3112
rect 14462 3106 14470 3140
rect 14504 3106 14510 3140
rect 14734 3239 14746 3273
rect 14734 3205 14780 3239
rect 14734 3171 14746 3205
rect 14734 3125 14780 3171
rect 14814 3273 14880 3285
rect 14814 3222 14830 3273
rect 14864 3222 14880 3273
rect 15150 3267 15184 3318
rect 14814 3205 14880 3222
rect 14814 3171 14830 3205
rect 14864 3171 14880 3205
rect 14814 3159 14880 3171
rect 15051 3233 15184 3267
rect 15239 3258 15275 3330
rect 15426 3326 15440 3360
rect 15474 3349 15492 3360
rect 15426 3315 15442 3326
rect 15476 3315 15492 3349
rect 15051 3212 15085 3233
rect 15223 3229 15275 3258
rect 15051 3157 15085 3178
rect 15121 3165 15137 3199
rect 15171 3165 15187 3199
rect 13872 3078 13882 3092
rect 10476 2948 10510 2982
rect 10476 2896 10510 2912
rect 11862 2972 11994 3008
rect 12166 3018 12200 3034
rect 12262 3018 12296 3034
rect 12200 2982 12201 2983
rect 11862 2924 11898 2972
rect 12166 2948 12201 2982
rect 12200 2946 12201 2948
rect 12262 2948 12296 2982
rect 12046 2924 12166 2946
rect 11862 2912 12166 2924
rect 12200 2912 12202 2946
rect 11862 2910 12202 2912
rect 11862 2888 12082 2910
rect 12166 2896 12200 2910
rect 12262 2896 12296 2912
rect 12358 3018 12392 3034
rect 13832 3008 13882 3078
rect 14182 3068 14198 3102
rect 14232 3068 14248 3102
rect 14462 3094 14510 3106
rect 14670 3091 14699 3125
rect 14733 3091 14791 3125
rect 14825 3091 14883 3125
rect 14917 3091 14946 3125
rect 15121 3123 15187 3165
rect 15257 3195 15275 3229
rect 15223 3157 15275 3195
rect 15426 3265 15472 3281
rect 15526 3277 15572 3397
rect 15710 3575 15744 3594
rect 15796 3585 16001 3594
rect 16035 3617 16244 3619
rect 16035 3585 16120 3617
rect 15796 3583 16120 3585
rect 16154 3594 16244 3617
rect 16484 3594 16518 3952
rect 17428 3926 17462 4137
rect 17659 3834 17693 4137
rect 17744 3918 17778 4532
rect 17944 4530 18010 4532
rect 18261 4537 18277 4571
rect 18311 4537 18327 4571
rect 18261 4503 18327 4537
rect 17816 4471 17850 4490
rect 17816 4403 17850 4405
rect 17816 4367 17850 4369
rect 17816 4282 17850 4301
rect 17912 4471 17946 4490
rect 17912 4403 17946 4405
rect 17912 4367 17946 4369
rect 17912 4282 17946 4301
rect 18008 4471 18042 4490
rect 18261 4469 18277 4503
rect 18311 4487 18327 4503
rect 18433 4639 18499 4681
rect 18467 4605 18499 4639
rect 18433 4571 18499 4605
rect 18467 4537 18499 4571
rect 18433 4503 18499 4537
rect 18311 4469 18397 4487
rect 18261 4453 18397 4469
rect 18467 4469 18499 4503
rect 18433 4453 18499 4469
rect 19335 4639 19401 4644
rect 19335 4605 19351 4639
rect 19385 4605 19401 4639
rect 19335 4571 19401 4605
rect 19335 4537 19351 4571
rect 19385 4537 19401 4571
rect 19335 4503 19401 4537
rect 19335 4469 19351 4503
rect 19385 4487 19401 4503
rect 19507 4639 19573 4681
rect 19541 4605 19573 4639
rect 19740 4675 20022 4681
rect 19740 4641 19779 4675
rect 19813 4673 20022 4675
rect 19813 4641 19898 4673
rect 19740 4639 19898 4641
rect 19932 4639 20022 4673
rect 19740 4606 20022 4639
rect 20149 4639 20215 4644
rect 19507 4571 19573 4605
rect 19541 4537 19573 4571
rect 20149 4605 20165 4639
rect 20199 4605 20215 4639
rect 20149 4571 20215 4605
rect 19507 4503 19573 4537
rect 19385 4469 19471 4487
rect 19335 4453 19471 4469
rect 19541 4469 19573 4503
rect 19507 4453 19573 4469
rect 19632 4567 19898 4568
rect 19632 4533 19848 4567
rect 19882 4533 19898 4567
rect 19632 4532 19898 4533
rect 18008 4403 18042 4405
rect 18259 4410 18329 4419
rect 18259 4376 18275 4410
rect 18309 4403 18329 4410
rect 18259 4369 18279 4376
rect 18313 4369 18329 4403
rect 18008 4367 18042 4369
rect 18363 4333 18397 4453
rect 18431 4410 18501 4419
rect 18431 4403 18449 4410
rect 18431 4369 18447 4403
rect 18483 4376 18501 4410
rect 18481 4369 18501 4376
rect 19333 4412 19403 4419
rect 19333 4378 19351 4412
rect 19385 4403 19403 4412
rect 19333 4369 19353 4378
rect 19387 4369 19403 4403
rect 19437 4333 19471 4453
rect 19505 4408 19575 4419
rect 19505 4403 19524 4408
rect 19505 4369 19521 4403
rect 19558 4374 19575 4408
rect 19555 4369 19575 4374
rect 18008 4282 18042 4301
rect 18263 4317 18311 4333
rect 18263 4283 18277 4317
rect 18263 4249 18311 4283
rect 17848 4205 17864 4239
rect 17898 4205 17914 4239
rect 18263 4215 18277 4249
rect 18263 4171 18311 4215
rect 18345 4317 18411 4333
rect 18345 4283 18361 4317
rect 18395 4287 18411 4317
rect 18345 4253 18363 4283
rect 18397 4253 18411 4287
rect 18345 4249 18411 4253
rect 18345 4215 18361 4249
rect 18395 4215 18411 4249
rect 18345 4205 18411 4215
rect 18445 4317 18499 4333
rect 18479 4283 18499 4317
rect 18445 4249 18499 4283
rect 18479 4215 18499 4249
rect 18445 4171 18499 4215
rect 19337 4317 19385 4333
rect 19337 4283 19351 4317
rect 19337 4249 19385 4283
rect 19337 4215 19351 4249
rect 19337 4171 19385 4215
rect 19419 4317 19485 4333
rect 19419 4292 19435 4317
rect 19419 4258 19433 4292
rect 19469 4283 19485 4317
rect 19467 4258 19485 4283
rect 19419 4249 19485 4258
rect 19419 4215 19435 4249
rect 19469 4215 19485 4249
rect 19419 4205 19485 4215
rect 19519 4317 19573 4333
rect 19553 4283 19573 4317
rect 19519 4249 19573 4283
rect 19553 4215 19573 4249
rect 19519 4171 19573 4215
rect 17960 4124 17976 4158
rect 18010 4124 18026 4158
rect 18242 4137 18271 4171
rect 18305 4137 18363 4171
rect 18397 4137 18455 4171
rect 18489 4137 18518 4171
rect 19316 4137 19345 4171
rect 19379 4137 19437 4171
rect 19471 4137 19529 4171
rect 19563 4137 19592 4171
rect 17832 4074 17866 4090
rect 17832 4004 17866 4038
rect 17832 3952 17866 3968
rect 17928 4074 17962 4090
rect 17928 4004 17962 4038
rect 17928 3952 17962 3968
rect 18024 4074 18058 4090
rect 18024 4004 18058 4038
rect 18058 3968 18406 3992
rect 18024 3952 18406 3968
rect 17744 3884 17880 3918
rect 17914 3884 17930 3918
rect 17659 3814 18054 3834
rect 17659 3809 17921 3814
rect 17659 3800 17800 3809
rect 17784 3775 17800 3800
rect 17834 3780 17921 3809
rect 17955 3790 18054 3814
rect 18226 3792 18272 3794
rect 18226 3790 18230 3792
rect 17955 3780 18230 3790
rect 17834 3775 18230 3780
rect 17784 3758 18230 3775
rect 18264 3758 18272 3792
rect 17784 3756 18272 3758
rect 18226 3750 18272 3756
rect 16558 3635 16587 3669
rect 16621 3635 16679 3669
rect 16713 3635 16771 3669
rect 16805 3635 16834 3669
rect 16154 3583 16390 3594
rect 15796 3575 16390 3583
rect 15796 3550 15798 3575
rect 15710 3507 15744 3509
rect 15710 3471 15744 3473
rect 15710 3386 15744 3405
rect 15832 3550 16356 3575
rect 16442 3575 16518 3594
rect 16442 3554 16444 3575
rect 15798 3507 15832 3509
rect 16054 3477 16070 3511
rect 16104 3477 16120 3511
rect 16356 3507 16390 3509
rect 15798 3471 15832 3473
rect 16356 3471 16390 3473
rect 15798 3386 15832 3405
rect 15926 3415 15960 3434
rect 15926 3347 15960 3349
rect 15738 3309 15754 3343
rect 15788 3309 15804 3343
rect 15926 3311 15960 3313
rect 15426 3231 15438 3265
rect 15426 3197 15472 3231
rect 15426 3163 15438 3197
rect 15016 3089 15045 3123
rect 15079 3089 15137 3123
rect 15171 3089 15229 3123
rect 15263 3089 15292 3123
rect 15426 3117 15472 3163
rect 15506 3265 15572 3277
rect 15506 3231 15522 3265
rect 15556 3231 15572 3265
rect 15506 3218 15572 3231
rect 15926 3226 15960 3245
rect 16022 3415 16056 3434
rect 16022 3347 16056 3349
rect 16022 3311 16056 3313
rect 16022 3226 16056 3245
rect 16118 3415 16152 3434
rect 16356 3386 16390 3405
rect 16478 3554 16518 3575
rect 16626 3593 16668 3635
rect 16904 3633 16933 3667
rect 16967 3633 17025 3667
rect 17059 3633 17117 3667
rect 17151 3633 17180 3667
rect 17325 3661 17359 3668
rect 16626 3559 16634 3593
rect 16444 3507 16478 3509
rect 16444 3471 16478 3473
rect 16626 3525 16668 3559
rect 16626 3491 16634 3525
rect 16626 3457 16668 3491
rect 16626 3423 16634 3457
rect 16626 3407 16668 3423
rect 16702 3593 16768 3601
rect 16702 3559 16718 3593
rect 16752 3559 16768 3593
rect 16702 3525 16768 3559
rect 16702 3491 16718 3525
rect 16752 3491 16768 3525
rect 16702 3457 16768 3491
rect 16702 3423 16718 3457
rect 16752 3423 16768 3457
rect 16702 3405 16768 3423
rect 16937 3583 16973 3599
rect 16937 3549 16939 3583
rect 16937 3515 16973 3549
rect 16937 3481 16939 3515
rect 17009 3583 17075 3633
rect 17250 3627 17279 3661
rect 17313 3627 17371 3661
rect 17405 3627 17463 3661
rect 17497 3627 17526 3661
rect 17626 3637 17642 3671
rect 17676 3637 17692 3671
rect 17850 3658 17964 3660
rect 17009 3549 17025 3583
rect 17059 3549 17075 3583
rect 17009 3515 17075 3549
rect 17009 3481 17025 3515
rect 17059 3481 17075 3515
rect 17109 3583 17163 3599
rect 17109 3549 17111 3583
rect 17145 3549 17163 3583
rect 17109 3502 17163 3549
rect 16937 3447 16973 3481
rect 17109 3468 17111 3502
rect 17145 3468 17163 3502
rect 16937 3413 17072 3447
rect 17109 3418 17163 3468
rect 16444 3386 16478 3405
rect 16118 3347 16152 3349
rect 16530 3371 16674 3372
rect 16530 3357 16688 3371
rect 16118 3311 16152 3313
rect 16384 3344 16450 3346
rect 16530 3344 16638 3357
rect 16384 3343 16638 3344
rect 16384 3309 16400 3343
rect 16434 3330 16638 3343
rect 16434 3310 16570 3330
rect 16622 3323 16638 3330
rect 16672 3323 16688 3357
rect 16434 3309 16450 3310
rect 16622 3273 16668 3289
rect 16722 3285 16768 3405
rect 17038 3384 17072 3413
rect 16925 3355 16993 3377
rect 16925 3354 16941 3355
rect 16925 3320 16939 3354
rect 16975 3321 16993 3355
rect 16973 3320 16993 3321
rect 16925 3303 16993 3320
rect 17038 3368 17093 3384
rect 17038 3334 17059 3368
rect 17038 3318 17093 3334
rect 17127 3368 17163 3418
rect 17318 3585 17360 3627
rect 17850 3619 18132 3658
rect 18272 3637 18288 3671
rect 18322 3637 18338 3671
rect 17850 3594 17889 3619
rect 17318 3551 17326 3585
rect 17318 3517 17360 3551
rect 17318 3483 17326 3517
rect 17318 3449 17360 3483
rect 17318 3415 17326 3449
rect 17318 3399 17360 3415
rect 17394 3585 17460 3593
rect 17394 3551 17410 3585
rect 17444 3551 17460 3585
rect 17394 3517 17460 3551
rect 17394 3483 17410 3517
rect 17444 3483 17460 3517
rect 17394 3449 17460 3483
rect 17394 3415 17410 3449
rect 17444 3415 17460 3449
rect 17394 3397 17460 3415
rect 17127 3366 17168 3368
rect 17127 3332 17132 3366
rect 17166 3332 17168 3366
rect 17127 3330 17168 3332
rect 17314 3360 17380 3363
rect 16152 3245 16398 3262
rect 16118 3228 16398 3245
rect 16118 3226 16152 3228
rect 15506 3197 15848 3218
rect 15506 3163 15522 3197
rect 15556 3186 15848 3197
rect 15556 3183 16024 3186
rect 15556 3182 15974 3183
rect 15556 3163 15578 3182
rect 15506 3158 15578 3163
rect 15506 3151 15572 3158
rect 15812 3150 15974 3182
rect 15958 3149 15974 3150
rect 16008 3149 16024 3183
rect 16350 3140 16398 3228
rect 15362 3083 15391 3117
rect 15425 3083 15483 3117
rect 15517 3083 15575 3117
rect 15609 3083 15638 3117
rect 15720 3112 15766 3122
rect 15720 3078 15726 3112
rect 15760 3092 15766 3112
rect 16350 3106 16358 3140
rect 16392 3106 16398 3140
rect 16622 3239 16634 3273
rect 16622 3205 16668 3239
rect 16622 3171 16634 3205
rect 16622 3125 16668 3171
rect 16702 3273 16768 3285
rect 16702 3222 16718 3273
rect 16752 3222 16768 3273
rect 17038 3267 17072 3318
rect 16702 3205 16768 3222
rect 16702 3171 16718 3205
rect 16752 3171 16768 3205
rect 16702 3159 16768 3171
rect 16939 3233 17072 3267
rect 17127 3258 17163 3330
rect 17314 3326 17328 3360
rect 17362 3349 17380 3360
rect 17314 3315 17330 3326
rect 17364 3315 17380 3349
rect 16939 3212 16973 3233
rect 17111 3229 17163 3258
rect 16939 3157 16973 3178
rect 17009 3165 17025 3199
rect 17059 3165 17075 3199
rect 15760 3078 15770 3092
rect 12358 2948 12392 2982
rect 12358 2896 12392 2912
rect 13750 2972 13882 3008
rect 14054 3018 14088 3034
rect 14150 3018 14184 3034
rect 14088 2982 14089 2983
rect 13750 2924 13786 2972
rect 14054 2948 14089 2982
rect 14088 2946 14089 2948
rect 14150 2948 14184 2982
rect 13934 2924 14054 2946
rect 13750 2912 14054 2924
rect 14088 2912 14090 2946
rect 13750 2910 14090 2912
rect 13750 2888 13970 2910
rect 14054 2896 14088 2910
rect 14150 2896 14184 2912
rect 14246 3018 14280 3034
rect 15720 3008 15770 3078
rect 16070 3068 16086 3102
rect 16120 3068 16136 3102
rect 16350 3094 16398 3106
rect 16558 3091 16587 3125
rect 16621 3091 16679 3125
rect 16713 3091 16771 3125
rect 16805 3091 16834 3125
rect 17009 3123 17075 3165
rect 17145 3195 17163 3229
rect 17111 3157 17163 3195
rect 17314 3265 17360 3281
rect 17414 3277 17460 3397
rect 17598 3575 17632 3594
rect 17684 3585 17889 3594
rect 17923 3617 18132 3619
rect 17923 3585 18008 3617
rect 17684 3583 18008 3585
rect 18042 3594 18132 3617
rect 18372 3594 18406 3952
rect 19316 3926 19350 4137
rect 19547 3834 19581 4137
rect 19632 3918 19666 4532
rect 19832 4530 19898 4532
rect 20149 4537 20165 4571
rect 20199 4537 20215 4571
rect 20149 4503 20215 4537
rect 19704 4471 19738 4490
rect 19704 4403 19738 4405
rect 19704 4367 19738 4369
rect 19704 4282 19738 4301
rect 19800 4471 19834 4490
rect 19800 4403 19834 4405
rect 19800 4367 19834 4369
rect 19800 4282 19834 4301
rect 19896 4471 19930 4490
rect 20149 4469 20165 4503
rect 20199 4487 20215 4503
rect 20321 4639 20387 4681
rect 20355 4605 20387 4639
rect 20321 4571 20387 4605
rect 20355 4537 20387 4571
rect 20321 4503 20387 4537
rect 20199 4469 20285 4487
rect 20149 4453 20285 4469
rect 20355 4469 20387 4503
rect 20321 4453 20387 4469
rect 21223 4639 21289 4644
rect 21223 4605 21239 4639
rect 21273 4605 21289 4639
rect 21223 4571 21289 4605
rect 21223 4537 21239 4571
rect 21273 4537 21289 4571
rect 21223 4503 21289 4537
rect 21223 4469 21239 4503
rect 21273 4487 21289 4503
rect 21395 4639 21461 4681
rect 21429 4605 21461 4639
rect 21628 4675 21910 4681
rect 21628 4641 21667 4675
rect 21701 4673 21910 4675
rect 21701 4641 21786 4673
rect 21628 4639 21786 4641
rect 21820 4639 21910 4673
rect 21628 4606 21910 4639
rect 22037 4639 22103 4644
rect 21395 4571 21461 4605
rect 21429 4537 21461 4571
rect 22037 4605 22053 4639
rect 22087 4605 22103 4639
rect 22037 4571 22103 4605
rect 21395 4503 21461 4537
rect 21273 4469 21359 4487
rect 21223 4453 21359 4469
rect 21429 4469 21461 4503
rect 21395 4453 21461 4469
rect 21520 4567 21786 4568
rect 21520 4533 21736 4567
rect 21770 4533 21786 4567
rect 21520 4532 21786 4533
rect 19896 4403 19930 4405
rect 20147 4410 20217 4419
rect 20147 4376 20163 4410
rect 20197 4403 20217 4410
rect 20147 4369 20167 4376
rect 20201 4369 20217 4403
rect 19896 4367 19930 4369
rect 20251 4333 20285 4453
rect 20319 4410 20389 4419
rect 20319 4403 20337 4410
rect 20319 4369 20335 4403
rect 20371 4376 20389 4410
rect 20369 4369 20389 4376
rect 21221 4412 21291 4419
rect 21221 4378 21239 4412
rect 21273 4403 21291 4412
rect 21221 4369 21241 4378
rect 21275 4369 21291 4403
rect 21325 4333 21359 4453
rect 21393 4408 21463 4419
rect 21393 4403 21412 4408
rect 21393 4369 21409 4403
rect 21446 4374 21463 4408
rect 21443 4369 21463 4374
rect 19896 4282 19930 4301
rect 20151 4317 20199 4333
rect 20151 4283 20165 4317
rect 20151 4249 20199 4283
rect 19736 4205 19752 4239
rect 19786 4205 19802 4239
rect 20151 4215 20165 4249
rect 20151 4171 20199 4215
rect 20233 4317 20299 4333
rect 20233 4283 20249 4317
rect 20283 4287 20299 4317
rect 20233 4253 20251 4283
rect 20285 4253 20299 4287
rect 20233 4249 20299 4253
rect 20233 4215 20249 4249
rect 20283 4215 20299 4249
rect 20233 4205 20299 4215
rect 20333 4317 20387 4333
rect 20367 4283 20387 4317
rect 20333 4249 20387 4283
rect 20367 4215 20387 4249
rect 20333 4171 20387 4215
rect 21225 4317 21273 4333
rect 21225 4283 21239 4317
rect 21225 4249 21273 4283
rect 21225 4215 21239 4249
rect 21225 4171 21273 4215
rect 21307 4317 21373 4333
rect 21307 4292 21323 4317
rect 21307 4258 21321 4292
rect 21357 4283 21373 4317
rect 21355 4258 21373 4283
rect 21307 4249 21373 4258
rect 21307 4215 21323 4249
rect 21357 4215 21373 4249
rect 21307 4205 21373 4215
rect 21407 4317 21461 4333
rect 21441 4283 21461 4317
rect 21407 4249 21461 4283
rect 21441 4215 21461 4249
rect 21407 4171 21461 4215
rect 19848 4124 19864 4158
rect 19898 4124 19914 4158
rect 20130 4137 20159 4171
rect 20193 4137 20251 4171
rect 20285 4137 20343 4171
rect 20377 4137 20406 4171
rect 21204 4137 21233 4171
rect 21267 4137 21325 4171
rect 21359 4137 21417 4171
rect 21451 4137 21480 4171
rect 19720 4074 19754 4090
rect 19720 4004 19754 4038
rect 19720 3952 19754 3968
rect 19816 4074 19850 4090
rect 19816 4004 19850 4038
rect 19816 3952 19850 3968
rect 19912 4074 19946 4090
rect 19912 4004 19946 4038
rect 19946 3968 20294 3992
rect 19912 3952 20294 3968
rect 19632 3884 19768 3918
rect 19802 3884 19818 3918
rect 19547 3814 19942 3834
rect 19547 3809 19809 3814
rect 19547 3800 19688 3809
rect 19672 3775 19688 3800
rect 19722 3780 19809 3809
rect 19843 3790 19942 3814
rect 20114 3792 20160 3794
rect 20114 3790 20118 3792
rect 19843 3780 20118 3790
rect 19722 3775 20118 3780
rect 19672 3758 20118 3775
rect 20152 3758 20160 3792
rect 19672 3756 20160 3758
rect 20114 3750 20160 3756
rect 18446 3635 18475 3669
rect 18509 3635 18567 3669
rect 18601 3635 18659 3669
rect 18693 3635 18722 3669
rect 18042 3583 18278 3594
rect 17684 3575 18278 3583
rect 17684 3550 17686 3575
rect 17598 3507 17632 3509
rect 17598 3471 17632 3473
rect 17598 3386 17632 3405
rect 17720 3550 18244 3575
rect 18330 3575 18406 3594
rect 18330 3554 18332 3575
rect 17686 3507 17720 3509
rect 17942 3477 17958 3511
rect 17992 3477 18008 3511
rect 18244 3507 18278 3509
rect 17686 3471 17720 3473
rect 18244 3471 18278 3473
rect 17686 3386 17720 3405
rect 17814 3415 17848 3434
rect 17814 3347 17848 3349
rect 17626 3309 17642 3343
rect 17676 3309 17692 3343
rect 17814 3311 17848 3313
rect 17314 3231 17326 3265
rect 17314 3197 17360 3231
rect 17314 3163 17326 3197
rect 16904 3089 16933 3123
rect 16967 3089 17025 3123
rect 17059 3089 17117 3123
rect 17151 3089 17180 3123
rect 17314 3117 17360 3163
rect 17394 3265 17460 3277
rect 17394 3231 17410 3265
rect 17444 3231 17460 3265
rect 17394 3218 17460 3231
rect 17814 3226 17848 3245
rect 17910 3415 17944 3434
rect 17910 3347 17944 3349
rect 17910 3311 17944 3313
rect 17910 3226 17944 3245
rect 18006 3415 18040 3434
rect 18244 3386 18278 3405
rect 18366 3554 18406 3575
rect 18514 3593 18556 3635
rect 18792 3633 18821 3667
rect 18855 3633 18913 3667
rect 18947 3633 19005 3667
rect 19039 3633 19068 3667
rect 19213 3661 19247 3668
rect 18514 3559 18522 3593
rect 18332 3507 18366 3509
rect 18332 3471 18366 3473
rect 18514 3525 18556 3559
rect 18514 3491 18522 3525
rect 18514 3457 18556 3491
rect 18514 3423 18522 3457
rect 18514 3407 18556 3423
rect 18590 3593 18656 3601
rect 18590 3559 18606 3593
rect 18640 3559 18656 3593
rect 18590 3525 18656 3559
rect 18590 3491 18606 3525
rect 18640 3491 18656 3525
rect 18590 3457 18656 3491
rect 18590 3423 18606 3457
rect 18640 3423 18656 3457
rect 18590 3405 18656 3423
rect 18825 3583 18861 3599
rect 18825 3549 18827 3583
rect 18825 3515 18861 3549
rect 18825 3481 18827 3515
rect 18897 3583 18963 3633
rect 19138 3627 19167 3661
rect 19201 3627 19259 3661
rect 19293 3627 19351 3661
rect 19385 3627 19414 3661
rect 19514 3637 19530 3671
rect 19564 3637 19580 3671
rect 19738 3658 19852 3660
rect 18897 3549 18913 3583
rect 18947 3549 18963 3583
rect 18897 3515 18963 3549
rect 18897 3481 18913 3515
rect 18947 3481 18963 3515
rect 18997 3583 19051 3599
rect 18997 3549 18999 3583
rect 19033 3549 19051 3583
rect 18997 3502 19051 3549
rect 18825 3447 18861 3481
rect 18997 3468 18999 3502
rect 19033 3468 19051 3502
rect 18825 3413 18960 3447
rect 18997 3418 19051 3468
rect 18332 3386 18366 3405
rect 18006 3347 18040 3349
rect 18418 3371 18562 3372
rect 18418 3357 18576 3371
rect 18006 3311 18040 3313
rect 18272 3344 18338 3346
rect 18418 3344 18526 3357
rect 18272 3343 18526 3344
rect 18272 3309 18288 3343
rect 18322 3330 18526 3343
rect 18322 3310 18458 3330
rect 18510 3323 18526 3330
rect 18560 3323 18576 3357
rect 18322 3309 18338 3310
rect 18510 3273 18556 3289
rect 18610 3285 18656 3405
rect 18926 3384 18960 3413
rect 18813 3355 18881 3377
rect 18813 3354 18829 3355
rect 18813 3320 18827 3354
rect 18863 3321 18881 3355
rect 18861 3320 18881 3321
rect 18813 3303 18881 3320
rect 18926 3368 18981 3384
rect 18926 3334 18947 3368
rect 18926 3318 18981 3334
rect 19015 3368 19051 3418
rect 19206 3585 19248 3627
rect 19738 3619 20020 3658
rect 20160 3637 20176 3671
rect 20210 3637 20226 3671
rect 19738 3594 19777 3619
rect 19206 3551 19214 3585
rect 19206 3517 19248 3551
rect 19206 3483 19214 3517
rect 19206 3449 19248 3483
rect 19206 3415 19214 3449
rect 19206 3399 19248 3415
rect 19282 3585 19348 3593
rect 19282 3551 19298 3585
rect 19332 3551 19348 3585
rect 19282 3517 19348 3551
rect 19282 3483 19298 3517
rect 19332 3483 19348 3517
rect 19282 3449 19348 3483
rect 19282 3415 19298 3449
rect 19332 3415 19348 3449
rect 19282 3397 19348 3415
rect 19015 3366 19056 3368
rect 19015 3332 19020 3366
rect 19054 3332 19056 3366
rect 19015 3330 19056 3332
rect 19202 3360 19268 3363
rect 18040 3245 18286 3262
rect 18006 3228 18286 3245
rect 18006 3226 18040 3228
rect 17394 3197 17736 3218
rect 17394 3163 17410 3197
rect 17444 3186 17736 3197
rect 17444 3183 17912 3186
rect 17444 3182 17862 3183
rect 17444 3163 17466 3182
rect 17394 3158 17466 3163
rect 17394 3151 17460 3158
rect 17700 3150 17862 3182
rect 17846 3149 17862 3150
rect 17896 3149 17912 3183
rect 18238 3140 18286 3228
rect 17250 3083 17279 3117
rect 17313 3083 17371 3117
rect 17405 3083 17463 3117
rect 17497 3083 17526 3117
rect 17608 3112 17654 3122
rect 17608 3078 17614 3112
rect 17648 3092 17654 3112
rect 18238 3106 18246 3140
rect 18280 3106 18286 3140
rect 18510 3239 18522 3273
rect 18510 3205 18556 3239
rect 18510 3171 18522 3205
rect 18510 3125 18556 3171
rect 18590 3273 18656 3285
rect 18590 3222 18606 3273
rect 18640 3222 18656 3273
rect 18926 3267 18960 3318
rect 18590 3205 18656 3222
rect 18590 3171 18606 3205
rect 18640 3171 18656 3205
rect 18590 3159 18656 3171
rect 18827 3233 18960 3267
rect 19015 3258 19051 3330
rect 19202 3326 19216 3360
rect 19250 3349 19268 3360
rect 19202 3315 19218 3326
rect 19252 3315 19268 3349
rect 18827 3212 18861 3233
rect 18999 3229 19051 3258
rect 18827 3157 18861 3178
rect 18897 3165 18913 3199
rect 18947 3165 18963 3199
rect 17648 3078 17658 3092
rect 14246 2948 14280 2982
rect 14246 2896 14280 2912
rect 15638 2972 15770 3008
rect 15942 3018 15976 3034
rect 16038 3018 16072 3034
rect 15976 2982 15977 2983
rect 15638 2924 15674 2972
rect 15942 2948 15977 2982
rect 15976 2946 15977 2948
rect 16038 2948 16072 2982
rect 15822 2924 15942 2946
rect 15638 2912 15942 2924
rect 15976 2912 15978 2946
rect 15638 2910 15978 2912
rect 15638 2888 15858 2910
rect 15942 2896 15976 2910
rect 16038 2896 16072 2912
rect 16134 3018 16168 3034
rect 17608 3008 17658 3078
rect 17958 3068 17974 3102
rect 18008 3068 18024 3102
rect 18238 3094 18286 3106
rect 18446 3091 18475 3125
rect 18509 3091 18567 3125
rect 18601 3091 18659 3125
rect 18693 3091 18722 3125
rect 18897 3123 18963 3165
rect 19033 3195 19051 3229
rect 18999 3157 19051 3195
rect 19202 3265 19248 3281
rect 19302 3277 19348 3397
rect 19486 3575 19520 3594
rect 19572 3585 19777 3594
rect 19811 3617 20020 3619
rect 19811 3585 19896 3617
rect 19572 3583 19896 3585
rect 19930 3594 20020 3617
rect 20260 3594 20294 3952
rect 21204 3926 21238 4137
rect 21435 3834 21469 4137
rect 21520 3918 21554 4532
rect 21720 4530 21786 4532
rect 22037 4537 22053 4571
rect 22087 4537 22103 4571
rect 22037 4503 22103 4537
rect 21592 4471 21626 4490
rect 21592 4403 21626 4405
rect 21592 4367 21626 4369
rect 21592 4282 21626 4301
rect 21688 4471 21722 4490
rect 21688 4403 21722 4405
rect 21688 4367 21722 4369
rect 21688 4282 21722 4301
rect 21784 4471 21818 4490
rect 22037 4469 22053 4503
rect 22087 4487 22103 4503
rect 22209 4639 22275 4681
rect 22243 4605 22275 4639
rect 22209 4571 22275 4605
rect 22243 4537 22275 4571
rect 22209 4503 22275 4537
rect 22087 4469 22173 4487
rect 22037 4453 22173 4469
rect 22243 4469 22275 4503
rect 22209 4453 22275 4469
rect 23111 4639 23177 4644
rect 23111 4605 23127 4639
rect 23161 4605 23177 4639
rect 23111 4571 23177 4605
rect 23111 4537 23127 4571
rect 23161 4537 23177 4571
rect 23111 4503 23177 4537
rect 23111 4469 23127 4503
rect 23161 4487 23177 4503
rect 23283 4639 23349 4681
rect 23317 4605 23349 4639
rect 23516 4675 23798 4681
rect 23516 4641 23555 4675
rect 23589 4673 23798 4675
rect 23589 4641 23674 4673
rect 23516 4639 23674 4641
rect 23708 4639 23798 4673
rect 23516 4606 23798 4639
rect 23925 4639 23991 4644
rect 23283 4571 23349 4605
rect 23317 4537 23349 4571
rect 23925 4605 23941 4639
rect 23975 4605 23991 4639
rect 23925 4571 23991 4605
rect 23283 4503 23349 4537
rect 23161 4469 23247 4487
rect 23111 4453 23247 4469
rect 23317 4469 23349 4503
rect 23283 4453 23349 4469
rect 23408 4567 23674 4568
rect 23408 4533 23624 4567
rect 23658 4533 23674 4567
rect 23408 4532 23674 4533
rect 21784 4403 21818 4405
rect 22035 4410 22105 4419
rect 22035 4376 22051 4410
rect 22085 4403 22105 4410
rect 22035 4369 22055 4376
rect 22089 4369 22105 4403
rect 21784 4367 21818 4369
rect 22139 4333 22173 4453
rect 22207 4410 22277 4419
rect 22207 4403 22225 4410
rect 22207 4369 22223 4403
rect 22259 4376 22277 4410
rect 22257 4369 22277 4376
rect 23109 4412 23179 4419
rect 23109 4378 23127 4412
rect 23161 4403 23179 4412
rect 23109 4369 23129 4378
rect 23163 4369 23179 4403
rect 23213 4333 23247 4453
rect 23281 4408 23351 4419
rect 23281 4403 23300 4408
rect 23281 4369 23297 4403
rect 23334 4374 23351 4408
rect 23331 4369 23351 4374
rect 21784 4282 21818 4301
rect 22039 4317 22087 4333
rect 22039 4283 22053 4317
rect 22039 4249 22087 4283
rect 21624 4205 21640 4239
rect 21674 4205 21690 4239
rect 22039 4215 22053 4249
rect 22039 4171 22087 4215
rect 22121 4317 22187 4333
rect 22121 4283 22137 4317
rect 22171 4287 22187 4317
rect 22121 4253 22139 4283
rect 22173 4253 22187 4287
rect 22121 4249 22187 4253
rect 22121 4215 22137 4249
rect 22171 4215 22187 4249
rect 22121 4205 22187 4215
rect 22221 4317 22275 4333
rect 22255 4283 22275 4317
rect 22221 4249 22275 4283
rect 22255 4215 22275 4249
rect 22221 4171 22275 4215
rect 23113 4317 23161 4333
rect 23113 4283 23127 4317
rect 23113 4249 23161 4283
rect 23113 4215 23127 4249
rect 23113 4171 23161 4215
rect 23195 4317 23261 4333
rect 23195 4292 23211 4317
rect 23195 4258 23209 4292
rect 23245 4283 23261 4317
rect 23243 4258 23261 4283
rect 23195 4249 23261 4258
rect 23195 4215 23211 4249
rect 23245 4215 23261 4249
rect 23195 4205 23261 4215
rect 23295 4317 23349 4333
rect 23329 4283 23349 4317
rect 23295 4249 23349 4283
rect 23329 4215 23349 4249
rect 23295 4171 23349 4215
rect 21736 4124 21752 4158
rect 21786 4124 21802 4158
rect 22018 4137 22047 4171
rect 22081 4137 22139 4171
rect 22173 4137 22231 4171
rect 22265 4137 22294 4171
rect 23092 4137 23121 4171
rect 23155 4137 23213 4171
rect 23247 4137 23305 4171
rect 23339 4137 23368 4171
rect 21608 4074 21642 4090
rect 21608 4004 21642 4038
rect 21608 3952 21642 3968
rect 21704 4074 21738 4090
rect 21704 4004 21738 4038
rect 21704 3952 21738 3968
rect 21800 4074 21834 4090
rect 21800 4004 21834 4038
rect 21834 3968 22182 3992
rect 21800 3952 22182 3968
rect 21520 3884 21656 3918
rect 21690 3884 21706 3918
rect 21435 3814 21830 3834
rect 21435 3809 21697 3814
rect 21435 3800 21576 3809
rect 21560 3775 21576 3800
rect 21610 3780 21697 3809
rect 21731 3790 21830 3814
rect 22002 3792 22048 3794
rect 22002 3790 22006 3792
rect 21731 3780 22006 3790
rect 21610 3775 22006 3780
rect 21560 3758 22006 3775
rect 22040 3758 22048 3792
rect 21560 3756 22048 3758
rect 22002 3750 22048 3756
rect 20334 3635 20363 3669
rect 20397 3635 20455 3669
rect 20489 3635 20547 3669
rect 20581 3635 20610 3669
rect 19930 3583 20166 3594
rect 19572 3575 20166 3583
rect 19572 3550 19574 3575
rect 19486 3507 19520 3509
rect 19486 3471 19520 3473
rect 19486 3386 19520 3405
rect 19608 3550 20132 3575
rect 20218 3575 20294 3594
rect 20218 3554 20220 3575
rect 19574 3507 19608 3509
rect 19830 3477 19846 3511
rect 19880 3477 19896 3511
rect 20132 3507 20166 3509
rect 19574 3471 19608 3473
rect 20132 3471 20166 3473
rect 19574 3386 19608 3405
rect 19702 3415 19736 3434
rect 19702 3347 19736 3349
rect 19514 3309 19530 3343
rect 19564 3309 19580 3343
rect 19702 3311 19736 3313
rect 19202 3231 19214 3265
rect 19202 3197 19248 3231
rect 19202 3163 19214 3197
rect 18792 3089 18821 3123
rect 18855 3089 18913 3123
rect 18947 3089 19005 3123
rect 19039 3089 19068 3123
rect 19202 3117 19248 3163
rect 19282 3265 19348 3277
rect 19282 3231 19298 3265
rect 19332 3231 19348 3265
rect 19282 3218 19348 3231
rect 19702 3226 19736 3245
rect 19798 3415 19832 3434
rect 19798 3347 19832 3349
rect 19798 3311 19832 3313
rect 19798 3226 19832 3245
rect 19894 3415 19928 3434
rect 20132 3386 20166 3405
rect 20254 3554 20294 3575
rect 20402 3593 20444 3635
rect 20680 3633 20709 3667
rect 20743 3633 20801 3667
rect 20835 3633 20893 3667
rect 20927 3633 20956 3667
rect 21101 3661 21135 3668
rect 20402 3559 20410 3593
rect 20220 3507 20254 3509
rect 20220 3471 20254 3473
rect 20402 3525 20444 3559
rect 20402 3491 20410 3525
rect 20402 3457 20444 3491
rect 20402 3423 20410 3457
rect 20402 3407 20444 3423
rect 20478 3593 20544 3601
rect 20478 3559 20494 3593
rect 20528 3559 20544 3593
rect 20478 3525 20544 3559
rect 20478 3491 20494 3525
rect 20528 3491 20544 3525
rect 20478 3457 20544 3491
rect 20478 3423 20494 3457
rect 20528 3423 20544 3457
rect 20478 3405 20544 3423
rect 20713 3583 20749 3599
rect 20713 3549 20715 3583
rect 20713 3515 20749 3549
rect 20713 3481 20715 3515
rect 20785 3583 20851 3633
rect 21026 3627 21055 3661
rect 21089 3627 21147 3661
rect 21181 3627 21239 3661
rect 21273 3627 21302 3661
rect 21402 3637 21418 3671
rect 21452 3637 21468 3671
rect 21626 3658 21740 3660
rect 20785 3549 20801 3583
rect 20835 3549 20851 3583
rect 20785 3515 20851 3549
rect 20785 3481 20801 3515
rect 20835 3481 20851 3515
rect 20885 3583 20939 3599
rect 20885 3549 20887 3583
rect 20921 3549 20939 3583
rect 20885 3502 20939 3549
rect 20713 3447 20749 3481
rect 20885 3468 20887 3502
rect 20921 3468 20939 3502
rect 20713 3413 20848 3447
rect 20885 3418 20939 3468
rect 20220 3386 20254 3405
rect 19894 3347 19928 3349
rect 20306 3371 20450 3372
rect 20306 3357 20464 3371
rect 19894 3311 19928 3313
rect 20160 3344 20226 3346
rect 20306 3344 20414 3357
rect 20160 3343 20414 3344
rect 20160 3309 20176 3343
rect 20210 3330 20414 3343
rect 20210 3310 20346 3330
rect 20398 3323 20414 3330
rect 20448 3323 20464 3357
rect 20210 3309 20226 3310
rect 20398 3273 20444 3289
rect 20498 3285 20544 3405
rect 20814 3384 20848 3413
rect 20701 3355 20769 3377
rect 20701 3354 20717 3355
rect 20701 3320 20715 3354
rect 20751 3321 20769 3355
rect 20749 3320 20769 3321
rect 20701 3303 20769 3320
rect 20814 3368 20869 3384
rect 20814 3334 20835 3368
rect 20814 3318 20869 3334
rect 20903 3368 20939 3418
rect 21094 3585 21136 3627
rect 21626 3619 21908 3658
rect 22048 3637 22064 3671
rect 22098 3637 22114 3671
rect 21626 3594 21665 3619
rect 21094 3551 21102 3585
rect 21094 3517 21136 3551
rect 21094 3483 21102 3517
rect 21094 3449 21136 3483
rect 21094 3415 21102 3449
rect 21094 3399 21136 3415
rect 21170 3585 21236 3593
rect 21170 3551 21186 3585
rect 21220 3551 21236 3585
rect 21170 3517 21236 3551
rect 21170 3483 21186 3517
rect 21220 3483 21236 3517
rect 21170 3449 21236 3483
rect 21170 3415 21186 3449
rect 21220 3415 21236 3449
rect 21170 3397 21236 3415
rect 20903 3366 20944 3368
rect 20903 3332 20908 3366
rect 20942 3332 20944 3366
rect 20903 3330 20944 3332
rect 21090 3360 21156 3363
rect 19928 3245 20174 3262
rect 19894 3228 20174 3245
rect 19894 3226 19928 3228
rect 19282 3197 19624 3218
rect 19282 3163 19298 3197
rect 19332 3186 19624 3197
rect 19332 3183 19800 3186
rect 19332 3182 19750 3183
rect 19332 3163 19354 3182
rect 19282 3158 19354 3163
rect 19282 3151 19348 3158
rect 19588 3150 19750 3182
rect 19734 3149 19750 3150
rect 19784 3149 19800 3183
rect 20126 3140 20174 3228
rect 19138 3083 19167 3117
rect 19201 3083 19259 3117
rect 19293 3083 19351 3117
rect 19385 3083 19414 3117
rect 19496 3112 19542 3122
rect 19496 3078 19502 3112
rect 19536 3092 19542 3112
rect 20126 3106 20134 3140
rect 20168 3106 20174 3140
rect 20398 3239 20410 3273
rect 20398 3205 20444 3239
rect 20398 3171 20410 3205
rect 20398 3125 20444 3171
rect 20478 3273 20544 3285
rect 20478 3222 20494 3273
rect 20528 3222 20544 3273
rect 20814 3267 20848 3318
rect 20478 3205 20544 3222
rect 20478 3171 20494 3205
rect 20528 3171 20544 3205
rect 20478 3159 20544 3171
rect 20715 3233 20848 3267
rect 20903 3258 20939 3330
rect 21090 3326 21104 3360
rect 21138 3349 21156 3360
rect 21090 3315 21106 3326
rect 21140 3315 21156 3349
rect 20715 3212 20749 3233
rect 20887 3229 20939 3258
rect 20715 3157 20749 3178
rect 20785 3165 20801 3199
rect 20835 3165 20851 3199
rect 19536 3078 19546 3092
rect 16134 2948 16168 2982
rect 16134 2896 16168 2912
rect 17526 2972 17658 3008
rect 17830 3018 17864 3034
rect 17926 3018 17960 3034
rect 17864 2982 17865 2983
rect 17526 2924 17562 2972
rect 17830 2948 17865 2982
rect 17864 2946 17865 2948
rect 17926 2948 17960 2982
rect 17710 2924 17830 2946
rect 17526 2912 17830 2924
rect 17864 2912 17866 2946
rect 17526 2910 17866 2912
rect 17526 2888 17746 2910
rect 17830 2896 17864 2910
rect 17926 2896 17960 2912
rect 18022 3018 18056 3034
rect 19496 3008 19546 3078
rect 19846 3068 19862 3102
rect 19896 3068 19912 3102
rect 20126 3094 20174 3106
rect 20334 3091 20363 3125
rect 20397 3091 20455 3125
rect 20489 3091 20547 3125
rect 20581 3091 20610 3125
rect 20785 3123 20851 3165
rect 20921 3195 20939 3229
rect 20887 3157 20939 3195
rect 21090 3265 21136 3281
rect 21190 3277 21236 3397
rect 21374 3575 21408 3594
rect 21460 3585 21665 3594
rect 21699 3617 21908 3619
rect 21699 3585 21784 3617
rect 21460 3583 21784 3585
rect 21818 3594 21908 3617
rect 22148 3594 22182 3952
rect 23092 3926 23126 4137
rect 23323 3834 23357 4137
rect 23408 3918 23442 4532
rect 23608 4530 23674 4532
rect 23925 4537 23941 4571
rect 23975 4537 23991 4571
rect 23925 4503 23991 4537
rect 23480 4471 23514 4490
rect 23480 4403 23514 4405
rect 23480 4367 23514 4369
rect 23480 4282 23514 4301
rect 23576 4471 23610 4490
rect 23576 4403 23610 4405
rect 23576 4367 23610 4369
rect 23576 4282 23610 4301
rect 23672 4471 23706 4490
rect 23925 4469 23941 4503
rect 23975 4487 23991 4503
rect 24097 4639 24163 4681
rect 24131 4605 24163 4639
rect 24097 4571 24163 4605
rect 24131 4537 24163 4571
rect 24097 4503 24163 4537
rect 23975 4469 24061 4487
rect 23925 4453 24061 4469
rect 24131 4469 24163 4503
rect 24097 4453 24163 4469
rect 24999 4639 25065 4644
rect 24999 4605 25015 4639
rect 25049 4605 25065 4639
rect 24999 4571 25065 4605
rect 24999 4537 25015 4571
rect 25049 4537 25065 4571
rect 24999 4503 25065 4537
rect 24999 4469 25015 4503
rect 25049 4487 25065 4503
rect 25171 4639 25237 4681
rect 25205 4605 25237 4639
rect 25404 4675 25686 4681
rect 25404 4641 25443 4675
rect 25477 4673 25686 4675
rect 25477 4641 25562 4673
rect 25404 4639 25562 4641
rect 25596 4639 25686 4673
rect 25404 4606 25686 4639
rect 25813 4639 25879 4644
rect 25171 4571 25237 4605
rect 25205 4537 25237 4571
rect 25813 4605 25829 4639
rect 25863 4605 25879 4639
rect 25813 4571 25879 4605
rect 25171 4503 25237 4537
rect 25049 4469 25135 4487
rect 24999 4453 25135 4469
rect 25205 4469 25237 4503
rect 25171 4453 25237 4469
rect 25296 4567 25562 4568
rect 25296 4533 25512 4567
rect 25546 4533 25562 4567
rect 25296 4532 25562 4533
rect 23672 4403 23706 4405
rect 23923 4410 23993 4419
rect 23923 4376 23939 4410
rect 23973 4403 23993 4410
rect 23923 4369 23943 4376
rect 23977 4369 23993 4403
rect 23672 4367 23706 4369
rect 24027 4333 24061 4453
rect 24095 4410 24165 4419
rect 24095 4403 24113 4410
rect 24095 4369 24111 4403
rect 24147 4376 24165 4410
rect 24145 4369 24165 4376
rect 24997 4412 25067 4419
rect 24997 4378 25015 4412
rect 25049 4403 25067 4412
rect 24997 4369 25017 4378
rect 25051 4369 25067 4403
rect 25101 4333 25135 4453
rect 25169 4408 25239 4419
rect 25169 4403 25188 4408
rect 25169 4369 25185 4403
rect 25222 4374 25239 4408
rect 25219 4369 25239 4374
rect 23672 4282 23706 4301
rect 23927 4317 23975 4333
rect 23927 4283 23941 4317
rect 23927 4249 23975 4283
rect 23512 4205 23528 4239
rect 23562 4205 23578 4239
rect 23927 4215 23941 4249
rect 23927 4171 23975 4215
rect 24009 4317 24075 4333
rect 24009 4283 24025 4317
rect 24059 4287 24075 4317
rect 24009 4253 24027 4283
rect 24061 4253 24075 4287
rect 24009 4249 24075 4253
rect 24009 4215 24025 4249
rect 24059 4215 24075 4249
rect 24009 4205 24075 4215
rect 24109 4317 24163 4333
rect 24143 4283 24163 4317
rect 24109 4249 24163 4283
rect 24143 4215 24163 4249
rect 24109 4171 24163 4215
rect 25001 4317 25049 4333
rect 25001 4283 25015 4317
rect 25001 4249 25049 4283
rect 25001 4215 25015 4249
rect 25001 4171 25049 4215
rect 25083 4317 25149 4333
rect 25083 4292 25099 4317
rect 25083 4258 25097 4292
rect 25133 4283 25149 4317
rect 25131 4258 25149 4283
rect 25083 4249 25149 4258
rect 25083 4215 25099 4249
rect 25133 4215 25149 4249
rect 25083 4205 25149 4215
rect 25183 4317 25237 4333
rect 25217 4283 25237 4317
rect 25183 4249 25237 4283
rect 25217 4215 25237 4249
rect 25183 4171 25237 4215
rect 23624 4124 23640 4158
rect 23674 4124 23690 4158
rect 23906 4137 23935 4171
rect 23969 4137 24027 4171
rect 24061 4137 24119 4171
rect 24153 4137 24182 4171
rect 24980 4137 25009 4171
rect 25043 4137 25101 4171
rect 25135 4137 25193 4171
rect 25227 4137 25256 4171
rect 23496 4074 23530 4090
rect 23496 4004 23530 4038
rect 23496 3952 23530 3968
rect 23592 4074 23626 4090
rect 23592 4004 23626 4038
rect 23592 3952 23626 3968
rect 23688 4074 23722 4090
rect 23688 4004 23722 4038
rect 23722 3968 24070 3992
rect 23688 3952 24070 3968
rect 23408 3884 23544 3918
rect 23578 3884 23594 3918
rect 23323 3814 23718 3834
rect 23323 3809 23585 3814
rect 23323 3800 23464 3809
rect 23448 3775 23464 3800
rect 23498 3780 23585 3809
rect 23619 3790 23718 3814
rect 23890 3792 23936 3794
rect 23890 3790 23894 3792
rect 23619 3780 23894 3790
rect 23498 3775 23894 3780
rect 23448 3758 23894 3775
rect 23928 3758 23936 3792
rect 23448 3756 23936 3758
rect 23890 3750 23936 3756
rect 22222 3635 22251 3669
rect 22285 3635 22343 3669
rect 22377 3635 22435 3669
rect 22469 3635 22498 3669
rect 21818 3583 22054 3594
rect 21460 3575 22054 3583
rect 21460 3550 21462 3575
rect 21374 3507 21408 3509
rect 21374 3471 21408 3473
rect 21374 3386 21408 3405
rect 21496 3550 22020 3575
rect 22106 3575 22182 3594
rect 22106 3554 22108 3575
rect 21462 3507 21496 3509
rect 21718 3477 21734 3511
rect 21768 3477 21784 3511
rect 22020 3507 22054 3509
rect 21462 3471 21496 3473
rect 22020 3471 22054 3473
rect 21462 3386 21496 3405
rect 21590 3415 21624 3434
rect 21590 3347 21624 3349
rect 21402 3309 21418 3343
rect 21452 3309 21468 3343
rect 21590 3311 21624 3313
rect 21090 3231 21102 3265
rect 21090 3197 21136 3231
rect 21090 3163 21102 3197
rect 20680 3089 20709 3123
rect 20743 3089 20801 3123
rect 20835 3089 20893 3123
rect 20927 3089 20956 3123
rect 21090 3117 21136 3163
rect 21170 3265 21236 3277
rect 21170 3231 21186 3265
rect 21220 3231 21236 3265
rect 21170 3218 21236 3231
rect 21590 3226 21624 3245
rect 21686 3415 21720 3434
rect 21686 3347 21720 3349
rect 21686 3311 21720 3313
rect 21686 3226 21720 3245
rect 21782 3415 21816 3434
rect 22020 3386 22054 3405
rect 22142 3554 22182 3575
rect 22290 3593 22332 3635
rect 22568 3633 22597 3667
rect 22631 3633 22689 3667
rect 22723 3633 22781 3667
rect 22815 3633 22844 3667
rect 22989 3661 23023 3668
rect 22290 3559 22298 3593
rect 22108 3507 22142 3509
rect 22108 3471 22142 3473
rect 22290 3525 22332 3559
rect 22290 3491 22298 3525
rect 22290 3457 22332 3491
rect 22290 3423 22298 3457
rect 22290 3407 22332 3423
rect 22366 3593 22432 3601
rect 22366 3559 22382 3593
rect 22416 3559 22432 3593
rect 22366 3525 22432 3559
rect 22366 3491 22382 3525
rect 22416 3491 22432 3525
rect 22366 3457 22432 3491
rect 22366 3423 22382 3457
rect 22416 3423 22432 3457
rect 22366 3405 22432 3423
rect 22601 3583 22637 3599
rect 22601 3549 22603 3583
rect 22601 3515 22637 3549
rect 22601 3481 22603 3515
rect 22673 3583 22739 3633
rect 22914 3627 22943 3661
rect 22977 3627 23035 3661
rect 23069 3627 23127 3661
rect 23161 3627 23190 3661
rect 23290 3637 23306 3671
rect 23340 3637 23356 3671
rect 23514 3658 23628 3660
rect 22673 3549 22689 3583
rect 22723 3549 22739 3583
rect 22673 3515 22739 3549
rect 22673 3481 22689 3515
rect 22723 3481 22739 3515
rect 22773 3583 22827 3599
rect 22773 3549 22775 3583
rect 22809 3549 22827 3583
rect 22773 3502 22827 3549
rect 22601 3447 22637 3481
rect 22773 3468 22775 3502
rect 22809 3468 22827 3502
rect 22601 3413 22736 3447
rect 22773 3418 22827 3468
rect 22108 3386 22142 3405
rect 21782 3347 21816 3349
rect 22194 3371 22338 3372
rect 22194 3357 22352 3371
rect 21782 3311 21816 3313
rect 22048 3344 22114 3346
rect 22194 3344 22302 3357
rect 22048 3343 22302 3344
rect 22048 3309 22064 3343
rect 22098 3330 22302 3343
rect 22098 3310 22234 3330
rect 22286 3323 22302 3330
rect 22336 3323 22352 3357
rect 22098 3309 22114 3310
rect 22286 3273 22332 3289
rect 22386 3285 22432 3405
rect 22702 3384 22736 3413
rect 22589 3355 22657 3377
rect 22589 3354 22605 3355
rect 22589 3320 22603 3354
rect 22639 3321 22657 3355
rect 22637 3320 22657 3321
rect 22589 3303 22657 3320
rect 22702 3368 22757 3384
rect 22702 3334 22723 3368
rect 22702 3318 22757 3334
rect 22791 3368 22827 3418
rect 22982 3585 23024 3627
rect 23514 3619 23796 3658
rect 23936 3637 23952 3671
rect 23986 3637 24002 3671
rect 23514 3594 23553 3619
rect 22982 3551 22990 3585
rect 22982 3517 23024 3551
rect 22982 3483 22990 3517
rect 22982 3449 23024 3483
rect 22982 3415 22990 3449
rect 22982 3399 23024 3415
rect 23058 3585 23124 3593
rect 23058 3551 23074 3585
rect 23108 3551 23124 3585
rect 23058 3517 23124 3551
rect 23058 3483 23074 3517
rect 23108 3483 23124 3517
rect 23058 3449 23124 3483
rect 23058 3415 23074 3449
rect 23108 3415 23124 3449
rect 23058 3397 23124 3415
rect 22791 3366 22832 3368
rect 22791 3332 22796 3366
rect 22830 3332 22832 3366
rect 22791 3330 22832 3332
rect 22978 3360 23044 3363
rect 21816 3245 22062 3262
rect 21782 3228 22062 3245
rect 21782 3226 21816 3228
rect 21170 3197 21512 3218
rect 21170 3163 21186 3197
rect 21220 3186 21512 3197
rect 21220 3183 21688 3186
rect 21220 3182 21638 3183
rect 21220 3163 21242 3182
rect 21170 3158 21242 3163
rect 21170 3151 21236 3158
rect 21476 3150 21638 3182
rect 21622 3149 21638 3150
rect 21672 3149 21688 3183
rect 22014 3140 22062 3228
rect 21026 3083 21055 3117
rect 21089 3083 21147 3117
rect 21181 3083 21239 3117
rect 21273 3083 21302 3117
rect 21384 3112 21430 3122
rect 21384 3078 21390 3112
rect 21424 3092 21430 3112
rect 22014 3106 22022 3140
rect 22056 3106 22062 3140
rect 22286 3239 22298 3273
rect 22286 3205 22332 3239
rect 22286 3171 22298 3205
rect 22286 3125 22332 3171
rect 22366 3273 22432 3285
rect 22366 3222 22382 3273
rect 22416 3222 22432 3273
rect 22702 3267 22736 3318
rect 22366 3205 22432 3222
rect 22366 3171 22382 3205
rect 22416 3171 22432 3205
rect 22366 3159 22432 3171
rect 22603 3233 22736 3267
rect 22791 3258 22827 3330
rect 22978 3326 22992 3360
rect 23026 3349 23044 3360
rect 22978 3315 22994 3326
rect 23028 3315 23044 3349
rect 22603 3212 22637 3233
rect 22775 3229 22827 3258
rect 22603 3157 22637 3178
rect 22673 3165 22689 3199
rect 22723 3165 22739 3199
rect 21424 3078 21434 3092
rect 18022 2948 18056 2982
rect 18022 2896 18056 2912
rect 19414 2972 19546 3008
rect 19718 3018 19752 3034
rect 19814 3018 19848 3034
rect 19752 2982 19753 2983
rect 19414 2924 19450 2972
rect 19718 2948 19753 2982
rect 19752 2946 19753 2948
rect 19814 2948 19848 2982
rect 19598 2924 19718 2946
rect 19414 2912 19718 2924
rect 19752 2912 19754 2946
rect 19414 2910 19754 2912
rect 19414 2888 19634 2910
rect 19718 2896 19752 2910
rect 19814 2896 19848 2912
rect 19910 3018 19944 3034
rect 21384 3008 21434 3078
rect 21734 3068 21750 3102
rect 21784 3068 21800 3102
rect 22014 3094 22062 3106
rect 22222 3091 22251 3125
rect 22285 3091 22343 3125
rect 22377 3091 22435 3125
rect 22469 3091 22498 3125
rect 22673 3123 22739 3165
rect 22809 3195 22827 3229
rect 22775 3157 22827 3195
rect 22978 3265 23024 3281
rect 23078 3277 23124 3397
rect 23262 3575 23296 3594
rect 23348 3585 23553 3594
rect 23587 3617 23796 3619
rect 23587 3585 23672 3617
rect 23348 3583 23672 3585
rect 23706 3594 23796 3617
rect 24036 3594 24070 3952
rect 24980 3926 25014 4137
rect 25211 3834 25245 4137
rect 25296 3918 25330 4532
rect 25496 4530 25562 4532
rect 25813 4537 25829 4571
rect 25863 4537 25879 4571
rect 25813 4503 25879 4537
rect 25368 4471 25402 4490
rect 25368 4403 25402 4405
rect 25368 4367 25402 4369
rect 25368 4282 25402 4301
rect 25464 4471 25498 4490
rect 25464 4403 25498 4405
rect 25464 4367 25498 4369
rect 25464 4282 25498 4301
rect 25560 4471 25594 4490
rect 25813 4469 25829 4503
rect 25863 4487 25879 4503
rect 25985 4639 26051 4681
rect 26019 4605 26051 4639
rect 25985 4571 26051 4605
rect 26019 4537 26051 4571
rect 25985 4503 26051 4537
rect 25863 4469 25949 4487
rect 25813 4453 25949 4469
rect 26019 4469 26051 4503
rect 25985 4453 26051 4469
rect 25560 4403 25594 4405
rect 25811 4410 25881 4419
rect 25811 4376 25827 4410
rect 25861 4403 25881 4410
rect 25811 4369 25831 4376
rect 25865 4369 25881 4403
rect 25560 4367 25594 4369
rect 25915 4333 25949 4453
rect 25983 4410 26053 4419
rect 25983 4403 26001 4410
rect 25983 4369 25999 4403
rect 26035 4376 26053 4410
rect 26033 4369 26053 4376
rect 25560 4282 25594 4301
rect 25815 4317 25863 4333
rect 25815 4283 25829 4317
rect 25815 4249 25863 4283
rect 25400 4205 25416 4239
rect 25450 4205 25466 4239
rect 25815 4215 25829 4249
rect 25815 4171 25863 4215
rect 25897 4317 25963 4333
rect 25897 4283 25913 4317
rect 25947 4287 25963 4317
rect 25897 4253 25915 4283
rect 25949 4253 25963 4287
rect 25897 4249 25963 4253
rect 25897 4215 25913 4249
rect 25947 4215 25963 4249
rect 25897 4205 25963 4215
rect 25997 4317 26051 4333
rect 26031 4283 26051 4317
rect 25997 4249 26051 4283
rect 26031 4215 26051 4249
rect 25997 4171 26051 4215
rect 25512 4124 25528 4158
rect 25562 4124 25578 4158
rect 25794 4137 25823 4171
rect 25857 4137 25915 4171
rect 25949 4137 26007 4171
rect 26041 4137 26070 4171
rect 25384 4074 25418 4090
rect 25384 4004 25418 4038
rect 25384 3952 25418 3968
rect 25480 4074 25514 4090
rect 25480 4004 25514 4038
rect 25480 3952 25514 3968
rect 25576 4074 25610 4090
rect 25576 4004 25610 4038
rect 25610 3968 25958 3992
rect 25576 3952 25958 3968
rect 25296 3884 25432 3918
rect 25466 3884 25482 3918
rect 25211 3814 25606 3834
rect 25211 3809 25473 3814
rect 25211 3800 25352 3809
rect 25336 3775 25352 3800
rect 25386 3780 25473 3809
rect 25507 3790 25606 3814
rect 25778 3792 25824 3794
rect 25778 3790 25782 3792
rect 25507 3780 25782 3790
rect 25386 3775 25782 3780
rect 25336 3758 25782 3775
rect 25816 3758 25824 3792
rect 25336 3756 25824 3758
rect 25778 3750 25824 3756
rect 24110 3635 24139 3669
rect 24173 3635 24231 3669
rect 24265 3635 24323 3669
rect 24357 3635 24386 3669
rect 23706 3583 23942 3594
rect 23348 3575 23942 3583
rect 23348 3550 23350 3575
rect 23262 3507 23296 3509
rect 23262 3471 23296 3473
rect 23262 3386 23296 3405
rect 23384 3550 23908 3575
rect 23994 3575 24070 3594
rect 23994 3554 23996 3575
rect 23350 3507 23384 3509
rect 23606 3477 23622 3511
rect 23656 3477 23672 3511
rect 23908 3507 23942 3509
rect 23350 3471 23384 3473
rect 23908 3471 23942 3473
rect 23350 3386 23384 3405
rect 23478 3415 23512 3434
rect 23478 3347 23512 3349
rect 23290 3309 23306 3343
rect 23340 3309 23356 3343
rect 23478 3311 23512 3313
rect 22978 3231 22990 3265
rect 22978 3197 23024 3231
rect 22978 3163 22990 3197
rect 22568 3089 22597 3123
rect 22631 3089 22689 3123
rect 22723 3089 22781 3123
rect 22815 3089 22844 3123
rect 22978 3117 23024 3163
rect 23058 3265 23124 3277
rect 23058 3231 23074 3265
rect 23108 3231 23124 3265
rect 23058 3218 23124 3231
rect 23478 3226 23512 3245
rect 23574 3415 23608 3434
rect 23574 3347 23608 3349
rect 23574 3311 23608 3313
rect 23574 3226 23608 3245
rect 23670 3415 23704 3434
rect 23908 3386 23942 3405
rect 24030 3554 24070 3575
rect 24178 3593 24220 3635
rect 24456 3633 24485 3667
rect 24519 3633 24577 3667
rect 24611 3633 24669 3667
rect 24703 3633 24732 3667
rect 24877 3661 24911 3668
rect 24178 3559 24186 3593
rect 23996 3507 24030 3509
rect 23996 3471 24030 3473
rect 24178 3525 24220 3559
rect 24178 3491 24186 3525
rect 24178 3457 24220 3491
rect 24178 3423 24186 3457
rect 24178 3407 24220 3423
rect 24254 3593 24320 3601
rect 24254 3559 24270 3593
rect 24304 3559 24320 3593
rect 24254 3525 24320 3559
rect 24254 3491 24270 3525
rect 24304 3491 24320 3525
rect 24254 3457 24320 3491
rect 24254 3423 24270 3457
rect 24304 3423 24320 3457
rect 24254 3405 24320 3423
rect 24489 3583 24525 3599
rect 24489 3549 24491 3583
rect 24489 3515 24525 3549
rect 24489 3481 24491 3515
rect 24561 3583 24627 3633
rect 24802 3627 24831 3661
rect 24865 3627 24923 3661
rect 24957 3627 25015 3661
rect 25049 3627 25078 3661
rect 25178 3637 25194 3671
rect 25228 3637 25244 3671
rect 25402 3658 25516 3660
rect 24561 3549 24577 3583
rect 24611 3549 24627 3583
rect 24561 3515 24627 3549
rect 24561 3481 24577 3515
rect 24611 3481 24627 3515
rect 24661 3583 24715 3599
rect 24661 3549 24663 3583
rect 24697 3549 24715 3583
rect 24661 3502 24715 3549
rect 24489 3447 24525 3481
rect 24661 3468 24663 3502
rect 24697 3468 24715 3502
rect 24489 3413 24624 3447
rect 24661 3418 24715 3468
rect 23996 3386 24030 3405
rect 23670 3347 23704 3349
rect 24082 3371 24226 3372
rect 24082 3357 24240 3371
rect 23670 3311 23704 3313
rect 23936 3344 24002 3346
rect 24082 3344 24190 3357
rect 23936 3343 24190 3344
rect 23936 3309 23952 3343
rect 23986 3330 24190 3343
rect 23986 3310 24122 3330
rect 24174 3323 24190 3330
rect 24224 3323 24240 3357
rect 23986 3309 24002 3310
rect 24174 3273 24220 3289
rect 24274 3285 24320 3405
rect 24590 3384 24624 3413
rect 24477 3355 24545 3377
rect 24477 3354 24493 3355
rect 24477 3320 24491 3354
rect 24527 3321 24545 3355
rect 24525 3320 24545 3321
rect 24477 3303 24545 3320
rect 24590 3368 24645 3384
rect 24590 3334 24611 3368
rect 24590 3318 24645 3334
rect 24679 3368 24715 3418
rect 24870 3585 24912 3627
rect 25402 3619 25684 3658
rect 25824 3637 25840 3671
rect 25874 3637 25890 3671
rect 25402 3594 25441 3619
rect 24870 3551 24878 3585
rect 24870 3517 24912 3551
rect 24870 3483 24878 3517
rect 24870 3449 24912 3483
rect 24870 3415 24878 3449
rect 24870 3399 24912 3415
rect 24946 3585 25012 3593
rect 24946 3551 24962 3585
rect 24996 3551 25012 3585
rect 24946 3517 25012 3551
rect 24946 3483 24962 3517
rect 24996 3483 25012 3517
rect 24946 3449 25012 3483
rect 24946 3415 24962 3449
rect 24996 3415 25012 3449
rect 24946 3397 25012 3415
rect 24679 3366 24720 3368
rect 24679 3332 24684 3366
rect 24718 3332 24720 3366
rect 24679 3330 24720 3332
rect 24866 3360 24932 3363
rect 23704 3245 23950 3262
rect 23670 3228 23950 3245
rect 23670 3226 23704 3228
rect 23058 3197 23400 3218
rect 23058 3163 23074 3197
rect 23108 3186 23400 3197
rect 23108 3183 23576 3186
rect 23108 3182 23526 3183
rect 23108 3163 23130 3182
rect 23058 3158 23130 3163
rect 23058 3151 23124 3158
rect 23364 3150 23526 3182
rect 23510 3149 23526 3150
rect 23560 3149 23576 3183
rect 23902 3140 23950 3228
rect 22914 3083 22943 3117
rect 22977 3083 23035 3117
rect 23069 3083 23127 3117
rect 23161 3083 23190 3117
rect 23272 3112 23318 3122
rect 23272 3078 23278 3112
rect 23312 3092 23318 3112
rect 23902 3106 23910 3140
rect 23944 3106 23950 3140
rect 24174 3239 24186 3273
rect 24174 3205 24220 3239
rect 24174 3171 24186 3205
rect 24174 3125 24220 3171
rect 24254 3273 24320 3285
rect 24254 3222 24270 3273
rect 24304 3222 24320 3273
rect 24590 3267 24624 3318
rect 24254 3205 24320 3222
rect 24254 3171 24270 3205
rect 24304 3171 24320 3205
rect 24254 3159 24320 3171
rect 24491 3233 24624 3267
rect 24679 3258 24715 3330
rect 24866 3326 24880 3360
rect 24914 3349 24932 3360
rect 24866 3315 24882 3326
rect 24916 3315 24932 3349
rect 24491 3212 24525 3233
rect 24663 3229 24715 3258
rect 24491 3157 24525 3178
rect 24561 3165 24577 3199
rect 24611 3165 24627 3199
rect 23312 3078 23322 3092
rect 19910 2948 19944 2982
rect 19910 2896 19944 2912
rect 21302 2972 21434 3008
rect 21606 3018 21640 3034
rect 21702 3018 21736 3034
rect 21640 2982 21641 2983
rect 21302 2924 21338 2972
rect 21606 2948 21641 2982
rect 21640 2946 21641 2948
rect 21702 2948 21736 2982
rect 21486 2924 21606 2946
rect 21302 2912 21606 2924
rect 21640 2912 21642 2946
rect 21302 2910 21642 2912
rect 21302 2888 21522 2910
rect 21606 2896 21640 2910
rect 21702 2896 21736 2912
rect 21798 3018 21832 3034
rect 23272 3008 23322 3078
rect 23622 3068 23638 3102
rect 23672 3068 23688 3102
rect 23902 3094 23950 3106
rect 24110 3091 24139 3125
rect 24173 3091 24231 3125
rect 24265 3091 24323 3125
rect 24357 3091 24386 3125
rect 24561 3123 24627 3165
rect 24697 3195 24715 3229
rect 24663 3157 24715 3195
rect 24866 3265 24912 3281
rect 24966 3277 25012 3397
rect 25150 3575 25184 3594
rect 25236 3585 25441 3594
rect 25475 3617 25684 3619
rect 25475 3585 25560 3617
rect 25236 3583 25560 3585
rect 25594 3594 25684 3617
rect 25924 3594 25958 3952
rect 25998 3635 26027 3669
rect 26061 3635 26119 3669
rect 26153 3635 26211 3669
rect 26245 3635 26274 3669
rect 25594 3583 25830 3594
rect 25236 3575 25830 3583
rect 25236 3550 25238 3575
rect 25150 3507 25184 3509
rect 25150 3471 25184 3473
rect 25150 3386 25184 3405
rect 25272 3550 25796 3575
rect 25882 3575 25958 3594
rect 25882 3554 25884 3575
rect 25238 3507 25272 3509
rect 25494 3477 25510 3511
rect 25544 3477 25560 3511
rect 25796 3507 25830 3509
rect 25238 3471 25272 3473
rect 25796 3471 25830 3473
rect 25238 3386 25272 3405
rect 25366 3415 25400 3434
rect 25366 3347 25400 3349
rect 25178 3309 25194 3343
rect 25228 3309 25244 3343
rect 25366 3311 25400 3313
rect 24866 3231 24878 3265
rect 24866 3197 24912 3231
rect 24866 3163 24878 3197
rect 24456 3089 24485 3123
rect 24519 3089 24577 3123
rect 24611 3089 24669 3123
rect 24703 3089 24732 3123
rect 24866 3117 24912 3163
rect 24946 3265 25012 3277
rect 24946 3231 24962 3265
rect 24996 3231 25012 3265
rect 24946 3218 25012 3231
rect 25366 3226 25400 3245
rect 25462 3415 25496 3434
rect 25462 3347 25496 3349
rect 25462 3311 25496 3313
rect 25462 3226 25496 3245
rect 25558 3415 25592 3434
rect 25796 3386 25830 3405
rect 25918 3554 25958 3575
rect 26066 3593 26108 3635
rect 26344 3633 26373 3667
rect 26407 3633 26465 3667
rect 26499 3633 26557 3667
rect 26591 3633 26620 3667
rect 26066 3559 26074 3593
rect 25884 3507 25918 3509
rect 25884 3471 25918 3473
rect 26066 3525 26108 3559
rect 26066 3491 26074 3525
rect 26066 3457 26108 3491
rect 26066 3423 26074 3457
rect 26066 3407 26108 3423
rect 26142 3593 26208 3601
rect 26142 3559 26158 3593
rect 26192 3559 26208 3593
rect 26142 3525 26208 3559
rect 26142 3491 26158 3525
rect 26192 3491 26208 3525
rect 26142 3457 26208 3491
rect 26142 3423 26158 3457
rect 26192 3423 26208 3457
rect 26142 3405 26208 3423
rect 26377 3583 26413 3599
rect 26377 3549 26379 3583
rect 26377 3515 26413 3549
rect 26377 3481 26379 3515
rect 26449 3583 26515 3633
rect 26449 3549 26465 3583
rect 26499 3549 26515 3583
rect 26449 3515 26515 3549
rect 26449 3481 26465 3515
rect 26499 3481 26515 3515
rect 26549 3583 26603 3599
rect 26549 3549 26551 3583
rect 26585 3549 26603 3583
rect 26549 3502 26603 3549
rect 26377 3447 26413 3481
rect 26549 3468 26551 3502
rect 26585 3468 26603 3502
rect 26377 3413 26512 3447
rect 26549 3418 26603 3468
rect 25884 3386 25918 3405
rect 25558 3347 25592 3349
rect 25970 3371 26114 3372
rect 25970 3357 26128 3371
rect 25558 3311 25592 3313
rect 25824 3344 25890 3346
rect 25970 3344 26078 3357
rect 25824 3343 26078 3344
rect 25824 3309 25840 3343
rect 25874 3330 26078 3343
rect 25874 3310 26010 3330
rect 26062 3323 26078 3330
rect 26112 3323 26128 3357
rect 25874 3309 25890 3310
rect 26062 3273 26108 3289
rect 26162 3285 26208 3405
rect 26478 3384 26512 3413
rect 26365 3355 26433 3377
rect 26365 3354 26381 3355
rect 26365 3320 26379 3354
rect 26415 3321 26433 3355
rect 26413 3320 26433 3321
rect 26365 3303 26433 3320
rect 26478 3368 26533 3384
rect 26478 3334 26499 3368
rect 26478 3318 26533 3334
rect 26567 3368 26603 3418
rect 26567 3366 26608 3368
rect 26567 3332 26572 3366
rect 26606 3332 26608 3366
rect 26567 3330 26608 3332
rect 25592 3245 25838 3262
rect 25558 3228 25838 3245
rect 25558 3226 25592 3228
rect 24946 3197 25288 3218
rect 24946 3163 24962 3197
rect 24996 3186 25288 3197
rect 24996 3183 25464 3186
rect 24996 3182 25414 3183
rect 24996 3163 25018 3182
rect 24946 3158 25018 3163
rect 24946 3151 25012 3158
rect 25252 3150 25414 3182
rect 25398 3149 25414 3150
rect 25448 3149 25464 3183
rect 25790 3140 25838 3228
rect 24802 3083 24831 3117
rect 24865 3083 24923 3117
rect 24957 3083 25015 3117
rect 25049 3083 25078 3117
rect 25160 3112 25206 3122
rect 25160 3078 25166 3112
rect 25200 3092 25206 3112
rect 25790 3106 25798 3140
rect 25832 3106 25838 3140
rect 26062 3239 26074 3273
rect 26062 3205 26108 3239
rect 26062 3171 26074 3205
rect 26062 3125 26108 3171
rect 26142 3273 26208 3285
rect 26142 3222 26158 3273
rect 26192 3222 26208 3273
rect 26478 3267 26512 3318
rect 26142 3205 26208 3222
rect 26142 3171 26158 3205
rect 26192 3171 26208 3205
rect 26142 3159 26208 3171
rect 26379 3233 26512 3267
rect 26567 3258 26603 3330
rect 26379 3212 26413 3233
rect 26551 3229 26603 3258
rect 26379 3157 26413 3178
rect 26449 3165 26465 3199
rect 26499 3165 26515 3199
rect 25200 3078 25210 3092
rect 21798 2948 21832 2982
rect 21798 2896 21832 2912
rect 23190 2972 23322 3008
rect 23494 3018 23528 3034
rect 23590 3018 23624 3034
rect 23528 2982 23529 2983
rect 23190 2924 23226 2972
rect 23494 2948 23529 2982
rect 23528 2946 23529 2948
rect 23590 2948 23624 2982
rect 23374 2924 23494 2946
rect 23190 2912 23494 2924
rect 23528 2912 23530 2946
rect 23190 2910 23530 2912
rect 23190 2888 23410 2910
rect 23494 2896 23528 2910
rect 23590 2896 23624 2912
rect 23686 3018 23720 3034
rect 25160 3008 25210 3078
rect 25510 3068 25526 3102
rect 25560 3068 25576 3102
rect 25790 3094 25838 3106
rect 25998 3091 26027 3125
rect 26061 3091 26119 3125
rect 26153 3091 26211 3125
rect 26245 3091 26274 3125
rect 26449 3123 26515 3165
rect 26585 3195 26603 3229
rect 26551 3157 26603 3195
rect 26344 3089 26373 3123
rect 26407 3089 26465 3123
rect 26499 3089 26557 3123
rect 26591 3089 26620 3123
rect 23686 2948 23720 2982
rect 23686 2896 23720 2912
rect 25078 2972 25210 3008
rect 25382 3018 25416 3034
rect 25478 3018 25512 3034
rect 25416 2982 25417 2983
rect 25078 2924 25114 2972
rect 25382 2948 25417 2982
rect 25416 2946 25417 2948
rect 25478 2948 25512 2982
rect 25262 2924 25382 2946
rect 25078 2912 25382 2924
rect 25416 2912 25418 2946
rect 25078 2910 25418 2912
rect 25078 2888 25298 2910
rect 25382 2896 25416 2910
rect 25478 2896 25512 2912
rect 25574 3018 25608 3034
rect 25574 2948 25608 2982
rect 25574 2896 25608 2912
rect -2900 2828 -2884 2862
rect -2850 2828 -2834 2862
rect -1012 2828 -996 2862
rect -962 2828 -946 2862
rect 876 2828 892 2862
rect 926 2828 942 2862
rect 2764 2828 2780 2862
rect 2814 2828 2830 2862
rect 4652 2828 4668 2862
rect 4702 2828 4718 2862
rect 6540 2828 6556 2862
rect 6590 2828 6606 2862
rect 8428 2828 8444 2862
rect 8478 2828 8494 2862
rect 10316 2828 10332 2862
rect 10366 2828 10382 2862
rect 12198 2828 12214 2862
rect 12248 2828 12264 2862
rect 14086 2828 14102 2862
rect 14136 2828 14152 2862
rect 15974 2828 15990 2862
rect 16024 2828 16040 2862
rect 17862 2828 17878 2862
rect 17912 2828 17928 2862
rect 19750 2828 19766 2862
rect 19800 2828 19816 2862
rect 21638 2828 21654 2862
rect 21688 2828 21704 2862
rect 23526 2828 23542 2862
rect 23576 2828 23592 2862
rect 25414 2828 25430 2862
rect 25464 2828 25480 2862
rect -2980 2758 -2710 2778
rect -2980 2753 -2843 2758
rect -2980 2719 -2964 2753
rect -2930 2724 -2843 2753
rect -2809 2724 -2710 2758
rect -2930 2719 -2710 2724
rect -2980 2700 -2710 2719
rect -1092 2758 -822 2778
rect -1092 2753 -955 2758
rect -1092 2719 -1076 2753
rect -1042 2724 -955 2753
rect -921 2724 -822 2758
rect -1042 2719 -822 2724
rect -1092 2700 -822 2719
rect 796 2758 1066 2778
rect 796 2753 933 2758
rect 796 2719 812 2753
rect 846 2724 933 2753
rect 967 2724 1066 2758
rect 846 2719 1066 2724
rect 796 2700 1066 2719
rect 2684 2758 2954 2778
rect 2684 2753 2821 2758
rect 2684 2719 2700 2753
rect 2734 2724 2821 2753
rect 2855 2724 2954 2758
rect 2734 2719 2954 2724
rect 2684 2700 2954 2719
rect 4572 2758 4842 2778
rect 4572 2753 4709 2758
rect 4572 2719 4588 2753
rect 4622 2724 4709 2753
rect 4743 2724 4842 2758
rect 4622 2719 4842 2724
rect 4572 2700 4842 2719
rect 6460 2758 6730 2778
rect 6460 2753 6597 2758
rect 6460 2719 6476 2753
rect 6510 2724 6597 2753
rect 6631 2724 6730 2758
rect 6510 2719 6730 2724
rect 6460 2700 6730 2719
rect 8348 2758 8618 2778
rect 8348 2753 8485 2758
rect 8348 2719 8364 2753
rect 8398 2724 8485 2753
rect 8519 2724 8618 2758
rect 8398 2719 8618 2724
rect 8348 2700 8618 2719
rect 10236 2758 10506 2778
rect 10236 2753 10373 2758
rect 10236 2719 10252 2753
rect 10286 2724 10373 2753
rect 10407 2724 10506 2758
rect 10286 2719 10506 2724
rect 10236 2700 10506 2719
rect 12118 2758 12388 2778
rect 12118 2753 12255 2758
rect 12118 2719 12134 2753
rect 12168 2724 12255 2753
rect 12289 2724 12388 2758
rect 12168 2719 12388 2724
rect 12118 2700 12388 2719
rect 14006 2758 14276 2778
rect 14006 2753 14143 2758
rect 14006 2719 14022 2753
rect 14056 2724 14143 2753
rect 14177 2724 14276 2758
rect 14056 2719 14276 2724
rect 14006 2700 14276 2719
rect 15894 2758 16164 2778
rect 15894 2753 16031 2758
rect 15894 2719 15910 2753
rect 15944 2724 16031 2753
rect 16065 2724 16164 2758
rect 15944 2719 16164 2724
rect 15894 2700 16164 2719
rect 17782 2758 18052 2778
rect 17782 2753 17919 2758
rect 17782 2719 17798 2753
rect 17832 2724 17919 2753
rect 17953 2724 18052 2758
rect 17832 2719 18052 2724
rect 17782 2700 18052 2719
rect 19670 2758 19940 2778
rect 19670 2753 19807 2758
rect 19670 2719 19686 2753
rect 19720 2724 19807 2753
rect 19841 2724 19940 2758
rect 19720 2719 19940 2724
rect 19670 2700 19940 2719
rect 21558 2758 21828 2778
rect 21558 2753 21695 2758
rect 21558 2719 21574 2753
rect 21608 2724 21695 2753
rect 21729 2724 21828 2758
rect 21608 2719 21828 2724
rect 21558 2700 21828 2719
rect 23446 2758 23716 2778
rect 23446 2753 23583 2758
rect 23446 2719 23462 2753
rect 23496 2724 23583 2753
rect 23617 2724 23716 2758
rect 23496 2719 23716 2724
rect 23446 2700 23716 2719
rect 25334 2758 25604 2778
rect 25334 2753 25471 2758
rect 25334 2719 25350 2753
rect 25384 2724 25471 2753
rect 25505 2724 25604 2758
rect 25384 2719 25604 2724
rect 25334 2700 25604 2719
<< viali >>
rect 2141 5305 2175 5339
rect 2233 5305 2267 5339
rect 2325 5305 2359 5339
rect 2417 5305 2451 5339
rect 2509 5305 2543 5339
rect 2601 5305 2635 5339
rect 2693 5305 2727 5339
rect 2785 5305 2819 5339
rect 2877 5305 2911 5339
rect 2969 5305 3003 5339
rect 3061 5305 3095 5339
rect 3153 5305 3187 5339
rect 3245 5305 3279 5339
rect 3337 5305 3371 5339
rect 3429 5305 3463 5339
rect 3521 5305 3555 5339
rect 4023 5303 4057 5337
rect 4115 5303 4149 5337
rect 4207 5303 4241 5337
rect 4299 5303 4333 5337
rect 4391 5303 4425 5337
rect 4483 5303 4517 5337
rect 4575 5303 4609 5337
rect 4667 5303 4701 5337
rect 4759 5303 4793 5337
rect 4851 5303 4885 5337
rect 4943 5303 4977 5337
rect 5035 5303 5069 5337
rect 5127 5303 5161 5337
rect 5219 5303 5253 5337
rect 5311 5303 5345 5337
rect 5403 5303 5437 5337
rect 17239 5305 17273 5339
rect 17331 5305 17365 5339
rect 17423 5305 17457 5339
rect 17515 5305 17549 5339
rect 17607 5305 17641 5339
rect 17699 5305 17733 5339
rect 17791 5305 17825 5339
rect 17883 5305 17917 5339
rect 17975 5305 18009 5339
rect 18067 5305 18101 5339
rect 18159 5305 18193 5339
rect 18251 5305 18285 5339
rect 18343 5305 18377 5339
rect 18435 5305 18469 5339
rect 18527 5305 18561 5339
rect 18619 5305 18653 5339
rect 2268 5068 2302 5102
rect 2381 5068 2415 5102
rect 2494 5073 2496 5102
rect 2496 5073 2528 5102
rect 2494 5068 2528 5073
rect 2607 5068 2641 5102
rect 2720 5068 2754 5102
rect 2833 5073 2866 5102
rect 2866 5073 2867 5102
rect 2833 5068 2867 5073
rect 2946 5068 2980 5102
rect 3062 5068 3096 5102
rect 3166 5073 3167 5102
rect 3167 5073 3200 5102
rect 3166 5068 3200 5073
rect 19121 5303 19155 5337
rect 19213 5303 19247 5337
rect 19305 5303 19339 5337
rect 19397 5303 19431 5337
rect 19489 5303 19523 5337
rect 19581 5303 19615 5337
rect 19673 5303 19707 5337
rect 19765 5303 19799 5337
rect 19857 5303 19891 5337
rect 19949 5303 19983 5337
rect 20041 5303 20075 5337
rect 20133 5303 20167 5337
rect 20225 5303 20259 5337
rect 20317 5303 20351 5337
rect 20409 5303 20443 5337
rect 20501 5303 20535 5337
rect 4022 5071 4036 5102
rect 4036 5071 4056 5102
rect 4022 5068 4056 5071
rect 4141 5068 4175 5102
rect 4260 5068 4294 5102
rect 4379 5071 4412 5102
rect 4412 5071 4413 5102
rect 4379 5068 4413 5071
rect 4498 5068 4532 5102
rect 4617 5068 4651 5102
rect 4736 5071 4748 5102
rect 4748 5071 4770 5102
rect 4736 5068 4770 5071
rect 2245 4975 2278 5007
rect 2278 4975 2279 5007
rect 2245 4973 2279 4975
rect 2411 4975 2412 5005
rect 2412 4975 2445 5005
rect 2411 4971 2445 4975
rect 2575 4975 2580 5003
rect 2580 4975 2609 5003
rect 2575 4969 2609 4975
rect 2746 4975 2748 5005
rect 2748 4975 2780 5005
rect 2746 4971 2780 4975
rect 2915 4975 2916 5001
rect 2916 4975 2949 5001
rect 2915 4967 2949 4975
rect 3084 4975 3118 5000
rect 3084 4966 3118 4975
rect 3250 4975 3252 5006
rect 3252 4975 3284 5006
rect 3250 4972 3284 4975
rect 3420 4975 3454 5008
rect 3420 4974 3454 4975
rect 17434 5073 17460 5102
rect 17460 5073 17468 5102
rect 17434 5068 17468 5073
rect 17531 5068 17565 5102
rect 17628 5068 17662 5102
rect 17725 5068 17759 5102
rect 17822 5068 17856 5102
rect 17919 5073 17930 5102
rect 17930 5073 17953 5102
rect 17919 5068 17953 5073
rect 18016 5068 18050 5102
rect 18113 5073 18132 5102
rect 18132 5073 18147 5102
rect 18113 5068 18147 5073
rect 18264 5073 18265 5102
rect 18265 5073 18298 5102
rect 18264 5068 18298 5073
rect 2141 4761 2175 4795
rect 2233 4761 2267 4795
rect 2325 4761 2359 4795
rect 2417 4761 2451 4795
rect 2509 4761 2543 4795
rect 2601 4761 2635 4795
rect 2693 4761 2727 4795
rect 2785 4761 2819 4795
rect 2877 4761 2911 4795
rect 2969 4761 3003 4795
rect 3061 4761 3095 4795
rect 3153 4761 3187 4795
rect 3245 4761 3279 4795
rect 3337 4761 3371 4795
rect 3429 4761 3463 4795
rect 3521 4761 3555 4795
rect 4630 5007 4664 5009
rect 4134 4973 4160 5005
rect 4160 4973 4168 5005
rect 4134 4971 4168 4973
rect 4294 4973 4328 5005
rect 4294 4971 4328 4973
rect 4461 4973 4462 4999
rect 4462 4973 4495 4999
rect 4461 4965 4495 4973
rect 4630 4975 4664 5007
rect 4794 4973 4798 4996
rect 4798 4973 4828 4996
rect 4794 4962 4828 4973
rect 4964 4973 4966 5002
rect 4966 4973 4998 5002
rect 4964 4968 4998 4973
rect 5134 4973 5168 5004
rect 5134 4970 5168 4973
rect 5293 4973 5302 5006
rect 5302 4973 5327 5006
rect 5293 4972 5327 4973
rect 19120 5071 19134 5102
rect 19134 5071 19154 5102
rect 19120 5068 19154 5071
rect 19228 5068 19262 5102
rect 19336 5071 19342 5102
rect 19342 5071 19370 5102
rect 19336 5068 19370 5071
rect 19444 5071 19476 5102
rect 19476 5071 19478 5102
rect 19444 5068 19478 5071
rect 19552 5068 19586 5102
rect 19660 5071 19679 5102
rect 19679 5071 19694 5102
rect 19660 5068 19694 5071
rect 19768 5068 19802 5102
rect 19876 5068 19910 5102
rect 17343 4975 17376 5001
rect 17376 4975 17377 5001
rect 17343 4967 17377 4975
rect 17506 4975 17510 4996
rect 17510 4975 17540 4996
rect 17506 4962 17540 4975
rect 17679 4975 17712 5000
rect 17712 4975 17713 5000
rect 17679 4966 17713 4975
rect 17844 4975 17846 5005
rect 17846 4975 17878 5005
rect 17844 4971 17878 4975
rect 18011 4975 18014 4992
rect 18014 4975 18045 4992
rect 18011 4958 18045 4975
rect 18179 4975 18182 4990
rect 18182 4975 18213 4990
rect 18179 4956 18213 4975
rect 18349 4975 18350 4999
rect 18350 4975 18383 4999
rect 18349 4965 18383 4975
rect 4023 4759 4057 4793
rect 4115 4759 4149 4793
rect 4207 4759 4241 4793
rect 4299 4759 4333 4793
rect 4391 4759 4425 4793
rect 4483 4759 4517 4793
rect 4575 4759 4609 4793
rect 4667 4759 4701 4793
rect 4759 4759 4793 4793
rect 4851 4759 4885 4793
rect 4943 4759 4977 4793
rect 5035 4759 5069 4793
rect 5127 4759 5161 4793
rect 5219 4759 5253 4793
rect 5311 4759 5345 4793
rect 5403 4759 5437 4793
rect 17239 4761 17273 4795
rect 17331 4761 17365 4795
rect 17423 4761 17457 4795
rect 17515 4761 17549 4795
rect 17607 4761 17641 4795
rect 17699 4761 17733 4795
rect 17791 4761 17825 4795
rect 17883 4761 17917 4795
rect 17975 4761 18009 4795
rect 18067 4761 18101 4795
rect 18159 4761 18193 4795
rect 18251 4761 18285 4795
rect 18343 4761 18377 4795
rect 18435 4761 18469 4795
rect 18527 4761 18561 4795
rect 18619 4761 18653 4795
rect 19728 5007 19762 5009
rect 19222 4973 19224 5000
rect 19224 4973 19256 5000
rect 19222 4966 19256 4973
rect 19395 4973 19426 5001
rect 19426 4973 19429 5001
rect 19395 4967 19429 4973
rect 19557 4973 19560 5006
rect 19560 4973 19591 5006
rect 19557 4972 19591 4973
rect 19728 4975 19762 5007
rect 19897 4973 19930 4995
rect 19930 4973 19931 4995
rect 19897 4961 19931 4973
rect 20062 4973 20064 4995
rect 20064 4973 20096 4995
rect 20062 4961 20096 4973
rect 20232 4973 20266 4993
rect 20232 4959 20266 4973
rect 20395 4973 20400 4997
rect 20400 4973 20429 4997
rect 20395 4963 20429 4973
rect 19121 4759 19155 4793
rect 19213 4759 19247 4793
rect 19305 4759 19339 4793
rect 19397 4759 19431 4793
rect 19489 4759 19523 4793
rect 19581 4759 19615 4793
rect 19673 4759 19707 4793
rect 19765 4759 19799 4793
rect 19857 4759 19891 4793
rect 19949 4759 19983 4793
rect 20041 4759 20075 4793
rect 20133 4759 20167 4793
rect 20225 4759 20259 4793
rect 20317 4759 20351 4793
rect 20409 4759 20443 4793
rect 20501 4759 20535 4793
rect -3305 4681 -3271 4715
rect -3213 4681 -3179 4715
rect -3121 4681 -3087 4715
rect -2491 4681 -2457 4715
rect -2399 4681 -2365 4715
rect -2307 4681 -2273 4715
rect -1417 4681 -1383 4715
rect -1325 4681 -1291 4715
rect -1233 4681 -1199 4715
rect -603 4681 -569 4715
rect -511 4681 -477 4715
rect -419 4681 -385 4715
rect 471 4681 505 4715
rect 563 4681 597 4715
rect 655 4681 689 4715
rect 1285 4681 1319 4715
rect 1377 4681 1411 4715
rect 1469 4681 1503 4715
rect 2359 4681 2393 4715
rect 2451 4681 2485 4715
rect 2543 4681 2577 4715
rect 3173 4681 3207 4715
rect 3265 4681 3299 4715
rect 3357 4681 3391 4715
rect 4247 4681 4281 4715
rect 4339 4681 4373 4715
rect 4431 4681 4465 4715
rect 5061 4681 5095 4715
rect 5153 4681 5187 4715
rect 5245 4681 5279 4715
rect 6135 4681 6169 4715
rect 6227 4681 6261 4715
rect 6319 4681 6353 4715
rect 6949 4681 6983 4715
rect 7041 4681 7075 4715
rect 7133 4681 7167 4715
rect 8023 4681 8057 4715
rect 8115 4681 8149 4715
rect 8207 4681 8241 4715
rect 8837 4681 8871 4715
rect 8929 4681 8963 4715
rect 9021 4681 9055 4715
rect 9911 4681 9945 4715
rect 10003 4681 10037 4715
rect 10095 4681 10129 4715
rect 10725 4681 10759 4715
rect 10817 4681 10851 4715
rect 10909 4681 10943 4715
rect 11793 4681 11827 4715
rect 11885 4681 11919 4715
rect 11977 4681 12011 4715
rect 12607 4681 12641 4715
rect 12699 4681 12733 4715
rect 12791 4681 12825 4715
rect 13681 4681 13715 4715
rect 13773 4681 13807 4715
rect 13865 4681 13899 4715
rect 14495 4681 14529 4715
rect 14587 4681 14621 4715
rect 14679 4681 14713 4715
rect 15569 4681 15603 4715
rect 15661 4681 15695 4715
rect 15753 4681 15787 4715
rect 16383 4681 16417 4715
rect 16475 4681 16509 4715
rect 16567 4681 16601 4715
rect 17457 4681 17491 4715
rect 17549 4681 17583 4715
rect 17641 4681 17675 4715
rect 18271 4681 18305 4715
rect 18363 4681 18397 4715
rect 18455 4681 18489 4715
rect 19345 4681 19379 4715
rect 19437 4681 19471 4715
rect 19529 4681 19563 4715
rect 20159 4681 20193 4715
rect 20251 4681 20285 4715
rect 20343 4681 20377 4715
rect 21233 4681 21267 4715
rect 21325 4681 21359 4715
rect 21417 4681 21451 4715
rect 22047 4681 22081 4715
rect 22139 4681 22173 4715
rect 22231 4681 22265 4715
rect 23121 4681 23155 4715
rect 23213 4681 23247 4715
rect 23305 4681 23339 4715
rect 23935 4681 23969 4715
rect 24027 4681 24061 4715
rect 24119 4681 24153 4715
rect 25009 4681 25043 4715
rect 25101 4681 25135 4715
rect 25193 4681 25227 4715
rect 25823 4681 25857 4715
rect 25915 4681 25949 4715
rect 26007 4681 26041 4715
rect -2871 4641 -2837 4675
rect -2802 4533 -2768 4567
rect -3299 4403 -3265 4412
rect -3299 4378 -3297 4403
rect -3297 4378 -3265 4403
rect -3126 4403 -3092 4408
rect -3126 4374 -3095 4403
rect -3095 4374 -3092 4403
rect -3217 4283 -3215 4292
rect -3215 4283 -3183 4292
rect -3217 4258 -3183 4283
rect -3305 4137 -3271 4171
rect -3213 4137 -3179 4171
rect -3121 4137 -3087 4171
rect -3334 3892 -3300 3926
rect -2946 4437 -2912 4439
rect -2946 4405 -2912 4437
rect -2946 4335 -2912 4367
rect -2946 4333 -2912 4335
rect -2850 4437 -2816 4439
rect -2850 4405 -2816 4437
rect -2850 4335 -2816 4367
rect -2850 4333 -2816 4335
rect -983 4641 -949 4675
rect -914 4533 -880 4567
rect -2754 4437 -2720 4439
rect -2754 4405 -2720 4437
rect -2487 4403 -2453 4410
rect -2487 4376 -2483 4403
rect -2483 4376 -2453 4403
rect -2754 4335 -2720 4367
rect -2754 4333 -2720 4335
rect -2313 4403 -2279 4410
rect -2313 4376 -2281 4403
rect -2281 4376 -2279 4403
rect -1411 4403 -1377 4412
rect -1411 4378 -1409 4403
rect -1409 4378 -1377 4403
rect -1238 4403 -1204 4408
rect -1238 4374 -1207 4403
rect -1207 4374 -1204 4403
rect -2898 4205 -2864 4239
rect -2399 4283 -2367 4287
rect -2367 4283 -2365 4287
rect -2399 4253 -2365 4283
rect -1329 4283 -1327 4292
rect -1327 4283 -1295 4292
rect -1329 4258 -1295 4283
rect -2786 4124 -2752 4158
rect -2491 4137 -2457 4171
rect -2399 4137 -2365 4171
rect -2307 4137 -2273 4171
rect -1417 4137 -1383 4171
rect -1325 4137 -1291 4171
rect -1233 4137 -1199 4171
rect -2930 4072 -2896 4074
rect -2930 4040 -2896 4072
rect -2930 3970 -2896 4002
rect -2930 3968 -2896 3970
rect -2834 4072 -2800 4074
rect -2834 4040 -2800 4072
rect -2834 3970 -2800 4002
rect -2834 3968 -2800 3970
rect -2738 4072 -2704 4074
rect -2738 4040 -2704 4072
rect -2738 3970 -2704 4002
rect -2738 3968 -2704 3970
rect -2882 3884 -2848 3918
rect -2962 3775 -2928 3809
rect -2532 3758 -2498 3792
rect -3483 3627 -3449 3661
rect -3391 3627 -3357 3661
rect -3299 3627 -3265 3661
rect -3120 3637 -3086 3671
rect -2474 3637 -2440 3671
rect -3434 3349 -3400 3360
rect -3434 3326 -3432 3349
rect -3432 3326 -3400 3349
rect -2873 3585 -2839 3619
rect -1446 3892 -1412 3926
rect -1058 4437 -1024 4439
rect -1058 4405 -1024 4437
rect -1058 4335 -1024 4367
rect -1058 4333 -1024 4335
rect -962 4437 -928 4439
rect -962 4405 -928 4437
rect -962 4335 -928 4367
rect -962 4333 -928 4335
rect 905 4641 939 4675
rect 974 4533 1008 4567
rect -866 4437 -832 4439
rect -866 4405 -832 4437
rect -599 4403 -565 4410
rect -599 4376 -595 4403
rect -595 4376 -565 4403
rect -866 4335 -832 4367
rect -866 4333 -832 4335
rect -425 4403 -391 4410
rect -425 4376 -393 4403
rect -393 4376 -391 4403
rect 477 4403 511 4412
rect 477 4378 479 4403
rect 479 4378 511 4403
rect 650 4403 684 4408
rect 650 4374 681 4403
rect 681 4374 684 4403
rect -1010 4205 -976 4239
rect -511 4283 -479 4287
rect -479 4283 -477 4287
rect -511 4253 -477 4283
rect 559 4283 561 4292
rect 561 4283 593 4292
rect 559 4258 593 4283
rect -898 4124 -864 4158
rect -603 4137 -569 4171
rect -511 4137 -477 4171
rect -419 4137 -385 4171
rect 471 4137 505 4171
rect 563 4137 597 4171
rect 655 4137 689 4171
rect -1042 4072 -1008 4074
rect -1042 4040 -1008 4072
rect -1042 3970 -1008 4002
rect -1042 3968 -1008 3970
rect -946 4072 -912 4074
rect -946 4040 -912 4072
rect -946 3970 -912 4002
rect -946 3968 -912 3970
rect -850 4072 -816 4074
rect -850 4040 -816 4072
rect -850 3970 -816 4002
rect -850 3968 -816 3970
rect -994 3884 -960 3918
rect -1074 3775 -1040 3809
rect -644 3758 -610 3792
rect -2287 3635 -2253 3669
rect -2195 3635 -2161 3669
rect -2103 3635 -2069 3669
rect -3164 3541 -3130 3543
rect -3164 3509 -3130 3541
rect -3164 3439 -3130 3471
rect -3164 3437 -3130 3439
rect -3076 3541 -3042 3543
rect -3076 3509 -3042 3541
rect -2518 3541 -2484 3543
rect -2804 3477 -2770 3511
rect -2518 3509 -2484 3541
rect -3076 3439 -3042 3471
rect -3076 3437 -3042 3439
rect -2518 3439 -2484 3471
rect -2518 3437 -2484 3439
rect -2948 3381 -2914 3383
rect -2948 3349 -2914 3381
rect -3120 3309 -3086 3343
rect -2948 3279 -2914 3311
rect -2948 3277 -2914 3279
rect -2852 3381 -2818 3383
rect -2852 3349 -2818 3381
rect -2852 3279 -2818 3311
rect -2852 3277 -2818 3279
rect -1941 3633 -1907 3667
rect -1849 3633 -1815 3667
rect -1757 3633 -1723 3667
rect -2430 3541 -2396 3543
rect -2430 3509 -2396 3541
rect -2430 3439 -2396 3471
rect -2430 3437 -2396 3439
rect -1595 3627 -1561 3661
rect -1503 3627 -1469 3661
rect -1411 3627 -1377 3661
rect -1232 3637 -1198 3671
rect -2756 3381 -2722 3383
rect -2756 3349 -2722 3381
rect -2756 3279 -2722 3311
rect -2474 3309 -2440 3343
rect -2756 3277 -2722 3279
rect -1935 3321 -1933 3354
rect -1933 3321 -1901 3354
rect -1935 3320 -1901 3321
rect -586 3637 -552 3671
rect -1742 3332 -1708 3366
rect -2900 3149 -2866 3183
rect -3483 3083 -3449 3117
rect -3391 3083 -3357 3117
rect -3299 3083 -3265 3117
rect -3148 3078 -3114 3112
rect -2516 3106 -2482 3140
rect -2156 3239 -2122 3256
rect -2156 3222 -2122 3239
rect -1546 3349 -1512 3360
rect -1546 3326 -1544 3349
rect -1544 3326 -1512 3349
rect -2788 3068 -2754 3102
rect -2287 3091 -2253 3125
rect -2195 3091 -2161 3125
rect -2103 3091 -2069 3125
rect -985 3585 -951 3619
rect 442 3892 476 3926
rect 830 4437 864 4439
rect 830 4405 864 4437
rect 830 4335 864 4367
rect 830 4333 864 4335
rect 926 4437 960 4439
rect 926 4405 960 4437
rect 926 4335 960 4367
rect 926 4333 960 4335
rect 2793 4641 2827 4675
rect 2862 4533 2896 4567
rect 1022 4437 1056 4439
rect 1022 4405 1056 4437
rect 1289 4403 1323 4410
rect 1289 4376 1293 4403
rect 1293 4376 1323 4403
rect 1022 4335 1056 4367
rect 1022 4333 1056 4335
rect 1463 4403 1497 4410
rect 1463 4376 1495 4403
rect 1495 4376 1497 4403
rect 2365 4403 2399 4412
rect 2365 4378 2367 4403
rect 2367 4378 2399 4403
rect 2538 4403 2572 4408
rect 2538 4374 2569 4403
rect 2569 4374 2572 4403
rect 878 4205 912 4239
rect 1377 4283 1409 4287
rect 1409 4283 1411 4287
rect 1377 4253 1411 4283
rect 2447 4283 2449 4292
rect 2449 4283 2481 4292
rect 2447 4258 2481 4283
rect 990 4124 1024 4158
rect 1285 4137 1319 4171
rect 1377 4137 1411 4171
rect 1469 4137 1503 4171
rect 2359 4137 2393 4171
rect 2451 4137 2485 4171
rect 2543 4137 2577 4171
rect 846 4072 880 4074
rect 846 4040 880 4072
rect 846 3970 880 4002
rect 846 3968 880 3970
rect 942 4072 976 4074
rect 942 4040 976 4072
rect 942 3970 976 4002
rect 942 3968 976 3970
rect 1038 4072 1072 4074
rect 1038 4040 1072 4072
rect 1038 3970 1072 4002
rect 1038 3968 1072 3970
rect 894 3884 928 3918
rect 814 3775 848 3809
rect 1244 3758 1278 3792
rect -399 3635 -365 3669
rect -307 3635 -273 3669
rect -215 3635 -181 3669
rect -1276 3541 -1242 3543
rect -1276 3509 -1242 3541
rect -1276 3439 -1242 3471
rect -1276 3437 -1242 3439
rect -1188 3541 -1154 3543
rect -1188 3509 -1154 3541
rect -630 3541 -596 3543
rect -916 3477 -882 3511
rect -630 3509 -596 3541
rect -1188 3439 -1154 3471
rect -1188 3437 -1154 3439
rect -630 3439 -596 3471
rect -630 3437 -596 3439
rect -1060 3381 -1026 3383
rect -1060 3349 -1026 3381
rect -1232 3309 -1198 3343
rect -1941 3089 -1907 3123
rect -1849 3089 -1815 3123
rect -1757 3089 -1723 3123
rect -1060 3279 -1026 3311
rect -1060 3277 -1026 3279
rect -964 3381 -930 3383
rect -964 3349 -930 3381
rect -964 3279 -930 3311
rect -964 3277 -930 3279
rect -53 3633 -19 3667
rect 39 3633 73 3667
rect 131 3633 165 3667
rect -542 3541 -508 3543
rect -542 3509 -508 3541
rect -542 3439 -508 3471
rect -542 3437 -508 3439
rect 293 3627 327 3661
rect 385 3627 419 3661
rect 477 3627 511 3661
rect 656 3637 690 3671
rect -868 3381 -834 3383
rect -868 3349 -834 3381
rect -868 3279 -834 3311
rect -586 3309 -552 3343
rect -868 3277 -834 3279
rect -47 3321 -45 3354
rect -45 3321 -13 3354
rect -47 3320 -13 3321
rect 1302 3637 1336 3671
rect 146 3332 180 3366
rect -1012 3149 -978 3183
rect -1595 3083 -1561 3117
rect -1503 3083 -1469 3117
rect -1411 3083 -1377 3117
rect -1260 3078 -1226 3112
rect -628 3106 -594 3140
rect -268 3239 -234 3256
rect -268 3222 -234 3239
rect 342 3349 376 3360
rect 342 3326 344 3349
rect 344 3326 376 3349
rect -2932 3016 -2898 3018
rect -2932 2984 -2898 3016
rect -2836 3016 -2802 3018
rect -2836 2984 -2802 3016
rect -2932 2914 -2898 2946
rect -2932 2912 -2898 2914
rect -2836 2914 -2802 2946
rect -2836 2912 -2802 2914
rect -2740 3016 -2706 3018
rect -2740 2984 -2706 3016
rect -900 3068 -866 3102
rect -399 3091 -365 3125
rect -307 3091 -273 3125
rect -215 3091 -181 3125
rect 903 3585 937 3619
rect 2330 3892 2364 3926
rect 2718 4437 2752 4439
rect 2718 4405 2752 4437
rect 2718 4335 2752 4367
rect 2718 4333 2752 4335
rect 2814 4437 2848 4439
rect 2814 4405 2848 4437
rect 2814 4335 2848 4367
rect 2814 4333 2848 4335
rect 4681 4641 4715 4675
rect 4750 4533 4784 4567
rect 2910 4437 2944 4439
rect 2910 4405 2944 4437
rect 3177 4403 3211 4410
rect 3177 4376 3181 4403
rect 3181 4376 3211 4403
rect 2910 4335 2944 4367
rect 2910 4333 2944 4335
rect 3351 4403 3385 4410
rect 3351 4376 3383 4403
rect 3383 4376 3385 4403
rect 4253 4403 4287 4412
rect 4253 4378 4255 4403
rect 4255 4378 4287 4403
rect 4426 4403 4460 4408
rect 4426 4374 4457 4403
rect 4457 4374 4460 4403
rect 2766 4205 2800 4239
rect 3265 4283 3297 4287
rect 3297 4283 3299 4287
rect 3265 4253 3299 4283
rect 4335 4283 4337 4292
rect 4337 4283 4369 4292
rect 4335 4258 4369 4283
rect 2878 4124 2912 4158
rect 3173 4137 3207 4171
rect 3265 4137 3299 4171
rect 3357 4137 3391 4171
rect 4247 4137 4281 4171
rect 4339 4137 4373 4171
rect 4431 4137 4465 4171
rect 2734 4072 2768 4074
rect 2734 4040 2768 4072
rect 2734 3970 2768 4002
rect 2734 3968 2768 3970
rect 2830 4072 2864 4074
rect 2830 4040 2864 4072
rect 2830 3970 2864 4002
rect 2830 3968 2864 3970
rect 2926 4072 2960 4074
rect 2926 4040 2960 4072
rect 2926 3970 2960 4002
rect 2926 3968 2960 3970
rect 2782 3884 2816 3918
rect 2702 3775 2736 3809
rect 3132 3758 3166 3792
rect 1489 3635 1523 3669
rect 1581 3635 1615 3669
rect 1673 3635 1707 3669
rect 612 3541 646 3543
rect 612 3509 646 3541
rect 612 3439 646 3471
rect 612 3437 646 3439
rect 700 3541 734 3543
rect 700 3509 734 3541
rect 1258 3541 1292 3543
rect 972 3477 1006 3511
rect 1258 3509 1292 3541
rect 700 3439 734 3471
rect 700 3437 734 3439
rect 1258 3439 1292 3471
rect 1258 3437 1292 3439
rect 828 3381 862 3383
rect 828 3349 862 3381
rect 656 3309 690 3343
rect -53 3089 -19 3123
rect 39 3089 73 3123
rect 131 3089 165 3123
rect 828 3279 862 3311
rect 828 3277 862 3279
rect 924 3381 958 3383
rect 924 3349 958 3381
rect 924 3279 958 3311
rect 924 3277 958 3279
rect 1835 3633 1869 3667
rect 1927 3633 1961 3667
rect 2019 3633 2053 3667
rect 1346 3541 1380 3543
rect 1346 3509 1380 3541
rect 1346 3439 1380 3471
rect 1346 3437 1380 3439
rect 2181 3627 2215 3661
rect 2273 3627 2307 3661
rect 2365 3627 2399 3661
rect 2544 3637 2578 3671
rect 1020 3381 1054 3383
rect 1020 3349 1054 3381
rect 1020 3279 1054 3311
rect 1302 3309 1336 3343
rect 1020 3277 1054 3279
rect 1841 3321 1843 3354
rect 1843 3321 1875 3354
rect 1841 3320 1875 3321
rect 3190 3637 3224 3671
rect 2034 3332 2068 3366
rect 876 3149 910 3183
rect 293 3083 327 3117
rect 385 3083 419 3117
rect 477 3083 511 3117
rect 628 3078 662 3112
rect 1260 3106 1294 3140
rect 1620 3239 1654 3256
rect 1620 3222 1654 3239
rect 2230 3349 2264 3360
rect 2230 3326 2232 3349
rect 2232 3326 2264 3349
rect -2740 2914 -2706 2946
rect -2740 2912 -2706 2914
rect -1044 3016 -1010 3018
rect -1044 2984 -1010 3016
rect -948 3016 -914 3018
rect -948 2984 -914 3016
rect -1044 2914 -1010 2946
rect -1044 2912 -1010 2914
rect -948 2914 -914 2946
rect -948 2912 -914 2914
rect -852 3016 -818 3018
rect -852 2984 -818 3016
rect 988 3068 1022 3102
rect 1489 3091 1523 3125
rect 1581 3091 1615 3125
rect 1673 3091 1707 3125
rect 2791 3585 2825 3619
rect 4218 3892 4252 3926
rect 4606 4437 4640 4439
rect 4606 4405 4640 4437
rect 4606 4335 4640 4367
rect 4606 4333 4640 4335
rect 4702 4437 4736 4439
rect 4702 4405 4736 4437
rect 4702 4335 4736 4367
rect 4702 4333 4736 4335
rect 6569 4641 6603 4675
rect 6638 4533 6672 4567
rect 4798 4437 4832 4439
rect 4798 4405 4832 4437
rect 5065 4403 5099 4410
rect 5065 4376 5069 4403
rect 5069 4376 5099 4403
rect 4798 4335 4832 4367
rect 4798 4333 4832 4335
rect 5239 4403 5273 4410
rect 5239 4376 5271 4403
rect 5271 4376 5273 4403
rect 6141 4403 6175 4412
rect 6141 4378 6143 4403
rect 6143 4378 6175 4403
rect 6314 4403 6348 4408
rect 6314 4374 6345 4403
rect 6345 4374 6348 4403
rect 4654 4205 4688 4239
rect 5153 4283 5185 4287
rect 5185 4283 5187 4287
rect 5153 4253 5187 4283
rect 6223 4283 6225 4292
rect 6225 4283 6257 4292
rect 6223 4258 6257 4283
rect 4766 4124 4800 4158
rect 5061 4137 5095 4171
rect 5153 4137 5187 4171
rect 5245 4137 5279 4171
rect 6135 4137 6169 4171
rect 6227 4137 6261 4171
rect 6319 4137 6353 4171
rect 4622 4072 4656 4074
rect 4622 4040 4656 4072
rect 4622 3970 4656 4002
rect 4622 3968 4656 3970
rect 4718 4072 4752 4074
rect 4718 4040 4752 4072
rect 4718 3970 4752 4002
rect 4718 3968 4752 3970
rect 4814 4072 4848 4074
rect 4814 4040 4848 4072
rect 4814 3970 4848 4002
rect 4814 3968 4848 3970
rect 4670 3884 4704 3918
rect 4590 3775 4624 3809
rect 5020 3758 5054 3792
rect 3377 3635 3411 3669
rect 3469 3635 3503 3669
rect 3561 3635 3595 3669
rect 2500 3541 2534 3543
rect 2500 3509 2534 3541
rect 2500 3439 2534 3471
rect 2500 3437 2534 3439
rect 2588 3541 2622 3543
rect 2588 3509 2622 3541
rect 3146 3541 3180 3543
rect 2860 3477 2894 3511
rect 3146 3509 3180 3541
rect 2588 3439 2622 3471
rect 2588 3437 2622 3439
rect 3146 3439 3180 3471
rect 3146 3437 3180 3439
rect 2716 3381 2750 3383
rect 2716 3349 2750 3381
rect 2544 3309 2578 3343
rect 1835 3089 1869 3123
rect 1927 3089 1961 3123
rect 2019 3089 2053 3123
rect 2716 3279 2750 3311
rect 2716 3277 2750 3279
rect 2812 3381 2846 3383
rect 2812 3349 2846 3381
rect 2812 3279 2846 3311
rect 2812 3277 2846 3279
rect 3723 3633 3757 3667
rect 3815 3633 3849 3667
rect 3907 3633 3941 3667
rect 3234 3541 3268 3543
rect 3234 3509 3268 3541
rect 3234 3439 3268 3471
rect 3234 3437 3268 3439
rect 4069 3627 4103 3661
rect 4161 3627 4195 3661
rect 4253 3627 4287 3661
rect 4432 3637 4466 3671
rect 2908 3381 2942 3383
rect 2908 3349 2942 3381
rect 2908 3279 2942 3311
rect 3190 3309 3224 3343
rect 2908 3277 2942 3279
rect 3729 3321 3731 3354
rect 3731 3321 3763 3354
rect 3729 3320 3763 3321
rect 5078 3637 5112 3671
rect 3922 3332 3956 3366
rect 2764 3149 2798 3183
rect 2181 3083 2215 3117
rect 2273 3083 2307 3117
rect 2365 3083 2399 3117
rect 2516 3078 2550 3112
rect 3148 3106 3182 3140
rect 3508 3239 3542 3256
rect 3508 3222 3542 3239
rect 4118 3349 4152 3360
rect 4118 3326 4120 3349
rect 4120 3326 4152 3349
rect -852 2914 -818 2946
rect -852 2912 -818 2914
rect 844 3016 878 3018
rect 844 2984 878 3016
rect 940 3016 974 3018
rect 940 2984 974 3016
rect 844 2914 878 2946
rect 844 2912 878 2914
rect 940 2914 974 2946
rect 940 2912 974 2914
rect 1036 3016 1070 3018
rect 1036 2984 1070 3016
rect 2876 3068 2910 3102
rect 3377 3091 3411 3125
rect 3469 3091 3503 3125
rect 3561 3091 3595 3125
rect 4679 3585 4713 3619
rect 6106 3892 6140 3926
rect 6494 4437 6528 4439
rect 6494 4405 6528 4437
rect 6494 4335 6528 4367
rect 6494 4333 6528 4335
rect 6590 4437 6624 4439
rect 6590 4405 6624 4437
rect 6590 4335 6624 4367
rect 6590 4333 6624 4335
rect 8457 4641 8491 4675
rect 8526 4533 8560 4567
rect 6686 4437 6720 4439
rect 6686 4405 6720 4437
rect 6953 4403 6987 4410
rect 6953 4376 6957 4403
rect 6957 4376 6987 4403
rect 6686 4335 6720 4367
rect 6686 4333 6720 4335
rect 7127 4403 7161 4410
rect 7127 4376 7159 4403
rect 7159 4376 7161 4403
rect 8029 4403 8063 4412
rect 8029 4378 8031 4403
rect 8031 4378 8063 4403
rect 8202 4403 8236 4408
rect 8202 4374 8233 4403
rect 8233 4374 8236 4403
rect 6542 4205 6576 4239
rect 7041 4283 7073 4287
rect 7073 4283 7075 4287
rect 7041 4253 7075 4283
rect 8111 4283 8113 4292
rect 8113 4283 8145 4292
rect 8111 4258 8145 4283
rect 6654 4124 6688 4158
rect 6949 4137 6983 4171
rect 7041 4137 7075 4171
rect 7133 4137 7167 4171
rect 8023 4137 8057 4171
rect 8115 4137 8149 4171
rect 8207 4137 8241 4171
rect 6510 4072 6544 4074
rect 6510 4040 6544 4072
rect 6510 3970 6544 4002
rect 6510 3968 6544 3970
rect 6606 4072 6640 4074
rect 6606 4040 6640 4072
rect 6606 3970 6640 4002
rect 6606 3968 6640 3970
rect 6702 4072 6736 4074
rect 6702 4040 6736 4072
rect 6702 3970 6736 4002
rect 6702 3968 6736 3970
rect 6558 3884 6592 3918
rect 6478 3775 6512 3809
rect 6908 3758 6942 3792
rect 5265 3635 5299 3669
rect 5357 3635 5391 3669
rect 5449 3635 5483 3669
rect 4388 3541 4422 3543
rect 4388 3509 4422 3541
rect 4388 3439 4422 3471
rect 4388 3437 4422 3439
rect 4476 3541 4510 3543
rect 4476 3509 4510 3541
rect 5034 3541 5068 3543
rect 4748 3477 4782 3511
rect 5034 3509 5068 3541
rect 4476 3439 4510 3471
rect 4476 3437 4510 3439
rect 5034 3439 5068 3471
rect 5034 3437 5068 3439
rect 4604 3381 4638 3383
rect 4604 3349 4638 3381
rect 4432 3309 4466 3343
rect 3723 3089 3757 3123
rect 3815 3089 3849 3123
rect 3907 3089 3941 3123
rect 4604 3279 4638 3311
rect 4604 3277 4638 3279
rect 4700 3381 4734 3383
rect 4700 3349 4734 3381
rect 4700 3279 4734 3311
rect 4700 3277 4734 3279
rect 5611 3633 5645 3667
rect 5703 3633 5737 3667
rect 5795 3633 5829 3667
rect 5122 3541 5156 3543
rect 5122 3509 5156 3541
rect 5122 3439 5156 3471
rect 5122 3437 5156 3439
rect 5957 3627 5991 3661
rect 6049 3627 6083 3661
rect 6141 3627 6175 3661
rect 6320 3637 6354 3671
rect 4796 3381 4830 3383
rect 4796 3349 4830 3381
rect 4796 3279 4830 3311
rect 5078 3309 5112 3343
rect 4796 3277 4830 3279
rect 5617 3321 5619 3354
rect 5619 3321 5651 3354
rect 5617 3320 5651 3321
rect 6966 3637 7000 3671
rect 5810 3332 5844 3366
rect 4652 3149 4686 3183
rect 4069 3083 4103 3117
rect 4161 3083 4195 3117
rect 4253 3083 4287 3117
rect 4404 3078 4438 3112
rect 5036 3106 5070 3140
rect 5396 3239 5430 3256
rect 5396 3222 5430 3239
rect 6006 3349 6040 3360
rect 6006 3326 6008 3349
rect 6008 3326 6040 3349
rect 1036 2914 1070 2946
rect 1036 2912 1070 2914
rect 2732 3016 2766 3018
rect 2732 2984 2766 3016
rect 2828 3016 2862 3018
rect 2828 2984 2862 3016
rect 2732 2914 2766 2946
rect 2732 2912 2766 2914
rect 2828 2914 2862 2946
rect 2828 2912 2862 2914
rect 2924 3016 2958 3018
rect 2924 2984 2958 3016
rect 4764 3068 4798 3102
rect 5265 3091 5299 3125
rect 5357 3091 5391 3125
rect 5449 3091 5483 3125
rect 6567 3585 6601 3619
rect 7994 3892 8028 3926
rect 8382 4437 8416 4439
rect 8382 4405 8416 4437
rect 8382 4335 8416 4367
rect 8382 4333 8416 4335
rect 8478 4437 8512 4439
rect 8478 4405 8512 4437
rect 8478 4335 8512 4367
rect 8478 4333 8512 4335
rect 10345 4641 10379 4675
rect 10414 4533 10448 4567
rect 8574 4437 8608 4439
rect 8574 4405 8608 4437
rect 8841 4403 8875 4410
rect 8841 4376 8845 4403
rect 8845 4376 8875 4403
rect 8574 4335 8608 4367
rect 8574 4333 8608 4335
rect 9015 4403 9049 4410
rect 9015 4376 9047 4403
rect 9047 4376 9049 4403
rect 9917 4403 9951 4412
rect 9917 4378 9919 4403
rect 9919 4378 9951 4403
rect 10090 4403 10124 4408
rect 10090 4374 10121 4403
rect 10121 4374 10124 4403
rect 8430 4205 8464 4239
rect 8929 4283 8961 4287
rect 8961 4283 8963 4287
rect 8929 4253 8963 4283
rect 9999 4283 10001 4292
rect 10001 4283 10033 4292
rect 9999 4258 10033 4283
rect 8542 4124 8576 4158
rect 8837 4137 8871 4171
rect 8929 4137 8963 4171
rect 9021 4137 9055 4171
rect 9911 4137 9945 4171
rect 10003 4137 10037 4171
rect 10095 4137 10129 4171
rect 8398 4072 8432 4074
rect 8398 4040 8432 4072
rect 8398 3970 8432 4002
rect 8398 3968 8432 3970
rect 8494 4072 8528 4074
rect 8494 4040 8528 4072
rect 8494 3970 8528 4002
rect 8494 3968 8528 3970
rect 8590 4072 8624 4074
rect 8590 4040 8624 4072
rect 8590 3970 8624 4002
rect 8590 3968 8624 3970
rect 8446 3884 8480 3918
rect 8366 3775 8400 3809
rect 8796 3758 8830 3792
rect 7153 3635 7187 3669
rect 7245 3635 7279 3669
rect 7337 3635 7371 3669
rect 6276 3541 6310 3543
rect 6276 3509 6310 3541
rect 6276 3439 6310 3471
rect 6276 3437 6310 3439
rect 6364 3541 6398 3543
rect 6364 3509 6398 3541
rect 6922 3541 6956 3543
rect 6636 3477 6670 3511
rect 6922 3509 6956 3541
rect 6364 3439 6398 3471
rect 6364 3437 6398 3439
rect 6922 3439 6956 3471
rect 6922 3437 6956 3439
rect 6492 3381 6526 3383
rect 6492 3349 6526 3381
rect 6320 3309 6354 3343
rect 5611 3089 5645 3123
rect 5703 3089 5737 3123
rect 5795 3089 5829 3123
rect 6492 3279 6526 3311
rect 6492 3277 6526 3279
rect 6588 3381 6622 3383
rect 6588 3349 6622 3381
rect 6588 3279 6622 3311
rect 6588 3277 6622 3279
rect 7499 3633 7533 3667
rect 7591 3633 7625 3667
rect 7683 3633 7717 3667
rect 7010 3541 7044 3543
rect 7010 3509 7044 3541
rect 7010 3439 7044 3471
rect 7010 3437 7044 3439
rect 7845 3627 7879 3661
rect 7937 3627 7971 3661
rect 8029 3627 8063 3661
rect 8208 3637 8242 3671
rect 6684 3381 6718 3383
rect 6684 3349 6718 3381
rect 6684 3279 6718 3311
rect 6966 3309 7000 3343
rect 6684 3277 6718 3279
rect 7505 3321 7507 3354
rect 7507 3321 7539 3354
rect 7505 3320 7539 3321
rect 8854 3637 8888 3671
rect 7698 3332 7732 3366
rect 6540 3149 6574 3183
rect 5957 3083 5991 3117
rect 6049 3083 6083 3117
rect 6141 3083 6175 3117
rect 6292 3078 6326 3112
rect 6924 3106 6958 3140
rect 7284 3239 7318 3256
rect 7284 3222 7318 3239
rect 7894 3349 7928 3360
rect 7894 3326 7896 3349
rect 7896 3326 7928 3349
rect 2924 2914 2958 2946
rect 2924 2912 2958 2914
rect 4620 3016 4654 3018
rect 4620 2984 4654 3016
rect 4716 3016 4750 3018
rect 4716 2984 4750 3016
rect 4620 2914 4654 2946
rect 4620 2912 4654 2914
rect 4716 2914 4750 2946
rect 4716 2912 4750 2914
rect 4812 3016 4846 3018
rect 4812 2984 4846 3016
rect 6652 3068 6686 3102
rect 7153 3091 7187 3125
rect 7245 3091 7279 3125
rect 7337 3091 7371 3125
rect 8455 3585 8489 3619
rect 9882 3892 9916 3926
rect 10270 4437 10304 4439
rect 10270 4405 10304 4437
rect 10270 4335 10304 4367
rect 10270 4333 10304 4335
rect 10366 4437 10400 4439
rect 10366 4405 10400 4437
rect 10366 4335 10400 4367
rect 10366 4333 10400 4335
rect 12227 4641 12261 4675
rect 12296 4533 12330 4567
rect 10462 4437 10496 4439
rect 10462 4405 10496 4437
rect 10729 4403 10763 4410
rect 10729 4376 10733 4403
rect 10733 4376 10763 4403
rect 10462 4335 10496 4367
rect 10462 4333 10496 4335
rect 10903 4403 10937 4410
rect 10903 4376 10935 4403
rect 10935 4376 10937 4403
rect 11799 4403 11833 4412
rect 11799 4378 11801 4403
rect 11801 4378 11833 4403
rect 11972 4403 12006 4408
rect 11972 4374 12003 4403
rect 12003 4374 12006 4403
rect 10318 4205 10352 4239
rect 10817 4283 10849 4287
rect 10849 4283 10851 4287
rect 10817 4253 10851 4283
rect 11881 4283 11883 4292
rect 11883 4283 11915 4292
rect 11881 4258 11915 4283
rect 10430 4124 10464 4158
rect 10725 4137 10759 4171
rect 10817 4137 10851 4171
rect 10909 4137 10943 4171
rect 11793 4137 11827 4171
rect 11885 4137 11919 4171
rect 11977 4137 12011 4171
rect 10286 4072 10320 4074
rect 10286 4040 10320 4072
rect 10286 3970 10320 4002
rect 10286 3968 10320 3970
rect 10382 4072 10416 4074
rect 10382 4040 10416 4072
rect 10382 3970 10416 4002
rect 10382 3968 10416 3970
rect 10478 4072 10512 4074
rect 10478 4040 10512 4072
rect 10478 3970 10512 4002
rect 10478 3968 10512 3970
rect 10334 3884 10368 3918
rect 10254 3775 10288 3809
rect 10684 3758 10718 3792
rect 9041 3635 9075 3669
rect 9133 3635 9167 3669
rect 9225 3635 9259 3669
rect 8164 3541 8198 3543
rect 8164 3509 8198 3541
rect 8164 3439 8198 3471
rect 8164 3437 8198 3439
rect 8252 3541 8286 3543
rect 8252 3509 8286 3541
rect 8810 3541 8844 3543
rect 8524 3477 8558 3511
rect 8810 3509 8844 3541
rect 8252 3439 8286 3471
rect 8252 3437 8286 3439
rect 8810 3439 8844 3471
rect 8810 3437 8844 3439
rect 8380 3381 8414 3383
rect 8380 3349 8414 3381
rect 8208 3309 8242 3343
rect 7499 3089 7533 3123
rect 7591 3089 7625 3123
rect 7683 3089 7717 3123
rect 8380 3279 8414 3311
rect 8380 3277 8414 3279
rect 8476 3381 8510 3383
rect 8476 3349 8510 3381
rect 8476 3279 8510 3311
rect 8476 3277 8510 3279
rect 9387 3633 9421 3667
rect 9479 3633 9513 3667
rect 9571 3633 9605 3667
rect 8898 3541 8932 3543
rect 8898 3509 8932 3541
rect 8898 3439 8932 3471
rect 8898 3437 8932 3439
rect 9733 3627 9767 3661
rect 9825 3627 9859 3661
rect 9917 3627 9951 3661
rect 10096 3637 10130 3671
rect 8572 3381 8606 3383
rect 8572 3349 8606 3381
rect 8572 3279 8606 3311
rect 8854 3309 8888 3343
rect 8572 3277 8606 3279
rect 9393 3321 9395 3354
rect 9395 3321 9427 3354
rect 9393 3320 9427 3321
rect 10742 3637 10776 3671
rect 9586 3332 9620 3366
rect 8428 3149 8462 3183
rect 7845 3083 7879 3117
rect 7937 3083 7971 3117
rect 8029 3083 8063 3117
rect 8180 3078 8214 3112
rect 8812 3106 8846 3140
rect 9172 3239 9206 3256
rect 9172 3222 9206 3239
rect 9782 3349 9816 3360
rect 9782 3326 9784 3349
rect 9784 3326 9816 3349
rect 4812 2914 4846 2946
rect 4812 2912 4846 2914
rect 6508 3016 6542 3018
rect 6508 2984 6542 3016
rect 6604 3016 6638 3018
rect 6604 2984 6638 3016
rect 6508 2914 6542 2946
rect 6508 2912 6542 2914
rect 6604 2914 6638 2946
rect 6604 2912 6638 2914
rect 6700 3016 6734 3018
rect 6700 2984 6734 3016
rect 8540 3068 8574 3102
rect 9041 3091 9075 3125
rect 9133 3091 9167 3125
rect 9225 3091 9259 3125
rect 10343 3585 10377 3619
rect 11764 3892 11798 3926
rect 12152 4437 12186 4439
rect 12152 4405 12186 4437
rect 12152 4335 12186 4367
rect 12152 4333 12186 4335
rect 12248 4437 12282 4439
rect 12248 4405 12282 4437
rect 12248 4335 12282 4367
rect 12248 4333 12282 4335
rect 14115 4641 14149 4675
rect 14184 4533 14218 4567
rect 12344 4437 12378 4439
rect 12344 4405 12378 4437
rect 12611 4403 12645 4410
rect 12611 4376 12615 4403
rect 12615 4376 12645 4403
rect 12344 4335 12378 4367
rect 12344 4333 12378 4335
rect 12785 4403 12819 4410
rect 12785 4376 12817 4403
rect 12817 4376 12819 4403
rect 13687 4403 13721 4412
rect 13687 4378 13689 4403
rect 13689 4378 13721 4403
rect 13860 4403 13894 4408
rect 13860 4374 13891 4403
rect 13891 4374 13894 4403
rect 12200 4205 12234 4239
rect 12699 4283 12731 4287
rect 12731 4283 12733 4287
rect 12699 4253 12733 4283
rect 13769 4283 13771 4292
rect 13771 4283 13803 4292
rect 13769 4258 13803 4283
rect 12312 4124 12346 4158
rect 12607 4137 12641 4171
rect 12699 4137 12733 4171
rect 12791 4137 12825 4171
rect 13681 4137 13715 4171
rect 13773 4137 13807 4171
rect 13865 4137 13899 4171
rect 12168 4072 12202 4074
rect 12168 4040 12202 4072
rect 12168 3970 12202 4002
rect 12168 3968 12202 3970
rect 12264 4072 12298 4074
rect 12264 4040 12298 4072
rect 12264 3970 12298 4002
rect 12264 3968 12298 3970
rect 12360 4072 12394 4074
rect 12360 4040 12394 4072
rect 12360 3970 12394 4002
rect 12360 3968 12394 3970
rect 12216 3884 12250 3918
rect 12136 3775 12170 3809
rect 12566 3758 12600 3792
rect 10929 3635 10963 3669
rect 11021 3635 11055 3669
rect 11113 3635 11147 3669
rect 10052 3541 10086 3543
rect 10052 3509 10086 3541
rect 10052 3439 10086 3471
rect 10052 3437 10086 3439
rect 10140 3541 10174 3543
rect 10140 3509 10174 3541
rect 10698 3541 10732 3543
rect 10412 3477 10446 3511
rect 10698 3509 10732 3541
rect 10140 3439 10174 3471
rect 10140 3437 10174 3439
rect 10698 3439 10732 3471
rect 10698 3437 10732 3439
rect 10268 3381 10302 3383
rect 10268 3349 10302 3381
rect 10096 3309 10130 3343
rect 9387 3089 9421 3123
rect 9479 3089 9513 3123
rect 9571 3089 9605 3123
rect 10268 3279 10302 3311
rect 10268 3277 10302 3279
rect 10364 3381 10398 3383
rect 10364 3349 10398 3381
rect 10364 3279 10398 3311
rect 10364 3277 10398 3279
rect 11275 3633 11309 3667
rect 11367 3633 11401 3667
rect 11459 3633 11493 3667
rect 10786 3541 10820 3543
rect 10786 3509 10820 3541
rect 10786 3439 10820 3471
rect 10786 3437 10820 3439
rect 11615 3627 11649 3661
rect 11707 3627 11741 3661
rect 11799 3627 11833 3661
rect 11978 3637 12012 3671
rect 10460 3381 10494 3383
rect 10460 3349 10494 3381
rect 10460 3279 10494 3311
rect 10742 3309 10776 3343
rect 10460 3277 10494 3279
rect 11281 3321 11283 3354
rect 11283 3321 11315 3354
rect 11281 3320 11315 3321
rect 12624 3637 12658 3671
rect 11474 3332 11508 3366
rect 10316 3149 10350 3183
rect 9733 3083 9767 3117
rect 9825 3083 9859 3117
rect 9917 3083 9951 3117
rect 10068 3078 10102 3112
rect 10700 3106 10734 3140
rect 11060 3239 11094 3256
rect 11060 3222 11094 3239
rect 11664 3349 11698 3360
rect 11664 3326 11666 3349
rect 11666 3326 11698 3349
rect 6700 2914 6734 2946
rect 6700 2912 6734 2914
rect 8396 3016 8430 3018
rect 8396 2984 8430 3016
rect 8492 3016 8526 3018
rect 8492 2984 8526 3016
rect 8396 2914 8430 2946
rect 8396 2912 8430 2914
rect 8492 2914 8526 2946
rect 8492 2912 8526 2914
rect 8588 3016 8622 3018
rect 8588 2984 8622 3016
rect 10428 3068 10462 3102
rect 10929 3091 10963 3125
rect 11021 3091 11055 3125
rect 11113 3091 11147 3125
rect 12225 3585 12259 3619
rect 13652 3892 13686 3926
rect 14040 4437 14074 4439
rect 14040 4405 14074 4437
rect 14040 4335 14074 4367
rect 14040 4333 14074 4335
rect 14136 4437 14170 4439
rect 14136 4405 14170 4437
rect 14136 4335 14170 4367
rect 14136 4333 14170 4335
rect 16003 4641 16037 4675
rect 16072 4533 16106 4567
rect 14232 4437 14266 4439
rect 14232 4405 14266 4437
rect 14499 4403 14533 4410
rect 14499 4376 14503 4403
rect 14503 4376 14533 4403
rect 14232 4335 14266 4367
rect 14232 4333 14266 4335
rect 14673 4403 14707 4410
rect 14673 4376 14705 4403
rect 14705 4376 14707 4403
rect 15575 4403 15609 4412
rect 15575 4378 15577 4403
rect 15577 4378 15609 4403
rect 15748 4403 15782 4408
rect 15748 4374 15779 4403
rect 15779 4374 15782 4403
rect 14088 4205 14122 4239
rect 14587 4283 14619 4287
rect 14619 4283 14621 4287
rect 14587 4253 14621 4283
rect 15657 4283 15659 4292
rect 15659 4283 15691 4292
rect 15657 4258 15691 4283
rect 14200 4124 14234 4158
rect 14495 4137 14529 4171
rect 14587 4137 14621 4171
rect 14679 4137 14713 4171
rect 15569 4137 15603 4171
rect 15661 4137 15695 4171
rect 15753 4137 15787 4171
rect 14056 4072 14090 4074
rect 14056 4040 14090 4072
rect 14056 3970 14090 4002
rect 14056 3968 14090 3970
rect 14152 4072 14186 4074
rect 14152 4040 14186 4072
rect 14152 3970 14186 4002
rect 14152 3968 14186 3970
rect 14248 4072 14282 4074
rect 14248 4040 14282 4072
rect 14248 3970 14282 4002
rect 14248 3968 14282 3970
rect 14104 3884 14138 3918
rect 14024 3775 14058 3809
rect 14454 3758 14488 3792
rect 12811 3635 12845 3669
rect 12903 3635 12937 3669
rect 12995 3635 13029 3669
rect 11934 3541 11968 3543
rect 11934 3509 11968 3541
rect 11934 3439 11968 3471
rect 11934 3437 11968 3439
rect 12022 3541 12056 3543
rect 12022 3509 12056 3541
rect 12580 3541 12614 3543
rect 12294 3477 12328 3511
rect 12580 3509 12614 3541
rect 12022 3439 12056 3471
rect 12022 3437 12056 3439
rect 12580 3439 12614 3471
rect 12580 3437 12614 3439
rect 12150 3381 12184 3383
rect 12150 3349 12184 3381
rect 11978 3309 12012 3343
rect 11275 3089 11309 3123
rect 11367 3089 11401 3123
rect 11459 3089 11493 3123
rect 12150 3279 12184 3311
rect 12150 3277 12184 3279
rect 12246 3381 12280 3383
rect 12246 3349 12280 3381
rect 12246 3279 12280 3311
rect 12246 3277 12280 3279
rect 13157 3633 13191 3667
rect 13249 3633 13283 3667
rect 13341 3633 13375 3667
rect 12668 3541 12702 3543
rect 12668 3509 12702 3541
rect 12668 3439 12702 3471
rect 12668 3437 12702 3439
rect 13503 3627 13537 3661
rect 13595 3627 13629 3661
rect 13687 3627 13721 3661
rect 13866 3637 13900 3671
rect 12342 3381 12376 3383
rect 12342 3349 12376 3381
rect 12342 3279 12376 3311
rect 12624 3309 12658 3343
rect 12342 3277 12376 3279
rect 13163 3321 13165 3354
rect 13165 3321 13197 3354
rect 13163 3320 13197 3321
rect 14512 3637 14546 3671
rect 13356 3332 13390 3366
rect 12198 3149 12232 3183
rect 11615 3083 11649 3117
rect 11707 3083 11741 3117
rect 11799 3083 11833 3117
rect 11950 3078 11984 3112
rect 12582 3106 12616 3140
rect 12942 3239 12976 3256
rect 12942 3222 12976 3239
rect 13552 3349 13586 3360
rect 13552 3326 13554 3349
rect 13554 3326 13586 3349
rect 8588 2914 8622 2946
rect 8588 2912 8622 2914
rect 10284 3016 10318 3018
rect 10284 2984 10318 3016
rect 10380 3016 10414 3018
rect 10380 2984 10414 3016
rect 10284 2914 10318 2946
rect 10284 2912 10318 2914
rect 10380 2914 10414 2946
rect 10380 2912 10414 2914
rect 10476 3016 10510 3018
rect 10476 2984 10510 3016
rect 12310 3068 12344 3102
rect 12811 3091 12845 3125
rect 12903 3091 12937 3125
rect 12995 3091 13029 3125
rect 14113 3585 14147 3619
rect 15540 3892 15574 3926
rect 15928 4437 15962 4439
rect 15928 4405 15962 4437
rect 15928 4335 15962 4367
rect 15928 4333 15962 4335
rect 16024 4437 16058 4439
rect 16024 4405 16058 4437
rect 16024 4335 16058 4367
rect 16024 4333 16058 4335
rect 17891 4641 17925 4675
rect 17960 4533 17994 4567
rect 16120 4437 16154 4439
rect 16120 4405 16154 4437
rect 16387 4403 16421 4410
rect 16387 4376 16391 4403
rect 16391 4376 16421 4403
rect 16120 4335 16154 4367
rect 16120 4333 16154 4335
rect 16561 4403 16595 4410
rect 16561 4376 16593 4403
rect 16593 4376 16595 4403
rect 17463 4403 17497 4412
rect 17463 4378 17465 4403
rect 17465 4378 17497 4403
rect 17636 4403 17670 4408
rect 17636 4374 17667 4403
rect 17667 4374 17670 4403
rect 15976 4205 16010 4239
rect 16475 4283 16507 4287
rect 16507 4283 16509 4287
rect 16475 4253 16509 4283
rect 17545 4283 17547 4292
rect 17547 4283 17579 4292
rect 17545 4258 17579 4283
rect 16088 4124 16122 4158
rect 16383 4137 16417 4171
rect 16475 4137 16509 4171
rect 16567 4137 16601 4171
rect 17457 4137 17491 4171
rect 17549 4137 17583 4171
rect 17641 4137 17675 4171
rect 15944 4072 15978 4074
rect 15944 4040 15978 4072
rect 15944 3970 15978 4002
rect 15944 3968 15978 3970
rect 16040 4072 16074 4074
rect 16040 4040 16074 4072
rect 16040 3970 16074 4002
rect 16040 3968 16074 3970
rect 16136 4072 16170 4074
rect 16136 4040 16170 4072
rect 16136 3970 16170 4002
rect 16136 3968 16170 3970
rect 15992 3884 16026 3918
rect 15912 3775 15946 3809
rect 16342 3758 16376 3792
rect 14699 3635 14733 3669
rect 14791 3635 14825 3669
rect 14883 3635 14917 3669
rect 13822 3541 13856 3543
rect 13822 3509 13856 3541
rect 13822 3439 13856 3471
rect 13822 3437 13856 3439
rect 13910 3541 13944 3543
rect 13910 3509 13944 3541
rect 14468 3541 14502 3543
rect 14182 3477 14216 3511
rect 14468 3509 14502 3541
rect 13910 3439 13944 3471
rect 13910 3437 13944 3439
rect 14468 3439 14502 3471
rect 14468 3437 14502 3439
rect 14038 3381 14072 3383
rect 14038 3349 14072 3381
rect 13866 3309 13900 3343
rect 13157 3089 13191 3123
rect 13249 3089 13283 3123
rect 13341 3089 13375 3123
rect 14038 3279 14072 3311
rect 14038 3277 14072 3279
rect 14134 3381 14168 3383
rect 14134 3349 14168 3381
rect 14134 3279 14168 3311
rect 14134 3277 14168 3279
rect 15045 3633 15079 3667
rect 15137 3633 15171 3667
rect 15229 3633 15263 3667
rect 14556 3541 14590 3543
rect 14556 3509 14590 3541
rect 14556 3439 14590 3471
rect 14556 3437 14590 3439
rect 15391 3627 15425 3661
rect 15483 3627 15517 3661
rect 15575 3627 15609 3661
rect 15754 3637 15788 3671
rect 14230 3381 14264 3383
rect 14230 3349 14264 3381
rect 14230 3279 14264 3311
rect 14512 3309 14546 3343
rect 14230 3277 14264 3279
rect 15051 3321 15053 3354
rect 15053 3321 15085 3354
rect 15051 3320 15085 3321
rect 16400 3637 16434 3671
rect 15244 3332 15278 3366
rect 14086 3149 14120 3183
rect 13503 3083 13537 3117
rect 13595 3083 13629 3117
rect 13687 3083 13721 3117
rect 13838 3078 13872 3112
rect 14470 3106 14504 3140
rect 14830 3239 14864 3256
rect 14830 3222 14864 3239
rect 15440 3349 15474 3360
rect 15440 3326 15442 3349
rect 15442 3326 15474 3349
rect 10476 2914 10510 2946
rect 10476 2912 10510 2914
rect 12166 3016 12200 3018
rect 12166 2984 12200 3016
rect 12262 3016 12296 3018
rect 12262 2984 12296 3016
rect 12166 2914 12200 2946
rect 12166 2912 12200 2914
rect 12262 2914 12296 2946
rect 12262 2912 12296 2914
rect 12358 3016 12392 3018
rect 12358 2984 12392 3016
rect 14198 3068 14232 3102
rect 14699 3091 14733 3125
rect 14791 3091 14825 3125
rect 14883 3091 14917 3125
rect 16001 3585 16035 3619
rect 17428 3892 17462 3926
rect 17816 4437 17850 4439
rect 17816 4405 17850 4437
rect 17816 4335 17850 4367
rect 17816 4333 17850 4335
rect 17912 4437 17946 4439
rect 17912 4405 17946 4437
rect 17912 4335 17946 4367
rect 17912 4333 17946 4335
rect 19779 4641 19813 4675
rect 19848 4533 19882 4567
rect 18008 4437 18042 4439
rect 18008 4405 18042 4437
rect 18275 4403 18309 4410
rect 18275 4376 18279 4403
rect 18279 4376 18309 4403
rect 18008 4335 18042 4367
rect 18008 4333 18042 4335
rect 18449 4403 18483 4410
rect 18449 4376 18481 4403
rect 18481 4376 18483 4403
rect 19351 4403 19385 4412
rect 19351 4378 19353 4403
rect 19353 4378 19385 4403
rect 19524 4403 19558 4408
rect 19524 4374 19555 4403
rect 19555 4374 19558 4403
rect 17864 4205 17898 4239
rect 18363 4283 18395 4287
rect 18395 4283 18397 4287
rect 18363 4253 18397 4283
rect 19433 4283 19435 4292
rect 19435 4283 19467 4292
rect 19433 4258 19467 4283
rect 17976 4124 18010 4158
rect 18271 4137 18305 4171
rect 18363 4137 18397 4171
rect 18455 4137 18489 4171
rect 19345 4137 19379 4171
rect 19437 4137 19471 4171
rect 19529 4137 19563 4171
rect 17832 4072 17866 4074
rect 17832 4040 17866 4072
rect 17832 3970 17866 4002
rect 17832 3968 17866 3970
rect 17928 4072 17962 4074
rect 17928 4040 17962 4072
rect 17928 3970 17962 4002
rect 17928 3968 17962 3970
rect 18024 4072 18058 4074
rect 18024 4040 18058 4072
rect 18024 3970 18058 4002
rect 18024 3968 18058 3970
rect 17880 3884 17914 3918
rect 17800 3775 17834 3809
rect 18230 3758 18264 3792
rect 16587 3635 16621 3669
rect 16679 3635 16713 3669
rect 16771 3635 16805 3669
rect 15710 3541 15744 3543
rect 15710 3509 15744 3541
rect 15710 3439 15744 3471
rect 15710 3437 15744 3439
rect 15798 3541 15832 3543
rect 15798 3509 15832 3541
rect 16356 3541 16390 3543
rect 16070 3477 16104 3511
rect 16356 3509 16390 3541
rect 15798 3439 15832 3471
rect 15798 3437 15832 3439
rect 16356 3439 16390 3471
rect 16356 3437 16390 3439
rect 15926 3381 15960 3383
rect 15926 3349 15960 3381
rect 15754 3309 15788 3343
rect 15045 3089 15079 3123
rect 15137 3089 15171 3123
rect 15229 3089 15263 3123
rect 15926 3279 15960 3311
rect 15926 3277 15960 3279
rect 16022 3381 16056 3383
rect 16022 3349 16056 3381
rect 16022 3279 16056 3311
rect 16022 3277 16056 3279
rect 16933 3633 16967 3667
rect 17025 3633 17059 3667
rect 17117 3633 17151 3667
rect 16444 3541 16478 3543
rect 16444 3509 16478 3541
rect 16444 3439 16478 3471
rect 16444 3437 16478 3439
rect 17279 3627 17313 3661
rect 17371 3627 17405 3661
rect 17463 3627 17497 3661
rect 17642 3637 17676 3671
rect 16118 3381 16152 3383
rect 16118 3349 16152 3381
rect 16118 3279 16152 3311
rect 16400 3309 16434 3343
rect 16118 3277 16152 3279
rect 16939 3321 16941 3354
rect 16941 3321 16973 3354
rect 16939 3320 16973 3321
rect 18288 3637 18322 3671
rect 17132 3332 17166 3366
rect 15974 3149 16008 3183
rect 15391 3083 15425 3117
rect 15483 3083 15517 3117
rect 15575 3083 15609 3117
rect 15726 3078 15760 3112
rect 16358 3106 16392 3140
rect 16718 3239 16752 3256
rect 16718 3222 16752 3239
rect 17328 3349 17362 3360
rect 17328 3326 17330 3349
rect 17330 3326 17362 3349
rect 12358 2914 12392 2946
rect 12358 2912 12392 2914
rect 14054 3016 14088 3018
rect 14054 2984 14088 3016
rect 14150 3016 14184 3018
rect 14150 2984 14184 3016
rect 14054 2914 14088 2946
rect 14054 2912 14088 2914
rect 14150 2914 14184 2946
rect 14150 2912 14184 2914
rect 14246 3016 14280 3018
rect 14246 2984 14280 3016
rect 16086 3068 16120 3102
rect 16587 3091 16621 3125
rect 16679 3091 16713 3125
rect 16771 3091 16805 3125
rect 17889 3585 17923 3619
rect 19316 3892 19350 3926
rect 19704 4437 19738 4439
rect 19704 4405 19738 4437
rect 19704 4335 19738 4367
rect 19704 4333 19738 4335
rect 19800 4437 19834 4439
rect 19800 4405 19834 4437
rect 19800 4335 19834 4367
rect 19800 4333 19834 4335
rect 21667 4641 21701 4675
rect 21736 4533 21770 4567
rect 19896 4437 19930 4439
rect 19896 4405 19930 4437
rect 20163 4403 20197 4410
rect 20163 4376 20167 4403
rect 20167 4376 20197 4403
rect 19896 4335 19930 4367
rect 19896 4333 19930 4335
rect 20337 4403 20371 4410
rect 20337 4376 20369 4403
rect 20369 4376 20371 4403
rect 21239 4403 21273 4412
rect 21239 4378 21241 4403
rect 21241 4378 21273 4403
rect 21412 4403 21446 4408
rect 21412 4374 21443 4403
rect 21443 4374 21446 4403
rect 19752 4205 19786 4239
rect 20251 4283 20283 4287
rect 20283 4283 20285 4287
rect 20251 4253 20285 4283
rect 21321 4283 21323 4292
rect 21323 4283 21355 4292
rect 21321 4258 21355 4283
rect 19864 4124 19898 4158
rect 20159 4137 20193 4171
rect 20251 4137 20285 4171
rect 20343 4137 20377 4171
rect 21233 4137 21267 4171
rect 21325 4137 21359 4171
rect 21417 4137 21451 4171
rect 19720 4072 19754 4074
rect 19720 4040 19754 4072
rect 19720 3970 19754 4002
rect 19720 3968 19754 3970
rect 19816 4072 19850 4074
rect 19816 4040 19850 4072
rect 19816 3970 19850 4002
rect 19816 3968 19850 3970
rect 19912 4072 19946 4074
rect 19912 4040 19946 4072
rect 19912 3970 19946 4002
rect 19912 3968 19946 3970
rect 19768 3884 19802 3918
rect 19688 3775 19722 3809
rect 20118 3758 20152 3792
rect 18475 3635 18509 3669
rect 18567 3635 18601 3669
rect 18659 3635 18693 3669
rect 17598 3541 17632 3543
rect 17598 3509 17632 3541
rect 17598 3439 17632 3471
rect 17598 3437 17632 3439
rect 17686 3541 17720 3543
rect 17686 3509 17720 3541
rect 18244 3541 18278 3543
rect 17958 3477 17992 3511
rect 18244 3509 18278 3541
rect 17686 3439 17720 3471
rect 17686 3437 17720 3439
rect 18244 3439 18278 3471
rect 18244 3437 18278 3439
rect 17814 3381 17848 3383
rect 17814 3349 17848 3381
rect 17642 3309 17676 3343
rect 16933 3089 16967 3123
rect 17025 3089 17059 3123
rect 17117 3089 17151 3123
rect 17814 3279 17848 3311
rect 17814 3277 17848 3279
rect 17910 3381 17944 3383
rect 17910 3349 17944 3381
rect 17910 3279 17944 3311
rect 17910 3277 17944 3279
rect 18821 3633 18855 3667
rect 18913 3633 18947 3667
rect 19005 3633 19039 3667
rect 18332 3541 18366 3543
rect 18332 3509 18366 3541
rect 18332 3439 18366 3471
rect 18332 3437 18366 3439
rect 19167 3627 19201 3661
rect 19259 3627 19293 3661
rect 19351 3627 19385 3661
rect 19530 3637 19564 3671
rect 18006 3381 18040 3383
rect 18006 3349 18040 3381
rect 18006 3279 18040 3311
rect 18288 3309 18322 3343
rect 18006 3277 18040 3279
rect 18827 3321 18829 3354
rect 18829 3321 18861 3354
rect 18827 3320 18861 3321
rect 20176 3637 20210 3671
rect 19020 3332 19054 3366
rect 17862 3149 17896 3183
rect 17279 3083 17313 3117
rect 17371 3083 17405 3117
rect 17463 3083 17497 3117
rect 17614 3078 17648 3112
rect 18246 3106 18280 3140
rect 18606 3239 18640 3256
rect 18606 3222 18640 3239
rect 19216 3349 19250 3360
rect 19216 3326 19218 3349
rect 19218 3326 19250 3349
rect 14246 2914 14280 2946
rect 14246 2912 14280 2914
rect 15942 3016 15976 3018
rect 15942 2984 15976 3016
rect 16038 3016 16072 3018
rect 16038 2984 16072 3016
rect 15942 2914 15976 2946
rect 15942 2912 15976 2914
rect 16038 2914 16072 2946
rect 16038 2912 16072 2914
rect 16134 3016 16168 3018
rect 16134 2984 16168 3016
rect 17974 3068 18008 3102
rect 18475 3091 18509 3125
rect 18567 3091 18601 3125
rect 18659 3091 18693 3125
rect 19777 3585 19811 3619
rect 21204 3892 21238 3926
rect 21592 4437 21626 4439
rect 21592 4405 21626 4437
rect 21592 4335 21626 4367
rect 21592 4333 21626 4335
rect 21688 4437 21722 4439
rect 21688 4405 21722 4437
rect 21688 4335 21722 4367
rect 21688 4333 21722 4335
rect 23555 4641 23589 4675
rect 23624 4533 23658 4567
rect 21784 4437 21818 4439
rect 21784 4405 21818 4437
rect 22051 4403 22085 4410
rect 22051 4376 22055 4403
rect 22055 4376 22085 4403
rect 21784 4335 21818 4367
rect 21784 4333 21818 4335
rect 22225 4403 22259 4410
rect 22225 4376 22257 4403
rect 22257 4376 22259 4403
rect 23127 4403 23161 4412
rect 23127 4378 23129 4403
rect 23129 4378 23161 4403
rect 23300 4403 23334 4408
rect 23300 4374 23331 4403
rect 23331 4374 23334 4403
rect 21640 4205 21674 4239
rect 22139 4283 22171 4287
rect 22171 4283 22173 4287
rect 22139 4253 22173 4283
rect 23209 4283 23211 4292
rect 23211 4283 23243 4292
rect 23209 4258 23243 4283
rect 21752 4124 21786 4158
rect 22047 4137 22081 4171
rect 22139 4137 22173 4171
rect 22231 4137 22265 4171
rect 23121 4137 23155 4171
rect 23213 4137 23247 4171
rect 23305 4137 23339 4171
rect 21608 4072 21642 4074
rect 21608 4040 21642 4072
rect 21608 3970 21642 4002
rect 21608 3968 21642 3970
rect 21704 4072 21738 4074
rect 21704 4040 21738 4072
rect 21704 3970 21738 4002
rect 21704 3968 21738 3970
rect 21800 4072 21834 4074
rect 21800 4040 21834 4072
rect 21800 3970 21834 4002
rect 21800 3968 21834 3970
rect 21656 3884 21690 3918
rect 21576 3775 21610 3809
rect 22006 3758 22040 3792
rect 20363 3635 20397 3669
rect 20455 3635 20489 3669
rect 20547 3635 20581 3669
rect 19486 3541 19520 3543
rect 19486 3509 19520 3541
rect 19486 3439 19520 3471
rect 19486 3437 19520 3439
rect 19574 3541 19608 3543
rect 19574 3509 19608 3541
rect 20132 3541 20166 3543
rect 19846 3477 19880 3511
rect 20132 3509 20166 3541
rect 19574 3439 19608 3471
rect 19574 3437 19608 3439
rect 20132 3439 20166 3471
rect 20132 3437 20166 3439
rect 19702 3381 19736 3383
rect 19702 3349 19736 3381
rect 19530 3309 19564 3343
rect 18821 3089 18855 3123
rect 18913 3089 18947 3123
rect 19005 3089 19039 3123
rect 19702 3279 19736 3311
rect 19702 3277 19736 3279
rect 19798 3381 19832 3383
rect 19798 3349 19832 3381
rect 19798 3279 19832 3311
rect 19798 3277 19832 3279
rect 20709 3633 20743 3667
rect 20801 3633 20835 3667
rect 20893 3633 20927 3667
rect 20220 3541 20254 3543
rect 20220 3509 20254 3541
rect 20220 3439 20254 3471
rect 20220 3437 20254 3439
rect 21055 3627 21089 3661
rect 21147 3627 21181 3661
rect 21239 3627 21273 3661
rect 21418 3637 21452 3671
rect 19894 3381 19928 3383
rect 19894 3349 19928 3381
rect 19894 3279 19928 3311
rect 20176 3309 20210 3343
rect 19894 3277 19928 3279
rect 20715 3321 20717 3354
rect 20717 3321 20749 3354
rect 20715 3320 20749 3321
rect 22064 3637 22098 3671
rect 20908 3332 20942 3366
rect 19750 3149 19784 3183
rect 19167 3083 19201 3117
rect 19259 3083 19293 3117
rect 19351 3083 19385 3117
rect 19502 3078 19536 3112
rect 20134 3106 20168 3140
rect 20494 3239 20528 3256
rect 20494 3222 20528 3239
rect 21104 3349 21138 3360
rect 21104 3326 21106 3349
rect 21106 3326 21138 3349
rect 16134 2914 16168 2946
rect 16134 2912 16168 2914
rect 17830 3016 17864 3018
rect 17830 2984 17864 3016
rect 17926 3016 17960 3018
rect 17926 2984 17960 3016
rect 17830 2914 17864 2946
rect 17830 2912 17864 2914
rect 17926 2914 17960 2946
rect 17926 2912 17960 2914
rect 18022 3016 18056 3018
rect 18022 2984 18056 3016
rect 19862 3068 19896 3102
rect 20363 3091 20397 3125
rect 20455 3091 20489 3125
rect 20547 3091 20581 3125
rect 21665 3585 21699 3619
rect 23092 3892 23126 3926
rect 23480 4437 23514 4439
rect 23480 4405 23514 4437
rect 23480 4335 23514 4367
rect 23480 4333 23514 4335
rect 23576 4437 23610 4439
rect 23576 4405 23610 4437
rect 23576 4335 23610 4367
rect 23576 4333 23610 4335
rect 25443 4641 25477 4675
rect 25512 4533 25546 4567
rect 23672 4437 23706 4439
rect 23672 4405 23706 4437
rect 23939 4403 23973 4410
rect 23939 4376 23943 4403
rect 23943 4376 23973 4403
rect 23672 4335 23706 4367
rect 23672 4333 23706 4335
rect 24113 4403 24147 4410
rect 24113 4376 24145 4403
rect 24145 4376 24147 4403
rect 25015 4403 25049 4412
rect 25015 4378 25017 4403
rect 25017 4378 25049 4403
rect 25188 4403 25222 4408
rect 25188 4374 25219 4403
rect 25219 4374 25222 4403
rect 23528 4205 23562 4239
rect 24027 4283 24059 4287
rect 24059 4283 24061 4287
rect 24027 4253 24061 4283
rect 25097 4283 25099 4292
rect 25099 4283 25131 4292
rect 25097 4258 25131 4283
rect 23640 4124 23674 4158
rect 23935 4137 23969 4171
rect 24027 4137 24061 4171
rect 24119 4137 24153 4171
rect 25009 4137 25043 4171
rect 25101 4137 25135 4171
rect 25193 4137 25227 4171
rect 23496 4072 23530 4074
rect 23496 4040 23530 4072
rect 23496 3970 23530 4002
rect 23496 3968 23530 3970
rect 23592 4072 23626 4074
rect 23592 4040 23626 4072
rect 23592 3970 23626 4002
rect 23592 3968 23626 3970
rect 23688 4072 23722 4074
rect 23688 4040 23722 4072
rect 23688 3970 23722 4002
rect 23688 3968 23722 3970
rect 23544 3884 23578 3918
rect 23464 3775 23498 3809
rect 23894 3758 23928 3792
rect 22251 3635 22285 3669
rect 22343 3635 22377 3669
rect 22435 3635 22469 3669
rect 21374 3541 21408 3543
rect 21374 3509 21408 3541
rect 21374 3439 21408 3471
rect 21374 3437 21408 3439
rect 21462 3541 21496 3543
rect 21462 3509 21496 3541
rect 22020 3541 22054 3543
rect 21734 3477 21768 3511
rect 22020 3509 22054 3541
rect 21462 3439 21496 3471
rect 21462 3437 21496 3439
rect 22020 3439 22054 3471
rect 22020 3437 22054 3439
rect 21590 3381 21624 3383
rect 21590 3349 21624 3381
rect 21418 3309 21452 3343
rect 20709 3089 20743 3123
rect 20801 3089 20835 3123
rect 20893 3089 20927 3123
rect 21590 3279 21624 3311
rect 21590 3277 21624 3279
rect 21686 3381 21720 3383
rect 21686 3349 21720 3381
rect 21686 3279 21720 3311
rect 21686 3277 21720 3279
rect 22597 3633 22631 3667
rect 22689 3633 22723 3667
rect 22781 3633 22815 3667
rect 22108 3541 22142 3543
rect 22108 3509 22142 3541
rect 22108 3439 22142 3471
rect 22108 3437 22142 3439
rect 22943 3627 22977 3661
rect 23035 3627 23069 3661
rect 23127 3627 23161 3661
rect 23306 3637 23340 3671
rect 21782 3381 21816 3383
rect 21782 3349 21816 3381
rect 21782 3279 21816 3311
rect 22064 3309 22098 3343
rect 21782 3277 21816 3279
rect 22603 3321 22605 3354
rect 22605 3321 22637 3354
rect 22603 3320 22637 3321
rect 23952 3637 23986 3671
rect 22796 3332 22830 3366
rect 21638 3149 21672 3183
rect 21055 3083 21089 3117
rect 21147 3083 21181 3117
rect 21239 3083 21273 3117
rect 21390 3078 21424 3112
rect 22022 3106 22056 3140
rect 22382 3239 22416 3256
rect 22382 3222 22416 3239
rect 22992 3349 23026 3360
rect 22992 3326 22994 3349
rect 22994 3326 23026 3349
rect 18022 2914 18056 2946
rect 18022 2912 18056 2914
rect 19718 3016 19752 3018
rect 19718 2984 19752 3016
rect 19814 3016 19848 3018
rect 19814 2984 19848 3016
rect 19718 2914 19752 2946
rect 19718 2912 19752 2914
rect 19814 2914 19848 2946
rect 19814 2912 19848 2914
rect 19910 3016 19944 3018
rect 19910 2984 19944 3016
rect 21750 3068 21784 3102
rect 22251 3091 22285 3125
rect 22343 3091 22377 3125
rect 22435 3091 22469 3125
rect 23553 3585 23587 3619
rect 24980 3892 25014 3926
rect 25368 4437 25402 4439
rect 25368 4405 25402 4437
rect 25368 4335 25402 4367
rect 25368 4333 25402 4335
rect 25464 4437 25498 4439
rect 25464 4405 25498 4437
rect 25464 4335 25498 4367
rect 25464 4333 25498 4335
rect 25560 4437 25594 4439
rect 25560 4405 25594 4437
rect 25827 4403 25861 4410
rect 25827 4376 25831 4403
rect 25831 4376 25861 4403
rect 25560 4335 25594 4367
rect 25560 4333 25594 4335
rect 26001 4403 26035 4410
rect 26001 4376 26033 4403
rect 26033 4376 26035 4403
rect 25416 4205 25450 4239
rect 25915 4283 25947 4287
rect 25947 4283 25949 4287
rect 25915 4253 25949 4283
rect 25528 4124 25562 4158
rect 25823 4137 25857 4171
rect 25915 4137 25949 4171
rect 26007 4137 26041 4171
rect 25384 4072 25418 4074
rect 25384 4040 25418 4072
rect 25384 3970 25418 4002
rect 25384 3968 25418 3970
rect 25480 4072 25514 4074
rect 25480 4040 25514 4072
rect 25480 3970 25514 4002
rect 25480 3968 25514 3970
rect 25576 4072 25610 4074
rect 25576 4040 25610 4072
rect 25576 3970 25610 4002
rect 25576 3968 25610 3970
rect 25432 3884 25466 3918
rect 25352 3775 25386 3809
rect 25782 3758 25816 3792
rect 24139 3635 24173 3669
rect 24231 3635 24265 3669
rect 24323 3635 24357 3669
rect 23262 3541 23296 3543
rect 23262 3509 23296 3541
rect 23262 3439 23296 3471
rect 23262 3437 23296 3439
rect 23350 3541 23384 3543
rect 23350 3509 23384 3541
rect 23908 3541 23942 3543
rect 23622 3477 23656 3511
rect 23908 3509 23942 3541
rect 23350 3439 23384 3471
rect 23350 3437 23384 3439
rect 23908 3439 23942 3471
rect 23908 3437 23942 3439
rect 23478 3381 23512 3383
rect 23478 3349 23512 3381
rect 23306 3309 23340 3343
rect 22597 3089 22631 3123
rect 22689 3089 22723 3123
rect 22781 3089 22815 3123
rect 23478 3279 23512 3311
rect 23478 3277 23512 3279
rect 23574 3381 23608 3383
rect 23574 3349 23608 3381
rect 23574 3279 23608 3311
rect 23574 3277 23608 3279
rect 24485 3633 24519 3667
rect 24577 3633 24611 3667
rect 24669 3633 24703 3667
rect 23996 3541 24030 3543
rect 23996 3509 24030 3541
rect 23996 3439 24030 3471
rect 23996 3437 24030 3439
rect 24831 3627 24865 3661
rect 24923 3627 24957 3661
rect 25015 3627 25049 3661
rect 25194 3637 25228 3671
rect 23670 3381 23704 3383
rect 23670 3349 23704 3381
rect 23670 3279 23704 3311
rect 23952 3309 23986 3343
rect 23670 3277 23704 3279
rect 24491 3321 24493 3354
rect 24493 3321 24525 3354
rect 24491 3320 24525 3321
rect 25840 3637 25874 3671
rect 24684 3332 24718 3366
rect 23526 3149 23560 3183
rect 22943 3083 22977 3117
rect 23035 3083 23069 3117
rect 23127 3083 23161 3117
rect 23278 3078 23312 3112
rect 23910 3106 23944 3140
rect 24270 3239 24304 3256
rect 24270 3222 24304 3239
rect 24880 3349 24914 3360
rect 24880 3326 24882 3349
rect 24882 3326 24914 3349
rect 19910 2914 19944 2946
rect 19910 2912 19944 2914
rect 21606 3016 21640 3018
rect 21606 2984 21640 3016
rect 21702 3016 21736 3018
rect 21702 2984 21736 3016
rect 21606 2914 21640 2946
rect 21606 2912 21640 2914
rect 21702 2914 21736 2946
rect 21702 2912 21736 2914
rect 21798 3016 21832 3018
rect 21798 2984 21832 3016
rect 23638 3068 23672 3102
rect 24139 3091 24173 3125
rect 24231 3091 24265 3125
rect 24323 3091 24357 3125
rect 25441 3585 25475 3619
rect 26027 3635 26061 3669
rect 26119 3635 26153 3669
rect 26211 3635 26245 3669
rect 25150 3541 25184 3543
rect 25150 3509 25184 3541
rect 25150 3439 25184 3471
rect 25150 3437 25184 3439
rect 25238 3541 25272 3543
rect 25238 3509 25272 3541
rect 25796 3541 25830 3543
rect 25510 3477 25544 3511
rect 25796 3509 25830 3541
rect 25238 3439 25272 3471
rect 25238 3437 25272 3439
rect 25796 3439 25830 3471
rect 25796 3437 25830 3439
rect 25366 3381 25400 3383
rect 25366 3349 25400 3381
rect 25194 3309 25228 3343
rect 24485 3089 24519 3123
rect 24577 3089 24611 3123
rect 24669 3089 24703 3123
rect 25366 3279 25400 3311
rect 25366 3277 25400 3279
rect 25462 3381 25496 3383
rect 25462 3349 25496 3381
rect 25462 3279 25496 3311
rect 25462 3277 25496 3279
rect 26373 3633 26407 3667
rect 26465 3633 26499 3667
rect 26557 3633 26591 3667
rect 25884 3541 25918 3543
rect 25884 3509 25918 3541
rect 25884 3439 25918 3471
rect 25884 3437 25918 3439
rect 25558 3381 25592 3383
rect 25558 3349 25592 3381
rect 25558 3279 25592 3311
rect 25840 3309 25874 3343
rect 25558 3277 25592 3279
rect 26379 3321 26381 3354
rect 26381 3321 26413 3354
rect 26379 3320 26413 3321
rect 26572 3332 26606 3366
rect 25414 3149 25448 3183
rect 24831 3083 24865 3117
rect 24923 3083 24957 3117
rect 25015 3083 25049 3117
rect 25166 3078 25200 3112
rect 25798 3106 25832 3140
rect 26158 3239 26192 3256
rect 26158 3222 26192 3239
rect 21798 2914 21832 2946
rect 21798 2912 21832 2914
rect 23494 3016 23528 3018
rect 23494 2984 23528 3016
rect 23590 3016 23624 3018
rect 23590 2984 23624 3016
rect 23494 2914 23528 2946
rect 23494 2912 23528 2914
rect 23590 2914 23624 2946
rect 23590 2912 23624 2914
rect 23686 3016 23720 3018
rect 23686 2984 23720 3016
rect 25526 3068 25560 3102
rect 26027 3091 26061 3125
rect 26119 3091 26153 3125
rect 26211 3091 26245 3125
rect 26373 3089 26407 3123
rect 26465 3089 26499 3123
rect 26557 3089 26591 3123
rect 23686 2914 23720 2946
rect 23686 2912 23720 2914
rect 25382 3016 25416 3018
rect 25382 2984 25416 3016
rect 25478 3016 25512 3018
rect 25478 2984 25512 3016
rect 25382 2914 25416 2946
rect 25382 2912 25416 2914
rect 25478 2914 25512 2946
rect 25478 2912 25512 2914
rect 25574 3016 25608 3018
rect 25574 2984 25608 3016
rect 25574 2914 25608 2946
rect 25574 2912 25608 2914
rect -2884 2828 -2850 2862
rect -996 2828 -962 2862
rect 892 2828 926 2862
rect 2780 2828 2814 2862
rect 4668 2828 4702 2862
rect 6556 2828 6590 2862
rect 8444 2828 8478 2862
rect 10332 2828 10366 2862
rect 12214 2828 12248 2862
rect 14102 2828 14136 2862
rect 15990 2828 16024 2862
rect 17878 2828 17912 2862
rect 19766 2828 19800 2862
rect 21654 2828 21688 2862
rect 23542 2828 23576 2862
rect 25430 2828 25464 2862
rect -2964 2719 -2930 2753
rect -1076 2719 -1042 2753
rect 812 2719 846 2753
rect 2700 2719 2734 2753
rect 4588 2719 4622 2753
rect 6476 2719 6510 2753
rect 8364 2719 8398 2753
rect 10252 2719 10286 2753
rect 12134 2719 12168 2753
rect 14022 2719 14056 2753
rect 15910 2719 15944 2753
rect 17798 2719 17832 2753
rect 19686 2719 19720 2753
rect 21574 2719 21608 2753
rect 23462 2719 23496 2753
rect 25350 2719 25384 2753
<< metal1 >>
rect 2112 5367 3584 5370
rect 3994 5367 5466 5368
rect 2112 5343 5466 5367
rect 2112 5339 4610 5343
rect 2112 5305 2141 5339
rect 2175 5305 2233 5339
rect 2267 5305 2325 5339
rect 2359 5305 2417 5339
rect 2451 5305 2509 5339
rect 2543 5305 2601 5339
rect 2635 5305 2693 5339
rect 2727 5305 2785 5339
rect 2819 5305 2877 5339
rect 2911 5305 2969 5339
rect 3003 5305 3061 5339
rect 3095 5305 3153 5339
rect 3187 5305 3245 5339
rect 3279 5305 3337 5339
rect 3371 5305 3429 5339
rect 3463 5305 3521 5339
rect 3555 5337 4610 5339
rect 4683 5337 5466 5343
rect 3555 5305 4023 5337
rect 2112 5303 4023 5305
rect 4057 5303 4115 5337
rect 4149 5303 4207 5337
rect 4241 5303 4299 5337
rect 4333 5303 4391 5337
rect 4425 5303 4483 5337
rect 4517 5303 4575 5337
rect 4609 5303 4610 5337
rect 4701 5303 4759 5337
rect 4793 5303 4851 5337
rect 4885 5303 4943 5337
rect 4977 5303 5035 5337
rect 5069 5303 5127 5337
rect 5161 5303 5219 5337
rect 5253 5303 5311 5337
rect 5345 5303 5403 5337
rect 5437 5303 5466 5337
rect 2112 5290 4610 5303
rect 4683 5290 5466 5303
rect 2112 5274 5466 5290
rect 17210 5365 18682 5370
rect 19092 5365 20564 5368
rect 17210 5343 20564 5365
rect 17210 5339 19704 5343
rect 17210 5305 17239 5339
rect 17273 5305 17331 5339
rect 17365 5305 17423 5339
rect 17457 5305 17515 5339
rect 17549 5305 17607 5339
rect 17641 5305 17699 5339
rect 17733 5305 17791 5339
rect 17825 5305 17883 5339
rect 17917 5305 17975 5339
rect 18009 5305 18067 5339
rect 18101 5305 18159 5339
rect 18193 5305 18251 5339
rect 18285 5305 18343 5339
rect 18377 5305 18435 5339
rect 18469 5305 18527 5339
rect 18561 5305 18619 5339
rect 18653 5337 19704 5339
rect 19780 5337 20564 5343
rect 18653 5305 19121 5337
rect 17210 5303 19121 5305
rect 19155 5303 19213 5337
rect 19247 5303 19305 5337
rect 19339 5303 19397 5337
rect 19431 5303 19489 5337
rect 19523 5303 19581 5337
rect 19615 5303 19673 5337
rect 19799 5303 19857 5337
rect 19891 5303 19949 5337
rect 19983 5303 20041 5337
rect 20075 5303 20133 5337
rect 20167 5303 20225 5337
rect 20259 5303 20317 5337
rect 20351 5303 20409 5337
rect 20443 5303 20501 5337
rect 20535 5303 20564 5337
rect 17210 5289 19704 5303
rect 19780 5289 20564 5303
rect 17210 5274 20564 5289
rect 3994 5272 5466 5274
rect 19092 5272 20564 5274
rect 3688 5108 3894 5220
rect 18800 5108 18998 5222
rect 2218 5102 5022 5108
rect 2218 5068 2268 5102
rect 2302 5068 2381 5102
rect 2415 5068 2494 5102
rect 2528 5068 2607 5102
rect 2641 5068 2720 5102
rect 2754 5068 2833 5102
rect 2867 5068 2946 5102
rect 2980 5068 3062 5102
rect 3096 5068 3166 5102
rect 3200 5068 4022 5102
rect 4056 5068 4141 5102
rect 4175 5068 4260 5102
rect 4294 5068 4379 5102
rect 4413 5068 4498 5102
rect 4532 5068 4617 5102
rect 4651 5068 4736 5102
rect 4770 5068 5022 5102
rect 2218 5062 5022 5068
rect 17369 5102 20060 5108
rect 17369 5068 17434 5102
rect 17468 5068 17531 5102
rect 17565 5068 17628 5102
rect 17662 5068 17725 5102
rect 17759 5068 17822 5102
rect 17856 5068 17919 5102
rect 17953 5068 18016 5102
rect 18050 5068 18113 5102
rect 18147 5068 18264 5102
rect 18298 5068 19120 5102
rect 19154 5068 19228 5102
rect 19262 5068 19336 5102
rect 19370 5068 19444 5102
rect 19478 5068 19552 5102
rect 19586 5068 19660 5102
rect 19694 5068 19768 5102
rect 19802 5068 19876 5102
rect 19910 5068 20060 5102
rect 17369 5062 20060 5068
rect 2230 5008 3467 5020
rect 2230 5007 3420 5008
rect 2230 4973 2245 5007
rect 2279 5006 3420 5007
rect 2279 5005 3250 5006
rect 2279 5002 2411 5005
rect 2445 5004 2746 5005
rect 2780 5004 3250 5005
rect 2445 5003 2740 5004
rect 2445 5002 2575 5003
rect 2279 4973 2282 5002
rect 2230 4950 2282 4973
rect 2334 4950 2389 5002
rect 2445 4971 2495 5002
rect 2441 4950 2495 4971
rect 2547 4969 2575 5002
rect 2609 5002 2740 5003
rect 2609 4969 2611 5002
rect 2547 4950 2611 4969
rect 2663 4952 2740 5002
rect 2792 5003 3250 5004
rect 3284 5003 3420 5006
rect 2792 4952 2874 5003
rect 2926 5001 2991 5003
rect 2949 4967 2991 5001
rect 2663 4951 2874 4952
rect 2926 4951 2991 4967
rect 3043 5000 3096 5003
rect 3043 4966 3084 5000
rect 3043 4951 3096 4966
rect 3148 4951 3202 5003
rect 3284 4972 3299 5003
rect 3254 4951 3299 4972
rect 3351 4951 3396 5003
rect 3454 4974 3467 5008
rect 3448 4951 3467 4974
rect 2663 4950 3467 4951
rect 2230 4936 3467 4950
rect 4120 5009 5346 5018
rect 4120 5005 4630 5009
rect 4120 4971 4134 5005
rect 4168 4999 4294 5005
rect 4328 5002 4630 5005
rect 4664 5006 5346 5009
rect 4664 5004 5293 5006
rect 4664 5002 5134 5004
rect 4328 4999 4622 5002
rect 4168 4971 4171 4999
rect 4120 4947 4171 4971
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4965 4461 4999
rect 4495 4965 4500 4999
rect 4436 4947 4500 4965
rect 4552 4950 4622 4999
rect 4674 5001 4964 5002
rect 4681 5000 4964 5001
rect 4998 5000 5134 5002
rect 5168 5000 5293 5004
rect 5327 5000 5346 5006
rect 4552 4949 4629 4950
rect 4681 4949 4763 5000
rect 4815 4996 4880 5000
rect 4828 4962 4880 4996
rect 4552 4948 4763 4949
rect 4815 4948 4880 4962
rect 4932 4968 4964 5000
rect 4932 4948 4985 4968
rect 5037 4948 5091 5000
rect 5168 4970 5188 5000
rect 5143 4948 5188 4970
rect 5240 4948 5285 5000
rect 5337 4948 5346 5000
rect 4552 4947 5346 4948
rect 4120 4934 5346 4947
rect 17321 5008 18588 5020
rect 17321 5001 17391 5008
rect 17321 4967 17343 5001
rect 17377 4967 17391 5001
rect 17321 4956 17391 4967
rect 17443 5006 18588 5008
rect 17443 4956 17503 5006
rect 17321 4954 17503 4956
rect 17555 4954 17610 5006
rect 17662 5000 17712 5006
rect 17764 5005 18588 5006
rect 17764 5004 17844 5005
rect 17878 5004 18588 5005
rect 17662 4966 17679 5000
rect 17662 4954 17712 4966
rect 17764 4954 17838 5004
rect 17321 4952 17838 4954
rect 17890 4952 17992 5004
rect 18044 4992 18129 5004
rect 18045 4958 18129 4992
rect 18181 4990 18226 5004
rect 18044 4952 18129 4958
rect 18213 4956 18226 4990
rect 18181 4952 18226 4956
rect 18278 4952 18326 5004
rect 18378 5003 18588 5004
rect 18378 4999 18415 5003
rect 18383 4965 18415 4999
rect 18378 4952 18415 4965
rect 17321 4951 18415 4952
rect 18467 4951 18511 5003
rect 18563 4951 18588 5003
rect 17321 4936 18588 4951
rect 19207 5009 20463 5018
rect 19207 5006 19728 5009
rect 19207 5002 19557 5006
rect 19591 5002 19728 5006
rect 19762 5002 20463 5009
rect 19207 5000 19225 5002
rect 19207 4966 19222 5000
rect 19207 4950 19225 4966
rect 19277 4950 19319 5002
rect 19371 5001 19418 5002
rect 19371 4967 19395 5001
rect 19371 4950 19418 4967
rect 19470 4950 19526 5002
rect 19591 4972 19622 5002
rect 19578 4950 19622 4972
rect 19674 4950 19720 5002
rect 19772 5001 20463 5002
rect 19772 4950 19839 5001
rect 19207 4949 19839 4950
rect 19891 4995 19953 5001
rect 19891 4961 19897 4995
rect 19931 4961 19953 4995
rect 19891 4949 19953 4961
rect 20005 4995 20070 5001
rect 20005 4961 20062 4995
rect 20005 4949 20070 4961
rect 20122 4949 20197 5001
rect 20249 4993 20312 5001
rect 20266 4959 20312 4993
rect 20249 4949 20312 4959
rect 20364 4997 20463 5001
rect 20364 4963 20395 4997
rect 20429 4963 20463 4997
rect 20364 4949 20463 4963
rect 19207 4934 20463 4949
rect -3552 4832 26658 4904
rect -3552 4716 -2017 4832
rect -1709 4716 -129 4832
rect 179 4716 1759 4832
rect 2067 4795 3647 4832
rect 2067 4761 2141 4795
rect 2175 4761 2233 4795
rect 2267 4761 2325 4795
rect 2359 4761 2417 4795
rect 2451 4761 2509 4795
rect 2543 4761 2601 4795
rect 2635 4761 2693 4795
rect 2727 4761 2785 4795
rect 2819 4761 2877 4795
rect 2911 4761 2969 4795
rect 3003 4761 3061 4795
rect 3095 4761 3153 4795
rect 3187 4761 3245 4795
rect 3279 4761 3337 4795
rect 3371 4761 3429 4795
rect 3463 4761 3521 4795
rect 3555 4761 3647 4795
rect 2067 4716 3647 4761
rect 3955 4793 5535 4832
rect 3955 4759 4023 4793
rect 4057 4759 4115 4793
rect 4149 4759 4207 4793
rect 4241 4759 4299 4793
rect 4333 4759 4391 4793
rect 4425 4759 4483 4793
rect 4517 4759 4575 4793
rect 4609 4759 4667 4793
rect 4701 4759 4759 4793
rect 4793 4759 4851 4793
rect 4885 4759 4943 4793
rect 4977 4759 5035 4793
rect 5069 4759 5127 4793
rect 5161 4759 5219 4793
rect 5253 4759 5311 4793
rect 5345 4759 5403 4793
rect 5437 4759 5535 4793
rect 3955 4716 5535 4759
rect 5843 4716 7423 4832
rect 7731 4716 9311 4832
rect 9619 4716 11199 4832
rect 11507 4716 13081 4832
rect 13389 4716 14969 4832
rect 15277 4716 16857 4832
rect 17165 4795 18745 4832
rect 17165 4761 17239 4795
rect 17273 4761 17331 4795
rect 17365 4761 17423 4795
rect 17457 4761 17515 4795
rect 17549 4761 17607 4795
rect 17641 4761 17699 4795
rect 17733 4761 17791 4795
rect 17825 4761 17883 4795
rect 17917 4761 17975 4795
rect 18009 4761 18067 4795
rect 18101 4761 18159 4795
rect 18193 4761 18251 4795
rect 18285 4761 18343 4795
rect 18377 4761 18435 4795
rect 18469 4761 18527 4795
rect 18561 4761 18619 4795
rect 18653 4761 18745 4795
rect 17165 4716 18745 4761
rect 19053 4793 20633 4832
rect 19053 4759 19121 4793
rect 19155 4759 19213 4793
rect 19247 4759 19305 4793
rect 19339 4759 19397 4793
rect 19431 4759 19489 4793
rect 19523 4759 19581 4793
rect 19615 4759 19673 4793
rect 19707 4759 19765 4793
rect 19799 4759 19857 4793
rect 19891 4759 19949 4793
rect 19983 4759 20041 4793
rect 20075 4759 20133 4793
rect 20167 4759 20225 4793
rect 20259 4759 20317 4793
rect 20351 4759 20409 4793
rect 20443 4759 20501 4793
rect 20535 4759 20633 4793
rect 19053 4716 20633 4759
rect 20941 4716 22521 4832
rect 22829 4716 24409 4832
rect 24717 4716 26297 4832
rect 26605 4716 26658 4832
rect -3552 4715 26658 4716
rect -3552 4681 -3305 4715
rect -3271 4681 -3213 4715
rect -3179 4681 -3121 4715
rect -3087 4681 -2491 4715
rect -2457 4681 -2399 4715
rect -2365 4681 -2307 4715
rect -2273 4681 -1417 4715
rect -1383 4681 -1325 4715
rect -1291 4681 -1233 4715
rect -1199 4681 -603 4715
rect -569 4681 -511 4715
rect -477 4681 -419 4715
rect -385 4681 471 4715
rect 505 4681 563 4715
rect 597 4681 655 4715
rect 689 4681 1285 4715
rect 1319 4681 1377 4715
rect 1411 4681 1469 4715
rect 1503 4681 2359 4715
rect 2393 4681 2451 4715
rect 2485 4681 2543 4715
rect 2577 4681 3173 4715
rect 3207 4681 3265 4715
rect 3299 4681 3357 4715
rect 3391 4681 4247 4715
rect 4281 4681 4339 4715
rect 4373 4681 4431 4715
rect 4465 4681 5061 4715
rect 5095 4681 5153 4715
rect 5187 4681 5245 4715
rect 5279 4681 6135 4715
rect 6169 4681 6227 4715
rect 6261 4681 6319 4715
rect 6353 4681 6949 4715
rect 6983 4681 7041 4715
rect 7075 4681 7133 4715
rect 7167 4681 8023 4715
rect 8057 4681 8115 4715
rect 8149 4681 8207 4715
rect 8241 4681 8837 4715
rect 8871 4681 8929 4715
rect 8963 4681 9021 4715
rect 9055 4681 9911 4715
rect 9945 4681 10003 4715
rect 10037 4681 10095 4715
rect 10129 4681 10725 4715
rect 10759 4681 10817 4715
rect 10851 4681 10909 4715
rect 10943 4681 11793 4715
rect 11827 4681 11885 4715
rect 11919 4681 11977 4715
rect 12011 4681 12607 4715
rect 12641 4681 12699 4715
rect 12733 4681 12791 4715
rect 12825 4681 13681 4715
rect 13715 4681 13773 4715
rect 13807 4681 13865 4715
rect 13899 4681 14495 4715
rect 14529 4681 14587 4715
rect 14621 4681 14679 4715
rect 14713 4681 15569 4715
rect 15603 4681 15661 4715
rect 15695 4681 15753 4715
rect 15787 4681 16383 4715
rect 16417 4681 16475 4715
rect 16509 4681 16567 4715
rect 16601 4681 17457 4715
rect 17491 4681 17549 4715
rect 17583 4681 17641 4715
rect 17675 4681 18271 4715
rect 18305 4681 18363 4715
rect 18397 4681 18455 4715
rect 18489 4681 19345 4715
rect 19379 4681 19437 4715
rect 19471 4681 19529 4715
rect 19563 4681 20159 4715
rect 20193 4681 20251 4715
rect 20285 4681 20343 4715
rect 20377 4681 21233 4715
rect 21267 4681 21325 4715
rect 21359 4681 21417 4715
rect 21451 4681 22047 4715
rect 22081 4681 22139 4715
rect 22173 4681 22231 4715
rect 22265 4681 23121 4715
rect 23155 4681 23213 4715
rect 23247 4681 23305 4715
rect 23339 4681 23935 4715
rect 23969 4681 24027 4715
rect 24061 4681 24119 4715
rect 24153 4681 25009 4715
rect 25043 4681 25101 4715
rect 25135 4681 25193 4715
rect 25227 4681 25823 4715
rect 25857 4681 25915 4715
rect 25949 4681 26007 4715
rect 26041 4681 26658 4715
rect -3552 4675 26658 4681
rect -3552 4650 -2871 4675
rect -3492 3692 -3414 4650
rect -2900 4641 -2871 4650
rect -2837 4650 -983 4675
rect -2837 4641 -2810 4650
rect -2900 4620 -2810 4641
rect -2814 4584 -2756 4586
rect -2814 4567 -2752 4584
rect -2814 4533 -2802 4567
rect -2768 4533 -2752 4567
rect -2814 4524 -2752 4533
rect -3314 4486 -2948 4490
rect -2866 4486 -2800 4494
rect -3314 4458 -2906 4486
rect -3314 4420 -3286 4458
rect -2992 4439 -2906 4458
rect -3314 4412 -3248 4420
rect -3314 4378 -3299 4412
rect -3265 4378 -3248 4412
rect -3314 4366 -3248 4378
rect -3142 4416 -3074 4422
rect -3142 4364 -3132 4416
rect -3080 4364 -3074 4416
rect -3142 4358 -3074 4364
rect -2992 4405 -2946 4439
rect -2912 4405 -2906 4439
rect -2866 4434 -2860 4486
rect -2808 4434 -2800 4486
rect -2866 4426 -2850 4434
rect -2992 4367 -2906 4405
rect -2992 4333 -2946 4367
rect -2912 4333 -2906 4367
rect -3232 4304 -3164 4310
rect -3232 4252 -3224 4304
rect -3172 4252 -3164 4304
rect -3232 4242 -3164 4252
rect -2992 4286 -2906 4333
rect -2856 4405 -2850 4426
rect -2816 4426 -2800 4434
rect -2760 4454 -2432 4486
rect -2760 4439 -2664 4454
rect -2816 4405 -2810 4426
rect -2856 4367 -2810 4405
rect -2856 4333 -2850 4367
rect -2816 4333 -2810 4367
rect -2856 4286 -2810 4333
rect -2760 4405 -2754 4439
rect -2720 4405 -2664 4439
rect -2460 4418 -2432 4454
rect -2760 4367 -2664 4405
rect -2760 4333 -2754 4367
rect -2720 4333 -2664 4367
rect -2502 4410 -2432 4418
rect -2502 4376 -2487 4410
rect -2453 4376 -2432 4410
rect -2502 4358 -2432 4376
rect -2326 4418 -2262 4424
rect -2326 4366 -2320 4418
rect -2268 4366 -2262 4418
rect -2326 4360 -2262 4366
rect -2760 4286 -2664 4333
rect -3334 4171 -3058 4202
rect -3334 4137 -3305 4171
rect -3271 4137 -3213 4171
rect -3179 4137 -3121 4171
rect -3087 4137 -3058 4171
rect -3334 4106 -3058 4137
rect -2992 4086 -2942 4286
rect -2910 4239 -2852 4254
rect -2910 4205 -2898 4239
rect -2864 4205 -2852 4239
rect -2910 4188 -2852 4205
rect -2798 4158 -2740 4176
rect -2798 4124 -2786 4158
rect -2752 4124 -2740 4158
rect -2798 4114 -2740 4124
rect -2710 4086 -2664 4286
rect -2414 4302 -2350 4308
rect -2414 4250 -2408 4302
rect -2356 4250 -2350 4302
rect -2414 4244 -2350 4250
rect -2520 4171 -2244 4202
rect -2520 4137 -2491 4171
rect -2457 4137 -2399 4171
rect -2365 4137 -2307 4171
rect -2273 4137 -2244 4171
rect -2520 4134 -2244 4137
rect -3352 4069 -3288 4076
rect -3352 4036 -3346 4069
rect -3294 4036 -3288 4069
rect -3176 4069 -3112 4076
rect -3176 4036 -3170 4069
rect -3294 4017 -3170 4036
rect -3118 4017 -3112 4069
rect -3346 4008 -3112 4017
rect -2992 4074 -2890 4086
rect -2992 4040 -2930 4074
rect -2896 4040 -2890 4074
rect -2992 4002 -2890 4040
rect -2840 4074 -2794 4086
rect -2840 4040 -2834 4074
rect -2800 4040 -2794 4074
rect -2840 4020 -2794 4040
rect -2744 4074 -2664 4086
rect -2744 4040 -2738 4074
rect -2704 4040 -2664 4074
rect -2992 3970 -2930 4002
rect -3196 3968 -2930 3970
rect -2896 3968 -2890 4002
rect -3196 3956 -2890 3968
rect -2850 4014 -2784 4020
rect -2850 3962 -2842 4014
rect -2790 3962 -2784 4014
rect -2850 3956 -2784 3962
rect -2744 4002 -2664 4040
rect -2744 3968 -2738 4002
rect -2704 3968 -2664 4002
rect -2548 4106 -2244 4134
rect -2744 3956 -2698 3968
rect -3196 3942 -2942 3956
rect -3352 3936 -3286 3942
rect -3352 3884 -3344 3936
rect -3292 3884 -3286 3936
rect -3352 3878 -3286 3884
rect -3512 3678 -3236 3692
rect -3512 3661 -3320 3678
rect -3268 3661 -3236 3678
rect -3512 3627 -3483 3661
rect -3449 3627 -3391 3661
rect -3357 3627 -3320 3661
rect -3265 3627 -3236 3661
rect -3512 3626 -3320 3627
rect -3268 3626 -3236 3627
rect -3512 3596 -3236 3626
rect -3196 3592 -3168 3942
rect -2896 3918 -2832 3928
rect -2896 3884 -2882 3918
rect -2848 3884 -2576 3918
rect -2896 3866 -2832 3884
rect -2980 3820 -2908 3832
rect -2980 3768 -2970 3820
rect -2918 3768 -2908 3820
rect -2980 3756 -2908 3768
rect -2610 3702 -2576 3884
rect -2548 3802 -2520 4106
rect -2548 3792 -2480 3802
rect -2548 3758 -2532 3792
rect -2498 3758 -2480 3792
rect -2548 3744 -2480 3758
rect -3136 3674 -2576 3702
rect -3136 3671 -3070 3674
rect -3136 3637 -3120 3671
rect -3086 3637 -3070 3671
rect -3136 3628 -3070 3637
rect -2902 3619 -2812 3640
rect -3196 3564 -3124 3592
rect -3170 3543 -3124 3564
rect -3170 3509 -3164 3543
rect -3130 3509 -3124 3543
rect -3170 3471 -3124 3509
rect -3170 3437 -3164 3471
rect -3130 3437 -3124 3471
rect -3170 3390 -3124 3437
rect -3082 3570 -3036 3590
rect -2902 3585 -2873 3619
rect -2839 3585 -2812 3619
rect -3082 3564 -3014 3570
rect -2902 3564 -2812 3585
rect -3082 3543 -3074 3564
rect -3082 3509 -3076 3543
rect -3022 3512 -3014 3564
rect -3042 3509 -3014 3512
rect -3082 3504 -3014 3509
rect -2816 3528 -2758 3530
rect -2610 3528 -2576 3674
rect -2490 3671 -2424 3682
rect -2490 3637 -2474 3671
rect -2440 3637 -2424 3671
rect -2490 3626 -2424 3637
rect -2316 3672 -1692 3704
rect -1604 3692 -1526 4650
rect -1012 4641 -983 4650
rect -949 4650 905 4675
rect -949 4641 -922 4650
rect -1012 4620 -922 4641
rect -926 4584 -868 4586
rect -926 4567 -864 4584
rect -926 4533 -914 4567
rect -880 4533 -864 4567
rect -926 4524 -864 4533
rect -1426 4486 -1060 4490
rect -978 4486 -912 4494
rect -1426 4458 -1018 4486
rect -1426 4420 -1398 4458
rect -1104 4439 -1018 4458
rect -1426 4412 -1360 4420
rect -1426 4378 -1411 4412
rect -1377 4378 -1360 4412
rect -1426 4366 -1360 4378
rect -1254 4416 -1186 4422
rect -1254 4364 -1244 4416
rect -1192 4364 -1186 4416
rect -1254 4358 -1186 4364
rect -1104 4405 -1058 4439
rect -1024 4405 -1018 4439
rect -978 4434 -972 4486
rect -920 4434 -912 4486
rect -978 4426 -962 4434
rect -1104 4367 -1018 4405
rect -1104 4333 -1058 4367
rect -1024 4333 -1018 4367
rect -1344 4304 -1276 4310
rect -1344 4252 -1336 4304
rect -1284 4252 -1276 4304
rect -1344 4242 -1276 4252
rect -1104 4286 -1018 4333
rect -968 4405 -962 4426
rect -928 4426 -912 4434
rect -872 4454 -544 4486
rect -872 4439 -776 4454
rect -928 4405 -922 4426
rect -968 4367 -922 4405
rect -968 4333 -962 4367
rect -928 4333 -922 4367
rect -968 4286 -922 4333
rect -872 4405 -866 4439
rect -832 4405 -776 4439
rect -572 4418 -544 4454
rect -872 4367 -776 4405
rect -872 4333 -866 4367
rect -832 4333 -776 4367
rect -614 4410 -544 4418
rect -614 4376 -599 4410
rect -565 4376 -544 4410
rect -614 4358 -544 4376
rect -438 4418 -374 4424
rect -438 4366 -432 4418
rect -380 4366 -374 4418
rect -438 4360 -374 4366
rect -872 4286 -776 4333
rect -1446 4171 -1170 4202
rect -1446 4137 -1417 4171
rect -1383 4137 -1325 4171
rect -1291 4137 -1233 4171
rect -1199 4137 -1170 4171
rect -1446 4106 -1170 4137
rect -1104 4086 -1054 4286
rect -1022 4239 -964 4254
rect -1022 4205 -1010 4239
rect -976 4205 -964 4239
rect -1022 4188 -964 4205
rect -910 4158 -852 4176
rect -910 4124 -898 4158
rect -864 4124 -852 4158
rect -910 4114 -852 4124
rect -822 4086 -776 4286
rect -526 4302 -462 4308
rect -526 4250 -520 4302
rect -468 4250 -462 4302
rect -526 4244 -462 4250
rect -632 4171 -356 4202
rect -632 4137 -603 4171
rect -569 4137 -511 4171
rect -477 4137 -419 4171
rect -385 4137 -356 4171
rect -632 4134 -356 4137
rect -1464 4069 -1400 4076
rect -1464 4036 -1458 4069
rect -1406 4036 -1400 4069
rect -1288 4069 -1224 4076
rect -1288 4036 -1282 4069
rect -1406 4017 -1282 4036
rect -1230 4017 -1224 4069
rect -1458 4008 -1224 4017
rect -1104 4074 -1002 4086
rect -1104 4040 -1042 4074
rect -1008 4040 -1002 4074
rect -1104 4002 -1002 4040
rect -952 4074 -906 4086
rect -952 4040 -946 4074
rect -912 4040 -906 4074
rect -952 4020 -906 4040
rect -856 4074 -776 4086
rect -856 4040 -850 4074
rect -816 4040 -776 4074
rect -1104 3970 -1042 4002
rect -1308 3968 -1042 3970
rect -1008 3968 -1002 4002
rect -1308 3956 -1002 3968
rect -962 4014 -896 4020
rect -962 3962 -954 4014
rect -902 3962 -896 4014
rect -962 3956 -896 3962
rect -856 4002 -776 4040
rect -856 3968 -850 4002
rect -816 3968 -776 4002
rect -660 4106 -356 4134
rect -856 3956 -810 3968
rect -1308 3942 -1054 3956
rect -1464 3936 -1398 3942
rect -1464 3884 -1456 3936
rect -1404 3884 -1398 3936
rect -1464 3878 -1398 3884
rect -2316 3669 -2286 3672
rect -2234 3669 -1692 3672
rect -2316 3635 -2287 3669
rect -2234 3635 -2195 3669
rect -2161 3635 -2103 3669
rect -2069 3667 -1692 3669
rect -2069 3635 -1941 3667
rect -2316 3620 -2286 3635
rect -2234 3633 -1941 3635
rect -1907 3633 -1849 3667
rect -1815 3633 -1757 3667
rect -1723 3633 -1692 3667
rect -2234 3620 -1692 3633
rect -2316 3602 -1692 3620
rect -1624 3678 -1348 3692
rect -1624 3661 -1432 3678
rect -1380 3661 -1348 3678
rect -1624 3627 -1595 3661
rect -1561 3627 -1503 3661
rect -1469 3627 -1432 3661
rect -1377 3627 -1348 3661
rect -1624 3626 -1432 3627
rect -1380 3626 -1348 3627
rect -1624 3596 -1348 3626
rect -1308 3592 -1280 3942
rect -1008 3918 -944 3928
rect -1008 3884 -994 3918
rect -960 3884 -688 3918
rect -1008 3866 -944 3884
rect -1092 3820 -1020 3832
rect -1092 3768 -1082 3820
rect -1030 3768 -1020 3820
rect -1092 3756 -1020 3768
rect -722 3702 -688 3884
rect -660 3802 -632 4106
rect -660 3792 -592 3802
rect -660 3758 -644 3792
rect -610 3758 -592 3792
rect -660 3744 -592 3758
rect -1248 3674 -688 3702
rect -1248 3671 -1182 3674
rect -1248 3637 -1232 3671
rect -1198 3637 -1182 3671
rect -1248 3628 -1182 3637
rect -1014 3619 -924 3640
rect -2816 3511 -2576 3528
rect -2532 3584 -2466 3590
rect -2532 3532 -2524 3584
rect -2472 3532 -2466 3584
rect -2532 3526 -2518 3532
rect -3082 3471 -3036 3504
rect -3082 3437 -3076 3471
rect -3042 3437 -3036 3471
rect -2816 3477 -2804 3511
rect -2770 3500 -2576 3511
rect -2524 3509 -2518 3526
rect -2484 3526 -2466 3532
rect -2436 3543 -2390 3590
rect -1308 3564 -1236 3592
rect -2484 3509 -2478 3526
rect -2770 3477 -2578 3500
rect -2816 3468 -2578 3477
rect -3082 3390 -3036 3437
rect -2868 3430 -2802 3438
rect -2954 3426 -2908 3430
rect -2994 3383 -2908 3426
rect -3532 3372 -3464 3378
rect -3532 3320 -3525 3372
rect -3473 3366 -3464 3372
rect -3473 3360 -3380 3366
rect -3473 3326 -3434 3360
rect -3400 3326 -3380 3360
rect -3473 3320 -3380 3326
rect -3532 3316 -3380 3320
rect -3136 3343 -3070 3354
rect -3532 3314 -3464 3316
rect -3136 3309 -3120 3343
rect -3086 3309 -3070 3343
rect -3136 3296 -3070 3309
rect -2994 3349 -2948 3383
rect -2914 3349 -2908 3383
rect -2868 3378 -2862 3430
rect -2810 3378 -2802 3430
rect -2868 3370 -2852 3378
rect -2994 3311 -2908 3349
rect -2994 3277 -2948 3311
rect -2914 3277 -2908 3311
rect -2994 3230 -2908 3277
rect -2858 3349 -2852 3370
rect -2818 3370 -2802 3378
rect -2762 3383 -2666 3430
rect -2818 3349 -2812 3370
rect -2858 3311 -2812 3349
rect -2858 3277 -2852 3311
rect -2818 3277 -2812 3311
rect -2858 3230 -2812 3277
rect -2762 3349 -2756 3383
rect -2722 3349 -2666 3383
rect -2762 3311 -2666 3349
rect -2762 3277 -2756 3311
rect -2722 3277 -2666 3311
rect -2762 3230 -2666 3277
rect -2994 3176 -2944 3230
rect -3512 3130 -3236 3148
rect -3512 3117 -3389 3130
rect -3337 3117 -3236 3130
rect -3160 3126 -3102 3134
rect -3512 3083 -3483 3117
rect -3449 3083 -3391 3117
rect -3337 3083 -3299 3117
rect -3265 3083 -3236 3117
rect -3512 3078 -3389 3083
rect -3337 3078 -3236 3083
rect -3512 3052 -3236 3078
rect -3168 3120 -3094 3126
rect -3168 3068 -3157 3120
rect -3105 3068 -3094 3120
rect -3014 3110 -2944 3176
rect -2912 3183 -2854 3198
rect -2912 3149 -2900 3183
rect -2866 3149 -2854 3183
rect -2912 3132 -2854 3149
rect -3168 3062 -3094 3068
rect -3160 3056 -3102 3062
rect -3444 2782 -3360 3052
rect -2994 3030 -2944 3110
rect -2800 3102 -2742 3120
rect -2800 3068 -2788 3102
rect -2754 3068 -2742 3102
rect -2800 3058 -2742 3068
rect -2712 3030 -2666 3230
rect -2994 3018 -2892 3030
rect -2994 2984 -2932 3018
rect -2898 2984 -2892 3018
rect -2994 2946 -2892 2984
rect -2842 3018 -2796 3030
rect -2842 2984 -2836 3018
rect -2802 2984 -2796 3018
rect -2842 2964 -2796 2984
rect -2746 3018 -2666 3030
rect -2746 2984 -2740 3018
rect -2706 2984 -2666 3018
rect -2994 2912 -2932 2946
rect -2898 2912 -2892 2946
rect -2994 2900 -2892 2912
rect -2852 2958 -2786 2964
rect -2852 2906 -2844 2958
rect -2792 2906 -2786 2958
rect -2852 2900 -2786 2906
rect -2746 2946 -2666 2984
rect -2746 2912 -2740 2946
rect -2706 2912 -2666 2946
rect -2638 3236 -2578 3468
rect -2524 3471 -2478 3509
rect -2524 3437 -2518 3471
rect -2484 3437 -2478 3471
rect -2524 3390 -2478 3437
rect -2436 3509 -2430 3543
rect -2396 3509 -2390 3543
rect -2436 3471 -2390 3509
rect -2436 3437 -2430 3471
rect -2396 3437 -2390 3471
rect -2436 3390 -2390 3437
rect -1282 3543 -1236 3564
rect -1282 3509 -1276 3543
rect -1242 3509 -1236 3543
rect -1282 3471 -1236 3509
rect -1282 3437 -1276 3471
rect -1242 3437 -1236 3471
rect -1282 3390 -1236 3437
rect -1194 3570 -1148 3590
rect -1014 3585 -985 3619
rect -951 3585 -924 3619
rect -1194 3564 -1126 3570
rect -1014 3564 -924 3585
rect -1194 3543 -1186 3564
rect -1194 3509 -1188 3543
rect -1134 3512 -1126 3564
rect -1154 3509 -1126 3512
rect -1194 3504 -1126 3509
rect -928 3528 -870 3530
rect -722 3528 -688 3674
rect -602 3671 -536 3682
rect -602 3637 -586 3671
rect -552 3637 -536 3671
rect -602 3626 -536 3637
rect -428 3672 196 3704
rect 284 3692 362 4650
rect 876 4641 905 4650
rect 939 4650 2793 4675
rect 939 4641 966 4650
rect 876 4620 966 4641
rect 962 4584 1020 4586
rect 962 4567 1024 4584
rect 962 4533 974 4567
rect 1008 4533 1024 4567
rect 962 4524 1024 4533
rect 462 4486 828 4490
rect 910 4486 976 4494
rect 462 4458 870 4486
rect 462 4420 490 4458
rect 784 4439 870 4458
rect 462 4412 528 4420
rect 462 4378 477 4412
rect 511 4378 528 4412
rect 462 4366 528 4378
rect 634 4416 702 4422
rect 634 4364 644 4416
rect 696 4364 702 4416
rect 634 4358 702 4364
rect 784 4405 830 4439
rect 864 4405 870 4439
rect 910 4434 916 4486
rect 968 4434 976 4486
rect 910 4426 926 4434
rect 784 4367 870 4405
rect 784 4333 830 4367
rect 864 4333 870 4367
rect 544 4304 612 4310
rect 544 4252 552 4304
rect 604 4252 612 4304
rect 544 4242 612 4252
rect 784 4286 870 4333
rect 920 4405 926 4426
rect 960 4426 976 4434
rect 1016 4454 1344 4486
rect 1016 4439 1112 4454
rect 960 4405 966 4426
rect 920 4367 966 4405
rect 920 4333 926 4367
rect 960 4333 966 4367
rect 920 4286 966 4333
rect 1016 4405 1022 4439
rect 1056 4405 1112 4439
rect 1316 4418 1344 4454
rect 1016 4367 1112 4405
rect 1016 4333 1022 4367
rect 1056 4333 1112 4367
rect 1274 4410 1344 4418
rect 1274 4376 1289 4410
rect 1323 4376 1344 4410
rect 1274 4358 1344 4376
rect 1450 4418 1514 4424
rect 1450 4366 1456 4418
rect 1508 4366 1514 4418
rect 1450 4360 1514 4366
rect 1016 4286 1112 4333
rect 442 4171 718 4202
rect 442 4137 471 4171
rect 505 4137 563 4171
rect 597 4137 655 4171
rect 689 4137 718 4171
rect 442 4106 718 4137
rect 784 4086 834 4286
rect 866 4239 924 4254
rect 866 4205 878 4239
rect 912 4205 924 4239
rect 866 4188 924 4205
rect 978 4158 1036 4176
rect 978 4124 990 4158
rect 1024 4124 1036 4158
rect 978 4114 1036 4124
rect 1066 4086 1112 4286
rect 1362 4302 1426 4308
rect 1362 4250 1368 4302
rect 1420 4250 1426 4302
rect 1362 4244 1426 4250
rect 1256 4171 1532 4202
rect 1256 4137 1285 4171
rect 1319 4137 1377 4171
rect 1411 4137 1469 4171
rect 1503 4137 1532 4171
rect 1256 4134 1532 4137
rect 424 4069 488 4076
rect 424 4036 430 4069
rect 482 4036 488 4069
rect 600 4069 664 4076
rect 600 4036 606 4069
rect 482 4017 606 4036
rect 658 4017 664 4069
rect 430 4008 664 4017
rect 784 4074 886 4086
rect 784 4040 846 4074
rect 880 4040 886 4074
rect 784 4002 886 4040
rect 936 4074 982 4086
rect 936 4040 942 4074
rect 976 4040 982 4074
rect 936 4020 982 4040
rect 1032 4074 1112 4086
rect 1032 4040 1038 4074
rect 1072 4040 1112 4074
rect 784 3970 846 4002
rect 580 3968 846 3970
rect 880 3968 886 4002
rect 580 3956 886 3968
rect 926 4014 992 4020
rect 926 3962 934 4014
rect 986 3962 992 4014
rect 926 3956 992 3962
rect 1032 4002 1112 4040
rect 1032 3968 1038 4002
rect 1072 3968 1112 4002
rect 1228 4106 1532 4134
rect 1032 3956 1078 3968
rect 580 3942 834 3956
rect 424 3936 490 3942
rect 424 3884 432 3936
rect 484 3884 490 3936
rect 424 3878 490 3884
rect -428 3669 -398 3672
rect -346 3669 196 3672
rect -428 3635 -399 3669
rect -346 3635 -307 3669
rect -273 3635 -215 3669
rect -181 3667 196 3669
rect -181 3635 -53 3667
rect -428 3620 -398 3635
rect -346 3633 -53 3635
rect -19 3633 39 3667
rect 73 3633 131 3667
rect 165 3633 196 3667
rect -346 3620 196 3633
rect -428 3602 196 3620
rect 264 3678 540 3692
rect 264 3661 456 3678
rect 508 3661 540 3678
rect 264 3627 293 3661
rect 327 3627 385 3661
rect 419 3627 456 3661
rect 511 3627 540 3661
rect 264 3626 456 3627
rect 508 3626 540 3627
rect 264 3596 540 3626
rect 580 3592 608 3942
rect 880 3918 944 3928
rect 880 3884 894 3918
rect 928 3884 1200 3918
rect 880 3866 944 3884
rect 796 3820 868 3832
rect 796 3768 806 3820
rect 858 3768 868 3820
rect 796 3756 868 3768
rect 1166 3702 1200 3884
rect 1228 3802 1256 4106
rect 1228 3792 1296 3802
rect 1228 3758 1244 3792
rect 1278 3758 1296 3792
rect 1228 3744 1296 3758
rect 640 3674 1200 3702
rect 640 3671 706 3674
rect 640 3637 656 3671
rect 690 3637 706 3671
rect 640 3628 706 3637
rect 874 3619 964 3640
rect -928 3511 -688 3528
rect -644 3584 -578 3590
rect -644 3532 -636 3584
rect -584 3532 -578 3584
rect -644 3526 -630 3532
rect -1194 3471 -1148 3504
rect -1194 3437 -1188 3471
rect -1154 3437 -1148 3471
rect -928 3477 -916 3511
rect -882 3500 -688 3511
rect -636 3509 -630 3526
rect -596 3526 -578 3532
rect -548 3543 -502 3590
rect 580 3564 652 3592
rect -596 3509 -590 3526
rect -882 3477 -690 3500
rect -928 3468 -690 3477
rect -1194 3390 -1148 3437
rect -980 3430 -914 3438
rect -1066 3426 -1020 3430
rect -1950 3368 -1878 3372
rect -2490 3343 -2424 3356
rect -2490 3309 -2474 3343
rect -2440 3309 -2424 3343
rect -2490 3300 -2424 3309
rect -1950 3316 -1941 3368
rect -1889 3316 -1878 3368
rect -1950 3304 -1878 3316
rect -1754 3366 -1680 3386
rect -1106 3383 -1020 3426
rect -1754 3332 -1742 3366
rect -1708 3332 -1680 3366
rect -1754 3308 -1680 3332
rect -1644 3372 -1576 3378
rect -1644 3320 -1637 3372
rect -1585 3366 -1576 3372
rect -1585 3360 -1492 3366
rect -1585 3326 -1546 3360
rect -1512 3326 -1492 3360
rect -1585 3320 -1492 3326
rect -1644 3316 -1492 3320
rect -1248 3343 -1182 3354
rect -1644 3314 -1576 3316
rect -1248 3309 -1232 3343
rect -1198 3309 -1182 3343
rect -1248 3296 -1182 3309
rect -1106 3349 -1060 3383
rect -1026 3349 -1020 3383
rect -980 3378 -974 3430
rect -922 3378 -914 3430
rect -980 3370 -964 3378
rect -1106 3311 -1020 3349
rect -1106 3277 -1060 3311
rect -1026 3277 -1020 3311
rect -2168 3256 -2110 3270
rect -2168 3236 -2156 3256
rect -2638 3222 -2156 3236
rect -2122 3222 -2110 3256
rect -2638 3202 -2110 3222
rect -1106 3230 -1020 3277
rect -970 3349 -964 3370
rect -930 3370 -914 3378
rect -874 3383 -778 3430
rect -930 3349 -924 3370
rect -970 3311 -924 3349
rect -970 3277 -964 3311
rect -930 3277 -924 3311
rect -970 3230 -924 3277
rect -874 3349 -868 3383
rect -834 3349 -778 3383
rect -874 3311 -778 3349
rect -874 3277 -868 3311
rect -834 3277 -778 3311
rect -874 3230 -778 3277
rect -2746 2900 -2700 2912
rect -2638 2872 -2578 3202
rect -1106 3176 -1056 3230
rect -2532 3152 -2456 3158
rect -2532 3100 -2524 3152
rect -2472 3100 -2456 3152
rect -2532 3094 -2456 3100
rect -2316 3125 -1694 3156
rect -2898 2862 -2578 2872
rect -2898 2828 -2884 2862
rect -2850 2828 -2578 2862
rect -2898 2810 -2578 2828
rect -2316 3091 -2287 3125
rect -2253 3091 -2195 3125
rect -2161 3091 -2103 3125
rect -2069 3123 -1694 3125
rect -2069 3091 -1941 3123
rect -2316 3089 -1941 3091
rect -1907 3089 -1849 3123
rect -1815 3089 -1757 3123
rect -1723 3089 -1694 3123
rect -2316 3058 -1694 3089
rect -1624 3130 -1348 3148
rect -1624 3117 -1501 3130
rect -1449 3117 -1348 3130
rect -1272 3126 -1214 3134
rect -1624 3083 -1595 3117
rect -1561 3083 -1503 3117
rect -1449 3083 -1411 3117
rect -1377 3083 -1348 3117
rect -1624 3078 -1501 3083
rect -1449 3078 -1348 3083
rect -2316 2782 -2218 3058
rect -1624 3052 -1348 3078
rect -1280 3120 -1206 3126
rect -1280 3068 -1269 3120
rect -1217 3068 -1206 3120
rect -1126 3110 -1056 3176
rect -1024 3183 -966 3198
rect -1024 3149 -1012 3183
rect -978 3149 -966 3183
rect -1024 3132 -966 3149
rect -1280 3062 -1206 3068
rect -1272 3056 -1214 3062
rect -1556 2782 -1472 3052
rect -1106 3030 -1056 3110
rect -912 3102 -854 3120
rect -912 3068 -900 3102
rect -866 3068 -854 3102
rect -912 3058 -854 3068
rect -824 3030 -778 3230
rect -1106 3018 -1004 3030
rect -1106 2984 -1044 3018
rect -1010 2984 -1004 3018
rect -1106 2946 -1004 2984
rect -954 3018 -908 3030
rect -954 2984 -948 3018
rect -914 2984 -908 3018
rect -954 2964 -908 2984
rect -858 3018 -778 3030
rect -858 2984 -852 3018
rect -818 2984 -778 3018
rect -1106 2912 -1044 2946
rect -1010 2912 -1004 2946
rect -1106 2900 -1004 2912
rect -964 2958 -898 2964
rect -964 2906 -956 2958
rect -904 2906 -898 2958
rect -964 2900 -898 2906
rect -858 2946 -778 2984
rect -858 2912 -852 2946
rect -818 2912 -778 2946
rect -750 3236 -690 3468
rect -636 3471 -590 3509
rect -636 3437 -630 3471
rect -596 3437 -590 3471
rect -636 3390 -590 3437
rect -548 3509 -542 3543
rect -508 3509 -502 3543
rect -548 3471 -502 3509
rect -548 3437 -542 3471
rect -508 3437 -502 3471
rect -548 3390 -502 3437
rect 606 3543 652 3564
rect 606 3509 612 3543
rect 646 3509 652 3543
rect 606 3471 652 3509
rect 606 3437 612 3471
rect 646 3437 652 3471
rect 606 3390 652 3437
rect 694 3570 740 3590
rect 874 3585 903 3619
rect 937 3585 964 3619
rect 694 3564 762 3570
rect 874 3564 964 3585
rect 694 3543 702 3564
rect 694 3509 700 3543
rect 754 3512 762 3564
rect 734 3509 762 3512
rect 694 3504 762 3509
rect 960 3528 1018 3530
rect 1166 3528 1200 3674
rect 1286 3671 1352 3682
rect 1286 3637 1302 3671
rect 1336 3637 1352 3671
rect 1286 3626 1352 3637
rect 1460 3672 2084 3704
rect 2172 3692 2250 4650
rect 2764 4641 2793 4650
rect 2827 4650 4681 4675
rect 2827 4641 2854 4650
rect 2764 4620 2854 4641
rect 2850 4584 2908 4586
rect 2850 4567 2912 4584
rect 2850 4533 2862 4567
rect 2896 4533 2912 4567
rect 2850 4524 2912 4533
rect 2350 4486 2716 4490
rect 2798 4486 2864 4494
rect 2350 4458 2758 4486
rect 2350 4420 2378 4458
rect 2672 4439 2758 4458
rect 2350 4412 2416 4420
rect 2350 4378 2365 4412
rect 2399 4378 2416 4412
rect 2350 4366 2416 4378
rect 2522 4416 2590 4422
rect 2522 4364 2532 4416
rect 2584 4364 2590 4416
rect 2522 4358 2590 4364
rect 2672 4405 2718 4439
rect 2752 4405 2758 4439
rect 2798 4434 2804 4486
rect 2856 4434 2864 4486
rect 2798 4426 2814 4434
rect 2672 4367 2758 4405
rect 2672 4333 2718 4367
rect 2752 4333 2758 4367
rect 2432 4304 2500 4310
rect 2432 4252 2440 4304
rect 2492 4252 2500 4304
rect 2432 4242 2500 4252
rect 2672 4286 2758 4333
rect 2808 4405 2814 4426
rect 2848 4426 2864 4434
rect 2904 4454 3232 4486
rect 2904 4439 3000 4454
rect 2848 4405 2854 4426
rect 2808 4367 2854 4405
rect 2808 4333 2814 4367
rect 2848 4333 2854 4367
rect 2808 4286 2854 4333
rect 2904 4405 2910 4439
rect 2944 4405 3000 4439
rect 3204 4418 3232 4454
rect 2904 4367 3000 4405
rect 2904 4333 2910 4367
rect 2944 4333 3000 4367
rect 3162 4410 3232 4418
rect 3162 4376 3177 4410
rect 3211 4376 3232 4410
rect 3162 4358 3232 4376
rect 3338 4418 3402 4424
rect 3338 4366 3344 4418
rect 3396 4366 3402 4418
rect 3338 4360 3402 4366
rect 2904 4286 3000 4333
rect 2330 4171 2606 4202
rect 2330 4137 2359 4171
rect 2393 4137 2451 4171
rect 2485 4137 2543 4171
rect 2577 4137 2606 4171
rect 2330 4106 2606 4137
rect 2672 4086 2722 4286
rect 2754 4239 2812 4254
rect 2754 4205 2766 4239
rect 2800 4205 2812 4239
rect 2754 4188 2812 4205
rect 2866 4158 2924 4176
rect 2866 4124 2878 4158
rect 2912 4124 2924 4158
rect 2866 4114 2924 4124
rect 2954 4086 3000 4286
rect 3250 4302 3314 4308
rect 3250 4250 3256 4302
rect 3308 4250 3314 4302
rect 3250 4244 3314 4250
rect 3144 4171 3420 4202
rect 3144 4137 3173 4171
rect 3207 4137 3265 4171
rect 3299 4137 3357 4171
rect 3391 4137 3420 4171
rect 3144 4134 3420 4137
rect 2312 4069 2376 4076
rect 2312 4036 2318 4069
rect 2370 4036 2376 4069
rect 2488 4069 2552 4076
rect 2488 4036 2494 4069
rect 2370 4017 2494 4036
rect 2546 4017 2552 4069
rect 2318 4008 2552 4017
rect 2672 4074 2774 4086
rect 2672 4040 2734 4074
rect 2768 4040 2774 4074
rect 2672 4002 2774 4040
rect 2824 4074 2870 4086
rect 2824 4040 2830 4074
rect 2864 4040 2870 4074
rect 2824 4020 2870 4040
rect 2920 4074 3000 4086
rect 2920 4040 2926 4074
rect 2960 4040 3000 4074
rect 2672 3970 2734 4002
rect 2468 3968 2734 3970
rect 2768 3968 2774 4002
rect 2468 3956 2774 3968
rect 2814 4014 2880 4020
rect 2814 3962 2822 4014
rect 2874 3962 2880 4014
rect 2814 3956 2880 3962
rect 2920 4002 3000 4040
rect 2920 3968 2926 4002
rect 2960 3968 3000 4002
rect 3116 4106 3420 4134
rect 2920 3956 2966 3968
rect 2468 3942 2722 3956
rect 2312 3936 2378 3942
rect 2312 3884 2320 3936
rect 2372 3884 2378 3936
rect 2312 3878 2378 3884
rect 1460 3669 1490 3672
rect 1542 3669 2084 3672
rect 1460 3635 1489 3669
rect 1542 3635 1581 3669
rect 1615 3635 1673 3669
rect 1707 3667 2084 3669
rect 1707 3635 1835 3667
rect 1460 3620 1490 3635
rect 1542 3633 1835 3635
rect 1869 3633 1927 3667
rect 1961 3633 2019 3667
rect 2053 3633 2084 3667
rect 1542 3620 2084 3633
rect 1460 3602 2084 3620
rect 2152 3678 2428 3692
rect 2152 3661 2344 3678
rect 2396 3661 2428 3678
rect 2152 3627 2181 3661
rect 2215 3627 2273 3661
rect 2307 3627 2344 3661
rect 2399 3627 2428 3661
rect 2152 3626 2344 3627
rect 2396 3626 2428 3627
rect 2152 3596 2428 3626
rect 2468 3592 2496 3942
rect 2768 3918 2832 3928
rect 2768 3884 2782 3918
rect 2816 3884 3088 3918
rect 2768 3866 2832 3884
rect 2684 3820 2756 3832
rect 2684 3768 2694 3820
rect 2746 3768 2756 3820
rect 2684 3756 2756 3768
rect 3054 3702 3088 3884
rect 3116 3802 3144 4106
rect 3116 3792 3184 3802
rect 3116 3758 3132 3792
rect 3166 3758 3184 3792
rect 3116 3744 3184 3758
rect 2528 3674 3088 3702
rect 2528 3671 2594 3674
rect 2528 3637 2544 3671
rect 2578 3637 2594 3671
rect 2528 3628 2594 3637
rect 2762 3619 2852 3640
rect 960 3511 1200 3528
rect 1244 3584 1310 3590
rect 1244 3532 1252 3584
rect 1304 3532 1310 3584
rect 1244 3526 1258 3532
rect 694 3471 740 3504
rect 694 3437 700 3471
rect 734 3437 740 3471
rect 960 3477 972 3511
rect 1006 3500 1200 3511
rect 1252 3509 1258 3526
rect 1292 3526 1310 3532
rect 1340 3543 1386 3590
rect 2468 3564 2540 3592
rect 1292 3509 1298 3526
rect 1006 3477 1198 3500
rect 960 3468 1198 3477
rect 694 3390 740 3437
rect 908 3430 974 3438
rect 822 3426 868 3430
rect -62 3368 10 3372
rect -602 3343 -536 3356
rect -602 3309 -586 3343
rect -552 3309 -536 3343
rect -602 3300 -536 3309
rect -62 3316 -53 3368
rect -1 3316 10 3368
rect -62 3304 10 3316
rect 134 3366 208 3386
rect 782 3383 868 3426
rect 134 3332 146 3366
rect 180 3332 208 3366
rect 134 3308 208 3332
rect 244 3372 312 3378
rect 244 3320 251 3372
rect 303 3366 312 3372
rect 303 3360 396 3366
rect 303 3326 342 3360
rect 376 3326 396 3360
rect 303 3320 396 3326
rect 244 3316 396 3320
rect 640 3343 706 3354
rect 244 3314 312 3316
rect 640 3309 656 3343
rect 690 3309 706 3343
rect 640 3296 706 3309
rect 782 3349 828 3383
rect 862 3349 868 3383
rect 908 3378 914 3430
rect 966 3378 974 3430
rect 908 3370 924 3378
rect 782 3311 868 3349
rect 782 3277 828 3311
rect 862 3277 868 3311
rect -280 3256 -222 3270
rect -280 3236 -268 3256
rect -750 3222 -268 3236
rect -234 3222 -222 3256
rect -750 3202 -222 3222
rect 782 3230 868 3277
rect 918 3349 924 3370
rect 958 3370 974 3378
rect 1014 3383 1110 3430
rect 958 3349 964 3370
rect 918 3311 964 3349
rect 918 3277 924 3311
rect 958 3277 964 3311
rect 918 3230 964 3277
rect 1014 3349 1020 3383
rect 1054 3349 1110 3383
rect 1014 3311 1110 3349
rect 1014 3277 1020 3311
rect 1054 3277 1110 3311
rect 1014 3230 1110 3277
rect -858 2900 -812 2912
rect -750 2872 -690 3202
rect 782 3176 832 3230
rect -644 3152 -568 3158
rect -644 3100 -636 3152
rect -584 3100 -568 3152
rect -644 3094 -568 3100
rect -428 3125 194 3156
rect -1010 2862 -690 2872
rect -1010 2828 -996 2862
rect -962 2828 -690 2862
rect -1010 2810 -690 2828
rect -428 3091 -399 3125
rect -365 3091 -307 3125
rect -273 3091 -215 3125
rect -181 3123 194 3125
rect -181 3091 -53 3123
rect -428 3089 -53 3091
rect -19 3089 39 3123
rect 73 3089 131 3123
rect 165 3089 194 3123
rect -428 3058 194 3089
rect 264 3130 540 3148
rect 264 3117 387 3130
rect 439 3117 540 3130
rect 616 3126 674 3134
rect 264 3083 293 3117
rect 327 3083 385 3117
rect 439 3083 477 3117
rect 511 3083 540 3117
rect 264 3078 387 3083
rect 439 3078 540 3083
rect -428 2782 -330 3058
rect 264 3052 540 3078
rect 608 3120 682 3126
rect 608 3068 619 3120
rect 671 3068 682 3120
rect 762 3110 832 3176
rect 864 3183 922 3198
rect 864 3149 876 3183
rect 910 3149 922 3183
rect 864 3132 922 3149
rect 608 3062 682 3068
rect 616 3056 674 3062
rect 332 2782 416 3052
rect 782 3030 832 3110
rect 976 3102 1034 3120
rect 976 3068 988 3102
rect 1022 3068 1034 3102
rect 976 3058 1034 3068
rect 1064 3030 1110 3230
rect 782 3018 884 3030
rect 782 2984 844 3018
rect 878 2984 884 3018
rect 782 2946 884 2984
rect 934 3018 980 3030
rect 934 2984 940 3018
rect 974 2984 980 3018
rect 934 2964 980 2984
rect 1030 3018 1110 3030
rect 1030 2984 1036 3018
rect 1070 2984 1110 3018
rect 782 2912 844 2946
rect 878 2912 884 2946
rect 782 2900 884 2912
rect 924 2958 990 2964
rect 924 2906 932 2958
rect 984 2906 990 2958
rect 924 2900 990 2906
rect 1030 2946 1110 2984
rect 1030 2912 1036 2946
rect 1070 2912 1110 2946
rect 1138 3236 1198 3468
rect 1252 3471 1298 3509
rect 1252 3437 1258 3471
rect 1292 3437 1298 3471
rect 1252 3390 1298 3437
rect 1340 3509 1346 3543
rect 1380 3509 1386 3543
rect 1340 3471 1386 3509
rect 1340 3437 1346 3471
rect 1380 3437 1386 3471
rect 1340 3390 1386 3437
rect 2494 3543 2540 3564
rect 2494 3509 2500 3543
rect 2534 3509 2540 3543
rect 2494 3471 2540 3509
rect 2494 3437 2500 3471
rect 2534 3437 2540 3471
rect 2494 3390 2540 3437
rect 2582 3570 2628 3590
rect 2762 3585 2791 3619
rect 2825 3585 2852 3619
rect 2582 3564 2650 3570
rect 2762 3564 2852 3585
rect 2582 3543 2590 3564
rect 2582 3509 2588 3543
rect 2642 3512 2650 3564
rect 2622 3509 2650 3512
rect 2582 3504 2650 3509
rect 2848 3528 2906 3530
rect 3054 3528 3088 3674
rect 3174 3671 3240 3682
rect 3174 3637 3190 3671
rect 3224 3637 3240 3671
rect 3174 3626 3240 3637
rect 3348 3672 3972 3704
rect 4060 3692 4138 4650
rect 4652 4641 4681 4650
rect 4715 4650 6569 4675
rect 4715 4641 4742 4650
rect 4652 4620 4742 4641
rect 4738 4584 4796 4586
rect 4738 4567 4800 4584
rect 4738 4533 4750 4567
rect 4784 4533 4800 4567
rect 4738 4524 4800 4533
rect 4238 4486 4604 4490
rect 4686 4486 4752 4494
rect 4238 4458 4646 4486
rect 4238 4420 4266 4458
rect 4560 4439 4646 4458
rect 4238 4412 4304 4420
rect 4238 4378 4253 4412
rect 4287 4378 4304 4412
rect 4238 4366 4304 4378
rect 4410 4416 4478 4422
rect 4410 4364 4420 4416
rect 4472 4364 4478 4416
rect 4410 4358 4478 4364
rect 4560 4405 4606 4439
rect 4640 4405 4646 4439
rect 4686 4434 4692 4486
rect 4744 4434 4752 4486
rect 4686 4426 4702 4434
rect 4560 4367 4646 4405
rect 4560 4333 4606 4367
rect 4640 4333 4646 4367
rect 4320 4304 4388 4310
rect 4320 4252 4328 4304
rect 4380 4252 4388 4304
rect 4320 4242 4388 4252
rect 4560 4286 4646 4333
rect 4696 4405 4702 4426
rect 4736 4426 4752 4434
rect 4792 4454 5120 4486
rect 4792 4439 4888 4454
rect 4736 4405 4742 4426
rect 4696 4367 4742 4405
rect 4696 4333 4702 4367
rect 4736 4333 4742 4367
rect 4696 4286 4742 4333
rect 4792 4405 4798 4439
rect 4832 4405 4888 4439
rect 5092 4418 5120 4454
rect 4792 4367 4888 4405
rect 4792 4333 4798 4367
rect 4832 4333 4888 4367
rect 5050 4410 5120 4418
rect 5050 4376 5065 4410
rect 5099 4376 5120 4410
rect 5050 4358 5120 4376
rect 5226 4418 5290 4424
rect 5226 4366 5232 4418
rect 5284 4366 5290 4418
rect 5226 4360 5290 4366
rect 4792 4286 4888 4333
rect 4218 4171 4494 4202
rect 4218 4137 4247 4171
rect 4281 4137 4339 4171
rect 4373 4137 4431 4171
rect 4465 4137 4494 4171
rect 4218 4106 4494 4137
rect 4560 4086 4610 4286
rect 4642 4239 4700 4254
rect 4642 4205 4654 4239
rect 4688 4205 4700 4239
rect 4642 4188 4700 4205
rect 4754 4158 4812 4176
rect 4754 4124 4766 4158
rect 4800 4124 4812 4158
rect 4754 4114 4812 4124
rect 4842 4086 4888 4286
rect 5138 4302 5202 4308
rect 5138 4250 5144 4302
rect 5196 4250 5202 4302
rect 5138 4244 5202 4250
rect 5032 4171 5308 4202
rect 5032 4137 5061 4171
rect 5095 4137 5153 4171
rect 5187 4137 5245 4171
rect 5279 4137 5308 4171
rect 5032 4134 5308 4137
rect 4200 4069 4264 4076
rect 4200 4036 4206 4069
rect 4258 4036 4264 4069
rect 4376 4069 4440 4076
rect 4376 4036 4382 4069
rect 4258 4017 4382 4036
rect 4434 4017 4440 4069
rect 4206 4008 4440 4017
rect 4560 4074 4662 4086
rect 4560 4040 4622 4074
rect 4656 4040 4662 4074
rect 4560 4002 4662 4040
rect 4712 4074 4758 4086
rect 4712 4040 4718 4074
rect 4752 4040 4758 4074
rect 4712 4020 4758 4040
rect 4808 4074 4888 4086
rect 4808 4040 4814 4074
rect 4848 4040 4888 4074
rect 4560 3970 4622 4002
rect 4356 3968 4622 3970
rect 4656 3968 4662 4002
rect 4356 3956 4662 3968
rect 4702 4014 4768 4020
rect 4702 3962 4710 4014
rect 4762 3962 4768 4014
rect 4702 3956 4768 3962
rect 4808 4002 4888 4040
rect 4808 3968 4814 4002
rect 4848 3968 4888 4002
rect 5004 4106 5308 4134
rect 4808 3956 4854 3968
rect 4356 3942 4610 3956
rect 4200 3936 4266 3942
rect 4200 3884 4208 3936
rect 4260 3884 4266 3936
rect 4200 3878 4266 3884
rect 3348 3669 3378 3672
rect 3430 3669 3972 3672
rect 3348 3635 3377 3669
rect 3430 3635 3469 3669
rect 3503 3635 3561 3669
rect 3595 3667 3972 3669
rect 3595 3635 3723 3667
rect 3348 3620 3378 3635
rect 3430 3633 3723 3635
rect 3757 3633 3815 3667
rect 3849 3633 3907 3667
rect 3941 3633 3972 3667
rect 3430 3620 3972 3633
rect 3348 3602 3972 3620
rect 4040 3678 4316 3692
rect 4040 3661 4232 3678
rect 4284 3661 4316 3678
rect 4040 3627 4069 3661
rect 4103 3627 4161 3661
rect 4195 3627 4232 3661
rect 4287 3627 4316 3661
rect 4040 3626 4232 3627
rect 4284 3626 4316 3627
rect 4040 3596 4316 3626
rect 4356 3592 4384 3942
rect 4656 3918 4720 3928
rect 4656 3884 4670 3918
rect 4704 3884 4976 3918
rect 4656 3866 4720 3884
rect 4572 3820 4644 3832
rect 4572 3768 4582 3820
rect 4634 3768 4644 3820
rect 4572 3756 4644 3768
rect 4942 3702 4976 3884
rect 5004 3802 5032 4106
rect 5004 3792 5072 3802
rect 5004 3758 5020 3792
rect 5054 3758 5072 3792
rect 5004 3744 5072 3758
rect 4416 3674 4976 3702
rect 4416 3671 4482 3674
rect 4416 3637 4432 3671
rect 4466 3637 4482 3671
rect 4416 3628 4482 3637
rect 4650 3619 4740 3640
rect 2848 3511 3088 3528
rect 3132 3584 3198 3590
rect 3132 3532 3140 3584
rect 3192 3532 3198 3584
rect 3132 3526 3146 3532
rect 2582 3471 2628 3504
rect 2582 3437 2588 3471
rect 2622 3437 2628 3471
rect 2848 3477 2860 3511
rect 2894 3500 3088 3511
rect 3140 3509 3146 3526
rect 3180 3526 3198 3532
rect 3228 3543 3274 3590
rect 4356 3564 4428 3592
rect 3180 3509 3186 3526
rect 2894 3477 3086 3500
rect 2848 3468 3086 3477
rect 2582 3390 2628 3437
rect 2796 3430 2862 3438
rect 2710 3426 2756 3430
rect 1826 3368 1898 3372
rect 1286 3343 1352 3356
rect 1286 3309 1302 3343
rect 1336 3309 1352 3343
rect 1286 3300 1352 3309
rect 1826 3316 1835 3368
rect 1887 3316 1898 3368
rect 1826 3304 1898 3316
rect 2022 3366 2096 3386
rect 2670 3383 2756 3426
rect 2022 3332 2034 3366
rect 2068 3332 2096 3366
rect 2022 3308 2096 3332
rect 2132 3372 2200 3378
rect 2132 3320 2139 3372
rect 2191 3366 2200 3372
rect 2191 3360 2284 3366
rect 2191 3326 2230 3360
rect 2264 3326 2284 3360
rect 2191 3320 2284 3326
rect 2132 3316 2284 3320
rect 2528 3343 2594 3354
rect 2132 3314 2200 3316
rect 2528 3309 2544 3343
rect 2578 3309 2594 3343
rect 2528 3296 2594 3309
rect 2670 3349 2716 3383
rect 2750 3349 2756 3383
rect 2796 3378 2802 3430
rect 2854 3378 2862 3430
rect 2796 3370 2812 3378
rect 2670 3311 2756 3349
rect 2670 3277 2716 3311
rect 2750 3277 2756 3311
rect 1608 3256 1666 3270
rect 1608 3236 1620 3256
rect 1138 3222 1620 3236
rect 1654 3222 1666 3256
rect 1138 3202 1666 3222
rect 2670 3230 2756 3277
rect 2806 3349 2812 3370
rect 2846 3370 2862 3378
rect 2902 3383 2998 3430
rect 2846 3349 2852 3370
rect 2806 3311 2852 3349
rect 2806 3277 2812 3311
rect 2846 3277 2852 3311
rect 2806 3230 2852 3277
rect 2902 3349 2908 3383
rect 2942 3349 2998 3383
rect 2902 3311 2998 3349
rect 2902 3277 2908 3311
rect 2942 3277 2998 3311
rect 2902 3230 2998 3277
rect 1030 2900 1076 2912
rect 1138 2872 1198 3202
rect 2670 3176 2720 3230
rect 1244 3152 1320 3158
rect 1244 3100 1252 3152
rect 1304 3100 1320 3152
rect 1244 3094 1320 3100
rect 1460 3125 2082 3156
rect 878 2862 1198 2872
rect 878 2828 892 2862
rect 926 2828 1198 2862
rect 878 2810 1198 2828
rect 1460 3091 1489 3125
rect 1523 3091 1581 3125
rect 1615 3091 1673 3125
rect 1707 3123 2082 3125
rect 1707 3091 1835 3123
rect 1460 3089 1835 3091
rect 1869 3089 1927 3123
rect 1961 3089 2019 3123
rect 2053 3089 2082 3123
rect 1460 3058 2082 3089
rect 2152 3130 2428 3148
rect 2152 3117 2275 3130
rect 2327 3117 2428 3130
rect 2504 3126 2562 3134
rect 2152 3083 2181 3117
rect 2215 3083 2273 3117
rect 2327 3083 2365 3117
rect 2399 3083 2428 3117
rect 2152 3078 2275 3083
rect 2327 3078 2428 3083
rect 1460 2782 1558 3058
rect 2152 3052 2428 3078
rect 2496 3120 2570 3126
rect 2496 3068 2507 3120
rect 2559 3068 2570 3120
rect 2650 3110 2720 3176
rect 2752 3183 2810 3198
rect 2752 3149 2764 3183
rect 2798 3149 2810 3183
rect 2752 3132 2810 3149
rect 2496 3062 2570 3068
rect 2504 3056 2562 3062
rect 2220 2782 2304 3052
rect 2670 3030 2720 3110
rect 2864 3102 2922 3120
rect 2864 3068 2876 3102
rect 2910 3068 2922 3102
rect 2864 3058 2922 3068
rect 2952 3030 2998 3230
rect 2670 3018 2772 3030
rect 2670 2984 2732 3018
rect 2766 2984 2772 3018
rect 2670 2946 2772 2984
rect 2822 3018 2868 3030
rect 2822 2984 2828 3018
rect 2862 2984 2868 3018
rect 2822 2964 2868 2984
rect 2918 3018 2998 3030
rect 2918 2984 2924 3018
rect 2958 2984 2998 3018
rect 2670 2912 2732 2946
rect 2766 2912 2772 2946
rect 2670 2900 2772 2912
rect 2812 2958 2878 2964
rect 2812 2906 2820 2958
rect 2872 2906 2878 2958
rect 2812 2900 2878 2906
rect 2918 2946 2998 2984
rect 2918 2912 2924 2946
rect 2958 2912 2998 2946
rect 3026 3236 3086 3468
rect 3140 3471 3186 3509
rect 3140 3437 3146 3471
rect 3180 3437 3186 3471
rect 3140 3390 3186 3437
rect 3228 3509 3234 3543
rect 3268 3509 3274 3543
rect 3228 3471 3274 3509
rect 3228 3437 3234 3471
rect 3268 3437 3274 3471
rect 3228 3390 3274 3437
rect 4382 3543 4428 3564
rect 4382 3509 4388 3543
rect 4422 3509 4428 3543
rect 4382 3471 4428 3509
rect 4382 3437 4388 3471
rect 4422 3437 4428 3471
rect 4382 3390 4428 3437
rect 4470 3570 4516 3590
rect 4650 3585 4679 3619
rect 4713 3585 4740 3619
rect 4470 3564 4538 3570
rect 4650 3564 4740 3585
rect 4470 3543 4478 3564
rect 4470 3509 4476 3543
rect 4530 3512 4538 3564
rect 4510 3509 4538 3512
rect 4470 3504 4538 3509
rect 4736 3528 4794 3530
rect 4942 3528 4976 3674
rect 5062 3671 5128 3682
rect 5062 3637 5078 3671
rect 5112 3637 5128 3671
rect 5062 3626 5128 3637
rect 5236 3672 5860 3704
rect 5948 3692 6026 4650
rect 6540 4641 6569 4650
rect 6603 4650 8457 4675
rect 6603 4641 6630 4650
rect 6540 4620 6630 4641
rect 6626 4584 6684 4586
rect 6626 4567 6688 4584
rect 6626 4533 6638 4567
rect 6672 4533 6688 4567
rect 6626 4524 6688 4533
rect 6126 4486 6492 4490
rect 6574 4486 6640 4494
rect 6126 4458 6534 4486
rect 6126 4420 6154 4458
rect 6448 4439 6534 4458
rect 6126 4412 6192 4420
rect 6126 4378 6141 4412
rect 6175 4378 6192 4412
rect 6126 4366 6192 4378
rect 6298 4416 6366 4422
rect 6298 4364 6308 4416
rect 6360 4364 6366 4416
rect 6298 4358 6366 4364
rect 6448 4405 6494 4439
rect 6528 4405 6534 4439
rect 6574 4434 6580 4486
rect 6632 4434 6640 4486
rect 6574 4426 6590 4434
rect 6448 4367 6534 4405
rect 6448 4333 6494 4367
rect 6528 4333 6534 4367
rect 6208 4304 6276 4310
rect 6208 4252 6216 4304
rect 6268 4252 6276 4304
rect 6208 4242 6276 4252
rect 6448 4286 6534 4333
rect 6584 4405 6590 4426
rect 6624 4426 6640 4434
rect 6680 4454 7008 4486
rect 6680 4439 6776 4454
rect 6624 4405 6630 4426
rect 6584 4367 6630 4405
rect 6584 4333 6590 4367
rect 6624 4333 6630 4367
rect 6584 4286 6630 4333
rect 6680 4405 6686 4439
rect 6720 4405 6776 4439
rect 6980 4418 7008 4454
rect 6680 4367 6776 4405
rect 6680 4333 6686 4367
rect 6720 4333 6776 4367
rect 6938 4410 7008 4418
rect 6938 4376 6953 4410
rect 6987 4376 7008 4410
rect 6938 4358 7008 4376
rect 7114 4418 7178 4424
rect 7114 4366 7120 4418
rect 7172 4366 7178 4418
rect 7114 4360 7178 4366
rect 6680 4286 6776 4333
rect 6106 4171 6382 4202
rect 6106 4137 6135 4171
rect 6169 4137 6227 4171
rect 6261 4137 6319 4171
rect 6353 4137 6382 4171
rect 6106 4106 6382 4137
rect 6448 4086 6498 4286
rect 6530 4239 6588 4254
rect 6530 4205 6542 4239
rect 6576 4205 6588 4239
rect 6530 4188 6588 4205
rect 6642 4158 6700 4176
rect 6642 4124 6654 4158
rect 6688 4124 6700 4158
rect 6642 4114 6700 4124
rect 6730 4086 6776 4286
rect 7026 4302 7090 4308
rect 7026 4250 7032 4302
rect 7084 4250 7090 4302
rect 7026 4244 7090 4250
rect 6920 4171 7196 4202
rect 6920 4137 6949 4171
rect 6983 4137 7041 4171
rect 7075 4137 7133 4171
rect 7167 4137 7196 4171
rect 6920 4134 7196 4137
rect 6088 4069 6152 4076
rect 6088 4036 6094 4069
rect 6146 4036 6152 4069
rect 6264 4069 6328 4076
rect 6264 4036 6270 4069
rect 6146 4017 6270 4036
rect 6322 4017 6328 4069
rect 6094 4008 6328 4017
rect 6448 4074 6550 4086
rect 6448 4040 6510 4074
rect 6544 4040 6550 4074
rect 6448 4002 6550 4040
rect 6600 4074 6646 4086
rect 6600 4040 6606 4074
rect 6640 4040 6646 4074
rect 6600 4020 6646 4040
rect 6696 4074 6776 4086
rect 6696 4040 6702 4074
rect 6736 4040 6776 4074
rect 6448 3970 6510 4002
rect 6244 3968 6510 3970
rect 6544 3968 6550 4002
rect 6244 3956 6550 3968
rect 6590 4014 6656 4020
rect 6590 3962 6598 4014
rect 6650 3962 6656 4014
rect 6590 3956 6656 3962
rect 6696 4002 6776 4040
rect 6696 3968 6702 4002
rect 6736 3968 6776 4002
rect 6892 4106 7196 4134
rect 6696 3956 6742 3968
rect 6244 3942 6498 3956
rect 6088 3936 6154 3942
rect 6088 3884 6096 3936
rect 6148 3884 6154 3936
rect 6088 3878 6154 3884
rect 5236 3669 5266 3672
rect 5318 3669 5860 3672
rect 5236 3635 5265 3669
rect 5318 3635 5357 3669
rect 5391 3635 5449 3669
rect 5483 3667 5860 3669
rect 5483 3635 5611 3667
rect 5236 3620 5266 3635
rect 5318 3633 5611 3635
rect 5645 3633 5703 3667
rect 5737 3633 5795 3667
rect 5829 3633 5860 3667
rect 5318 3620 5860 3633
rect 5236 3602 5860 3620
rect 5928 3678 6204 3692
rect 5928 3661 6120 3678
rect 6172 3661 6204 3678
rect 5928 3627 5957 3661
rect 5991 3627 6049 3661
rect 6083 3627 6120 3661
rect 6175 3627 6204 3661
rect 5928 3626 6120 3627
rect 6172 3626 6204 3627
rect 5928 3596 6204 3626
rect 6244 3592 6272 3942
rect 6544 3918 6608 3928
rect 6544 3884 6558 3918
rect 6592 3884 6864 3918
rect 6544 3866 6608 3884
rect 6460 3820 6532 3832
rect 6460 3768 6470 3820
rect 6522 3768 6532 3820
rect 6460 3756 6532 3768
rect 6830 3702 6864 3884
rect 6892 3802 6920 4106
rect 6892 3792 6960 3802
rect 6892 3758 6908 3792
rect 6942 3758 6960 3792
rect 6892 3744 6960 3758
rect 6304 3674 6864 3702
rect 6304 3671 6370 3674
rect 6304 3637 6320 3671
rect 6354 3637 6370 3671
rect 6304 3628 6370 3637
rect 6538 3619 6628 3640
rect 4736 3511 4976 3528
rect 5020 3584 5086 3590
rect 5020 3532 5028 3584
rect 5080 3532 5086 3584
rect 5020 3526 5034 3532
rect 4470 3471 4516 3504
rect 4470 3437 4476 3471
rect 4510 3437 4516 3471
rect 4736 3477 4748 3511
rect 4782 3500 4976 3511
rect 5028 3509 5034 3526
rect 5068 3526 5086 3532
rect 5116 3543 5162 3590
rect 6244 3564 6316 3592
rect 5068 3509 5074 3526
rect 4782 3477 4974 3500
rect 4736 3468 4974 3477
rect 4470 3390 4516 3437
rect 4684 3430 4750 3438
rect 4598 3426 4644 3430
rect 3714 3368 3786 3372
rect 3174 3343 3240 3356
rect 3174 3309 3190 3343
rect 3224 3309 3240 3343
rect 3174 3300 3240 3309
rect 3714 3316 3723 3368
rect 3775 3316 3786 3368
rect 3714 3304 3786 3316
rect 3910 3366 3984 3386
rect 4558 3383 4644 3426
rect 3910 3332 3922 3366
rect 3956 3332 3984 3366
rect 3910 3308 3984 3332
rect 4020 3372 4088 3378
rect 4020 3320 4027 3372
rect 4079 3366 4088 3372
rect 4079 3360 4172 3366
rect 4079 3326 4118 3360
rect 4152 3326 4172 3360
rect 4079 3320 4172 3326
rect 4020 3316 4172 3320
rect 4416 3343 4482 3354
rect 4020 3314 4088 3316
rect 4416 3309 4432 3343
rect 4466 3309 4482 3343
rect 4416 3296 4482 3309
rect 4558 3349 4604 3383
rect 4638 3349 4644 3383
rect 4684 3378 4690 3430
rect 4742 3378 4750 3430
rect 4684 3370 4700 3378
rect 4558 3311 4644 3349
rect 4558 3277 4604 3311
rect 4638 3277 4644 3311
rect 3496 3256 3554 3270
rect 3496 3236 3508 3256
rect 3026 3222 3508 3236
rect 3542 3222 3554 3256
rect 3026 3202 3554 3222
rect 4558 3230 4644 3277
rect 4694 3349 4700 3370
rect 4734 3370 4750 3378
rect 4790 3383 4886 3430
rect 4734 3349 4740 3370
rect 4694 3311 4740 3349
rect 4694 3277 4700 3311
rect 4734 3277 4740 3311
rect 4694 3230 4740 3277
rect 4790 3349 4796 3383
rect 4830 3349 4886 3383
rect 4790 3311 4886 3349
rect 4790 3277 4796 3311
rect 4830 3277 4886 3311
rect 4790 3230 4886 3277
rect 2918 2900 2964 2912
rect 3026 2872 3086 3202
rect 4558 3176 4608 3230
rect 3132 3152 3208 3158
rect 3132 3100 3140 3152
rect 3192 3100 3208 3152
rect 3132 3094 3208 3100
rect 3348 3125 3970 3156
rect 2766 2862 3086 2872
rect 2766 2828 2780 2862
rect 2814 2828 3086 2862
rect 2766 2810 3086 2828
rect 3348 3091 3377 3125
rect 3411 3091 3469 3125
rect 3503 3091 3561 3125
rect 3595 3123 3970 3125
rect 3595 3091 3723 3123
rect 3348 3089 3723 3091
rect 3757 3089 3815 3123
rect 3849 3089 3907 3123
rect 3941 3089 3970 3123
rect 3348 3058 3970 3089
rect 4040 3130 4316 3148
rect 4040 3117 4163 3130
rect 4215 3117 4316 3130
rect 4392 3126 4450 3134
rect 4040 3083 4069 3117
rect 4103 3083 4161 3117
rect 4215 3083 4253 3117
rect 4287 3083 4316 3117
rect 4040 3078 4163 3083
rect 4215 3078 4316 3083
rect 3348 2782 3446 3058
rect 4040 3052 4316 3078
rect 4384 3120 4458 3126
rect 4384 3068 4395 3120
rect 4447 3068 4458 3120
rect 4538 3110 4608 3176
rect 4640 3183 4698 3198
rect 4640 3149 4652 3183
rect 4686 3149 4698 3183
rect 4640 3132 4698 3149
rect 4384 3062 4458 3068
rect 4392 3056 4450 3062
rect 4108 2782 4192 3052
rect 4558 3030 4608 3110
rect 4752 3102 4810 3120
rect 4752 3068 4764 3102
rect 4798 3068 4810 3102
rect 4752 3058 4810 3068
rect 4840 3030 4886 3230
rect 4558 3018 4660 3030
rect 4558 2984 4620 3018
rect 4654 2984 4660 3018
rect 4558 2946 4660 2984
rect 4710 3018 4756 3030
rect 4710 2984 4716 3018
rect 4750 2984 4756 3018
rect 4710 2964 4756 2984
rect 4806 3018 4886 3030
rect 4806 2984 4812 3018
rect 4846 2984 4886 3018
rect 4558 2912 4620 2946
rect 4654 2912 4660 2946
rect 4558 2900 4660 2912
rect 4700 2958 4766 2964
rect 4700 2906 4708 2958
rect 4760 2906 4766 2958
rect 4700 2900 4766 2906
rect 4806 2946 4886 2984
rect 4806 2912 4812 2946
rect 4846 2912 4886 2946
rect 4914 3236 4974 3468
rect 5028 3471 5074 3509
rect 5028 3437 5034 3471
rect 5068 3437 5074 3471
rect 5028 3390 5074 3437
rect 5116 3509 5122 3543
rect 5156 3509 5162 3543
rect 5116 3471 5162 3509
rect 5116 3437 5122 3471
rect 5156 3437 5162 3471
rect 5116 3390 5162 3437
rect 6270 3543 6316 3564
rect 6270 3509 6276 3543
rect 6310 3509 6316 3543
rect 6270 3471 6316 3509
rect 6270 3437 6276 3471
rect 6310 3437 6316 3471
rect 6270 3390 6316 3437
rect 6358 3570 6404 3590
rect 6538 3585 6567 3619
rect 6601 3585 6628 3619
rect 6358 3564 6426 3570
rect 6538 3564 6628 3585
rect 6358 3543 6366 3564
rect 6358 3509 6364 3543
rect 6418 3512 6426 3564
rect 6398 3509 6426 3512
rect 6358 3504 6426 3509
rect 6624 3528 6682 3530
rect 6830 3528 6864 3674
rect 6950 3671 7016 3682
rect 6950 3637 6966 3671
rect 7000 3637 7016 3671
rect 6950 3626 7016 3637
rect 7124 3672 7748 3704
rect 7836 3692 7914 4650
rect 8428 4641 8457 4650
rect 8491 4650 10345 4675
rect 8491 4641 8518 4650
rect 8428 4620 8518 4641
rect 8514 4584 8572 4586
rect 8514 4567 8576 4584
rect 8514 4533 8526 4567
rect 8560 4533 8576 4567
rect 8514 4524 8576 4533
rect 8014 4486 8380 4490
rect 8462 4486 8528 4494
rect 8014 4458 8422 4486
rect 8014 4420 8042 4458
rect 8336 4439 8422 4458
rect 8014 4412 8080 4420
rect 8014 4378 8029 4412
rect 8063 4378 8080 4412
rect 8014 4366 8080 4378
rect 8186 4416 8254 4422
rect 8186 4364 8196 4416
rect 8248 4364 8254 4416
rect 8186 4358 8254 4364
rect 8336 4405 8382 4439
rect 8416 4405 8422 4439
rect 8462 4434 8468 4486
rect 8520 4434 8528 4486
rect 8462 4426 8478 4434
rect 8336 4367 8422 4405
rect 8336 4333 8382 4367
rect 8416 4333 8422 4367
rect 8096 4304 8164 4310
rect 8096 4252 8104 4304
rect 8156 4252 8164 4304
rect 8096 4242 8164 4252
rect 8336 4286 8422 4333
rect 8472 4405 8478 4426
rect 8512 4426 8528 4434
rect 8568 4454 8896 4486
rect 8568 4439 8664 4454
rect 8512 4405 8518 4426
rect 8472 4367 8518 4405
rect 8472 4333 8478 4367
rect 8512 4333 8518 4367
rect 8472 4286 8518 4333
rect 8568 4405 8574 4439
rect 8608 4405 8664 4439
rect 8868 4418 8896 4454
rect 8568 4367 8664 4405
rect 8568 4333 8574 4367
rect 8608 4333 8664 4367
rect 8826 4410 8896 4418
rect 8826 4376 8841 4410
rect 8875 4376 8896 4410
rect 8826 4358 8896 4376
rect 9002 4418 9066 4424
rect 9002 4366 9008 4418
rect 9060 4366 9066 4418
rect 9002 4360 9066 4366
rect 8568 4286 8664 4333
rect 7994 4171 8270 4202
rect 7994 4137 8023 4171
rect 8057 4137 8115 4171
rect 8149 4137 8207 4171
rect 8241 4137 8270 4171
rect 7994 4106 8270 4137
rect 8336 4086 8386 4286
rect 8418 4239 8476 4254
rect 8418 4205 8430 4239
rect 8464 4205 8476 4239
rect 8418 4188 8476 4205
rect 8530 4158 8588 4176
rect 8530 4124 8542 4158
rect 8576 4124 8588 4158
rect 8530 4114 8588 4124
rect 8618 4086 8664 4286
rect 8914 4302 8978 4308
rect 8914 4250 8920 4302
rect 8972 4250 8978 4302
rect 8914 4244 8978 4250
rect 8808 4171 9084 4202
rect 8808 4137 8837 4171
rect 8871 4137 8929 4171
rect 8963 4137 9021 4171
rect 9055 4137 9084 4171
rect 8808 4134 9084 4137
rect 7976 4069 8040 4076
rect 7976 4036 7982 4069
rect 8034 4036 8040 4069
rect 8152 4069 8216 4076
rect 8152 4036 8158 4069
rect 8034 4017 8158 4036
rect 8210 4017 8216 4069
rect 7982 4008 8216 4017
rect 8336 4074 8438 4086
rect 8336 4040 8398 4074
rect 8432 4040 8438 4074
rect 8336 4002 8438 4040
rect 8488 4074 8534 4086
rect 8488 4040 8494 4074
rect 8528 4040 8534 4074
rect 8488 4020 8534 4040
rect 8584 4074 8664 4086
rect 8584 4040 8590 4074
rect 8624 4040 8664 4074
rect 8336 3970 8398 4002
rect 8132 3968 8398 3970
rect 8432 3968 8438 4002
rect 8132 3956 8438 3968
rect 8478 4014 8544 4020
rect 8478 3962 8486 4014
rect 8538 3962 8544 4014
rect 8478 3956 8544 3962
rect 8584 4002 8664 4040
rect 8584 3968 8590 4002
rect 8624 3968 8664 4002
rect 8780 4106 9084 4134
rect 8584 3956 8630 3968
rect 8132 3942 8386 3956
rect 7976 3936 8042 3942
rect 7976 3884 7984 3936
rect 8036 3884 8042 3936
rect 7976 3878 8042 3884
rect 7124 3669 7154 3672
rect 7206 3669 7748 3672
rect 7124 3635 7153 3669
rect 7206 3635 7245 3669
rect 7279 3635 7337 3669
rect 7371 3667 7748 3669
rect 7371 3635 7499 3667
rect 7124 3620 7154 3635
rect 7206 3633 7499 3635
rect 7533 3633 7591 3667
rect 7625 3633 7683 3667
rect 7717 3633 7748 3667
rect 7206 3620 7748 3633
rect 7124 3602 7748 3620
rect 7816 3678 8092 3692
rect 7816 3661 8008 3678
rect 8060 3661 8092 3678
rect 7816 3627 7845 3661
rect 7879 3627 7937 3661
rect 7971 3627 8008 3661
rect 8063 3627 8092 3661
rect 7816 3626 8008 3627
rect 8060 3626 8092 3627
rect 7816 3596 8092 3626
rect 8132 3592 8160 3942
rect 8432 3918 8496 3928
rect 8432 3884 8446 3918
rect 8480 3884 8752 3918
rect 8432 3866 8496 3884
rect 8348 3820 8420 3832
rect 8348 3768 8358 3820
rect 8410 3768 8420 3820
rect 8348 3756 8420 3768
rect 8718 3702 8752 3884
rect 8780 3802 8808 4106
rect 8780 3792 8848 3802
rect 8780 3758 8796 3792
rect 8830 3758 8848 3792
rect 8780 3744 8848 3758
rect 8192 3674 8752 3702
rect 8192 3671 8258 3674
rect 8192 3637 8208 3671
rect 8242 3637 8258 3671
rect 8192 3628 8258 3637
rect 8426 3619 8516 3640
rect 6624 3511 6864 3528
rect 6908 3584 6974 3590
rect 6908 3532 6916 3584
rect 6968 3532 6974 3584
rect 6908 3526 6922 3532
rect 6358 3471 6404 3504
rect 6358 3437 6364 3471
rect 6398 3437 6404 3471
rect 6624 3477 6636 3511
rect 6670 3500 6864 3511
rect 6916 3509 6922 3526
rect 6956 3526 6974 3532
rect 7004 3543 7050 3590
rect 8132 3564 8204 3592
rect 6956 3509 6962 3526
rect 6670 3477 6862 3500
rect 6624 3468 6862 3477
rect 6358 3390 6404 3437
rect 6572 3430 6638 3438
rect 6486 3426 6532 3430
rect 5602 3368 5674 3372
rect 5062 3343 5128 3356
rect 5062 3309 5078 3343
rect 5112 3309 5128 3343
rect 5062 3300 5128 3309
rect 5602 3316 5611 3368
rect 5663 3316 5674 3368
rect 5602 3304 5674 3316
rect 5798 3366 5872 3386
rect 6446 3383 6532 3426
rect 5798 3332 5810 3366
rect 5844 3332 5872 3366
rect 5798 3308 5872 3332
rect 5908 3372 5976 3378
rect 5908 3320 5915 3372
rect 5967 3366 5976 3372
rect 5967 3360 6060 3366
rect 5967 3326 6006 3360
rect 6040 3326 6060 3360
rect 5967 3320 6060 3326
rect 5908 3316 6060 3320
rect 6304 3343 6370 3354
rect 5908 3314 5976 3316
rect 6304 3309 6320 3343
rect 6354 3309 6370 3343
rect 6304 3296 6370 3309
rect 6446 3349 6492 3383
rect 6526 3349 6532 3383
rect 6572 3378 6578 3430
rect 6630 3378 6638 3430
rect 6572 3370 6588 3378
rect 6446 3311 6532 3349
rect 6446 3277 6492 3311
rect 6526 3277 6532 3311
rect 5384 3256 5442 3270
rect 5384 3236 5396 3256
rect 4914 3222 5396 3236
rect 5430 3222 5442 3256
rect 4914 3202 5442 3222
rect 6446 3230 6532 3277
rect 6582 3349 6588 3370
rect 6622 3370 6638 3378
rect 6678 3383 6774 3430
rect 6622 3349 6628 3370
rect 6582 3311 6628 3349
rect 6582 3277 6588 3311
rect 6622 3277 6628 3311
rect 6582 3230 6628 3277
rect 6678 3349 6684 3383
rect 6718 3349 6774 3383
rect 6678 3311 6774 3349
rect 6678 3277 6684 3311
rect 6718 3277 6774 3311
rect 6678 3230 6774 3277
rect 4806 2900 4852 2912
rect 4914 2872 4974 3202
rect 6446 3176 6496 3230
rect 5020 3152 5096 3158
rect 5020 3100 5028 3152
rect 5080 3100 5096 3152
rect 5020 3094 5096 3100
rect 5236 3125 5858 3156
rect 4654 2862 4974 2872
rect 4654 2828 4668 2862
rect 4702 2828 4974 2862
rect 4654 2810 4974 2828
rect 5236 3091 5265 3125
rect 5299 3091 5357 3125
rect 5391 3091 5449 3125
rect 5483 3123 5858 3125
rect 5483 3091 5611 3123
rect 5236 3089 5611 3091
rect 5645 3089 5703 3123
rect 5737 3089 5795 3123
rect 5829 3089 5858 3123
rect 5236 3058 5858 3089
rect 5928 3130 6204 3148
rect 5928 3117 6051 3130
rect 6103 3117 6204 3130
rect 6280 3126 6338 3134
rect 5928 3083 5957 3117
rect 5991 3083 6049 3117
rect 6103 3083 6141 3117
rect 6175 3083 6204 3117
rect 5928 3078 6051 3083
rect 6103 3078 6204 3083
rect 5236 2782 5334 3058
rect 5928 3052 6204 3078
rect 6272 3120 6346 3126
rect 6272 3068 6283 3120
rect 6335 3068 6346 3120
rect 6426 3110 6496 3176
rect 6528 3183 6586 3198
rect 6528 3149 6540 3183
rect 6574 3149 6586 3183
rect 6528 3132 6586 3149
rect 6272 3062 6346 3068
rect 6280 3056 6338 3062
rect 5996 2782 6080 3052
rect 6446 3030 6496 3110
rect 6640 3102 6698 3120
rect 6640 3068 6652 3102
rect 6686 3068 6698 3102
rect 6640 3058 6698 3068
rect 6728 3030 6774 3230
rect 6446 3018 6548 3030
rect 6446 2984 6508 3018
rect 6542 2984 6548 3018
rect 6446 2946 6548 2984
rect 6598 3018 6644 3030
rect 6598 2984 6604 3018
rect 6638 2984 6644 3018
rect 6598 2964 6644 2984
rect 6694 3018 6774 3030
rect 6694 2984 6700 3018
rect 6734 2984 6774 3018
rect 6446 2912 6508 2946
rect 6542 2912 6548 2946
rect 6446 2900 6548 2912
rect 6588 2958 6654 2964
rect 6588 2906 6596 2958
rect 6648 2906 6654 2958
rect 6588 2900 6654 2906
rect 6694 2946 6774 2984
rect 6694 2912 6700 2946
rect 6734 2912 6774 2946
rect 6802 3236 6862 3468
rect 6916 3471 6962 3509
rect 6916 3437 6922 3471
rect 6956 3437 6962 3471
rect 6916 3390 6962 3437
rect 7004 3509 7010 3543
rect 7044 3509 7050 3543
rect 7004 3471 7050 3509
rect 7004 3437 7010 3471
rect 7044 3437 7050 3471
rect 7004 3390 7050 3437
rect 8158 3543 8204 3564
rect 8158 3509 8164 3543
rect 8198 3509 8204 3543
rect 8158 3471 8204 3509
rect 8158 3437 8164 3471
rect 8198 3437 8204 3471
rect 8158 3390 8204 3437
rect 8246 3570 8292 3590
rect 8426 3585 8455 3619
rect 8489 3585 8516 3619
rect 8246 3564 8314 3570
rect 8426 3564 8516 3585
rect 8246 3543 8254 3564
rect 8246 3509 8252 3543
rect 8306 3512 8314 3564
rect 8286 3509 8314 3512
rect 8246 3504 8314 3509
rect 8512 3528 8570 3530
rect 8718 3528 8752 3674
rect 8838 3671 8904 3682
rect 8838 3637 8854 3671
rect 8888 3637 8904 3671
rect 8838 3626 8904 3637
rect 9012 3672 9636 3704
rect 9724 3692 9802 4650
rect 10316 4641 10345 4650
rect 10379 4650 12227 4675
rect 10379 4641 10406 4650
rect 10316 4620 10406 4641
rect 10402 4584 10460 4586
rect 10402 4567 10464 4584
rect 10402 4533 10414 4567
rect 10448 4533 10464 4567
rect 10402 4524 10464 4533
rect 9902 4486 10268 4490
rect 10350 4486 10416 4494
rect 9902 4458 10310 4486
rect 9902 4420 9930 4458
rect 10224 4439 10310 4458
rect 9902 4412 9968 4420
rect 9902 4378 9917 4412
rect 9951 4378 9968 4412
rect 9902 4366 9968 4378
rect 10074 4416 10142 4422
rect 10074 4364 10084 4416
rect 10136 4364 10142 4416
rect 10074 4358 10142 4364
rect 10224 4405 10270 4439
rect 10304 4405 10310 4439
rect 10350 4434 10356 4486
rect 10408 4434 10416 4486
rect 10350 4426 10366 4434
rect 10224 4367 10310 4405
rect 10224 4333 10270 4367
rect 10304 4333 10310 4367
rect 9984 4304 10052 4310
rect 9984 4252 9992 4304
rect 10044 4252 10052 4304
rect 9984 4242 10052 4252
rect 10224 4286 10310 4333
rect 10360 4405 10366 4426
rect 10400 4426 10416 4434
rect 10456 4454 10784 4486
rect 10456 4439 10552 4454
rect 10400 4405 10406 4426
rect 10360 4367 10406 4405
rect 10360 4333 10366 4367
rect 10400 4333 10406 4367
rect 10360 4286 10406 4333
rect 10456 4405 10462 4439
rect 10496 4405 10552 4439
rect 10756 4418 10784 4454
rect 10456 4367 10552 4405
rect 10456 4333 10462 4367
rect 10496 4333 10552 4367
rect 10714 4410 10784 4418
rect 10714 4376 10729 4410
rect 10763 4376 10784 4410
rect 10714 4358 10784 4376
rect 10890 4418 10954 4424
rect 10890 4366 10896 4418
rect 10948 4366 10954 4418
rect 10890 4360 10954 4366
rect 10456 4286 10552 4333
rect 9882 4171 10158 4202
rect 9882 4137 9911 4171
rect 9945 4137 10003 4171
rect 10037 4137 10095 4171
rect 10129 4137 10158 4171
rect 9882 4106 10158 4137
rect 10224 4086 10274 4286
rect 10306 4239 10364 4254
rect 10306 4205 10318 4239
rect 10352 4205 10364 4239
rect 10306 4188 10364 4205
rect 10418 4158 10476 4176
rect 10418 4124 10430 4158
rect 10464 4124 10476 4158
rect 10418 4114 10476 4124
rect 10506 4086 10552 4286
rect 10802 4302 10866 4308
rect 10802 4250 10808 4302
rect 10860 4250 10866 4302
rect 10802 4244 10866 4250
rect 10696 4171 10972 4202
rect 10696 4137 10725 4171
rect 10759 4137 10817 4171
rect 10851 4137 10909 4171
rect 10943 4137 10972 4171
rect 10696 4134 10972 4137
rect 9864 4069 9928 4076
rect 9864 4036 9870 4069
rect 9922 4036 9928 4069
rect 10040 4069 10104 4076
rect 10040 4036 10046 4069
rect 9922 4017 10046 4036
rect 10098 4017 10104 4069
rect 9870 4008 10104 4017
rect 10224 4074 10326 4086
rect 10224 4040 10286 4074
rect 10320 4040 10326 4074
rect 10224 4002 10326 4040
rect 10376 4074 10422 4086
rect 10376 4040 10382 4074
rect 10416 4040 10422 4074
rect 10376 4020 10422 4040
rect 10472 4074 10552 4086
rect 10472 4040 10478 4074
rect 10512 4040 10552 4074
rect 10224 3970 10286 4002
rect 10020 3968 10286 3970
rect 10320 3968 10326 4002
rect 10020 3956 10326 3968
rect 10366 4014 10432 4020
rect 10366 3962 10374 4014
rect 10426 3962 10432 4014
rect 10366 3956 10432 3962
rect 10472 4002 10552 4040
rect 10472 3968 10478 4002
rect 10512 3968 10552 4002
rect 10668 4106 10972 4134
rect 10472 3956 10518 3968
rect 10020 3942 10274 3956
rect 9864 3936 9930 3942
rect 9864 3884 9872 3936
rect 9924 3884 9930 3936
rect 9864 3878 9930 3884
rect 9012 3669 9042 3672
rect 9094 3669 9636 3672
rect 9012 3635 9041 3669
rect 9094 3635 9133 3669
rect 9167 3635 9225 3669
rect 9259 3667 9636 3669
rect 9259 3635 9387 3667
rect 9012 3620 9042 3635
rect 9094 3633 9387 3635
rect 9421 3633 9479 3667
rect 9513 3633 9571 3667
rect 9605 3633 9636 3667
rect 9094 3620 9636 3633
rect 9012 3602 9636 3620
rect 9704 3678 9980 3692
rect 9704 3661 9896 3678
rect 9948 3661 9980 3678
rect 9704 3627 9733 3661
rect 9767 3627 9825 3661
rect 9859 3627 9896 3661
rect 9951 3627 9980 3661
rect 9704 3626 9896 3627
rect 9948 3626 9980 3627
rect 9704 3596 9980 3626
rect 10020 3592 10048 3942
rect 10320 3918 10384 3928
rect 10320 3884 10334 3918
rect 10368 3884 10640 3918
rect 10320 3866 10384 3884
rect 10236 3820 10308 3832
rect 10236 3768 10246 3820
rect 10298 3768 10308 3820
rect 10236 3756 10308 3768
rect 10606 3702 10640 3884
rect 10668 3802 10696 4106
rect 10668 3792 10736 3802
rect 10668 3758 10684 3792
rect 10718 3758 10736 3792
rect 10668 3744 10736 3758
rect 10080 3674 10640 3702
rect 10080 3671 10146 3674
rect 10080 3637 10096 3671
rect 10130 3637 10146 3671
rect 10080 3628 10146 3637
rect 10314 3619 10404 3640
rect 8512 3511 8752 3528
rect 8796 3584 8862 3590
rect 8796 3532 8804 3584
rect 8856 3532 8862 3584
rect 8796 3526 8810 3532
rect 8246 3471 8292 3504
rect 8246 3437 8252 3471
rect 8286 3437 8292 3471
rect 8512 3477 8524 3511
rect 8558 3500 8752 3511
rect 8804 3509 8810 3526
rect 8844 3526 8862 3532
rect 8892 3543 8938 3590
rect 10020 3564 10092 3592
rect 8844 3509 8850 3526
rect 8558 3477 8750 3500
rect 8512 3468 8750 3477
rect 8246 3390 8292 3437
rect 8460 3430 8526 3438
rect 8374 3426 8420 3430
rect 7490 3368 7562 3372
rect 6950 3343 7016 3356
rect 6950 3309 6966 3343
rect 7000 3309 7016 3343
rect 6950 3300 7016 3309
rect 7490 3316 7499 3368
rect 7551 3316 7562 3368
rect 7490 3304 7562 3316
rect 7686 3366 7760 3386
rect 8334 3383 8420 3426
rect 7686 3332 7698 3366
rect 7732 3332 7760 3366
rect 7686 3308 7760 3332
rect 7796 3372 7864 3378
rect 7796 3320 7803 3372
rect 7855 3366 7864 3372
rect 7855 3360 7948 3366
rect 7855 3326 7894 3360
rect 7928 3326 7948 3360
rect 7855 3320 7948 3326
rect 7796 3316 7948 3320
rect 8192 3343 8258 3354
rect 7796 3314 7864 3316
rect 8192 3309 8208 3343
rect 8242 3309 8258 3343
rect 8192 3296 8258 3309
rect 8334 3349 8380 3383
rect 8414 3349 8420 3383
rect 8460 3378 8466 3430
rect 8518 3378 8526 3430
rect 8460 3370 8476 3378
rect 8334 3311 8420 3349
rect 8334 3277 8380 3311
rect 8414 3277 8420 3311
rect 7272 3256 7330 3270
rect 7272 3236 7284 3256
rect 6802 3222 7284 3236
rect 7318 3222 7330 3256
rect 6802 3202 7330 3222
rect 8334 3230 8420 3277
rect 8470 3349 8476 3370
rect 8510 3370 8526 3378
rect 8566 3383 8662 3430
rect 8510 3349 8516 3370
rect 8470 3311 8516 3349
rect 8470 3277 8476 3311
rect 8510 3277 8516 3311
rect 8470 3230 8516 3277
rect 8566 3349 8572 3383
rect 8606 3349 8662 3383
rect 8566 3311 8662 3349
rect 8566 3277 8572 3311
rect 8606 3277 8662 3311
rect 8566 3230 8662 3277
rect 6694 2900 6740 2912
rect 6802 2872 6862 3202
rect 8334 3176 8384 3230
rect 6908 3152 6984 3158
rect 6908 3100 6916 3152
rect 6968 3100 6984 3152
rect 6908 3094 6984 3100
rect 7124 3125 7746 3156
rect 6542 2862 6862 2872
rect 6542 2828 6556 2862
rect 6590 2828 6862 2862
rect 6542 2810 6862 2828
rect 7124 3091 7153 3125
rect 7187 3091 7245 3125
rect 7279 3091 7337 3125
rect 7371 3123 7746 3125
rect 7371 3091 7499 3123
rect 7124 3089 7499 3091
rect 7533 3089 7591 3123
rect 7625 3089 7683 3123
rect 7717 3089 7746 3123
rect 7124 3058 7746 3089
rect 7816 3130 8092 3148
rect 7816 3117 7939 3130
rect 7991 3117 8092 3130
rect 8168 3126 8226 3134
rect 7816 3083 7845 3117
rect 7879 3083 7937 3117
rect 7991 3083 8029 3117
rect 8063 3083 8092 3117
rect 7816 3078 7939 3083
rect 7991 3078 8092 3083
rect 7124 2782 7222 3058
rect 7816 3052 8092 3078
rect 8160 3120 8234 3126
rect 8160 3068 8171 3120
rect 8223 3068 8234 3120
rect 8314 3110 8384 3176
rect 8416 3183 8474 3198
rect 8416 3149 8428 3183
rect 8462 3149 8474 3183
rect 8416 3132 8474 3149
rect 8160 3062 8234 3068
rect 8168 3056 8226 3062
rect 7884 2782 7968 3052
rect 8334 3030 8384 3110
rect 8528 3102 8586 3120
rect 8528 3068 8540 3102
rect 8574 3068 8586 3102
rect 8528 3058 8586 3068
rect 8616 3030 8662 3230
rect 8334 3018 8436 3030
rect 8334 2984 8396 3018
rect 8430 2984 8436 3018
rect 8334 2946 8436 2984
rect 8486 3018 8532 3030
rect 8486 2984 8492 3018
rect 8526 2984 8532 3018
rect 8486 2964 8532 2984
rect 8582 3018 8662 3030
rect 8582 2984 8588 3018
rect 8622 2984 8662 3018
rect 8334 2912 8396 2946
rect 8430 2912 8436 2946
rect 8334 2900 8436 2912
rect 8476 2958 8542 2964
rect 8476 2906 8484 2958
rect 8536 2906 8542 2958
rect 8476 2900 8542 2906
rect 8582 2946 8662 2984
rect 8582 2912 8588 2946
rect 8622 2912 8662 2946
rect 8690 3236 8750 3468
rect 8804 3471 8850 3509
rect 8804 3437 8810 3471
rect 8844 3437 8850 3471
rect 8804 3390 8850 3437
rect 8892 3509 8898 3543
rect 8932 3509 8938 3543
rect 8892 3471 8938 3509
rect 8892 3437 8898 3471
rect 8932 3437 8938 3471
rect 8892 3390 8938 3437
rect 10046 3543 10092 3564
rect 10046 3509 10052 3543
rect 10086 3509 10092 3543
rect 10046 3471 10092 3509
rect 10046 3437 10052 3471
rect 10086 3437 10092 3471
rect 10046 3390 10092 3437
rect 10134 3570 10180 3590
rect 10314 3585 10343 3619
rect 10377 3585 10404 3619
rect 10134 3564 10202 3570
rect 10314 3564 10404 3585
rect 10134 3543 10142 3564
rect 10134 3509 10140 3543
rect 10194 3512 10202 3564
rect 10174 3509 10202 3512
rect 10134 3504 10202 3509
rect 10400 3528 10458 3530
rect 10606 3528 10640 3674
rect 10726 3671 10792 3682
rect 10726 3637 10742 3671
rect 10776 3637 10792 3671
rect 10726 3626 10792 3637
rect 10900 3672 11524 3704
rect 11606 3692 11684 4650
rect 12198 4641 12227 4650
rect 12261 4650 14115 4675
rect 12261 4641 12288 4650
rect 12198 4620 12288 4641
rect 12284 4584 12342 4586
rect 12284 4567 12346 4584
rect 12284 4533 12296 4567
rect 12330 4533 12346 4567
rect 12284 4524 12346 4533
rect 11784 4486 12150 4490
rect 12232 4486 12298 4494
rect 11784 4458 12192 4486
rect 11784 4420 11812 4458
rect 12106 4439 12192 4458
rect 11784 4412 11850 4420
rect 11784 4378 11799 4412
rect 11833 4378 11850 4412
rect 11784 4366 11850 4378
rect 11956 4416 12024 4422
rect 11956 4364 11966 4416
rect 12018 4364 12024 4416
rect 11956 4358 12024 4364
rect 12106 4405 12152 4439
rect 12186 4405 12192 4439
rect 12232 4434 12238 4486
rect 12290 4434 12298 4486
rect 12232 4426 12248 4434
rect 12106 4367 12192 4405
rect 12106 4333 12152 4367
rect 12186 4333 12192 4367
rect 11866 4304 11934 4310
rect 11866 4252 11874 4304
rect 11926 4252 11934 4304
rect 11866 4242 11934 4252
rect 12106 4286 12192 4333
rect 12242 4405 12248 4426
rect 12282 4426 12298 4434
rect 12338 4454 12666 4486
rect 12338 4439 12434 4454
rect 12282 4405 12288 4426
rect 12242 4367 12288 4405
rect 12242 4333 12248 4367
rect 12282 4333 12288 4367
rect 12242 4286 12288 4333
rect 12338 4405 12344 4439
rect 12378 4405 12434 4439
rect 12638 4418 12666 4454
rect 12338 4367 12434 4405
rect 12338 4333 12344 4367
rect 12378 4333 12434 4367
rect 12596 4410 12666 4418
rect 12596 4376 12611 4410
rect 12645 4376 12666 4410
rect 12596 4358 12666 4376
rect 12772 4418 12836 4424
rect 12772 4366 12778 4418
rect 12830 4366 12836 4418
rect 12772 4360 12836 4366
rect 12338 4286 12434 4333
rect 11764 4171 12040 4202
rect 11764 4137 11793 4171
rect 11827 4137 11885 4171
rect 11919 4137 11977 4171
rect 12011 4137 12040 4171
rect 11764 4106 12040 4137
rect 12106 4086 12156 4286
rect 12188 4239 12246 4254
rect 12188 4205 12200 4239
rect 12234 4205 12246 4239
rect 12188 4188 12246 4205
rect 12300 4158 12358 4176
rect 12300 4124 12312 4158
rect 12346 4124 12358 4158
rect 12300 4114 12358 4124
rect 12388 4086 12434 4286
rect 12684 4302 12748 4308
rect 12684 4250 12690 4302
rect 12742 4250 12748 4302
rect 12684 4244 12748 4250
rect 12578 4171 12854 4202
rect 12578 4137 12607 4171
rect 12641 4137 12699 4171
rect 12733 4137 12791 4171
rect 12825 4137 12854 4171
rect 12578 4134 12854 4137
rect 11746 4069 11810 4076
rect 11746 4036 11752 4069
rect 11804 4036 11810 4069
rect 11922 4069 11986 4076
rect 11922 4036 11928 4069
rect 11804 4017 11928 4036
rect 11980 4017 11986 4069
rect 11752 4008 11986 4017
rect 12106 4074 12208 4086
rect 12106 4040 12168 4074
rect 12202 4040 12208 4074
rect 12106 4002 12208 4040
rect 12258 4074 12304 4086
rect 12258 4040 12264 4074
rect 12298 4040 12304 4074
rect 12258 4020 12304 4040
rect 12354 4074 12434 4086
rect 12354 4040 12360 4074
rect 12394 4040 12434 4074
rect 12106 3970 12168 4002
rect 11902 3968 12168 3970
rect 12202 3968 12208 4002
rect 11902 3956 12208 3968
rect 12248 4014 12314 4020
rect 12248 3962 12256 4014
rect 12308 3962 12314 4014
rect 12248 3956 12314 3962
rect 12354 4002 12434 4040
rect 12354 3968 12360 4002
rect 12394 3968 12434 4002
rect 12550 4106 12854 4134
rect 12354 3956 12400 3968
rect 11902 3942 12156 3956
rect 11746 3936 11812 3942
rect 11746 3884 11754 3936
rect 11806 3884 11812 3936
rect 11746 3878 11812 3884
rect 10900 3669 10930 3672
rect 10982 3669 11524 3672
rect 10900 3635 10929 3669
rect 10982 3635 11021 3669
rect 11055 3635 11113 3669
rect 11147 3667 11524 3669
rect 11147 3635 11275 3667
rect 10900 3620 10930 3635
rect 10982 3633 11275 3635
rect 11309 3633 11367 3667
rect 11401 3633 11459 3667
rect 11493 3633 11524 3667
rect 10982 3620 11524 3633
rect 10900 3602 11524 3620
rect 11586 3678 11862 3692
rect 11586 3661 11778 3678
rect 11830 3661 11862 3678
rect 11586 3627 11615 3661
rect 11649 3627 11707 3661
rect 11741 3627 11778 3661
rect 11833 3627 11862 3661
rect 11586 3626 11778 3627
rect 11830 3626 11862 3627
rect 11586 3596 11862 3626
rect 11902 3592 11930 3942
rect 12202 3918 12266 3928
rect 12202 3884 12216 3918
rect 12250 3884 12522 3918
rect 12202 3866 12266 3884
rect 12118 3820 12190 3832
rect 12118 3768 12128 3820
rect 12180 3768 12190 3820
rect 12118 3756 12190 3768
rect 12488 3702 12522 3884
rect 12550 3802 12578 4106
rect 12550 3792 12618 3802
rect 12550 3758 12566 3792
rect 12600 3758 12618 3792
rect 12550 3744 12618 3758
rect 11962 3674 12522 3702
rect 11962 3671 12028 3674
rect 11962 3637 11978 3671
rect 12012 3637 12028 3671
rect 11962 3628 12028 3637
rect 12196 3619 12286 3640
rect 10400 3511 10640 3528
rect 10684 3584 10750 3590
rect 10684 3532 10692 3584
rect 10744 3532 10750 3584
rect 10684 3526 10698 3532
rect 10134 3471 10180 3504
rect 10134 3437 10140 3471
rect 10174 3437 10180 3471
rect 10400 3477 10412 3511
rect 10446 3500 10640 3511
rect 10692 3509 10698 3526
rect 10732 3526 10750 3532
rect 10780 3543 10826 3590
rect 11902 3564 11974 3592
rect 10732 3509 10738 3526
rect 10446 3477 10638 3500
rect 10400 3468 10638 3477
rect 10134 3390 10180 3437
rect 10348 3430 10414 3438
rect 10262 3426 10308 3430
rect 9378 3368 9450 3372
rect 8838 3343 8904 3356
rect 8838 3309 8854 3343
rect 8888 3309 8904 3343
rect 8838 3300 8904 3309
rect 9378 3316 9387 3368
rect 9439 3316 9450 3368
rect 9378 3304 9450 3316
rect 9574 3366 9648 3386
rect 10222 3383 10308 3426
rect 9574 3332 9586 3366
rect 9620 3332 9648 3366
rect 9574 3308 9648 3332
rect 9684 3372 9752 3378
rect 9684 3320 9691 3372
rect 9743 3366 9752 3372
rect 9743 3360 9836 3366
rect 9743 3326 9782 3360
rect 9816 3326 9836 3360
rect 9743 3320 9836 3326
rect 9684 3316 9836 3320
rect 10080 3343 10146 3354
rect 9684 3314 9752 3316
rect 10080 3309 10096 3343
rect 10130 3309 10146 3343
rect 10080 3296 10146 3309
rect 10222 3349 10268 3383
rect 10302 3349 10308 3383
rect 10348 3378 10354 3430
rect 10406 3378 10414 3430
rect 10348 3370 10364 3378
rect 10222 3311 10308 3349
rect 10222 3277 10268 3311
rect 10302 3277 10308 3311
rect 9160 3256 9218 3270
rect 9160 3236 9172 3256
rect 8690 3222 9172 3236
rect 9206 3222 9218 3256
rect 8690 3202 9218 3222
rect 10222 3230 10308 3277
rect 10358 3349 10364 3370
rect 10398 3370 10414 3378
rect 10454 3383 10550 3430
rect 10398 3349 10404 3370
rect 10358 3311 10404 3349
rect 10358 3277 10364 3311
rect 10398 3277 10404 3311
rect 10358 3230 10404 3277
rect 10454 3349 10460 3383
rect 10494 3349 10550 3383
rect 10454 3311 10550 3349
rect 10454 3277 10460 3311
rect 10494 3277 10550 3311
rect 10454 3230 10550 3277
rect 8582 2900 8628 2912
rect 8690 2872 8750 3202
rect 10222 3176 10272 3230
rect 8796 3152 8872 3158
rect 8796 3100 8804 3152
rect 8856 3100 8872 3152
rect 8796 3094 8872 3100
rect 9012 3125 9634 3156
rect 8430 2862 8750 2872
rect 8430 2828 8444 2862
rect 8478 2828 8750 2862
rect 8430 2810 8750 2828
rect 9012 3091 9041 3125
rect 9075 3091 9133 3125
rect 9167 3091 9225 3125
rect 9259 3123 9634 3125
rect 9259 3091 9387 3123
rect 9012 3089 9387 3091
rect 9421 3089 9479 3123
rect 9513 3089 9571 3123
rect 9605 3089 9634 3123
rect 9012 3058 9634 3089
rect 9704 3130 9980 3148
rect 9704 3117 9827 3130
rect 9879 3117 9980 3130
rect 10056 3126 10114 3134
rect 9704 3083 9733 3117
rect 9767 3083 9825 3117
rect 9879 3083 9917 3117
rect 9951 3083 9980 3117
rect 9704 3078 9827 3083
rect 9879 3078 9980 3083
rect 9012 2782 9110 3058
rect 9704 3052 9980 3078
rect 10048 3120 10122 3126
rect 10048 3068 10059 3120
rect 10111 3068 10122 3120
rect 10202 3110 10272 3176
rect 10304 3183 10362 3198
rect 10304 3149 10316 3183
rect 10350 3149 10362 3183
rect 10304 3132 10362 3149
rect 10048 3062 10122 3068
rect 10056 3056 10114 3062
rect 9772 2782 9856 3052
rect 10222 3030 10272 3110
rect 10416 3102 10474 3120
rect 10416 3068 10428 3102
rect 10462 3068 10474 3102
rect 10416 3058 10474 3068
rect 10504 3030 10550 3230
rect 10222 3018 10324 3030
rect 10222 2984 10284 3018
rect 10318 2984 10324 3018
rect 10222 2946 10324 2984
rect 10374 3018 10420 3030
rect 10374 2984 10380 3018
rect 10414 2984 10420 3018
rect 10374 2964 10420 2984
rect 10470 3018 10550 3030
rect 10470 2984 10476 3018
rect 10510 2984 10550 3018
rect 10222 2912 10284 2946
rect 10318 2912 10324 2946
rect 10222 2900 10324 2912
rect 10364 2958 10430 2964
rect 10364 2906 10372 2958
rect 10424 2906 10430 2958
rect 10364 2900 10430 2906
rect 10470 2946 10550 2984
rect 10470 2912 10476 2946
rect 10510 2912 10550 2946
rect 10578 3236 10638 3468
rect 10692 3471 10738 3509
rect 10692 3437 10698 3471
rect 10732 3437 10738 3471
rect 10692 3390 10738 3437
rect 10780 3509 10786 3543
rect 10820 3509 10826 3543
rect 10780 3471 10826 3509
rect 10780 3437 10786 3471
rect 10820 3437 10826 3471
rect 10780 3390 10826 3437
rect 11928 3543 11974 3564
rect 11928 3509 11934 3543
rect 11968 3509 11974 3543
rect 11928 3471 11974 3509
rect 11928 3437 11934 3471
rect 11968 3437 11974 3471
rect 11928 3390 11974 3437
rect 12016 3570 12062 3590
rect 12196 3585 12225 3619
rect 12259 3585 12286 3619
rect 12016 3564 12084 3570
rect 12196 3564 12286 3585
rect 12016 3543 12024 3564
rect 12016 3509 12022 3543
rect 12076 3512 12084 3564
rect 12056 3509 12084 3512
rect 12016 3504 12084 3509
rect 12282 3528 12340 3530
rect 12488 3528 12522 3674
rect 12608 3671 12674 3682
rect 12608 3637 12624 3671
rect 12658 3637 12674 3671
rect 12608 3626 12674 3637
rect 12782 3672 13406 3704
rect 13494 3692 13572 4650
rect 14086 4641 14115 4650
rect 14149 4650 16003 4675
rect 14149 4641 14176 4650
rect 14086 4620 14176 4641
rect 14172 4584 14230 4586
rect 14172 4567 14234 4584
rect 14172 4533 14184 4567
rect 14218 4533 14234 4567
rect 14172 4524 14234 4533
rect 13672 4486 14038 4490
rect 14120 4486 14186 4494
rect 13672 4458 14080 4486
rect 13672 4420 13700 4458
rect 13994 4439 14080 4458
rect 13672 4412 13738 4420
rect 13672 4378 13687 4412
rect 13721 4378 13738 4412
rect 13672 4366 13738 4378
rect 13844 4416 13912 4422
rect 13844 4364 13854 4416
rect 13906 4364 13912 4416
rect 13844 4358 13912 4364
rect 13994 4405 14040 4439
rect 14074 4405 14080 4439
rect 14120 4434 14126 4486
rect 14178 4434 14186 4486
rect 14120 4426 14136 4434
rect 13994 4367 14080 4405
rect 13994 4333 14040 4367
rect 14074 4333 14080 4367
rect 13754 4304 13822 4310
rect 13754 4252 13762 4304
rect 13814 4252 13822 4304
rect 13754 4242 13822 4252
rect 13994 4286 14080 4333
rect 14130 4405 14136 4426
rect 14170 4426 14186 4434
rect 14226 4454 14554 4486
rect 14226 4439 14322 4454
rect 14170 4405 14176 4426
rect 14130 4367 14176 4405
rect 14130 4333 14136 4367
rect 14170 4333 14176 4367
rect 14130 4286 14176 4333
rect 14226 4405 14232 4439
rect 14266 4405 14322 4439
rect 14526 4418 14554 4454
rect 14226 4367 14322 4405
rect 14226 4333 14232 4367
rect 14266 4333 14322 4367
rect 14484 4410 14554 4418
rect 14484 4376 14499 4410
rect 14533 4376 14554 4410
rect 14484 4358 14554 4376
rect 14660 4418 14724 4424
rect 14660 4366 14666 4418
rect 14718 4366 14724 4418
rect 14660 4360 14724 4366
rect 14226 4286 14322 4333
rect 13652 4171 13928 4202
rect 13652 4137 13681 4171
rect 13715 4137 13773 4171
rect 13807 4137 13865 4171
rect 13899 4137 13928 4171
rect 13652 4106 13928 4137
rect 13994 4086 14044 4286
rect 14076 4239 14134 4254
rect 14076 4205 14088 4239
rect 14122 4205 14134 4239
rect 14076 4188 14134 4205
rect 14188 4158 14246 4176
rect 14188 4124 14200 4158
rect 14234 4124 14246 4158
rect 14188 4114 14246 4124
rect 14276 4086 14322 4286
rect 14572 4302 14636 4308
rect 14572 4250 14578 4302
rect 14630 4250 14636 4302
rect 14572 4244 14636 4250
rect 14466 4171 14742 4202
rect 14466 4137 14495 4171
rect 14529 4137 14587 4171
rect 14621 4137 14679 4171
rect 14713 4137 14742 4171
rect 14466 4134 14742 4137
rect 13634 4069 13698 4076
rect 13634 4036 13640 4069
rect 13692 4036 13698 4069
rect 13810 4069 13874 4076
rect 13810 4036 13816 4069
rect 13692 4017 13816 4036
rect 13868 4017 13874 4069
rect 13640 4008 13874 4017
rect 13994 4074 14096 4086
rect 13994 4040 14056 4074
rect 14090 4040 14096 4074
rect 13994 4002 14096 4040
rect 14146 4074 14192 4086
rect 14146 4040 14152 4074
rect 14186 4040 14192 4074
rect 14146 4020 14192 4040
rect 14242 4074 14322 4086
rect 14242 4040 14248 4074
rect 14282 4040 14322 4074
rect 13994 3970 14056 4002
rect 13790 3968 14056 3970
rect 14090 3968 14096 4002
rect 13790 3956 14096 3968
rect 14136 4014 14202 4020
rect 14136 3962 14144 4014
rect 14196 3962 14202 4014
rect 14136 3956 14202 3962
rect 14242 4002 14322 4040
rect 14242 3968 14248 4002
rect 14282 3968 14322 4002
rect 14438 4106 14742 4134
rect 14242 3956 14288 3968
rect 13790 3942 14044 3956
rect 13634 3936 13700 3942
rect 13634 3884 13642 3936
rect 13694 3884 13700 3936
rect 13634 3878 13700 3884
rect 12782 3669 12812 3672
rect 12864 3669 13406 3672
rect 12782 3635 12811 3669
rect 12864 3635 12903 3669
rect 12937 3635 12995 3669
rect 13029 3667 13406 3669
rect 13029 3635 13157 3667
rect 12782 3620 12812 3635
rect 12864 3633 13157 3635
rect 13191 3633 13249 3667
rect 13283 3633 13341 3667
rect 13375 3633 13406 3667
rect 12864 3620 13406 3633
rect 12782 3602 13406 3620
rect 13474 3678 13750 3692
rect 13474 3661 13666 3678
rect 13718 3661 13750 3678
rect 13474 3627 13503 3661
rect 13537 3627 13595 3661
rect 13629 3627 13666 3661
rect 13721 3627 13750 3661
rect 13474 3626 13666 3627
rect 13718 3626 13750 3627
rect 13474 3596 13750 3626
rect 13790 3592 13818 3942
rect 14090 3918 14154 3928
rect 14090 3884 14104 3918
rect 14138 3884 14410 3918
rect 14090 3866 14154 3884
rect 14006 3820 14078 3832
rect 14006 3768 14016 3820
rect 14068 3768 14078 3820
rect 14006 3756 14078 3768
rect 14376 3702 14410 3884
rect 14438 3802 14466 4106
rect 14438 3792 14506 3802
rect 14438 3758 14454 3792
rect 14488 3758 14506 3792
rect 14438 3744 14506 3758
rect 13850 3674 14410 3702
rect 13850 3671 13916 3674
rect 13850 3637 13866 3671
rect 13900 3637 13916 3671
rect 13850 3628 13916 3637
rect 14084 3619 14174 3640
rect 12282 3511 12522 3528
rect 12566 3584 12632 3590
rect 12566 3532 12574 3584
rect 12626 3532 12632 3584
rect 12566 3526 12580 3532
rect 12016 3471 12062 3504
rect 12016 3437 12022 3471
rect 12056 3437 12062 3471
rect 12282 3477 12294 3511
rect 12328 3500 12522 3511
rect 12574 3509 12580 3526
rect 12614 3526 12632 3532
rect 12662 3543 12708 3590
rect 13790 3564 13862 3592
rect 12614 3509 12620 3526
rect 12328 3477 12520 3500
rect 12282 3468 12520 3477
rect 12016 3390 12062 3437
rect 12230 3430 12296 3438
rect 12144 3426 12190 3430
rect 11266 3368 11338 3372
rect 10726 3343 10792 3356
rect 10726 3309 10742 3343
rect 10776 3309 10792 3343
rect 10726 3300 10792 3309
rect 11266 3316 11275 3368
rect 11327 3316 11338 3368
rect 11266 3304 11338 3316
rect 11462 3366 11536 3386
rect 12104 3383 12190 3426
rect 11462 3332 11474 3366
rect 11508 3332 11536 3366
rect 11462 3308 11536 3332
rect 11566 3372 11634 3378
rect 11566 3320 11573 3372
rect 11625 3366 11634 3372
rect 11625 3360 11718 3366
rect 11625 3326 11664 3360
rect 11698 3326 11718 3360
rect 11625 3320 11718 3326
rect 11566 3316 11718 3320
rect 11962 3343 12028 3354
rect 11566 3314 11634 3316
rect 11962 3309 11978 3343
rect 12012 3309 12028 3343
rect 11962 3296 12028 3309
rect 12104 3349 12150 3383
rect 12184 3349 12190 3383
rect 12230 3378 12236 3430
rect 12288 3378 12296 3430
rect 12230 3370 12246 3378
rect 12104 3311 12190 3349
rect 12104 3277 12150 3311
rect 12184 3277 12190 3311
rect 11048 3256 11106 3270
rect 11048 3236 11060 3256
rect 10578 3222 11060 3236
rect 11094 3222 11106 3256
rect 10578 3202 11106 3222
rect 12104 3230 12190 3277
rect 12240 3349 12246 3370
rect 12280 3370 12296 3378
rect 12336 3383 12432 3430
rect 12280 3349 12286 3370
rect 12240 3311 12286 3349
rect 12240 3277 12246 3311
rect 12280 3277 12286 3311
rect 12240 3230 12286 3277
rect 12336 3349 12342 3383
rect 12376 3349 12432 3383
rect 12336 3311 12432 3349
rect 12336 3277 12342 3311
rect 12376 3277 12432 3311
rect 12336 3230 12432 3277
rect 10470 2900 10516 2912
rect 10578 2872 10638 3202
rect 12104 3176 12154 3230
rect 10684 3152 10760 3158
rect 10684 3100 10692 3152
rect 10744 3100 10760 3152
rect 10684 3094 10760 3100
rect 10900 3125 11522 3156
rect 10318 2862 10638 2872
rect 10318 2828 10332 2862
rect 10366 2828 10638 2862
rect 10318 2810 10638 2828
rect 10900 3091 10929 3125
rect 10963 3091 11021 3125
rect 11055 3091 11113 3125
rect 11147 3123 11522 3125
rect 11147 3091 11275 3123
rect 10900 3089 11275 3091
rect 11309 3089 11367 3123
rect 11401 3089 11459 3123
rect 11493 3089 11522 3123
rect 10900 3058 11522 3089
rect 11586 3130 11862 3148
rect 11586 3117 11709 3130
rect 11761 3117 11862 3130
rect 11938 3126 11996 3134
rect 11586 3083 11615 3117
rect 11649 3083 11707 3117
rect 11761 3083 11799 3117
rect 11833 3083 11862 3117
rect 11586 3078 11709 3083
rect 11761 3078 11862 3083
rect 10900 2782 10998 3058
rect 11586 3052 11862 3078
rect 11930 3120 12004 3126
rect 11930 3068 11941 3120
rect 11993 3068 12004 3120
rect 12084 3110 12154 3176
rect 12186 3183 12244 3198
rect 12186 3149 12198 3183
rect 12232 3149 12244 3183
rect 12186 3132 12244 3149
rect 11930 3062 12004 3068
rect 11938 3056 11996 3062
rect 11654 2782 11738 3052
rect 12104 3030 12154 3110
rect 12298 3102 12356 3120
rect 12298 3068 12310 3102
rect 12344 3068 12356 3102
rect 12298 3058 12356 3068
rect 12386 3030 12432 3230
rect 12104 3018 12206 3030
rect 12104 2984 12166 3018
rect 12200 2984 12206 3018
rect 12104 2946 12206 2984
rect 12256 3018 12302 3030
rect 12256 2984 12262 3018
rect 12296 2984 12302 3018
rect 12256 2964 12302 2984
rect 12352 3018 12432 3030
rect 12352 2984 12358 3018
rect 12392 2984 12432 3018
rect 12104 2912 12166 2946
rect 12200 2912 12206 2946
rect 12104 2900 12206 2912
rect 12246 2958 12312 2964
rect 12246 2906 12254 2958
rect 12306 2906 12312 2958
rect 12246 2900 12312 2906
rect 12352 2946 12432 2984
rect 12352 2912 12358 2946
rect 12392 2912 12432 2946
rect 12460 3236 12520 3468
rect 12574 3471 12620 3509
rect 12574 3437 12580 3471
rect 12614 3437 12620 3471
rect 12574 3390 12620 3437
rect 12662 3509 12668 3543
rect 12702 3509 12708 3543
rect 12662 3471 12708 3509
rect 12662 3437 12668 3471
rect 12702 3437 12708 3471
rect 12662 3390 12708 3437
rect 13816 3543 13862 3564
rect 13816 3509 13822 3543
rect 13856 3509 13862 3543
rect 13816 3471 13862 3509
rect 13816 3437 13822 3471
rect 13856 3437 13862 3471
rect 13816 3390 13862 3437
rect 13904 3570 13950 3590
rect 14084 3585 14113 3619
rect 14147 3585 14174 3619
rect 13904 3564 13972 3570
rect 14084 3564 14174 3585
rect 13904 3543 13912 3564
rect 13904 3509 13910 3543
rect 13964 3512 13972 3564
rect 13944 3509 13972 3512
rect 13904 3504 13972 3509
rect 14170 3528 14228 3530
rect 14376 3528 14410 3674
rect 14496 3671 14562 3682
rect 14496 3637 14512 3671
rect 14546 3637 14562 3671
rect 14496 3626 14562 3637
rect 14670 3672 15294 3704
rect 15382 3692 15460 4650
rect 15974 4641 16003 4650
rect 16037 4650 17891 4675
rect 16037 4641 16064 4650
rect 15974 4620 16064 4641
rect 16060 4584 16118 4586
rect 16060 4567 16122 4584
rect 16060 4533 16072 4567
rect 16106 4533 16122 4567
rect 16060 4524 16122 4533
rect 15560 4486 15926 4490
rect 16008 4486 16074 4494
rect 15560 4458 15968 4486
rect 15560 4420 15588 4458
rect 15882 4439 15968 4458
rect 15560 4412 15626 4420
rect 15560 4378 15575 4412
rect 15609 4378 15626 4412
rect 15560 4366 15626 4378
rect 15732 4416 15800 4422
rect 15732 4364 15742 4416
rect 15794 4364 15800 4416
rect 15732 4358 15800 4364
rect 15882 4405 15928 4439
rect 15962 4405 15968 4439
rect 16008 4434 16014 4486
rect 16066 4434 16074 4486
rect 16008 4426 16024 4434
rect 15882 4367 15968 4405
rect 15882 4333 15928 4367
rect 15962 4333 15968 4367
rect 15642 4304 15710 4310
rect 15642 4252 15650 4304
rect 15702 4252 15710 4304
rect 15642 4242 15710 4252
rect 15882 4286 15968 4333
rect 16018 4405 16024 4426
rect 16058 4426 16074 4434
rect 16114 4454 16442 4486
rect 16114 4439 16210 4454
rect 16058 4405 16064 4426
rect 16018 4367 16064 4405
rect 16018 4333 16024 4367
rect 16058 4333 16064 4367
rect 16018 4286 16064 4333
rect 16114 4405 16120 4439
rect 16154 4405 16210 4439
rect 16414 4418 16442 4454
rect 16114 4367 16210 4405
rect 16114 4333 16120 4367
rect 16154 4333 16210 4367
rect 16372 4410 16442 4418
rect 16372 4376 16387 4410
rect 16421 4376 16442 4410
rect 16372 4358 16442 4376
rect 16548 4418 16612 4424
rect 16548 4366 16554 4418
rect 16606 4366 16612 4418
rect 16548 4360 16612 4366
rect 16114 4286 16210 4333
rect 15540 4171 15816 4202
rect 15540 4137 15569 4171
rect 15603 4137 15661 4171
rect 15695 4137 15753 4171
rect 15787 4137 15816 4171
rect 15540 4106 15816 4137
rect 15882 4086 15932 4286
rect 15964 4239 16022 4254
rect 15964 4205 15976 4239
rect 16010 4205 16022 4239
rect 15964 4188 16022 4205
rect 16076 4158 16134 4176
rect 16076 4124 16088 4158
rect 16122 4124 16134 4158
rect 16076 4114 16134 4124
rect 16164 4086 16210 4286
rect 16460 4302 16524 4308
rect 16460 4250 16466 4302
rect 16518 4250 16524 4302
rect 16460 4244 16524 4250
rect 16354 4171 16630 4202
rect 16354 4137 16383 4171
rect 16417 4137 16475 4171
rect 16509 4137 16567 4171
rect 16601 4137 16630 4171
rect 16354 4134 16630 4137
rect 15522 4069 15586 4076
rect 15522 4036 15528 4069
rect 15580 4036 15586 4069
rect 15698 4069 15762 4076
rect 15698 4036 15704 4069
rect 15580 4017 15704 4036
rect 15756 4017 15762 4069
rect 15528 4008 15762 4017
rect 15882 4074 15984 4086
rect 15882 4040 15944 4074
rect 15978 4040 15984 4074
rect 15882 4002 15984 4040
rect 16034 4074 16080 4086
rect 16034 4040 16040 4074
rect 16074 4040 16080 4074
rect 16034 4020 16080 4040
rect 16130 4074 16210 4086
rect 16130 4040 16136 4074
rect 16170 4040 16210 4074
rect 15882 3970 15944 4002
rect 15678 3968 15944 3970
rect 15978 3968 15984 4002
rect 15678 3956 15984 3968
rect 16024 4014 16090 4020
rect 16024 3962 16032 4014
rect 16084 3962 16090 4014
rect 16024 3956 16090 3962
rect 16130 4002 16210 4040
rect 16130 3968 16136 4002
rect 16170 3968 16210 4002
rect 16326 4106 16630 4134
rect 16130 3956 16176 3968
rect 15678 3942 15932 3956
rect 15522 3936 15588 3942
rect 15522 3884 15530 3936
rect 15582 3884 15588 3936
rect 15522 3878 15588 3884
rect 14670 3669 14700 3672
rect 14752 3669 15294 3672
rect 14670 3635 14699 3669
rect 14752 3635 14791 3669
rect 14825 3635 14883 3669
rect 14917 3667 15294 3669
rect 14917 3635 15045 3667
rect 14670 3620 14700 3635
rect 14752 3633 15045 3635
rect 15079 3633 15137 3667
rect 15171 3633 15229 3667
rect 15263 3633 15294 3667
rect 14752 3620 15294 3633
rect 14670 3602 15294 3620
rect 15362 3678 15638 3692
rect 15362 3661 15554 3678
rect 15606 3661 15638 3678
rect 15362 3627 15391 3661
rect 15425 3627 15483 3661
rect 15517 3627 15554 3661
rect 15609 3627 15638 3661
rect 15362 3626 15554 3627
rect 15606 3626 15638 3627
rect 15362 3596 15638 3626
rect 15678 3592 15706 3942
rect 15978 3918 16042 3928
rect 15978 3884 15992 3918
rect 16026 3884 16298 3918
rect 15978 3866 16042 3884
rect 15894 3820 15966 3832
rect 15894 3768 15904 3820
rect 15956 3768 15966 3820
rect 15894 3756 15966 3768
rect 16264 3702 16298 3884
rect 16326 3802 16354 4106
rect 16326 3792 16394 3802
rect 16326 3758 16342 3792
rect 16376 3758 16394 3792
rect 16326 3744 16394 3758
rect 15738 3674 16298 3702
rect 15738 3671 15804 3674
rect 15738 3637 15754 3671
rect 15788 3637 15804 3671
rect 15738 3628 15804 3637
rect 15972 3619 16062 3640
rect 14170 3511 14410 3528
rect 14454 3584 14520 3590
rect 14454 3532 14462 3584
rect 14514 3532 14520 3584
rect 14454 3526 14468 3532
rect 13904 3471 13950 3504
rect 13904 3437 13910 3471
rect 13944 3437 13950 3471
rect 14170 3477 14182 3511
rect 14216 3500 14410 3511
rect 14462 3509 14468 3526
rect 14502 3526 14520 3532
rect 14550 3543 14596 3590
rect 15678 3564 15750 3592
rect 14502 3509 14508 3526
rect 14216 3477 14408 3500
rect 14170 3468 14408 3477
rect 13904 3390 13950 3437
rect 14118 3430 14184 3438
rect 14032 3426 14078 3430
rect 13148 3368 13220 3372
rect 12608 3343 12674 3356
rect 12608 3309 12624 3343
rect 12658 3309 12674 3343
rect 12608 3300 12674 3309
rect 13148 3316 13157 3368
rect 13209 3316 13220 3368
rect 13148 3304 13220 3316
rect 13344 3366 13418 3386
rect 13992 3383 14078 3426
rect 13344 3332 13356 3366
rect 13390 3332 13418 3366
rect 13344 3308 13418 3332
rect 13454 3372 13522 3378
rect 13454 3320 13461 3372
rect 13513 3366 13522 3372
rect 13513 3360 13606 3366
rect 13513 3326 13552 3360
rect 13586 3326 13606 3360
rect 13513 3320 13606 3326
rect 13454 3316 13606 3320
rect 13850 3343 13916 3354
rect 13454 3314 13522 3316
rect 13850 3309 13866 3343
rect 13900 3309 13916 3343
rect 13850 3296 13916 3309
rect 13992 3349 14038 3383
rect 14072 3349 14078 3383
rect 14118 3378 14124 3430
rect 14176 3378 14184 3430
rect 14118 3370 14134 3378
rect 13992 3311 14078 3349
rect 13992 3277 14038 3311
rect 14072 3277 14078 3311
rect 12930 3256 12988 3270
rect 12930 3236 12942 3256
rect 12460 3222 12942 3236
rect 12976 3222 12988 3256
rect 12460 3202 12988 3222
rect 13992 3230 14078 3277
rect 14128 3349 14134 3370
rect 14168 3370 14184 3378
rect 14224 3383 14320 3430
rect 14168 3349 14174 3370
rect 14128 3311 14174 3349
rect 14128 3277 14134 3311
rect 14168 3277 14174 3311
rect 14128 3230 14174 3277
rect 14224 3349 14230 3383
rect 14264 3349 14320 3383
rect 14224 3311 14320 3349
rect 14224 3277 14230 3311
rect 14264 3277 14320 3311
rect 14224 3230 14320 3277
rect 12352 2900 12398 2912
rect 12460 2872 12520 3202
rect 13992 3176 14042 3230
rect 12566 3152 12642 3158
rect 12566 3100 12574 3152
rect 12626 3100 12642 3152
rect 12566 3094 12642 3100
rect 12782 3125 13404 3156
rect 12200 2862 12520 2872
rect 12200 2828 12214 2862
rect 12248 2828 12520 2862
rect 12200 2810 12520 2828
rect 12782 3091 12811 3125
rect 12845 3091 12903 3125
rect 12937 3091 12995 3125
rect 13029 3123 13404 3125
rect 13029 3091 13157 3123
rect 12782 3089 13157 3091
rect 13191 3089 13249 3123
rect 13283 3089 13341 3123
rect 13375 3089 13404 3123
rect 12782 3058 13404 3089
rect 13474 3130 13750 3148
rect 13474 3117 13597 3130
rect 13649 3117 13750 3130
rect 13826 3126 13884 3134
rect 13474 3083 13503 3117
rect 13537 3083 13595 3117
rect 13649 3083 13687 3117
rect 13721 3083 13750 3117
rect 13474 3078 13597 3083
rect 13649 3078 13750 3083
rect 12782 2782 12880 3058
rect 13474 3052 13750 3078
rect 13818 3120 13892 3126
rect 13818 3068 13829 3120
rect 13881 3068 13892 3120
rect 13972 3110 14042 3176
rect 14074 3183 14132 3198
rect 14074 3149 14086 3183
rect 14120 3149 14132 3183
rect 14074 3132 14132 3149
rect 13818 3062 13892 3068
rect 13826 3056 13884 3062
rect 13542 2782 13626 3052
rect 13992 3030 14042 3110
rect 14186 3102 14244 3120
rect 14186 3068 14198 3102
rect 14232 3068 14244 3102
rect 14186 3058 14244 3068
rect 14274 3030 14320 3230
rect 13992 3018 14094 3030
rect 13992 2984 14054 3018
rect 14088 2984 14094 3018
rect 13992 2946 14094 2984
rect 14144 3018 14190 3030
rect 14144 2984 14150 3018
rect 14184 2984 14190 3018
rect 14144 2964 14190 2984
rect 14240 3018 14320 3030
rect 14240 2984 14246 3018
rect 14280 2984 14320 3018
rect 13992 2912 14054 2946
rect 14088 2912 14094 2946
rect 13992 2900 14094 2912
rect 14134 2958 14200 2964
rect 14134 2906 14142 2958
rect 14194 2906 14200 2958
rect 14134 2900 14200 2906
rect 14240 2946 14320 2984
rect 14240 2912 14246 2946
rect 14280 2912 14320 2946
rect 14348 3236 14408 3468
rect 14462 3471 14508 3509
rect 14462 3437 14468 3471
rect 14502 3437 14508 3471
rect 14462 3390 14508 3437
rect 14550 3509 14556 3543
rect 14590 3509 14596 3543
rect 14550 3471 14596 3509
rect 14550 3437 14556 3471
rect 14590 3437 14596 3471
rect 14550 3390 14596 3437
rect 15704 3543 15750 3564
rect 15704 3509 15710 3543
rect 15744 3509 15750 3543
rect 15704 3471 15750 3509
rect 15704 3437 15710 3471
rect 15744 3437 15750 3471
rect 15704 3390 15750 3437
rect 15792 3570 15838 3590
rect 15972 3585 16001 3619
rect 16035 3585 16062 3619
rect 15792 3564 15860 3570
rect 15972 3564 16062 3585
rect 15792 3543 15800 3564
rect 15792 3509 15798 3543
rect 15852 3512 15860 3564
rect 15832 3509 15860 3512
rect 15792 3504 15860 3509
rect 16058 3528 16116 3530
rect 16264 3528 16298 3674
rect 16384 3671 16450 3682
rect 16384 3637 16400 3671
rect 16434 3637 16450 3671
rect 16384 3626 16450 3637
rect 16558 3672 17182 3704
rect 17270 3692 17348 4650
rect 17862 4641 17891 4650
rect 17925 4650 19779 4675
rect 17925 4641 17952 4650
rect 17862 4620 17952 4641
rect 17948 4584 18006 4586
rect 17948 4567 18010 4584
rect 17948 4533 17960 4567
rect 17994 4533 18010 4567
rect 17948 4524 18010 4533
rect 17448 4486 17814 4490
rect 17896 4486 17962 4494
rect 17448 4458 17856 4486
rect 17448 4420 17476 4458
rect 17770 4439 17856 4458
rect 17448 4412 17514 4420
rect 17448 4378 17463 4412
rect 17497 4378 17514 4412
rect 17448 4366 17514 4378
rect 17620 4416 17688 4422
rect 17620 4364 17630 4416
rect 17682 4364 17688 4416
rect 17620 4358 17688 4364
rect 17770 4405 17816 4439
rect 17850 4405 17856 4439
rect 17896 4434 17902 4486
rect 17954 4434 17962 4486
rect 17896 4426 17912 4434
rect 17770 4367 17856 4405
rect 17770 4333 17816 4367
rect 17850 4333 17856 4367
rect 17530 4304 17598 4310
rect 17530 4252 17538 4304
rect 17590 4252 17598 4304
rect 17530 4242 17598 4252
rect 17770 4286 17856 4333
rect 17906 4405 17912 4426
rect 17946 4426 17962 4434
rect 18002 4454 18330 4486
rect 18002 4439 18098 4454
rect 17946 4405 17952 4426
rect 17906 4367 17952 4405
rect 17906 4333 17912 4367
rect 17946 4333 17952 4367
rect 17906 4286 17952 4333
rect 18002 4405 18008 4439
rect 18042 4405 18098 4439
rect 18302 4418 18330 4454
rect 18002 4367 18098 4405
rect 18002 4333 18008 4367
rect 18042 4333 18098 4367
rect 18260 4410 18330 4418
rect 18260 4376 18275 4410
rect 18309 4376 18330 4410
rect 18260 4358 18330 4376
rect 18436 4418 18500 4424
rect 18436 4366 18442 4418
rect 18494 4366 18500 4418
rect 18436 4360 18500 4366
rect 18002 4286 18098 4333
rect 17428 4171 17704 4202
rect 17428 4137 17457 4171
rect 17491 4137 17549 4171
rect 17583 4137 17641 4171
rect 17675 4137 17704 4171
rect 17428 4106 17704 4137
rect 17770 4086 17820 4286
rect 17852 4239 17910 4254
rect 17852 4205 17864 4239
rect 17898 4205 17910 4239
rect 17852 4188 17910 4205
rect 17964 4158 18022 4176
rect 17964 4124 17976 4158
rect 18010 4124 18022 4158
rect 17964 4114 18022 4124
rect 18052 4086 18098 4286
rect 18348 4302 18412 4308
rect 18348 4250 18354 4302
rect 18406 4250 18412 4302
rect 18348 4244 18412 4250
rect 18242 4171 18518 4202
rect 18242 4137 18271 4171
rect 18305 4137 18363 4171
rect 18397 4137 18455 4171
rect 18489 4137 18518 4171
rect 18242 4134 18518 4137
rect 17410 4069 17474 4076
rect 17410 4036 17416 4069
rect 17468 4036 17474 4069
rect 17586 4069 17650 4076
rect 17586 4036 17592 4069
rect 17468 4017 17592 4036
rect 17644 4017 17650 4069
rect 17416 4008 17650 4017
rect 17770 4074 17872 4086
rect 17770 4040 17832 4074
rect 17866 4040 17872 4074
rect 17770 4002 17872 4040
rect 17922 4074 17968 4086
rect 17922 4040 17928 4074
rect 17962 4040 17968 4074
rect 17922 4020 17968 4040
rect 18018 4074 18098 4086
rect 18018 4040 18024 4074
rect 18058 4040 18098 4074
rect 17770 3970 17832 4002
rect 17566 3968 17832 3970
rect 17866 3968 17872 4002
rect 17566 3956 17872 3968
rect 17912 4014 17978 4020
rect 17912 3962 17920 4014
rect 17972 3962 17978 4014
rect 17912 3956 17978 3962
rect 18018 4002 18098 4040
rect 18018 3968 18024 4002
rect 18058 3968 18098 4002
rect 18214 4106 18518 4134
rect 18018 3956 18064 3968
rect 17566 3942 17820 3956
rect 17410 3936 17476 3942
rect 17410 3884 17418 3936
rect 17470 3884 17476 3936
rect 17410 3878 17476 3884
rect 16558 3669 16588 3672
rect 16640 3669 17182 3672
rect 16558 3635 16587 3669
rect 16640 3635 16679 3669
rect 16713 3635 16771 3669
rect 16805 3667 17182 3669
rect 16805 3635 16933 3667
rect 16558 3620 16588 3635
rect 16640 3633 16933 3635
rect 16967 3633 17025 3667
rect 17059 3633 17117 3667
rect 17151 3633 17182 3667
rect 16640 3620 17182 3633
rect 16558 3602 17182 3620
rect 17250 3678 17526 3692
rect 17250 3661 17442 3678
rect 17494 3661 17526 3678
rect 17250 3627 17279 3661
rect 17313 3627 17371 3661
rect 17405 3627 17442 3661
rect 17497 3627 17526 3661
rect 17250 3626 17442 3627
rect 17494 3626 17526 3627
rect 17250 3596 17526 3626
rect 17566 3592 17594 3942
rect 17866 3918 17930 3928
rect 17866 3884 17880 3918
rect 17914 3884 18186 3918
rect 17866 3866 17930 3884
rect 17782 3820 17854 3832
rect 17782 3768 17792 3820
rect 17844 3768 17854 3820
rect 17782 3756 17854 3768
rect 18152 3702 18186 3884
rect 18214 3802 18242 4106
rect 18214 3792 18282 3802
rect 18214 3758 18230 3792
rect 18264 3758 18282 3792
rect 18214 3744 18282 3758
rect 17626 3674 18186 3702
rect 17626 3671 17692 3674
rect 17626 3637 17642 3671
rect 17676 3637 17692 3671
rect 17626 3628 17692 3637
rect 17860 3619 17950 3640
rect 16058 3511 16298 3528
rect 16342 3584 16408 3590
rect 16342 3532 16350 3584
rect 16402 3532 16408 3584
rect 16342 3526 16356 3532
rect 15792 3471 15838 3504
rect 15792 3437 15798 3471
rect 15832 3437 15838 3471
rect 16058 3477 16070 3511
rect 16104 3500 16298 3511
rect 16350 3509 16356 3526
rect 16390 3526 16408 3532
rect 16438 3543 16484 3590
rect 17566 3564 17638 3592
rect 16390 3509 16396 3526
rect 16104 3477 16296 3500
rect 16058 3468 16296 3477
rect 15792 3390 15838 3437
rect 16006 3430 16072 3438
rect 15920 3426 15966 3430
rect 15036 3368 15108 3372
rect 14496 3343 14562 3356
rect 14496 3309 14512 3343
rect 14546 3309 14562 3343
rect 14496 3300 14562 3309
rect 15036 3316 15045 3368
rect 15097 3316 15108 3368
rect 15036 3304 15108 3316
rect 15232 3366 15306 3386
rect 15880 3383 15966 3426
rect 15232 3332 15244 3366
rect 15278 3332 15306 3366
rect 15232 3308 15306 3332
rect 15342 3372 15410 3378
rect 15342 3320 15349 3372
rect 15401 3366 15410 3372
rect 15401 3360 15494 3366
rect 15401 3326 15440 3360
rect 15474 3326 15494 3360
rect 15401 3320 15494 3326
rect 15342 3316 15494 3320
rect 15738 3343 15804 3354
rect 15342 3314 15410 3316
rect 15738 3309 15754 3343
rect 15788 3309 15804 3343
rect 15738 3296 15804 3309
rect 15880 3349 15926 3383
rect 15960 3349 15966 3383
rect 16006 3378 16012 3430
rect 16064 3378 16072 3430
rect 16006 3370 16022 3378
rect 15880 3311 15966 3349
rect 15880 3277 15926 3311
rect 15960 3277 15966 3311
rect 14818 3256 14876 3270
rect 14818 3236 14830 3256
rect 14348 3222 14830 3236
rect 14864 3222 14876 3256
rect 14348 3202 14876 3222
rect 15880 3230 15966 3277
rect 16016 3349 16022 3370
rect 16056 3370 16072 3378
rect 16112 3383 16208 3430
rect 16056 3349 16062 3370
rect 16016 3311 16062 3349
rect 16016 3277 16022 3311
rect 16056 3277 16062 3311
rect 16016 3230 16062 3277
rect 16112 3349 16118 3383
rect 16152 3349 16208 3383
rect 16112 3311 16208 3349
rect 16112 3277 16118 3311
rect 16152 3277 16208 3311
rect 16112 3230 16208 3277
rect 14240 2900 14286 2912
rect 14348 2872 14408 3202
rect 15880 3176 15930 3230
rect 14454 3152 14530 3158
rect 14454 3100 14462 3152
rect 14514 3100 14530 3152
rect 14454 3094 14530 3100
rect 14670 3125 15292 3156
rect 14088 2862 14408 2872
rect 14088 2828 14102 2862
rect 14136 2828 14408 2862
rect 14088 2810 14408 2828
rect 14670 3091 14699 3125
rect 14733 3091 14791 3125
rect 14825 3091 14883 3125
rect 14917 3123 15292 3125
rect 14917 3091 15045 3123
rect 14670 3089 15045 3091
rect 15079 3089 15137 3123
rect 15171 3089 15229 3123
rect 15263 3089 15292 3123
rect 14670 3058 15292 3089
rect 15362 3130 15638 3148
rect 15362 3117 15485 3130
rect 15537 3117 15638 3130
rect 15714 3126 15772 3134
rect 15362 3083 15391 3117
rect 15425 3083 15483 3117
rect 15537 3083 15575 3117
rect 15609 3083 15638 3117
rect 15362 3078 15485 3083
rect 15537 3078 15638 3083
rect 14670 2782 14768 3058
rect 15362 3052 15638 3078
rect 15706 3120 15780 3126
rect 15706 3068 15717 3120
rect 15769 3068 15780 3120
rect 15860 3110 15930 3176
rect 15962 3183 16020 3198
rect 15962 3149 15974 3183
rect 16008 3149 16020 3183
rect 15962 3132 16020 3149
rect 15706 3062 15780 3068
rect 15714 3056 15772 3062
rect 15430 2782 15514 3052
rect 15880 3030 15930 3110
rect 16074 3102 16132 3120
rect 16074 3068 16086 3102
rect 16120 3068 16132 3102
rect 16074 3058 16132 3068
rect 16162 3030 16208 3230
rect 15880 3018 15982 3030
rect 15880 2984 15942 3018
rect 15976 2984 15982 3018
rect 15880 2946 15982 2984
rect 16032 3018 16078 3030
rect 16032 2984 16038 3018
rect 16072 2984 16078 3018
rect 16032 2964 16078 2984
rect 16128 3018 16208 3030
rect 16128 2984 16134 3018
rect 16168 2984 16208 3018
rect 15880 2912 15942 2946
rect 15976 2912 15982 2946
rect 15880 2900 15982 2912
rect 16022 2958 16088 2964
rect 16022 2906 16030 2958
rect 16082 2906 16088 2958
rect 16022 2900 16088 2906
rect 16128 2946 16208 2984
rect 16128 2912 16134 2946
rect 16168 2912 16208 2946
rect 16236 3236 16296 3468
rect 16350 3471 16396 3509
rect 16350 3437 16356 3471
rect 16390 3437 16396 3471
rect 16350 3390 16396 3437
rect 16438 3509 16444 3543
rect 16478 3509 16484 3543
rect 16438 3471 16484 3509
rect 16438 3437 16444 3471
rect 16478 3437 16484 3471
rect 16438 3390 16484 3437
rect 17592 3543 17638 3564
rect 17592 3509 17598 3543
rect 17632 3509 17638 3543
rect 17592 3471 17638 3509
rect 17592 3437 17598 3471
rect 17632 3437 17638 3471
rect 17592 3390 17638 3437
rect 17680 3570 17726 3590
rect 17860 3585 17889 3619
rect 17923 3585 17950 3619
rect 17680 3564 17748 3570
rect 17860 3564 17950 3585
rect 17680 3543 17688 3564
rect 17680 3509 17686 3543
rect 17740 3512 17748 3564
rect 17720 3509 17748 3512
rect 17680 3504 17748 3509
rect 17946 3528 18004 3530
rect 18152 3528 18186 3674
rect 18272 3671 18338 3682
rect 18272 3637 18288 3671
rect 18322 3637 18338 3671
rect 18272 3626 18338 3637
rect 18446 3672 19070 3704
rect 19158 3692 19236 4650
rect 19750 4641 19779 4650
rect 19813 4650 21667 4675
rect 19813 4641 19840 4650
rect 19750 4620 19840 4641
rect 19836 4584 19894 4586
rect 19836 4567 19898 4584
rect 19836 4533 19848 4567
rect 19882 4533 19898 4567
rect 19836 4524 19898 4533
rect 19336 4486 19702 4490
rect 19784 4486 19850 4494
rect 19336 4458 19744 4486
rect 19336 4420 19364 4458
rect 19658 4439 19744 4458
rect 19336 4412 19402 4420
rect 19336 4378 19351 4412
rect 19385 4378 19402 4412
rect 19336 4366 19402 4378
rect 19508 4416 19576 4422
rect 19508 4364 19518 4416
rect 19570 4364 19576 4416
rect 19508 4358 19576 4364
rect 19658 4405 19704 4439
rect 19738 4405 19744 4439
rect 19784 4434 19790 4486
rect 19842 4434 19850 4486
rect 19784 4426 19800 4434
rect 19658 4367 19744 4405
rect 19658 4333 19704 4367
rect 19738 4333 19744 4367
rect 19418 4304 19486 4310
rect 19418 4252 19426 4304
rect 19478 4252 19486 4304
rect 19418 4242 19486 4252
rect 19658 4286 19744 4333
rect 19794 4405 19800 4426
rect 19834 4426 19850 4434
rect 19890 4454 20218 4486
rect 19890 4439 19986 4454
rect 19834 4405 19840 4426
rect 19794 4367 19840 4405
rect 19794 4333 19800 4367
rect 19834 4333 19840 4367
rect 19794 4286 19840 4333
rect 19890 4405 19896 4439
rect 19930 4405 19986 4439
rect 20190 4418 20218 4454
rect 19890 4367 19986 4405
rect 19890 4333 19896 4367
rect 19930 4333 19986 4367
rect 20148 4410 20218 4418
rect 20148 4376 20163 4410
rect 20197 4376 20218 4410
rect 20148 4358 20218 4376
rect 20324 4418 20388 4424
rect 20324 4366 20330 4418
rect 20382 4366 20388 4418
rect 20324 4360 20388 4366
rect 19890 4286 19986 4333
rect 19316 4171 19592 4202
rect 19316 4137 19345 4171
rect 19379 4137 19437 4171
rect 19471 4137 19529 4171
rect 19563 4137 19592 4171
rect 19316 4106 19592 4137
rect 19658 4086 19708 4286
rect 19740 4239 19798 4254
rect 19740 4205 19752 4239
rect 19786 4205 19798 4239
rect 19740 4188 19798 4205
rect 19852 4158 19910 4176
rect 19852 4124 19864 4158
rect 19898 4124 19910 4158
rect 19852 4114 19910 4124
rect 19940 4086 19986 4286
rect 20236 4302 20300 4308
rect 20236 4250 20242 4302
rect 20294 4250 20300 4302
rect 20236 4244 20300 4250
rect 20130 4171 20406 4202
rect 20130 4137 20159 4171
rect 20193 4137 20251 4171
rect 20285 4137 20343 4171
rect 20377 4137 20406 4171
rect 20130 4134 20406 4137
rect 19298 4069 19362 4076
rect 19298 4036 19304 4069
rect 19356 4036 19362 4069
rect 19474 4069 19538 4076
rect 19474 4036 19480 4069
rect 19356 4017 19480 4036
rect 19532 4017 19538 4069
rect 19304 4008 19538 4017
rect 19658 4074 19760 4086
rect 19658 4040 19720 4074
rect 19754 4040 19760 4074
rect 19658 4002 19760 4040
rect 19810 4074 19856 4086
rect 19810 4040 19816 4074
rect 19850 4040 19856 4074
rect 19810 4020 19856 4040
rect 19906 4074 19986 4086
rect 19906 4040 19912 4074
rect 19946 4040 19986 4074
rect 19658 3970 19720 4002
rect 19454 3968 19720 3970
rect 19754 3968 19760 4002
rect 19454 3956 19760 3968
rect 19800 4014 19866 4020
rect 19800 3962 19808 4014
rect 19860 3962 19866 4014
rect 19800 3956 19866 3962
rect 19906 4002 19986 4040
rect 19906 3968 19912 4002
rect 19946 3968 19986 4002
rect 20102 4106 20406 4134
rect 19906 3956 19952 3968
rect 19454 3942 19708 3956
rect 19298 3936 19364 3942
rect 19298 3884 19306 3936
rect 19358 3884 19364 3936
rect 19298 3878 19364 3884
rect 18446 3669 18476 3672
rect 18528 3669 19070 3672
rect 18446 3635 18475 3669
rect 18528 3635 18567 3669
rect 18601 3635 18659 3669
rect 18693 3667 19070 3669
rect 18693 3635 18821 3667
rect 18446 3620 18476 3635
rect 18528 3633 18821 3635
rect 18855 3633 18913 3667
rect 18947 3633 19005 3667
rect 19039 3633 19070 3667
rect 18528 3620 19070 3633
rect 18446 3602 19070 3620
rect 19138 3678 19414 3692
rect 19138 3661 19330 3678
rect 19382 3661 19414 3678
rect 19138 3627 19167 3661
rect 19201 3627 19259 3661
rect 19293 3627 19330 3661
rect 19385 3627 19414 3661
rect 19138 3626 19330 3627
rect 19382 3626 19414 3627
rect 19138 3596 19414 3626
rect 19454 3592 19482 3942
rect 19754 3918 19818 3928
rect 19754 3884 19768 3918
rect 19802 3884 20074 3918
rect 19754 3866 19818 3884
rect 19670 3820 19742 3832
rect 19670 3768 19680 3820
rect 19732 3768 19742 3820
rect 19670 3756 19742 3768
rect 20040 3702 20074 3884
rect 20102 3802 20130 4106
rect 20102 3792 20170 3802
rect 20102 3758 20118 3792
rect 20152 3758 20170 3792
rect 20102 3744 20170 3758
rect 19514 3674 20074 3702
rect 19514 3671 19580 3674
rect 19514 3637 19530 3671
rect 19564 3637 19580 3671
rect 19514 3628 19580 3637
rect 19748 3619 19838 3640
rect 17946 3511 18186 3528
rect 18230 3584 18296 3590
rect 18230 3532 18238 3584
rect 18290 3532 18296 3584
rect 18230 3526 18244 3532
rect 17680 3471 17726 3504
rect 17680 3437 17686 3471
rect 17720 3437 17726 3471
rect 17946 3477 17958 3511
rect 17992 3500 18186 3511
rect 18238 3509 18244 3526
rect 18278 3526 18296 3532
rect 18326 3543 18372 3590
rect 19454 3564 19526 3592
rect 18278 3509 18284 3526
rect 17992 3477 18184 3500
rect 17946 3468 18184 3477
rect 17680 3390 17726 3437
rect 17894 3430 17960 3438
rect 17808 3426 17854 3430
rect 16924 3368 16996 3372
rect 16384 3343 16450 3356
rect 16384 3309 16400 3343
rect 16434 3309 16450 3343
rect 16384 3300 16450 3309
rect 16924 3316 16933 3368
rect 16985 3316 16996 3368
rect 16924 3304 16996 3316
rect 17120 3366 17194 3386
rect 17768 3383 17854 3426
rect 17120 3332 17132 3366
rect 17166 3332 17194 3366
rect 17120 3308 17194 3332
rect 17230 3372 17298 3378
rect 17230 3320 17237 3372
rect 17289 3366 17298 3372
rect 17289 3360 17382 3366
rect 17289 3326 17328 3360
rect 17362 3326 17382 3360
rect 17289 3320 17382 3326
rect 17230 3316 17382 3320
rect 17626 3343 17692 3354
rect 17230 3314 17298 3316
rect 17626 3309 17642 3343
rect 17676 3309 17692 3343
rect 17626 3296 17692 3309
rect 17768 3349 17814 3383
rect 17848 3349 17854 3383
rect 17894 3378 17900 3430
rect 17952 3378 17960 3430
rect 17894 3370 17910 3378
rect 17768 3311 17854 3349
rect 17768 3277 17814 3311
rect 17848 3277 17854 3311
rect 16706 3256 16764 3270
rect 16706 3236 16718 3256
rect 16236 3222 16718 3236
rect 16752 3222 16764 3256
rect 16236 3202 16764 3222
rect 17768 3230 17854 3277
rect 17904 3349 17910 3370
rect 17944 3370 17960 3378
rect 18000 3383 18096 3430
rect 17944 3349 17950 3370
rect 17904 3311 17950 3349
rect 17904 3277 17910 3311
rect 17944 3277 17950 3311
rect 17904 3230 17950 3277
rect 18000 3349 18006 3383
rect 18040 3349 18096 3383
rect 18000 3311 18096 3349
rect 18000 3277 18006 3311
rect 18040 3277 18096 3311
rect 18000 3230 18096 3277
rect 16128 2900 16174 2912
rect 16236 2872 16296 3202
rect 17768 3176 17818 3230
rect 16342 3152 16418 3158
rect 16342 3100 16350 3152
rect 16402 3100 16418 3152
rect 16342 3094 16418 3100
rect 16558 3125 17180 3156
rect 15976 2862 16296 2872
rect 15976 2828 15990 2862
rect 16024 2828 16296 2862
rect 15976 2810 16296 2828
rect 16558 3091 16587 3125
rect 16621 3091 16679 3125
rect 16713 3091 16771 3125
rect 16805 3123 17180 3125
rect 16805 3091 16933 3123
rect 16558 3089 16933 3091
rect 16967 3089 17025 3123
rect 17059 3089 17117 3123
rect 17151 3089 17180 3123
rect 16558 3058 17180 3089
rect 17250 3130 17526 3148
rect 17250 3117 17373 3130
rect 17425 3117 17526 3130
rect 17602 3126 17660 3134
rect 17250 3083 17279 3117
rect 17313 3083 17371 3117
rect 17425 3083 17463 3117
rect 17497 3083 17526 3117
rect 17250 3078 17373 3083
rect 17425 3078 17526 3083
rect 16558 2782 16656 3058
rect 17250 3052 17526 3078
rect 17594 3120 17668 3126
rect 17594 3068 17605 3120
rect 17657 3068 17668 3120
rect 17748 3110 17818 3176
rect 17850 3183 17908 3198
rect 17850 3149 17862 3183
rect 17896 3149 17908 3183
rect 17850 3132 17908 3149
rect 17594 3062 17668 3068
rect 17602 3056 17660 3062
rect 17318 2782 17402 3052
rect 17768 3030 17818 3110
rect 17962 3102 18020 3120
rect 17962 3068 17974 3102
rect 18008 3068 18020 3102
rect 17962 3058 18020 3068
rect 18050 3030 18096 3230
rect 17768 3018 17870 3030
rect 17768 2984 17830 3018
rect 17864 2984 17870 3018
rect 17768 2946 17870 2984
rect 17920 3018 17966 3030
rect 17920 2984 17926 3018
rect 17960 2984 17966 3018
rect 17920 2964 17966 2984
rect 18016 3018 18096 3030
rect 18016 2984 18022 3018
rect 18056 2984 18096 3018
rect 17768 2912 17830 2946
rect 17864 2912 17870 2946
rect 17768 2900 17870 2912
rect 17910 2958 17976 2964
rect 17910 2906 17918 2958
rect 17970 2906 17976 2958
rect 17910 2900 17976 2906
rect 18016 2946 18096 2984
rect 18016 2912 18022 2946
rect 18056 2912 18096 2946
rect 18124 3236 18184 3468
rect 18238 3471 18284 3509
rect 18238 3437 18244 3471
rect 18278 3437 18284 3471
rect 18238 3390 18284 3437
rect 18326 3509 18332 3543
rect 18366 3509 18372 3543
rect 18326 3471 18372 3509
rect 18326 3437 18332 3471
rect 18366 3437 18372 3471
rect 18326 3390 18372 3437
rect 19480 3543 19526 3564
rect 19480 3509 19486 3543
rect 19520 3509 19526 3543
rect 19480 3471 19526 3509
rect 19480 3437 19486 3471
rect 19520 3437 19526 3471
rect 19480 3390 19526 3437
rect 19568 3570 19614 3590
rect 19748 3585 19777 3619
rect 19811 3585 19838 3619
rect 19568 3564 19636 3570
rect 19748 3564 19838 3585
rect 19568 3543 19576 3564
rect 19568 3509 19574 3543
rect 19628 3512 19636 3564
rect 19608 3509 19636 3512
rect 19568 3504 19636 3509
rect 19834 3528 19892 3530
rect 20040 3528 20074 3674
rect 20160 3671 20226 3682
rect 20160 3637 20176 3671
rect 20210 3637 20226 3671
rect 20160 3626 20226 3637
rect 20334 3672 20958 3704
rect 21046 3692 21124 4650
rect 21638 4641 21667 4650
rect 21701 4650 23555 4675
rect 21701 4641 21728 4650
rect 21638 4620 21728 4641
rect 21724 4584 21782 4586
rect 21724 4567 21786 4584
rect 21724 4533 21736 4567
rect 21770 4533 21786 4567
rect 21724 4524 21786 4533
rect 21224 4486 21590 4490
rect 21672 4486 21738 4494
rect 21224 4458 21632 4486
rect 21224 4420 21252 4458
rect 21546 4439 21632 4458
rect 21224 4412 21290 4420
rect 21224 4378 21239 4412
rect 21273 4378 21290 4412
rect 21224 4366 21290 4378
rect 21396 4416 21464 4422
rect 21396 4364 21406 4416
rect 21458 4364 21464 4416
rect 21396 4358 21464 4364
rect 21546 4405 21592 4439
rect 21626 4405 21632 4439
rect 21672 4434 21678 4486
rect 21730 4434 21738 4486
rect 21672 4426 21688 4434
rect 21546 4367 21632 4405
rect 21546 4333 21592 4367
rect 21626 4333 21632 4367
rect 21306 4304 21374 4310
rect 21306 4252 21314 4304
rect 21366 4252 21374 4304
rect 21306 4242 21374 4252
rect 21546 4286 21632 4333
rect 21682 4405 21688 4426
rect 21722 4426 21738 4434
rect 21778 4454 22106 4486
rect 21778 4439 21874 4454
rect 21722 4405 21728 4426
rect 21682 4367 21728 4405
rect 21682 4333 21688 4367
rect 21722 4333 21728 4367
rect 21682 4286 21728 4333
rect 21778 4405 21784 4439
rect 21818 4405 21874 4439
rect 22078 4418 22106 4454
rect 21778 4367 21874 4405
rect 21778 4333 21784 4367
rect 21818 4333 21874 4367
rect 22036 4410 22106 4418
rect 22036 4376 22051 4410
rect 22085 4376 22106 4410
rect 22036 4358 22106 4376
rect 22212 4418 22276 4424
rect 22212 4366 22218 4418
rect 22270 4366 22276 4418
rect 22212 4360 22276 4366
rect 21778 4286 21874 4333
rect 21204 4171 21480 4202
rect 21204 4137 21233 4171
rect 21267 4137 21325 4171
rect 21359 4137 21417 4171
rect 21451 4137 21480 4171
rect 21204 4106 21480 4137
rect 21546 4086 21596 4286
rect 21628 4239 21686 4254
rect 21628 4205 21640 4239
rect 21674 4205 21686 4239
rect 21628 4188 21686 4205
rect 21740 4158 21798 4176
rect 21740 4124 21752 4158
rect 21786 4124 21798 4158
rect 21740 4114 21798 4124
rect 21828 4086 21874 4286
rect 22124 4302 22188 4308
rect 22124 4250 22130 4302
rect 22182 4250 22188 4302
rect 22124 4244 22188 4250
rect 22018 4171 22294 4202
rect 22018 4137 22047 4171
rect 22081 4137 22139 4171
rect 22173 4137 22231 4171
rect 22265 4137 22294 4171
rect 22018 4134 22294 4137
rect 21186 4069 21250 4076
rect 21186 4036 21192 4069
rect 21244 4036 21250 4069
rect 21362 4069 21426 4076
rect 21362 4036 21368 4069
rect 21244 4017 21368 4036
rect 21420 4017 21426 4069
rect 21192 4008 21426 4017
rect 21546 4074 21648 4086
rect 21546 4040 21608 4074
rect 21642 4040 21648 4074
rect 21546 4002 21648 4040
rect 21698 4074 21744 4086
rect 21698 4040 21704 4074
rect 21738 4040 21744 4074
rect 21698 4020 21744 4040
rect 21794 4074 21874 4086
rect 21794 4040 21800 4074
rect 21834 4040 21874 4074
rect 21546 3970 21608 4002
rect 21342 3968 21608 3970
rect 21642 3968 21648 4002
rect 21342 3956 21648 3968
rect 21688 4014 21754 4020
rect 21688 3962 21696 4014
rect 21748 3962 21754 4014
rect 21688 3956 21754 3962
rect 21794 4002 21874 4040
rect 21794 3968 21800 4002
rect 21834 3968 21874 4002
rect 21990 4106 22294 4134
rect 21794 3956 21840 3968
rect 21342 3942 21596 3956
rect 21186 3936 21252 3942
rect 21186 3884 21194 3936
rect 21246 3884 21252 3936
rect 21186 3878 21252 3884
rect 20334 3669 20364 3672
rect 20416 3669 20958 3672
rect 20334 3635 20363 3669
rect 20416 3635 20455 3669
rect 20489 3635 20547 3669
rect 20581 3667 20958 3669
rect 20581 3635 20709 3667
rect 20334 3620 20364 3635
rect 20416 3633 20709 3635
rect 20743 3633 20801 3667
rect 20835 3633 20893 3667
rect 20927 3633 20958 3667
rect 20416 3620 20958 3633
rect 20334 3602 20958 3620
rect 21026 3678 21302 3692
rect 21026 3661 21218 3678
rect 21270 3661 21302 3678
rect 21026 3627 21055 3661
rect 21089 3627 21147 3661
rect 21181 3627 21218 3661
rect 21273 3627 21302 3661
rect 21026 3626 21218 3627
rect 21270 3626 21302 3627
rect 21026 3596 21302 3626
rect 21342 3592 21370 3942
rect 21642 3918 21706 3928
rect 21642 3884 21656 3918
rect 21690 3884 21962 3918
rect 21642 3866 21706 3884
rect 21558 3820 21630 3832
rect 21558 3768 21568 3820
rect 21620 3768 21630 3820
rect 21558 3756 21630 3768
rect 21928 3702 21962 3884
rect 21990 3802 22018 4106
rect 21990 3792 22058 3802
rect 21990 3758 22006 3792
rect 22040 3758 22058 3792
rect 21990 3744 22058 3758
rect 21402 3674 21962 3702
rect 21402 3671 21468 3674
rect 21402 3637 21418 3671
rect 21452 3637 21468 3671
rect 21402 3628 21468 3637
rect 21636 3619 21726 3640
rect 19834 3511 20074 3528
rect 20118 3584 20184 3590
rect 20118 3532 20126 3584
rect 20178 3532 20184 3584
rect 20118 3526 20132 3532
rect 19568 3471 19614 3504
rect 19568 3437 19574 3471
rect 19608 3437 19614 3471
rect 19834 3477 19846 3511
rect 19880 3500 20074 3511
rect 20126 3509 20132 3526
rect 20166 3526 20184 3532
rect 20214 3543 20260 3590
rect 21342 3564 21414 3592
rect 20166 3509 20172 3526
rect 19880 3477 20072 3500
rect 19834 3468 20072 3477
rect 19568 3390 19614 3437
rect 19782 3430 19848 3438
rect 19696 3426 19742 3430
rect 18812 3368 18884 3372
rect 18272 3343 18338 3356
rect 18272 3309 18288 3343
rect 18322 3309 18338 3343
rect 18272 3300 18338 3309
rect 18812 3316 18821 3368
rect 18873 3316 18884 3368
rect 18812 3304 18884 3316
rect 19008 3366 19082 3386
rect 19656 3383 19742 3426
rect 19008 3332 19020 3366
rect 19054 3332 19082 3366
rect 19008 3308 19082 3332
rect 19118 3372 19186 3378
rect 19118 3320 19125 3372
rect 19177 3366 19186 3372
rect 19177 3360 19270 3366
rect 19177 3326 19216 3360
rect 19250 3326 19270 3360
rect 19177 3320 19270 3326
rect 19118 3316 19270 3320
rect 19514 3343 19580 3354
rect 19118 3314 19186 3316
rect 19514 3309 19530 3343
rect 19564 3309 19580 3343
rect 19514 3296 19580 3309
rect 19656 3349 19702 3383
rect 19736 3349 19742 3383
rect 19782 3378 19788 3430
rect 19840 3378 19848 3430
rect 19782 3370 19798 3378
rect 19656 3311 19742 3349
rect 19656 3277 19702 3311
rect 19736 3277 19742 3311
rect 18594 3256 18652 3270
rect 18594 3236 18606 3256
rect 18124 3222 18606 3236
rect 18640 3222 18652 3256
rect 18124 3202 18652 3222
rect 19656 3230 19742 3277
rect 19792 3349 19798 3370
rect 19832 3370 19848 3378
rect 19888 3383 19984 3430
rect 19832 3349 19838 3370
rect 19792 3311 19838 3349
rect 19792 3277 19798 3311
rect 19832 3277 19838 3311
rect 19792 3230 19838 3277
rect 19888 3349 19894 3383
rect 19928 3349 19984 3383
rect 19888 3311 19984 3349
rect 19888 3277 19894 3311
rect 19928 3277 19984 3311
rect 19888 3230 19984 3277
rect 18016 2900 18062 2912
rect 18124 2872 18184 3202
rect 19656 3176 19706 3230
rect 18230 3152 18306 3158
rect 18230 3100 18238 3152
rect 18290 3100 18306 3152
rect 18230 3094 18306 3100
rect 18446 3125 19068 3156
rect 17864 2862 18184 2872
rect 17864 2828 17878 2862
rect 17912 2828 18184 2862
rect 17864 2810 18184 2828
rect 18446 3091 18475 3125
rect 18509 3091 18567 3125
rect 18601 3091 18659 3125
rect 18693 3123 19068 3125
rect 18693 3091 18821 3123
rect 18446 3089 18821 3091
rect 18855 3089 18913 3123
rect 18947 3089 19005 3123
rect 19039 3089 19068 3123
rect 18446 3058 19068 3089
rect 19138 3130 19414 3148
rect 19138 3117 19261 3130
rect 19313 3117 19414 3130
rect 19490 3126 19548 3134
rect 19138 3083 19167 3117
rect 19201 3083 19259 3117
rect 19313 3083 19351 3117
rect 19385 3083 19414 3117
rect 19138 3078 19261 3083
rect 19313 3078 19414 3083
rect 18446 2782 18544 3058
rect 19138 3052 19414 3078
rect 19482 3120 19556 3126
rect 19482 3068 19493 3120
rect 19545 3068 19556 3120
rect 19636 3110 19706 3176
rect 19738 3183 19796 3198
rect 19738 3149 19750 3183
rect 19784 3149 19796 3183
rect 19738 3132 19796 3149
rect 19482 3062 19556 3068
rect 19490 3056 19548 3062
rect 19206 2782 19290 3052
rect 19656 3030 19706 3110
rect 19850 3102 19908 3120
rect 19850 3068 19862 3102
rect 19896 3068 19908 3102
rect 19850 3058 19908 3068
rect 19938 3030 19984 3230
rect 19656 3018 19758 3030
rect 19656 2984 19718 3018
rect 19752 2984 19758 3018
rect 19656 2946 19758 2984
rect 19808 3018 19854 3030
rect 19808 2984 19814 3018
rect 19848 2984 19854 3018
rect 19808 2964 19854 2984
rect 19904 3018 19984 3030
rect 19904 2984 19910 3018
rect 19944 2984 19984 3018
rect 19656 2912 19718 2946
rect 19752 2912 19758 2946
rect 19656 2900 19758 2912
rect 19798 2958 19864 2964
rect 19798 2906 19806 2958
rect 19858 2906 19864 2958
rect 19798 2900 19864 2906
rect 19904 2946 19984 2984
rect 19904 2912 19910 2946
rect 19944 2912 19984 2946
rect 20012 3236 20072 3468
rect 20126 3471 20172 3509
rect 20126 3437 20132 3471
rect 20166 3437 20172 3471
rect 20126 3390 20172 3437
rect 20214 3509 20220 3543
rect 20254 3509 20260 3543
rect 20214 3471 20260 3509
rect 20214 3437 20220 3471
rect 20254 3437 20260 3471
rect 20214 3390 20260 3437
rect 21368 3543 21414 3564
rect 21368 3509 21374 3543
rect 21408 3509 21414 3543
rect 21368 3471 21414 3509
rect 21368 3437 21374 3471
rect 21408 3437 21414 3471
rect 21368 3390 21414 3437
rect 21456 3570 21502 3590
rect 21636 3585 21665 3619
rect 21699 3585 21726 3619
rect 21456 3564 21524 3570
rect 21636 3564 21726 3585
rect 21456 3543 21464 3564
rect 21456 3509 21462 3543
rect 21516 3512 21524 3564
rect 21496 3509 21524 3512
rect 21456 3504 21524 3509
rect 21722 3528 21780 3530
rect 21928 3528 21962 3674
rect 22048 3671 22114 3682
rect 22048 3637 22064 3671
rect 22098 3637 22114 3671
rect 22048 3626 22114 3637
rect 22222 3672 22846 3704
rect 22934 3692 23012 4650
rect 23526 4641 23555 4650
rect 23589 4650 25443 4675
rect 23589 4641 23616 4650
rect 23526 4620 23616 4641
rect 23612 4584 23670 4586
rect 23612 4567 23674 4584
rect 23612 4533 23624 4567
rect 23658 4533 23674 4567
rect 23612 4524 23674 4533
rect 23112 4486 23478 4490
rect 23560 4486 23626 4494
rect 23112 4458 23520 4486
rect 23112 4420 23140 4458
rect 23434 4439 23520 4458
rect 23112 4412 23178 4420
rect 23112 4378 23127 4412
rect 23161 4378 23178 4412
rect 23112 4366 23178 4378
rect 23284 4416 23352 4422
rect 23284 4364 23294 4416
rect 23346 4364 23352 4416
rect 23284 4358 23352 4364
rect 23434 4405 23480 4439
rect 23514 4405 23520 4439
rect 23560 4434 23566 4486
rect 23618 4434 23626 4486
rect 23560 4426 23576 4434
rect 23434 4367 23520 4405
rect 23434 4333 23480 4367
rect 23514 4333 23520 4367
rect 23194 4304 23262 4310
rect 23194 4252 23202 4304
rect 23254 4252 23262 4304
rect 23194 4242 23262 4252
rect 23434 4286 23520 4333
rect 23570 4405 23576 4426
rect 23610 4426 23626 4434
rect 23666 4454 23994 4486
rect 23666 4439 23762 4454
rect 23610 4405 23616 4426
rect 23570 4367 23616 4405
rect 23570 4333 23576 4367
rect 23610 4333 23616 4367
rect 23570 4286 23616 4333
rect 23666 4405 23672 4439
rect 23706 4405 23762 4439
rect 23966 4418 23994 4454
rect 23666 4367 23762 4405
rect 23666 4333 23672 4367
rect 23706 4333 23762 4367
rect 23924 4410 23994 4418
rect 23924 4376 23939 4410
rect 23973 4376 23994 4410
rect 23924 4358 23994 4376
rect 24100 4418 24164 4424
rect 24100 4366 24106 4418
rect 24158 4366 24164 4418
rect 24100 4360 24164 4366
rect 23666 4286 23762 4333
rect 23092 4171 23368 4202
rect 23092 4137 23121 4171
rect 23155 4137 23213 4171
rect 23247 4137 23305 4171
rect 23339 4137 23368 4171
rect 23092 4106 23368 4137
rect 23434 4086 23484 4286
rect 23516 4239 23574 4254
rect 23516 4205 23528 4239
rect 23562 4205 23574 4239
rect 23516 4188 23574 4205
rect 23628 4158 23686 4176
rect 23628 4124 23640 4158
rect 23674 4124 23686 4158
rect 23628 4114 23686 4124
rect 23716 4086 23762 4286
rect 24012 4302 24076 4308
rect 24012 4250 24018 4302
rect 24070 4250 24076 4302
rect 24012 4244 24076 4250
rect 23906 4171 24182 4202
rect 23906 4137 23935 4171
rect 23969 4137 24027 4171
rect 24061 4137 24119 4171
rect 24153 4137 24182 4171
rect 23906 4134 24182 4137
rect 23074 4069 23138 4076
rect 23074 4036 23080 4069
rect 23132 4036 23138 4069
rect 23250 4069 23314 4076
rect 23250 4036 23256 4069
rect 23132 4017 23256 4036
rect 23308 4017 23314 4069
rect 23080 4008 23314 4017
rect 23434 4074 23536 4086
rect 23434 4040 23496 4074
rect 23530 4040 23536 4074
rect 23434 4002 23536 4040
rect 23586 4074 23632 4086
rect 23586 4040 23592 4074
rect 23626 4040 23632 4074
rect 23586 4020 23632 4040
rect 23682 4074 23762 4086
rect 23682 4040 23688 4074
rect 23722 4040 23762 4074
rect 23434 3970 23496 4002
rect 23230 3968 23496 3970
rect 23530 3968 23536 4002
rect 23230 3956 23536 3968
rect 23576 4014 23642 4020
rect 23576 3962 23584 4014
rect 23636 3962 23642 4014
rect 23576 3956 23642 3962
rect 23682 4002 23762 4040
rect 23682 3968 23688 4002
rect 23722 3968 23762 4002
rect 23878 4106 24182 4134
rect 23682 3956 23728 3968
rect 23230 3942 23484 3956
rect 23074 3936 23140 3942
rect 23074 3884 23082 3936
rect 23134 3884 23140 3936
rect 23074 3878 23140 3884
rect 22222 3669 22252 3672
rect 22304 3669 22846 3672
rect 22222 3635 22251 3669
rect 22304 3635 22343 3669
rect 22377 3635 22435 3669
rect 22469 3667 22846 3669
rect 22469 3635 22597 3667
rect 22222 3620 22252 3635
rect 22304 3633 22597 3635
rect 22631 3633 22689 3667
rect 22723 3633 22781 3667
rect 22815 3633 22846 3667
rect 22304 3620 22846 3633
rect 22222 3602 22846 3620
rect 22914 3678 23190 3692
rect 22914 3661 23106 3678
rect 23158 3661 23190 3678
rect 22914 3627 22943 3661
rect 22977 3627 23035 3661
rect 23069 3627 23106 3661
rect 23161 3627 23190 3661
rect 22914 3626 23106 3627
rect 23158 3626 23190 3627
rect 22914 3596 23190 3626
rect 23230 3592 23258 3942
rect 23530 3918 23594 3928
rect 23530 3884 23544 3918
rect 23578 3884 23850 3918
rect 23530 3866 23594 3884
rect 23446 3820 23518 3832
rect 23446 3768 23456 3820
rect 23508 3768 23518 3820
rect 23446 3756 23518 3768
rect 23816 3702 23850 3884
rect 23878 3802 23906 4106
rect 23878 3792 23946 3802
rect 23878 3758 23894 3792
rect 23928 3758 23946 3792
rect 23878 3744 23946 3758
rect 23290 3674 23850 3702
rect 23290 3671 23356 3674
rect 23290 3637 23306 3671
rect 23340 3637 23356 3671
rect 23290 3628 23356 3637
rect 23524 3619 23614 3640
rect 21722 3511 21962 3528
rect 22006 3584 22072 3590
rect 22006 3532 22014 3584
rect 22066 3532 22072 3584
rect 22006 3526 22020 3532
rect 21456 3471 21502 3504
rect 21456 3437 21462 3471
rect 21496 3437 21502 3471
rect 21722 3477 21734 3511
rect 21768 3500 21962 3511
rect 22014 3509 22020 3526
rect 22054 3526 22072 3532
rect 22102 3543 22148 3590
rect 23230 3564 23302 3592
rect 22054 3509 22060 3526
rect 21768 3477 21960 3500
rect 21722 3468 21960 3477
rect 21456 3390 21502 3437
rect 21670 3430 21736 3438
rect 21584 3426 21630 3430
rect 20700 3368 20772 3372
rect 20160 3343 20226 3356
rect 20160 3309 20176 3343
rect 20210 3309 20226 3343
rect 20160 3300 20226 3309
rect 20700 3316 20709 3368
rect 20761 3316 20772 3368
rect 20700 3304 20772 3316
rect 20896 3366 20970 3386
rect 21544 3383 21630 3426
rect 20896 3332 20908 3366
rect 20942 3332 20970 3366
rect 20896 3308 20970 3332
rect 21006 3372 21074 3378
rect 21006 3320 21013 3372
rect 21065 3366 21074 3372
rect 21065 3360 21158 3366
rect 21065 3326 21104 3360
rect 21138 3326 21158 3360
rect 21065 3320 21158 3326
rect 21006 3316 21158 3320
rect 21402 3343 21468 3354
rect 21006 3314 21074 3316
rect 21402 3309 21418 3343
rect 21452 3309 21468 3343
rect 21402 3296 21468 3309
rect 21544 3349 21590 3383
rect 21624 3349 21630 3383
rect 21670 3378 21676 3430
rect 21728 3378 21736 3430
rect 21670 3370 21686 3378
rect 21544 3311 21630 3349
rect 21544 3277 21590 3311
rect 21624 3277 21630 3311
rect 20482 3256 20540 3270
rect 20482 3236 20494 3256
rect 20012 3222 20494 3236
rect 20528 3222 20540 3256
rect 20012 3202 20540 3222
rect 21544 3230 21630 3277
rect 21680 3349 21686 3370
rect 21720 3370 21736 3378
rect 21776 3383 21872 3430
rect 21720 3349 21726 3370
rect 21680 3311 21726 3349
rect 21680 3277 21686 3311
rect 21720 3277 21726 3311
rect 21680 3230 21726 3277
rect 21776 3349 21782 3383
rect 21816 3349 21872 3383
rect 21776 3311 21872 3349
rect 21776 3277 21782 3311
rect 21816 3277 21872 3311
rect 21776 3230 21872 3277
rect 19904 2900 19950 2912
rect 20012 2872 20072 3202
rect 21544 3176 21594 3230
rect 20118 3152 20194 3158
rect 20118 3100 20126 3152
rect 20178 3100 20194 3152
rect 20118 3094 20194 3100
rect 20334 3125 20956 3156
rect 19752 2862 20072 2872
rect 19752 2828 19766 2862
rect 19800 2828 20072 2862
rect 19752 2810 20072 2828
rect 20334 3091 20363 3125
rect 20397 3091 20455 3125
rect 20489 3091 20547 3125
rect 20581 3123 20956 3125
rect 20581 3091 20709 3123
rect 20334 3089 20709 3091
rect 20743 3089 20801 3123
rect 20835 3089 20893 3123
rect 20927 3089 20956 3123
rect 20334 3058 20956 3089
rect 21026 3130 21302 3148
rect 21026 3117 21149 3130
rect 21201 3117 21302 3130
rect 21378 3126 21436 3134
rect 21026 3083 21055 3117
rect 21089 3083 21147 3117
rect 21201 3083 21239 3117
rect 21273 3083 21302 3117
rect 21026 3078 21149 3083
rect 21201 3078 21302 3083
rect 20334 2782 20432 3058
rect 21026 3052 21302 3078
rect 21370 3120 21444 3126
rect 21370 3068 21381 3120
rect 21433 3068 21444 3120
rect 21524 3110 21594 3176
rect 21626 3183 21684 3198
rect 21626 3149 21638 3183
rect 21672 3149 21684 3183
rect 21626 3132 21684 3149
rect 21370 3062 21444 3068
rect 21378 3056 21436 3062
rect 21094 2782 21178 3052
rect 21544 3030 21594 3110
rect 21738 3102 21796 3120
rect 21738 3068 21750 3102
rect 21784 3068 21796 3102
rect 21738 3058 21796 3068
rect 21826 3030 21872 3230
rect 21544 3018 21646 3030
rect 21544 2984 21606 3018
rect 21640 2984 21646 3018
rect 21544 2946 21646 2984
rect 21696 3018 21742 3030
rect 21696 2984 21702 3018
rect 21736 2984 21742 3018
rect 21696 2964 21742 2984
rect 21792 3018 21872 3030
rect 21792 2984 21798 3018
rect 21832 2984 21872 3018
rect 21544 2912 21606 2946
rect 21640 2912 21646 2946
rect 21544 2900 21646 2912
rect 21686 2958 21752 2964
rect 21686 2906 21694 2958
rect 21746 2906 21752 2958
rect 21686 2900 21752 2906
rect 21792 2946 21872 2984
rect 21792 2912 21798 2946
rect 21832 2912 21872 2946
rect 21900 3236 21960 3468
rect 22014 3471 22060 3509
rect 22014 3437 22020 3471
rect 22054 3437 22060 3471
rect 22014 3390 22060 3437
rect 22102 3509 22108 3543
rect 22142 3509 22148 3543
rect 22102 3471 22148 3509
rect 22102 3437 22108 3471
rect 22142 3437 22148 3471
rect 22102 3390 22148 3437
rect 23256 3543 23302 3564
rect 23256 3509 23262 3543
rect 23296 3509 23302 3543
rect 23256 3471 23302 3509
rect 23256 3437 23262 3471
rect 23296 3437 23302 3471
rect 23256 3390 23302 3437
rect 23344 3570 23390 3590
rect 23524 3585 23553 3619
rect 23587 3585 23614 3619
rect 23344 3564 23412 3570
rect 23524 3564 23614 3585
rect 23344 3543 23352 3564
rect 23344 3509 23350 3543
rect 23404 3512 23412 3564
rect 23384 3509 23412 3512
rect 23344 3504 23412 3509
rect 23610 3528 23668 3530
rect 23816 3528 23850 3674
rect 23936 3671 24002 3682
rect 23936 3637 23952 3671
rect 23986 3637 24002 3671
rect 23936 3626 24002 3637
rect 24110 3672 24734 3704
rect 24822 3692 24900 4650
rect 25414 4641 25443 4650
rect 25477 4650 26658 4675
rect 25477 4641 25504 4650
rect 25414 4620 25504 4641
rect 25500 4584 25558 4586
rect 25500 4567 25562 4584
rect 25500 4533 25512 4567
rect 25546 4533 25562 4567
rect 25500 4524 25562 4533
rect 25000 4486 25366 4490
rect 25448 4486 25514 4494
rect 25000 4458 25408 4486
rect 25000 4420 25028 4458
rect 25322 4439 25408 4458
rect 25000 4412 25066 4420
rect 25000 4378 25015 4412
rect 25049 4378 25066 4412
rect 25000 4366 25066 4378
rect 25172 4416 25240 4422
rect 25172 4364 25182 4416
rect 25234 4364 25240 4416
rect 25172 4358 25240 4364
rect 25322 4405 25368 4439
rect 25402 4405 25408 4439
rect 25448 4434 25454 4486
rect 25506 4434 25514 4486
rect 25448 4426 25464 4434
rect 25322 4367 25408 4405
rect 25322 4333 25368 4367
rect 25402 4333 25408 4367
rect 25082 4304 25150 4310
rect 25082 4252 25090 4304
rect 25142 4252 25150 4304
rect 25082 4242 25150 4252
rect 25322 4286 25408 4333
rect 25458 4405 25464 4426
rect 25498 4426 25514 4434
rect 25554 4454 25882 4486
rect 25554 4439 25650 4454
rect 25498 4405 25504 4426
rect 25458 4367 25504 4405
rect 25458 4333 25464 4367
rect 25498 4333 25504 4367
rect 25458 4286 25504 4333
rect 25554 4405 25560 4439
rect 25594 4405 25650 4439
rect 25854 4418 25882 4454
rect 25554 4367 25650 4405
rect 25554 4333 25560 4367
rect 25594 4333 25650 4367
rect 25812 4410 25882 4418
rect 25812 4376 25827 4410
rect 25861 4376 25882 4410
rect 25812 4358 25882 4376
rect 25988 4418 26052 4424
rect 25988 4366 25994 4418
rect 26046 4366 26052 4418
rect 25988 4360 26052 4366
rect 25554 4286 25650 4333
rect 24980 4171 25256 4202
rect 24980 4137 25009 4171
rect 25043 4137 25101 4171
rect 25135 4137 25193 4171
rect 25227 4137 25256 4171
rect 24980 4106 25256 4137
rect 25322 4086 25372 4286
rect 25404 4239 25462 4254
rect 25404 4205 25416 4239
rect 25450 4205 25462 4239
rect 25404 4188 25462 4205
rect 25516 4158 25574 4176
rect 25516 4124 25528 4158
rect 25562 4124 25574 4158
rect 25516 4114 25574 4124
rect 25604 4086 25650 4286
rect 25900 4302 25964 4308
rect 25900 4250 25906 4302
rect 25958 4250 25964 4302
rect 25900 4244 25964 4250
rect 25794 4171 26070 4202
rect 25794 4137 25823 4171
rect 25857 4137 25915 4171
rect 25949 4137 26007 4171
rect 26041 4137 26070 4171
rect 25794 4134 26070 4137
rect 24962 4069 25026 4076
rect 24962 4036 24968 4069
rect 25020 4036 25026 4069
rect 25138 4069 25202 4076
rect 25138 4036 25144 4069
rect 25020 4017 25144 4036
rect 25196 4017 25202 4069
rect 24968 4008 25202 4017
rect 25322 4074 25424 4086
rect 25322 4040 25384 4074
rect 25418 4040 25424 4074
rect 25322 4002 25424 4040
rect 25474 4074 25520 4086
rect 25474 4040 25480 4074
rect 25514 4040 25520 4074
rect 25474 4020 25520 4040
rect 25570 4074 25650 4086
rect 25570 4040 25576 4074
rect 25610 4040 25650 4074
rect 25322 3970 25384 4002
rect 25118 3968 25384 3970
rect 25418 3968 25424 4002
rect 25118 3956 25424 3968
rect 25464 4014 25530 4020
rect 25464 3962 25472 4014
rect 25524 3962 25530 4014
rect 25464 3956 25530 3962
rect 25570 4002 25650 4040
rect 25570 3968 25576 4002
rect 25610 3968 25650 4002
rect 25766 4106 26070 4134
rect 25570 3956 25616 3968
rect 25118 3942 25372 3956
rect 24962 3936 25028 3942
rect 24962 3884 24970 3936
rect 25022 3884 25028 3936
rect 24962 3878 25028 3884
rect 24110 3669 24140 3672
rect 24192 3669 24734 3672
rect 24110 3635 24139 3669
rect 24192 3635 24231 3669
rect 24265 3635 24323 3669
rect 24357 3667 24734 3669
rect 24357 3635 24485 3667
rect 24110 3620 24140 3635
rect 24192 3633 24485 3635
rect 24519 3633 24577 3667
rect 24611 3633 24669 3667
rect 24703 3633 24734 3667
rect 24192 3620 24734 3633
rect 24110 3602 24734 3620
rect 24802 3678 25078 3692
rect 24802 3661 24994 3678
rect 25046 3661 25078 3678
rect 24802 3627 24831 3661
rect 24865 3627 24923 3661
rect 24957 3627 24994 3661
rect 25049 3627 25078 3661
rect 24802 3626 24994 3627
rect 25046 3626 25078 3627
rect 24802 3596 25078 3626
rect 25118 3592 25146 3942
rect 25418 3918 25482 3928
rect 25418 3884 25432 3918
rect 25466 3884 25738 3918
rect 25418 3866 25482 3884
rect 25334 3820 25406 3832
rect 25334 3768 25344 3820
rect 25396 3768 25406 3820
rect 25334 3756 25406 3768
rect 25704 3702 25738 3884
rect 25766 3802 25794 4106
rect 25766 3792 25834 3802
rect 25766 3758 25782 3792
rect 25816 3758 25834 3792
rect 25766 3744 25834 3758
rect 25178 3674 25738 3702
rect 25178 3671 25244 3674
rect 25178 3637 25194 3671
rect 25228 3637 25244 3671
rect 25178 3628 25244 3637
rect 25412 3619 25502 3640
rect 23610 3511 23850 3528
rect 23894 3584 23960 3590
rect 23894 3532 23902 3584
rect 23954 3532 23960 3584
rect 23894 3526 23908 3532
rect 23344 3471 23390 3504
rect 23344 3437 23350 3471
rect 23384 3437 23390 3471
rect 23610 3477 23622 3511
rect 23656 3500 23850 3511
rect 23902 3509 23908 3526
rect 23942 3526 23960 3532
rect 23990 3543 24036 3590
rect 25118 3564 25190 3592
rect 23942 3509 23948 3526
rect 23656 3477 23848 3500
rect 23610 3468 23848 3477
rect 23344 3390 23390 3437
rect 23558 3430 23624 3438
rect 23472 3426 23518 3430
rect 22588 3368 22660 3372
rect 22048 3343 22114 3356
rect 22048 3309 22064 3343
rect 22098 3309 22114 3343
rect 22048 3300 22114 3309
rect 22588 3316 22597 3368
rect 22649 3316 22660 3368
rect 22588 3304 22660 3316
rect 22784 3366 22858 3386
rect 23432 3383 23518 3426
rect 22784 3332 22796 3366
rect 22830 3332 22858 3366
rect 22784 3308 22858 3332
rect 22894 3372 22962 3378
rect 22894 3320 22901 3372
rect 22953 3366 22962 3372
rect 22953 3360 23046 3366
rect 22953 3326 22992 3360
rect 23026 3326 23046 3360
rect 22953 3320 23046 3326
rect 22894 3316 23046 3320
rect 23290 3343 23356 3354
rect 22894 3314 22962 3316
rect 23290 3309 23306 3343
rect 23340 3309 23356 3343
rect 23290 3296 23356 3309
rect 23432 3349 23478 3383
rect 23512 3349 23518 3383
rect 23558 3378 23564 3430
rect 23616 3378 23624 3430
rect 23558 3370 23574 3378
rect 23432 3311 23518 3349
rect 23432 3277 23478 3311
rect 23512 3277 23518 3311
rect 22370 3256 22428 3270
rect 22370 3236 22382 3256
rect 21900 3222 22382 3236
rect 22416 3222 22428 3256
rect 21900 3202 22428 3222
rect 23432 3230 23518 3277
rect 23568 3349 23574 3370
rect 23608 3370 23624 3378
rect 23664 3383 23760 3430
rect 23608 3349 23614 3370
rect 23568 3311 23614 3349
rect 23568 3277 23574 3311
rect 23608 3277 23614 3311
rect 23568 3230 23614 3277
rect 23664 3349 23670 3383
rect 23704 3349 23760 3383
rect 23664 3311 23760 3349
rect 23664 3277 23670 3311
rect 23704 3277 23760 3311
rect 23664 3230 23760 3277
rect 21792 2900 21838 2912
rect 21900 2872 21960 3202
rect 23432 3176 23482 3230
rect 22006 3152 22082 3158
rect 22006 3100 22014 3152
rect 22066 3100 22082 3152
rect 22006 3094 22082 3100
rect 22222 3125 22844 3156
rect 21640 2862 21960 2872
rect 21640 2828 21654 2862
rect 21688 2828 21960 2862
rect 21640 2810 21960 2828
rect 22222 3091 22251 3125
rect 22285 3091 22343 3125
rect 22377 3091 22435 3125
rect 22469 3123 22844 3125
rect 22469 3091 22597 3123
rect 22222 3089 22597 3091
rect 22631 3089 22689 3123
rect 22723 3089 22781 3123
rect 22815 3089 22844 3123
rect 22222 3058 22844 3089
rect 22914 3130 23190 3148
rect 22914 3117 23037 3130
rect 23089 3117 23190 3130
rect 23266 3126 23324 3134
rect 22914 3083 22943 3117
rect 22977 3083 23035 3117
rect 23089 3083 23127 3117
rect 23161 3083 23190 3117
rect 22914 3078 23037 3083
rect 23089 3078 23190 3083
rect 22222 2782 22320 3058
rect 22914 3052 23190 3078
rect 23258 3120 23332 3126
rect 23258 3068 23269 3120
rect 23321 3068 23332 3120
rect 23412 3110 23482 3176
rect 23514 3183 23572 3198
rect 23514 3149 23526 3183
rect 23560 3149 23572 3183
rect 23514 3132 23572 3149
rect 23258 3062 23332 3068
rect 23266 3056 23324 3062
rect 22982 2782 23066 3052
rect 23432 3030 23482 3110
rect 23626 3102 23684 3120
rect 23626 3068 23638 3102
rect 23672 3068 23684 3102
rect 23626 3058 23684 3068
rect 23714 3030 23760 3230
rect 23432 3018 23534 3030
rect 23432 2984 23494 3018
rect 23528 2984 23534 3018
rect 23432 2946 23534 2984
rect 23584 3018 23630 3030
rect 23584 2984 23590 3018
rect 23624 2984 23630 3018
rect 23584 2964 23630 2984
rect 23680 3018 23760 3030
rect 23680 2984 23686 3018
rect 23720 2984 23760 3018
rect 23432 2912 23494 2946
rect 23528 2912 23534 2946
rect 23432 2900 23534 2912
rect 23574 2958 23640 2964
rect 23574 2906 23582 2958
rect 23634 2906 23640 2958
rect 23574 2900 23640 2906
rect 23680 2946 23760 2984
rect 23680 2912 23686 2946
rect 23720 2912 23760 2946
rect 23788 3236 23848 3468
rect 23902 3471 23948 3509
rect 23902 3437 23908 3471
rect 23942 3437 23948 3471
rect 23902 3390 23948 3437
rect 23990 3509 23996 3543
rect 24030 3509 24036 3543
rect 23990 3471 24036 3509
rect 23990 3437 23996 3471
rect 24030 3437 24036 3471
rect 23990 3390 24036 3437
rect 25144 3543 25190 3564
rect 25144 3509 25150 3543
rect 25184 3509 25190 3543
rect 25144 3471 25190 3509
rect 25144 3437 25150 3471
rect 25184 3437 25190 3471
rect 25144 3390 25190 3437
rect 25232 3570 25278 3590
rect 25412 3585 25441 3619
rect 25475 3585 25502 3619
rect 25232 3564 25300 3570
rect 25412 3564 25502 3585
rect 25232 3543 25240 3564
rect 25232 3509 25238 3543
rect 25292 3512 25300 3564
rect 25272 3509 25300 3512
rect 25232 3504 25300 3509
rect 25498 3528 25556 3530
rect 25704 3528 25738 3674
rect 25824 3671 25890 3682
rect 25824 3637 25840 3671
rect 25874 3637 25890 3671
rect 25824 3626 25890 3637
rect 25998 3672 26622 3704
rect 25998 3669 26028 3672
rect 26080 3669 26622 3672
rect 25998 3635 26027 3669
rect 26080 3635 26119 3669
rect 26153 3635 26211 3669
rect 26245 3667 26622 3669
rect 26245 3635 26373 3667
rect 25998 3620 26028 3635
rect 26080 3633 26373 3635
rect 26407 3633 26465 3667
rect 26499 3633 26557 3667
rect 26591 3633 26622 3667
rect 26080 3620 26622 3633
rect 25998 3602 26622 3620
rect 25498 3511 25738 3528
rect 25782 3584 25848 3590
rect 25782 3532 25790 3584
rect 25842 3532 25848 3584
rect 25782 3526 25796 3532
rect 25232 3471 25278 3504
rect 25232 3437 25238 3471
rect 25272 3437 25278 3471
rect 25498 3477 25510 3511
rect 25544 3500 25738 3511
rect 25790 3509 25796 3526
rect 25830 3526 25848 3532
rect 25878 3543 25924 3590
rect 25830 3509 25836 3526
rect 25544 3477 25736 3500
rect 25498 3468 25736 3477
rect 25232 3390 25278 3437
rect 25446 3430 25512 3438
rect 25360 3426 25406 3430
rect 24476 3368 24548 3372
rect 23936 3343 24002 3356
rect 23936 3309 23952 3343
rect 23986 3309 24002 3343
rect 23936 3300 24002 3309
rect 24476 3316 24485 3368
rect 24537 3316 24548 3368
rect 24476 3304 24548 3316
rect 24672 3366 24746 3386
rect 25320 3383 25406 3426
rect 24672 3332 24684 3366
rect 24718 3332 24746 3366
rect 24672 3308 24746 3332
rect 24782 3372 24850 3378
rect 24782 3320 24789 3372
rect 24841 3366 24850 3372
rect 24841 3360 24934 3366
rect 24841 3326 24880 3360
rect 24914 3326 24934 3360
rect 24841 3320 24934 3326
rect 24782 3316 24934 3320
rect 25178 3343 25244 3354
rect 24782 3314 24850 3316
rect 25178 3309 25194 3343
rect 25228 3309 25244 3343
rect 25178 3296 25244 3309
rect 25320 3349 25366 3383
rect 25400 3349 25406 3383
rect 25446 3378 25452 3430
rect 25504 3378 25512 3430
rect 25446 3370 25462 3378
rect 25320 3311 25406 3349
rect 25320 3277 25366 3311
rect 25400 3277 25406 3311
rect 24258 3256 24316 3270
rect 24258 3236 24270 3256
rect 23788 3222 24270 3236
rect 24304 3222 24316 3256
rect 23788 3202 24316 3222
rect 25320 3230 25406 3277
rect 25456 3349 25462 3370
rect 25496 3370 25512 3378
rect 25552 3383 25648 3430
rect 25496 3349 25502 3370
rect 25456 3311 25502 3349
rect 25456 3277 25462 3311
rect 25496 3277 25502 3311
rect 25456 3230 25502 3277
rect 25552 3349 25558 3383
rect 25592 3349 25648 3383
rect 25552 3311 25648 3349
rect 25552 3277 25558 3311
rect 25592 3277 25648 3311
rect 25552 3230 25648 3277
rect 23680 2900 23726 2912
rect 23788 2872 23848 3202
rect 25320 3176 25370 3230
rect 23894 3152 23970 3158
rect 23894 3100 23902 3152
rect 23954 3100 23970 3152
rect 23894 3094 23970 3100
rect 24110 3125 24732 3156
rect 23528 2862 23848 2872
rect 23528 2828 23542 2862
rect 23576 2828 23848 2862
rect 23528 2810 23848 2828
rect 24110 3091 24139 3125
rect 24173 3091 24231 3125
rect 24265 3091 24323 3125
rect 24357 3123 24732 3125
rect 24357 3091 24485 3123
rect 24110 3089 24485 3091
rect 24519 3089 24577 3123
rect 24611 3089 24669 3123
rect 24703 3089 24732 3123
rect 24110 3058 24732 3089
rect 24802 3130 25078 3148
rect 24802 3117 24925 3130
rect 24977 3117 25078 3130
rect 25154 3126 25212 3134
rect 24802 3083 24831 3117
rect 24865 3083 24923 3117
rect 24977 3083 25015 3117
rect 25049 3083 25078 3117
rect 24802 3078 24925 3083
rect 24977 3078 25078 3083
rect 24110 2782 24208 3058
rect 24802 3052 25078 3078
rect 25146 3120 25220 3126
rect 25146 3068 25157 3120
rect 25209 3068 25220 3120
rect 25300 3110 25370 3176
rect 25402 3183 25460 3198
rect 25402 3149 25414 3183
rect 25448 3149 25460 3183
rect 25402 3132 25460 3149
rect 25146 3062 25220 3068
rect 25154 3056 25212 3062
rect 24870 2782 24954 3052
rect 25320 3030 25370 3110
rect 25514 3102 25572 3120
rect 25514 3068 25526 3102
rect 25560 3068 25572 3102
rect 25514 3058 25572 3068
rect 25602 3030 25648 3230
rect 25320 3018 25422 3030
rect 25320 2984 25382 3018
rect 25416 2984 25422 3018
rect 25320 2946 25422 2984
rect 25472 3018 25518 3030
rect 25472 2984 25478 3018
rect 25512 2984 25518 3018
rect 25472 2964 25518 2984
rect 25568 3018 25648 3030
rect 25568 2984 25574 3018
rect 25608 2984 25648 3018
rect 25320 2912 25382 2946
rect 25416 2912 25422 2946
rect 25320 2900 25422 2912
rect 25462 2958 25528 2964
rect 25462 2906 25470 2958
rect 25522 2906 25528 2958
rect 25462 2900 25528 2906
rect 25568 2946 25648 2984
rect 25568 2912 25574 2946
rect 25608 2912 25648 2946
rect 25676 3236 25736 3468
rect 25790 3471 25836 3509
rect 25790 3437 25796 3471
rect 25830 3437 25836 3471
rect 25790 3390 25836 3437
rect 25878 3509 25884 3543
rect 25918 3509 25924 3543
rect 25878 3471 25924 3509
rect 25878 3437 25884 3471
rect 25918 3437 25924 3471
rect 25878 3390 25924 3437
rect 26364 3368 26436 3372
rect 25824 3343 25890 3356
rect 25824 3309 25840 3343
rect 25874 3309 25890 3343
rect 25824 3300 25890 3309
rect 26364 3316 26373 3368
rect 26425 3316 26436 3368
rect 26364 3304 26436 3316
rect 26560 3366 26744 3386
rect 26560 3332 26572 3366
rect 26606 3332 26744 3366
rect 26560 3308 26744 3332
rect 26146 3256 26204 3270
rect 26146 3236 26158 3256
rect 25676 3222 26158 3236
rect 26192 3222 26204 3256
rect 25676 3202 26204 3222
rect 25568 2900 25614 2912
rect 25676 2872 25736 3202
rect 25782 3152 25858 3158
rect 25782 3100 25790 3152
rect 25842 3100 25858 3152
rect 25782 3094 25858 3100
rect 25998 3125 26620 3156
rect 25416 2862 25736 2872
rect 25416 2828 25430 2862
rect 25464 2828 25736 2862
rect 25416 2810 25736 2828
rect 25998 3091 26027 3125
rect 26061 3091 26119 3125
rect 26153 3091 26211 3125
rect 26245 3123 26620 3125
rect 26245 3091 26373 3123
rect 25998 3089 26373 3091
rect 26407 3089 26465 3123
rect 26499 3089 26557 3123
rect 26591 3089 26620 3123
rect 25998 3058 26620 3089
rect 25998 2782 26096 3058
rect -3544 2753 26658 2782
rect -3544 2719 -2964 2753
rect -2930 2719 -1076 2753
rect -1042 2719 812 2753
rect 846 2719 2700 2753
rect 2734 2719 4588 2753
rect 4622 2719 6476 2753
rect 6510 2719 8364 2753
rect 8398 2719 10252 2753
rect 10286 2719 12134 2753
rect 12168 2719 14022 2753
rect 14056 2719 15910 2753
rect 15944 2719 17798 2753
rect 17832 2719 19686 2753
rect 19720 2719 21574 2753
rect 21608 2719 23462 2753
rect 23496 2719 25350 2753
rect 25384 2719 26658 2753
rect -3544 2708 26658 2719
rect -3544 2592 -2017 2708
rect -1709 2592 -129 2708
rect 179 2592 1759 2708
rect 2067 2592 3647 2708
rect 3955 2592 5535 2708
rect 5843 2592 7423 2708
rect 7731 2592 9311 2708
rect 9619 2592 11199 2708
rect 11507 2592 13081 2708
rect 13389 2592 14969 2708
rect 15277 2592 16857 2708
rect 17165 2592 18745 2708
rect 19053 2592 20633 2708
rect 20941 2592 22521 2708
rect 22829 2592 24409 2708
rect 24717 2592 26297 2708
rect 26605 2592 26658 2708
rect -3544 2528 26658 2592
<< via1 >>
rect 4610 5337 4683 5343
rect 4610 5303 4667 5337
rect 4667 5303 4683 5337
rect 4610 5290 4683 5303
rect 19704 5337 19780 5343
rect 19704 5303 19707 5337
rect 19707 5303 19765 5337
rect 19765 5303 19780 5337
rect 19704 5289 19780 5303
rect 2282 4950 2334 5002
rect 2389 4971 2411 5002
rect 2411 4971 2441 5002
rect 2389 4950 2441 4971
rect 2495 4950 2547 5002
rect 2611 4950 2663 5002
rect 2740 4971 2746 5004
rect 2746 4971 2780 5004
rect 2780 4971 2792 5004
rect 2740 4952 2792 4971
rect 2874 5001 2926 5003
rect 2874 4967 2915 5001
rect 2915 4967 2926 5001
rect 2874 4951 2926 4967
rect 2991 4951 3043 5003
rect 3096 5000 3148 5003
rect 3096 4966 3118 5000
rect 3118 4966 3148 5000
rect 3096 4951 3148 4966
rect 3202 4972 3250 5003
rect 3250 4972 3254 5003
rect 3202 4951 3254 4972
rect 3299 4951 3351 5003
rect 3396 4974 3420 5003
rect 3420 4974 3448 5003
rect 3396 4951 3448 4974
rect 4171 4947 4223 4999
rect 4278 4971 4294 4999
rect 4294 4971 4328 4999
rect 4328 4971 4330 4999
rect 4278 4947 4330 4971
rect 4384 4947 4436 4999
rect 4500 4947 4552 4999
rect 4622 4975 4630 5002
rect 4630 4975 4664 5002
rect 4664 5001 4674 5002
rect 4664 4975 4681 5001
rect 4622 4950 4681 4975
rect 4629 4949 4681 4950
rect 4763 4996 4815 5000
rect 4763 4962 4794 4996
rect 4794 4962 4815 4996
rect 4763 4948 4815 4962
rect 4880 4948 4932 5000
rect 4985 4968 4998 5000
rect 4998 4968 5037 5000
rect 4985 4948 5037 4968
rect 5091 4970 5134 5000
rect 5134 4970 5143 5000
rect 5091 4948 5143 4970
rect 5188 4948 5240 5000
rect 5285 4972 5293 5000
rect 5293 4972 5327 5000
rect 5327 4972 5337 5000
rect 5285 4948 5337 4972
rect 17391 4956 17443 5008
rect 17503 4996 17555 5006
rect 17503 4962 17506 4996
rect 17506 4962 17540 4996
rect 17540 4962 17555 4996
rect 17503 4954 17555 4962
rect 17610 4954 17662 5006
rect 17712 5000 17764 5006
rect 17712 4966 17713 5000
rect 17713 4966 17764 5000
rect 17712 4954 17764 4966
rect 17838 4971 17844 5004
rect 17844 4971 17878 5004
rect 17878 4971 17890 5004
rect 17838 4952 17890 4971
rect 17992 4992 18044 5004
rect 17992 4958 18011 4992
rect 18011 4958 18044 4992
rect 18129 4990 18181 5004
rect 17992 4952 18044 4958
rect 18129 4956 18179 4990
rect 18179 4956 18181 4990
rect 18129 4952 18181 4956
rect 18226 4952 18278 5004
rect 18326 4999 18378 5004
rect 18326 4965 18349 4999
rect 18349 4965 18378 4999
rect 18326 4952 18378 4965
rect 18415 4951 18467 5003
rect 18511 4951 18563 5003
rect 19225 5000 19277 5002
rect 19225 4966 19256 5000
rect 19256 4966 19277 5000
rect 19225 4950 19277 4966
rect 19319 4950 19371 5002
rect 19418 5001 19470 5002
rect 19418 4967 19429 5001
rect 19429 4967 19470 5001
rect 19418 4950 19470 4967
rect 19526 4972 19557 5002
rect 19557 4972 19578 5002
rect 19526 4950 19578 4972
rect 19622 4950 19674 5002
rect 19720 4975 19728 5002
rect 19728 4975 19762 5002
rect 19762 4975 19772 5002
rect 19720 4950 19772 4975
rect 19839 4949 19891 5001
rect 19953 4949 20005 5001
rect 20070 4995 20122 5001
rect 20070 4961 20096 4995
rect 20096 4961 20122 4995
rect 20070 4949 20122 4961
rect 20197 4993 20249 5001
rect 20197 4959 20232 4993
rect 20232 4959 20249 4993
rect 20197 4949 20249 4959
rect 20312 4949 20364 5001
rect -2017 4716 -1709 4832
rect -129 4716 179 4832
rect 1759 4716 2067 4832
rect 3647 4716 3955 4832
rect 5535 4716 5843 4832
rect 7423 4716 7731 4832
rect 9311 4716 9619 4832
rect 11199 4716 11507 4832
rect 13081 4716 13389 4832
rect 14969 4716 15277 4832
rect 16857 4716 17165 4832
rect 18745 4716 19053 4832
rect 20633 4716 20941 4832
rect 22521 4716 22829 4832
rect 24409 4716 24717 4832
rect 26297 4716 26605 4832
rect -3132 4408 -3080 4416
rect -3132 4374 -3126 4408
rect -3126 4374 -3092 4408
rect -3092 4374 -3080 4408
rect -3132 4364 -3080 4374
rect -2860 4439 -2808 4486
rect -2860 4434 -2850 4439
rect -2850 4434 -2816 4439
rect -2816 4434 -2808 4439
rect -3224 4292 -3172 4304
rect -3224 4258 -3217 4292
rect -3217 4258 -3183 4292
rect -3183 4258 -3172 4292
rect -3224 4252 -3172 4258
rect -2320 4410 -2268 4418
rect -2320 4376 -2313 4410
rect -2313 4376 -2279 4410
rect -2279 4376 -2268 4410
rect -2320 4366 -2268 4376
rect -2408 4287 -2356 4302
rect -2408 4253 -2399 4287
rect -2399 4253 -2365 4287
rect -2365 4253 -2356 4287
rect -2408 4250 -2356 4253
rect -3346 4017 -3294 4069
rect -3170 4017 -3118 4069
rect -2842 4002 -2790 4014
rect -2842 3968 -2834 4002
rect -2834 3968 -2800 4002
rect -2800 3968 -2790 4002
rect -2842 3962 -2790 3968
rect -3344 3926 -3292 3936
rect -3344 3892 -3334 3926
rect -3334 3892 -3300 3926
rect -3300 3892 -3292 3926
rect -3344 3884 -3292 3892
rect -3320 3661 -3268 3678
rect -3320 3627 -3299 3661
rect -3299 3627 -3268 3661
rect -3320 3626 -3268 3627
rect -2970 3809 -2918 3820
rect -2970 3775 -2962 3809
rect -2962 3775 -2928 3809
rect -2928 3775 -2918 3809
rect -2970 3768 -2918 3775
rect -3074 3543 -3022 3564
rect -3074 3512 -3042 3543
rect -3042 3512 -3022 3543
rect -1244 4408 -1192 4416
rect -1244 4374 -1238 4408
rect -1238 4374 -1204 4408
rect -1204 4374 -1192 4408
rect -1244 4364 -1192 4374
rect -972 4439 -920 4486
rect -972 4434 -962 4439
rect -962 4434 -928 4439
rect -928 4434 -920 4439
rect -1336 4292 -1284 4304
rect -1336 4258 -1329 4292
rect -1329 4258 -1295 4292
rect -1295 4258 -1284 4292
rect -1336 4252 -1284 4258
rect -432 4410 -380 4418
rect -432 4376 -425 4410
rect -425 4376 -391 4410
rect -391 4376 -380 4410
rect -432 4366 -380 4376
rect -520 4287 -468 4302
rect -520 4253 -511 4287
rect -511 4253 -477 4287
rect -477 4253 -468 4287
rect -520 4250 -468 4253
rect -1458 4017 -1406 4069
rect -1282 4017 -1230 4069
rect -954 4002 -902 4014
rect -954 3968 -946 4002
rect -946 3968 -912 4002
rect -912 3968 -902 4002
rect -954 3962 -902 3968
rect -1456 3926 -1404 3936
rect -1456 3892 -1446 3926
rect -1446 3892 -1412 3926
rect -1412 3892 -1404 3926
rect -1456 3884 -1404 3892
rect -2286 3669 -2234 3672
rect -2286 3635 -2253 3669
rect -2253 3635 -2234 3669
rect -2286 3620 -2234 3635
rect -1432 3661 -1380 3678
rect -1432 3627 -1411 3661
rect -1411 3627 -1380 3661
rect -1432 3626 -1380 3627
rect -1082 3809 -1030 3820
rect -1082 3775 -1074 3809
rect -1074 3775 -1040 3809
rect -1040 3775 -1030 3809
rect -1082 3768 -1030 3775
rect -2524 3543 -2472 3584
rect -2524 3532 -2518 3543
rect -2518 3532 -2484 3543
rect -2484 3532 -2472 3543
rect -3525 3320 -3473 3372
rect -2862 3383 -2810 3430
rect -2862 3378 -2852 3383
rect -2852 3378 -2818 3383
rect -2818 3378 -2810 3383
rect -3389 3117 -3337 3130
rect -3389 3083 -3357 3117
rect -3357 3083 -3337 3117
rect -3389 3078 -3337 3083
rect -3157 3112 -3105 3120
rect -3157 3078 -3148 3112
rect -3148 3078 -3114 3112
rect -3114 3078 -3105 3112
rect -3157 3068 -3105 3078
rect -2844 2946 -2792 2958
rect -2844 2912 -2836 2946
rect -2836 2912 -2802 2946
rect -2802 2912 -2792 2946
rect -2844 2906 -2792 2912
rect -1186 3543 -1134 3564
rect -1186 3512 -1154 3543
rect -1154 3512 -1134 3543
rect 644 4408 696 4416
rect 644 4374 650 4408
rect 650 4374 684 4408
rect 684 4374 696 4408
rect 644 4364 696 4374
rect 916 4439 968 4486
rect 916 4434 926 4439
rect 926 4434 960 4439
rect 960 4434 968 4439
rect 552 4292 604 4304
rect 552 4258 559 4292
rect 559 4258 593 4292
rect 593 4258 604 4292
rect 552 4252 604 4258
rect 1456 4410 1508 4418
rect 1456 4376 1463 4410
rect 1463 4376 1497 4410
rect 1497 4376 1508 4410
rect 1456 4366 1508 4376
rect 1368 4287 1420 4302
rect 1368 4253 1377 4287
rect 1377 4253 1411 4287
rect 1411 4253 1420 4287
rect 1368 4250 1420 4253
rect 430 4017 482 4069
rect 606 4017 658 4069
rect 934 4002 986 4014
rect 934 3968 942 4002
rect 942 3968 976 4002
rect 976 3968 986 4002
rect 934 3962 986 3968
rect 432 3926 484 3936
rect 432 3892 442 3926
rect 442 3892 476 3926
rect 476 3892 484 3926
rect 432 3884 484 3892
rect -398 3669 -346 3672
rect -398 3635 -365 3669
rect -365 3635 -346 3669
rect -398 3620 -346 3635
rect 456 3661 508 3678
rect 456 3627 477 3661
rect 477 3627 508 3661
rect 456 3626 508 3627
rect 806 3809 858 3820
rect 806 3775 814 3809
rect 814 3775 848 3809
rect 848 3775 858 3809
rect 806 3768 858 3775
rect -636 3543 -584 3584
rect -636 3532 -630 3543
rect -630 3532 -596 3543
rect -596 3532 -584 3543
rect -1941 3354 -1889 3368
rect -1941 3320 -1935 3354
rect -1935 3320 -1901 3354
rect -1901 3320 -1889 3354
rect -1941 3316 -1889 3320
rect -1637 3320 -1585 3372
rect -974 3383 -922 3430
rect -974 3378 -964 3383
rect -964 3378 -930 3383
rect -930 3378 -922 3383
rect -2524 3140 -2472 3152
rect -2524 3106 -2516 3140
rect -2516 3106 -2482 3140
rect -2482 3106 -2472 3140
rect -2524 3100 -2472 3106
rect -1501 3117 -1449 3130
rect -1501 3083 -1469 3117
rect -1469 3083 -1449 3117
rect -1501 3078 -1449 3083
rect -1269 3112 -1217 3120
rect -1269 3078 -1260 3112
rect -1260 3078 -1226 3112
rect -1226 3078 -1217 3112
rect -1269 3068 -1217 3078
rect -956 2946 -904 2958
rect -956 2912 -948 2946
rect -948 2912 -914 2946
rect -914 2912 -904 2946
rect -956 2906 -904 2912
rect 702 3543 754 3564
rect 702 3512 734 3543
rect 734 3512 754 3543
rect 2532 4408 2584 4416
rect 2532 4374 2538 4408
rect 2538 4374 2572 4408
rect 2572 4374 2584 4408
rect 2532 4364 2584 4374
rect 2804 4439 2856 4486
rect 2804 4434 2814 4439
rect 2814 4434 2848 4439
rect 2848 4434 2856 4439
rect 2440 4292 2492 4304
rect 2440 4258 2447 4292
rect 2447 4258 2481 4292
rect 2481 4258 2492 4292
rect 2440 4252 2492 4258
rect 3344 4410 3396 4418
rect 3344 4376 3351 4410
rect 3351 4376 3385 4410
rect 3385 4376 3396 4410
rect 3344 4366 3396 4376
rect 3256 4287 3308 4302
rect 3256 4253 3265 4287
rect 3265 4253 3299 4287
rect 3299 4253 3308 4287
rect 3256 4250 3308 4253
rect 2318 4017 2370 4069
rect 2494 4017 2546 4069
rect 2822 4002 2874 4014
rect 2822 3968 2830 4002
rect 2830 3968 2864 4002
rect 2864 3968 2874 4002
rect 2822 3962 2874 3968
rect 2320 3926 2372 3936
rect 2320 3892 2330 3926
rect 2330 3892 2364 3926
rect 2364 3892 2372 3926
rect 2320 3884 2372 3892
rect 1490 3669 1542 3672
rect 1490 3635 1523 3669
rect 1523 3635 1542 3669
rect 1490 3620 1542 3635
rect 2344 3661 2396 3678
rect 2344 3627 2365 3661
rect 2365 3627 2396 3661
rect 2344 3626 2396 3627
rect 2694 3809 2746 3820
rect 2694 3775 2702 3809
rect 2702 3775 2736 3809
rect 2736 3775 2746 3809
rect 2694 3768 2746 3775
rect 1252 3543 1304 3584
rect 1252 3532 1258 3543
rect 1258 3532 1292 3543
rect 1292 3532 1304 3543
rect -53 3354 -1 3368
rect -53 3320 -47 3354
rect -47 3320 -13 3354
rect -13 3320 -1 3354
rect -53 3316 -1 3320
rect 251 3320 303 3372
rect 914 3383 966 3430
rect 914 3378 924 3383
rect 924 3378 958 3383
rect 958 3378 966 3383
rect -636 3140 -584 3152
rect -636 3106 -628 3140
rect -628 3106 -594 3140
rect -594 3106 -584 3140
rect -636 3100 -584 3106
rect 387 3117 439 3130
rect 387 3083 419 3117
rect 419 3083 439 3117
rect 387 3078 439 3083
rect 619 3112 671 3120
rect 619 3078 628 3112
rect 628 3078 662 3112
rect 662 3078 671 3112
rect 619 3068 671 3078
rect 932 2946 984 2958
rect 932 2912 940 2946
rect 940 2912 974 2946
rect 974 2912 984 2946
rect 932 2906 984 2912
rect 2590 3543 2642 3564
rect 2590 3512 2622 3543
rect 2622 3512 2642 3543
rect 4420 4408 4472 4416
rect 4420 4374 4426 4408
rect 4426 4374 4460 4408
rect 4460 4374 4472 4408
rect 4420 4364 4472 4374
rect 4692 4439 4744 4486
rect 4692 4434 4702 4439
rect 4702 4434 4736 4439
rect 4736 4434 4744 4439
rect 4328 4292 4380 4304
rect 4328 4258 4335 4292
rect 4335 4258 4369 4292
rect 4369 4258 4380 4292
rect 4328 4252 4380 4258
rect 5232 4410 5284 4418
rect 5232 4376 5239 4410
rect 5239 4376 5273 4410
rect 5273 4376 5284 4410
rect 5232 4366 5284 4376
rect 5144 4287 5196 4302
rect 5144 4253 5153 4287
rect 5153 4253 5187 4287
rect 5187 4253 5196 4287
rect 5144 4250 5196 4253
rect 4206 4017 4258 4069
rect 4382 4017 4434 4069
rect 4710 4002 4762 4014
rect 4710 3968 4718 4002
rect 4718 3968 4752 4002
rect 4752 3968 4762 4002
rect 4710 3962 4762 3968
rect 4208 3926 4260 3936
rect 4208 3892 4218 3926
rect 4218 3892 4252 3926
rect 4252 3892 4260 3926
rect 4208 3884 4260 3892
rect 3378 3669 3430 3672
rect 3378 3635 3411 3669
rect 3411 3635 3430 3669
rect 3378 3620 3430 3635
rect 4232 3661 4284 3678
rect 4232 3627 4253 3661
rect 4253 3627 4284 3661
rect 4232 3626 4284 3627
rect 4582 3809 4634 3820
rect 4582 3775 4590 3809
rect 4590 3775 4624 3809
rect 4624 3775 4634 3809
rect 4582 3768 4634 3775
rect 3140 3543 3192 3584
rect 3140 3532 3146 3543
rect 3146 3532 3180 3543
rect 3180 3532 3192 3543
rect 1835 3354 1887 3368
rect 1835 3320 1841 3354
rect 1841 3320 1875 3354
rect 1875 3320 1887 3354
rect 1835 3316 1887 3320
rect 2139 3320 2191 3372
rect 2802 3383 2854 3430
rect 2802 3378 2812 3383
rect 2812 3378 2846 3383
rect 2846 3378 2854 3383
rect 1252 3140 1304 3152
rect 1252 3106 1260 3140
rect 1260 3106 1294 3140
rect 1294 3106 1304 3140
rect 1252 3100 1304 3106
rect 2275 3117 2327 3130
rect 2275 3083 2307 3117
rect 2307 3083 2327 3117
rect 2275 3078 2327 3083
rect 2507 3112 2559 3120
rect 2507 3078 2516 3112
rect 2516 3078 2550 3112
rect 2550 3078 2559 3112
rect 2507 3068 2559 3078
rect 2820 2946 2872 2958
rect 2820 2912 2828 2946
rect 2828 2912 2862 2946
rect 2862 2912 2872 2946
rect 2820 2906 2872 2912
rect 4478 3543 4530 3564
rect 4478 3512 4510 3543
rect 4510 3512 4530 3543
rect 6308 4408 6360 4416
rect 6308 4374 6314 4408
rect 6314 4374 6348 4408
rect 6348 4374 6360 4408
rect 6308 4364 6360 4374
rect 6580 4439 6632 4486
rect 6580 4434 6590 4439
rect 6590 4434 6624 4439
rect 6624 4434 6632 4439
rect 6216 4292 6268 4304
rect 6216 4258 6223 4292
rect 6223 4258 6257 4292
rect 6257 4258 6268 4292
rect 6216 4252 6268 4258
rect 7120 4410 7172 4418
rect 7120 4376 7127 4410
rect 7127 4376 7161 4410
rect 7161 4376 7172 4410
rect 7120 4366 7172 4376
rect 7032 4287 7084 4302
rect 7032 4253 7041 4287
rect 7041 4253 7075 4287
rect 7075 4253 7084 4287
rect 7032 4250 7084 4253
rect 6094 4017 6146 4069
rect 6270 4017 6322 4069
rect 6598 4002 6650 4014
rect 6598 3968 6606 4002
rect 6606 3968 6640 4002
rect 6640 3968 6650 4002
rect 6598 3962 6650 3968
rect 6096 3926 6148 3936
rect 6096 3892 6106 3926
rect 6106 3892 6140 3926
rect 6140 3892 6148 3926
rect 6096 3884 6148 3892
rect 5266 3669 5318 3672
rect 5266 3635 5299 3669
rect 5299 3635 5318 3669
rect 5266 3620 5318 3635
rect 6120 3661 6172 3678
rect 6120 3627 6141 3661
rect 6141 3627 6172 3661
rect 6120 3626 6172 3627
rect 6470 3809 6522 3820
rect 6470 3775 6478 3809
rect 6478 3775 6512 3809
rect 6512 3775 6522 3809
rect 6470 3768 6522 3775
rect 5028 3543 5080 3584
rect 5028 3532 5034 3543
rect 5034 3532 5068 3543
rect 5068 3532 5080 3543
rect 3723 3354 3775 3368
rect 3723 3320 3729 3354
rect 3729 3320 3763 3354
rect 3763 3320 3775 3354
rect 3723 3316 3775 3320
rect 4027 3320 4079 3372
rect 4690 3383 4742 3430
rect 4690 3378 4700 3383
rect 4700 3378 4734 3383
rect 4734 3378 4742 3383
rect 3140 3140 3192 3152
rect 3140 3106 3148 3140
rect 3148 3106 3182 3140
rect 3182 3106 3192 3140
rect 3140 3100 3192 3106
rect 4163 3117 4215 3130
rect 4163 3083 4195 3117
rect 4195 3083 4215 3117
rect 4163 3078 4215 3083
rect 4395 3112 4447 3120
rect 4395 3078 4404 3112
rect 4404 3078 4438 3112
rect 4438 3078 4447 3112
rect 4395 3068 4447 3078
rect 4708 2946 4760 2958
rect 4708 2912 4716 2946
rect 4716 2912 4750 2946
rect 4750 2912 4760 2946
rect 4708 2906 4760 2912
rect 6366 3543 6418 3564
rect 6366 3512 6398 3543
rect 6398 3512 6418 3543
rect 8196 4408 8248 4416
rect 8196 4374 8202 4408
rect 8202 4374 8236 4408
rect 8236 4374 8248 4408
rect 8196 4364 8248 4374
rect 8468 4439 8520 4486
rect 8468 4434 8478 4439
rect 8478 4434 8512 4439
rect 8512 4434 8520 4439
rect 8104 4292 8156 4304
rect 8104 4258 8111 4292
rect 8111 4258 8145 4292
rect 8145 4258 8156 4292
rect 8104 4252 8156 4258
rect 9008 4410 9060 4418
rect 9008 4376 9015 4410
rect 9015 4376 9049 4410
rect 9049 4376 9060 4410
rect 9008 4366 9060 4376
rect 8920 4287 8972 4302
rect 8920 4253 8929 4287
rect 8929 4253 8963 4287
rect 8963 4253 8972 4287
rect 8920 4250 8972 4253
rect 7982 4017 8034 4069
rect 8158 4017 8210 4069
rect 8486 4002 8538 4014
rect 8486 3968 8494 4002
rect 8494 3968 8528 4002
rect 8528 3968 8538 4002
rect 8486 3962 8538 3968
rect 7984 3926 8036 3936
rect 7984 3892 7994 3926
rect 7994 3892 8028 3926
rect 8028 3892 8036 3926
rect 7984 3884 8036 3892
rect 7154 3669 7206 3672
rect 7154 3635 7187 3669
rect 7187 3635 7206 3669
rect 7154 3620 7206 3635
rect 8008 3661 8060 3678
rect 8008 3627 8029 3661
rect 8029 3627 8060 3661
rect 8008 3626 8060 3627
rect 8358 3809 8410 3820
rect 8358 3775 8366 3809
rect 8366 3775 8400 3809
rect 8400 3775 8410 3809
rect 8358 3768 8410 3775
rect 6916 3543 6968 3584
rect 6916 3532 6922 3543
rect 6922 3532 6956 3543
rect 6956 3532 6968 3543
rect 5611 3354 5663 3368
rect 5611 3320 5617 3354
rect 5617 3320 5651 3354
rect 5651 3320 5663 3354
rect 5611 3316 5663 3320
rect 5915 3320 5967 3372
rect 6578 3383 6630 3430
rect 6578 3378 6588 3383
rect 6588 3378 6622 3383
rect 6622 3378 6630 3383
rect 5028 3140 5080 3152
rect 5028 3106 5036 3140
rect 5036 3106 5070 3140
rect 5070 3106 5080 3140
rect 5028 3100 5080 3106
rect 6051 3117 6103 3130
rect 6051 3083 6083 3117
rect 6083 3083 6103 3117
rect 6051 3078 6103 3083
rect 6283 3112 6335 3120
rect 6283 3078 6292 3112
rect 6292 3078 6326 3112
rect 6326 3078 6335 3112
rect 6283 3068 6335 3078
rect 6596 2946 6648 2958
rect 6596 2912 6604 2946
rect 6604 2912 6638 2946
rect 6638 2912 6648 2946
rect 6596 2906 6648 2912
rect 8254 3543 8306 3564
rect 8254 3512 8286 3543
rect 8286 3512 8306 3543
rect 10084 4408 10136 4416
rect 10084 4374 10090 4408
rect 10090 4374 10124 4408
rect 10124 4374 10136 4408
rect 10084 4364 10136 4374
rect 10356 4439 10408 4486
rect 10356 4434 10366 4439
rect 10366 4434 10400 4439
rect 10400 4434 10408 4439
rect 9992 4292 10044 4304
rect 9992 4258 9999 4292
rect 9999 4258 10033 4292
rect 10033 4258 10044 4292
rect 9992 4252 10044 4258
rect 10896 4410 10948 4418
rect 10896 4376 10903 4410
rect 10903 4376 10937 4410
rect 10937 4376 10948 4410
rect 10896 4366 10948 4376
rect 10808 4287 10860 4302
rect 10808 4253 10817 4287
rect 10817 4253 10851 4287
rect 10851 4253 10860 4287
rect 10808 4250 10860 4253
rect 9870 4017 9922 4069
rect 10046 4017 10098 4069
rect 10374 4002 10426 4014
rect 10374 3968 10382 4002
rect 10382 3968 10416 4002
rect 10416 3968 10426 4002
rect 10374 3962 10426 3968
rect 9872 3926 9924 3936
rect 9872 3892 9882 3926
rect 9882 3892 9916 3926
rect 9916 3892 9924 3926
rect 9872 3884 9924 3892
rect 9042 3669 9094 3672
rect 9042 3635 9075 3669
rect 9075 3635 9094 3669
rect 9042 3620 9094 3635
rect 9896 3661 9948 3678
rect 9896 3627 9917 3661
rect 9917 3627 9948 3661
rect 9896 3626 9948 3627
rect 10246 3809 10298 3820
rect 10246 3775 10254 3809
rect 10254 3775 10288 3809
rect 10288 3775 10298 3809
rect 10246 3768 10298 3775
rect 8804 3543 8856 3584
rect 8804 3532 8810 3543
rect 8810 3532 8844 3543
rect 8844 3532 8856 3543
rect 7499 3354 7551 3368
rect 7499 3320 7505 3354
rect 7505 3320 7539 3354
rect 7539 3320 7551 3354
rect 7499 3316 7551 3320
rect 7803 3320 7855 3372
rect 8466 3383 8518 3430
rect 8466 3378 8476 3383
rect 8476 3378 8510 3383
rect 8510 3378 8518 3383
rect 6916 3140 6968 3152
rect 6916 3106 6924 3140
rect 6924 3106 6958 3140
rect 6958 3106 6968 3140
rect 6916 3100 6968 3106
rect 7939 3117 7991 3130
rect 7939 3083 7971 3117
rect 7971 3083 7991 3117
rect 7939 3078 7991 3083
rect 8171 3112 8223 3120
rect 8171 3078 8180 3112
rect 8180 3078 8214 3112
rect 8214 3078 8223 3112
rect 8171 3068 8223 3078
rect 8484 2946 8536 2958
rect 8484 2912 8492 2946
rect 8492 2912 8526 2946
rect 8526 2912 8536 2946
rect 8484 2906 8536 2912
rect 10142 3543 10194 3564
rect 10142 3512 10174 3543
rect 10174 3512 10194 3543
rect 11966 4408 12018 4416
rect 11966 4374 11972 4408
rect 11972 4374 12006 4408
rect 12006 4374 12018 4408
rect 11966 4364 12018 4374
rect 12238 4439 12290 4486
rect 12238 4434 12248 4439
rect 12248 4434 12282 4439
rect 12282 4434 12290 4439
rect 11874 4292 11926 4304
rect 11874 4258 11881 4292
rect 11881 4258 11915 4292
rect 11915 4258 11926 4292
rect 11874 4252 11926 4258
rect 12778 4410 12830 4418
rect 12778 4376 12785 4410
rect 12785 4376 12819 4410
rect 12819 4376 12830 4410
rect 12778 4366 12830 4376
rect 12690 4287 12742 4302
rect 12690 4253 12699 4287
rect 12699 4253 12733 4287
rect 12733 4253 12742 4287
rect 12690 4250 12742 4253
rect 11752 4017 11804 4069
rect 11928 4017 11980 4069
rect 12256 4002 12308 4014
rect 12256 3968 12264 4002
rect 12264 3968 12298 4002
rect 12298 3968 12308 4002
rect 12256 3962 12308 3968
rect 11754 3926 11806 3936
rect 11754 3892 11764 3926
rect 11764 3892 11798 3926
rect 11798 3892 11806 3926
rect 11754 3884 11806 3892
rect 10930 3669 10982 3672
rect 10930 3635 10963 3669
rect 10963 3635 10982 3669
rect 10930 3620 10982 3635
rect 11778 3661 11830 3678
rect 11778 3627 11799 3661
rect 11799 3627 11830 3661
rect 11778 3626 11830 3627
rect 12128 3809 12180 3820
rect 12128 3775 12136 3809
rect 12136 3775 12170 3809
rect 12170 3775 12180 3809
rect 12128 3768 12180 3775
rect 10692 3543 10744 3584
rect 10692 3532 10698 3543
rect 10698 3532 10732 3543
rect 10732 3532 10744 3543
rect 9387 3354 9439 3368
rect 9387 3320 9393 3354
rect 9393 3320 9427 3354
rect 9427 3320 9439 3354
rect 9387 3316 9439 3320
rect 9691 3320 9743 3372
rect 10354 3383 10406 3430
rect 10354 3378 10364 3383
rect 10364 3378 10398 3383
rect 10398 3378 10406 3383
rect 8804 3140 8856 3152
rect 8804 3106 8812 3140
rect 8812 3106 8846 3140
rect 8846 3106 8856 3140
rect 8804 3100 8856 3106
rect 9827 3117 9879 3130
rect 9827 3083 9859 3117
rect 9859 3083 9879 3117
rect 9827 3078 9879 3083
rect 10059 3112 10111 3120
rect 10059 3078 10068 3112
rect 10068 3078 10102 3112
rect 10102 3078 10111 3112
rect 10059 3068 10111 3078
rect 10372 2946 10424 2958
rect 10372 2912 10380 2946
rect 10380 2912 10414 2946
rect 10414 2912 10424 2946
rect 10372 2906 10424 2912
rect 12024 3543 12076 3564
rect 12024 3512 12056 3543
rect 12056 3512 12076 3543
rect 13854 4408 13906 4416
rect 13854 4374 13860 4408
rect 13860 4374 13894 4408
rect 13894 4374 13906 4408
rect 13854 4364 13906 4374
rect 14126 4439 14178 4486
rect 14126 4434 14136 4439
rect 14136 4434 14170 4439
rect 14170 4434 14178 4439
rect 13762 4292 13814 4304
rect 13762 4258 13769 4292
rect 13769 4258 13803 4292
rect 13803 4258 13814 4292
rect 13762 4252 13814 4258
rect 14666 4410 14718 4418
rect 14666 4376 14673 4410
rect 14673 4376 14707 4410
rect 14707 4376 14718 4410
rect 14666 4366 14718 4376
rect 14578 4287 14630 4302
rect 14578 4253 14587 4287
rect 14587 4253 14621 4287
rect 14621 4253 14630 4287
rect 14578 4250 14630 4253
rect 13640 4017 13692 4069
rect 13816 4017 13868 4069
rect 14144 4002 14196 4014
rect 14144 3968 14152 4002
rect 14152 3968 14186 4002
rect 14186 3968 14196 4002
rect 14144 3962 14196 3968
rect 13642 3926 13694 3936
rect 13642 3892 13652 3926
rect 13652 3892 13686 3926
rect 13686 3892 13694 3926
rect 13642 3884 13694 3892
rect 12812 3669 12864 3672
rect 12812 3635 12845 3669
rect 12845 3635 12864 3669
rect 12812 3620 12864 3635
rect 13666 3661 13718 3678
rect 13666 3627 13687 3661
rect 13687 3627 13718 3661
rect 13666 3626 13718 3627
rect 14016 3809 14068 3820
rect 14016 3775 14024 3809
rect 14024 3775 14058 3809
rect 14058 3775 14068 3809
rect 14016 3768 14068 3775
rect 12574 3543 12626 3584
rect 12574 3532 12580 3543
rect 12580 3532 12614 3543
rect 12614 3532 12626 3543
rect 11275 3354 11327 3368
rect 11275 3320 11281 3354
rect 11281 3320 11315 3354
rect 11315 3320 11327 3354
rect 11275 3316 11327 3320
rect 11573 3320 11625 3372
rect 12236 3383 12288 3430
rect 12236 3378 12246 3383
rect 12246 3378 12280 3383
rect 12280 3378 12288 3383
rect 10692 3140 10744 3152
rect 10692 3106 10700 3140
rect 10700 3106 10734 3140
rect 10734 3106 10744 3140
rect 10692 3100 10744 3106
rect 11709 3117 11761 3130
rect 11709 3083 11741 3117
rect 11741 3083 11761 3117
rect 11709 3078 11761 3083
rect 11941 3112 11993 3120
rect 11941 3078 11950 3112
rect 11950 3078 11984 3112
rect 11984 3078 11993 3112
rect 11941 3068 11993 3078
rect 12254 2946 12306 2958
rect 12254 2912 12262 2946
rect 12262 2912 12296 2946
rect 12296 2912 12306 2946
rect 12254 2906 12306 2912
rect 13912 3543 13964 3564
rect 13912 3512 13944 3543
rect 13944 3512 13964 3543
rect 15742 4408 15794 4416
rect 15742 4374 15748 4408
rect 15748 4374 15782 4408
rect 15782 4374 15794 4408
rect 15742 4364 15794 4374
rect 16014 4439 16066 4486
rect 16014 4434 16024 4439
rect 16024 4434 16058 4439
rect 16058 4434 16066 4439
rect 15650 4292 15702 4304
rect 15650 4258 15657 4292
rect 15657 4258 15691 4292
rect 15691 4258 15702 4292
rect 15650 4252 15702 4258
rect 16554 4410 16606 4418
rect 16554 4376 16561 4410
rect 16561 4376 16595 4410
rect 16595 4376 16606 4410
rect 16554 4366 16606 4376
rect 16466 4287 16518 4302
rect 16466 4253 16475 4287
rect 16475 4253 16509 4287
rect 16509 4253 16518 4287
rect 16466 4250 16518 4253
rect 15528 4017 15580 4069
rect 15704 4017 15756 4069
rect 16032 4002 16084 4014
rect 16032 3968 16040 4002
rect 16040 3968 16074 4002
rect 16074 3968 16084 4002
rect 16032 3962 16084 3968
rect 15530 3926 15582 3936
rect 15530 3892 15540 3926
rect 15540 3892 15574 3926
rect 15574 3892 15582 3926
rect 15530 3884 15582 3892
rect 14700 3669 14752 3672
rect 14700 3635 14733 3669
rect 14733 3635 14752 3669
rect 14700 3620 14752 3635
rect 15554 3661 15606 3678
rect 15554 3627 15575 3661
rect 15575 3627 15606 3661
rect 15554 3626 15606 3627
rect 15904 3809 15956 3820
rect 15904 3775 15912 3809
rect 15912 3775 15946 3809
rect 15946 3775 15956 3809
rect 15904 3768 15956 3775
rect 14462 3543 14514 3584
rect 14462 3532 14468 3543
rect 14468 3532 14502 3543
rect 14502 3532 14514 3543
rect 13157 3354 13209 3368
rect 13157 3320 13163 3354
rect 13163 3320 13197 3354
rect 13197 3320 13209 3354
rect 13157 3316 13209 3320
rect 13461 3320 13513 3372
rect 14124 3383 14176 3430
rect 14124 3378 14134 3383
rect 14134 3378 14168 3383
rect 14168 3378 14176 3383
rect 12574 3140 12626 3152
rect 12574 3106 12582 3140
rect 12582 3106 12616 3140
rect 12616 3106 12626 3140
rect 12574 3100 12626 3106
rect 13597 3117 13649 3130
rect 13597 3083 13629 3117
rect 13629 3083 13649 3117
rect 13597 3078 13649 3083
rect 13829 3112 13881 3120
rect 13829 3078 13838 3112
rect 13838 3078 13872 3112
rect 13872 3078 13881 3112
rect 13829 3068 13881 3078
rect 14142 2946 14194 2958
rect 14142 2912 14150 2946
rect 14150 2912 14184 2946
rect 14184 2912 14194 2946
rect 14142 2906 14194 2912
rect 15800 3543 15852 3564
rect 15800 3512 15832 3543
rect 15832 3512 15852 3543
rect 17630 4408 17682 4416
rect 17630 4374 17636 4408
rect 17636 4374 17670 4408
rect 17670 4374 17682 4408
rect 17630 4364 17682 4374
rect 17902 4439 17954 4486
rect 17902 4434 17912 4439
rect 17912 4434 17946 4439
rect 17946 4434 17954 4439
rect 17538 4292 17590 4304
rect 17538 4258 17545 4292
rect 17545 4258 17579 4292
rect 17579 4258 17590 4292
rect 17538 4252 17590 4258
rect 18442 4410 18494 4418
rect 18442 4376 18449 4410
rect 18449 4376 18483 4410
rect 18483 4376 18494 4410
rect 18442 4366 18494 4376
rect 18354 4287 18406 4302
rect 18354 4253 18363 4287
rect 18363 4253 18397 4287
rect 18397 4253 18406 4287
rect 18354 4250 18406 4253
rect 17416 4017 17468 4069
rect 17592 4017 17644 4069
rect 17920 4002 17972 4014
rect 17920 3968 17928 4002
rect 17928 3968 17962 4002
rect 17962 3968 17972 4002
rect 17920 3962 17972 3968
rect 17418 3926 17470 3936
rect 17418 3892 17428 3926
rect 17428 3892 17462 3926
rect 17462 3892 17470 3926
rect 17418 3884 17470 3892
rect 16588 3669 16640 3672
rect 16588 3635 16621 3669
rect 16621 3635 16640 3669
rect 16588 3620 16640 3635
rect 17442 3661 17494 3678
rect 17442 3627 17463 3661
rect 17463 3627 17494 3661
rect 17442 3626 17494 3627
rect 17792 3809 17844 3820
rect 17792 3775 17800 3809
rect 17800 3775 17834 3809
rect 17834 3775 17844 3809
rect 17792 3768 17844 3775
rect 16350 3543 16402 3584
rect 16350 3532 16356 3543
rect 16356 3532 16390 3543
rect 16390 3532 16402 3543
rect 15045 3354 15097 3368
rect 15045 3320 15051 3354
rect 15051 3320 15085 3354
rect 15085 3320 15097 3354
rect 15045 3316 15097 3320
rect 15349 3320 15401 3372
rect 16012 3383 16064 3430
rect 16012 3378 16022 3383
rect 16022 3378 16056 3383
rect 16056 3378 16064 3383
rect 14462 3140 14514 3152
rect 14462 3106 14470 3140
rect 14470 3106 14504 3140
rect 14504 3106 14514 3140
rect 14462 3100 14514 3106
rect 15485 3117 15537 3130
rect 15485 3083 15517 3117
rect 15517 3083 15537 3117
rect 15485 3078 15537 3083
rect 15717 3112 15769 3120
rect 15717 3078 15726 3112
rect 15726 3078 15760 3112
rect 15760 3078 15769 3112
rect 15717 3068 15769 3078
rect 16030 2946 16082 2958
rect 16030 2912 16038 2946
rect 16038 2912 16072 2946
rect 16072 2912 16082 2946
rect 16030 2906 16082 2912
rect 17688 3543 17740 3564
rect 17688 3512 17720 3543
rect 17720 3512 17740 3543
rect 19518 4408 19570 4416
rect 19518 4374 19524 4408
rect 19524 4374 19558 4408
rect 19558 4374 19570 4408
rect 19518 4364 19570 4374
rect 19790 4439 19842 4486
rect 19790 4434 19800 4439
rect 19800 4434 19834 4439
rect 19834 4434 19842 4439
rect 19426 4292 19478 4304
rect 19426 4258 19433 4292
rect 19433 4258 19467 4292
rect 19467 4258 19478 4292
rect 19426 4252 19478 4258
rect 20330 4410 20382 4418
rect 20330 4376 20337 4410
rect 20337 4376 20371 4410
rect 20371 4376 20382 4410
rect 20330 4366 20382 4376
rect 20242 4287 20294 4302
rect 20242 4253 20251 4287
rect 20251 4253 20285 4287
rect 20285 4253 20294 4287
rect 20242 4250 20294 4253
rect 19304 4017 19356 4069
rect 19480 4017 19532 4069
rect 19808 4002 19860 4014
rect 19808 3968 19816 4002
rect 19816 3968 19850 4002
rect 19850 3968 19860 4002
rect 19808 3962 19860 3968
rect 19306 3926 19358 3936
rect 19306 3892 19316 3926
rect 19316 3892 19350 3926
rect 19350 3892 19358 3926
rect 19306 3884 19358 3892
rect 18476 3669 18528 3672
rect 18476 3635 18509 3669
rect 18509 3635 18528 3669
rect 18476 3620 18528 3635
rect 19330 3661 19382 3678
rect 19330 3627 19351 3661
rect 19351 3627 19382 3661
rect 19330 3626 19382 3627
rect 19680 3809 19732 3820
rect 19680 3775 19688 3809
rect 19688 3775 19722 3809
rect 19722 3775 19732 3809
rect 19680 3768 19732 3775
rect 18238 3543 18290 3584
rect 18238 3532 18244 3543
rect 18244 3532 18278 3543
rect 18278 3532 18290 3543
rect 16933 3354 16985 3368
rect 16933 3320 16939 3354
rect 16939 3320 16973 3354
rect 16973 3320 16985 3354
rect 16933 3316 16985 3320
rect 17237 3320 17289 3372
rect 17900 3383 17952 3430
rect 17900 3378 17910 3383
rect 17910 3378 17944 3383
rect 17944 3378 17952 3383
rect 16350 3140 16402 3152
rect 16350 3106 16358 3140
rect 16358 3106 16392 3140
rect 16392 3106 16402 3140
rect 16350 3100 16402 3106
rect 17373 3117 17425 3130
rect 17373 3083 17405 3117
rect 17405 3083 17425 3117
rect 17373 3078 17425 3083
rect 17605 3112 17657 3120
rect 17605 3078 17614 3112
rect 17614 3078 17648 3112
rect 17648 3078 17657 3112
rect 17605 3068 17657 3078
rect 17918 2946 17970 2958
rect 17918 2912 17926 2946
rect 17926 2912 17960 2946
rect 17960 2912 17970 2946
rect 17918 2906 17970 2912
rect 19576 3543 19628 3564
rect 19576 3512 19608 3543
rect 19608 3512 19628 3543
rect 21406 4408 21458 4416
rect 21406 4374 21412 4408
rect 21412 4374 21446 4408
rect 21446 4374 21458 4408
rect 21406 4364 21458 4374
rect 21678 4439 21730 4486
rect 21678 4434 21688 4439
rect 21688 4434 21722 4439
rect 21722 4434 21730 4439
rect 21314 4292 21366 4304
rect 21314 4258 21321 4292
rect 21321 4258 21355 4292
rect 21355 4258 21366 4292
rect 21314 4252 21366 4258
rect 22218 4410 22270 4418
rect 22218 4376 22225 4410
rect 22225 4376 22259 4410
rect 22259 4376 22270 4410
rect 22218 4366 22270 4376
rect 22130 4287 22182 4302
rect 22130 4253 22139 4287
rect 22139 4253 22173 4287
rect 22173 4253 22182 4287
rect 22130 4250 22182 4253
rect 21192 4017 21244 4069
rect 21368 4017 21420 4069
rect 21696 4002 21748 4014
rect 21696 3968 21704 4002
rect 21704 3968 21738 4002
rect 21738 3968 21748 4002
rect 21696 3962 21748 3968
rect 21194 3926 21246 3936
rect 21194 3892 21204 3926
rect 21204 3892 21238 3926
rect 21238 3892 21246 3926
rect 21194 3884 21246 3892
rect 20364 3669 20416 3672
rect 20364 3635 20397 3669
rect 20397 3635 20416 3669
rect 20364 3620 20416 3635
rect 21218 3661 21270 3678
rect 21218 3627 21239 3661
rect 21239 3627 21270 3661
rect 21218 3626 21270 3627
rect 21568 3809 21620 3820
rect 21568 3775 21576 3809
rect 21576 3775 21610 3809
rect 21610 3775 21620 3809
rect 21568 3768 21620 3775
rect 20126 3543 20178 3584
rect 20126 3532 20132 3543
rect 20132 3532 20166 3543
rect 20166 3532 20178 3543
rect 18821 3354 18873 3368
rect 18821 3320 18827 3354
rect 18827 3320 18861 3354
rect 18861 3320 18873 3354
rect 18821 3316 18873 3320
rect 19125 3320 19177 3372
rect 19788 3383 19840 3430
rect 19788 3378 19798 3383
rect 19798 3378 19832 3383
rect 19832 3378 19840 3383
rect 18238 3140 18290 3152
rect 18238 3106 18246 3140
rect 18246 3106 18280 3140
rect 18280 3106 18290 3140
rect 18238 3100 18290 3106
rect 19261 3117 19313 3130
rect 19261 3083 19293 3117
rect 19293 3083 19313 3117
rect 19261 3078 19313 3083
rect 19493 3112 19545 3120
rect 19493 3078 19502 3112
rect 19502 3078 19536 3112
rect 19536 3078 19545 3112
rect 19493 3068 19545 3078
rect 19806 2946 19858 2958
rect 19806 2912 19814 2946
rect 19814 2912 19848 2946
rect 19848 2912 19858 2946
rect 19806 2906 19858 2912
rect 21464 3543 21516 3564
rect 21464 3512 21496 3543
rect 21496 3512 21516 3543
rect 23294 4408 23346 4416
rect 23294 4374 23300 4408
rect 23300 4374 23334 4408
rect 23334 4374 23346 4408
rect 23294 4364 23346 4374
rect 23566 4439 23618 4486
rect 23566 4434 23576 4439
rect 23576 4434 23610 4439
rect 23610 4434 23618 4439
rect 23202 4292 23254 4304
rect 23202 4258 23209 4292
rect 23209 4258 23243 4292
rect 23243 4258 23254 4292
rect 23202 4252 23254 4258
rect 24106 4410 24158 4418
rect 24106 4376 24113 4410
rect 24113 4376 24147 4410
rect 24147 4376 24158 4410
rect 24106 4366 24158 4376
rect 24018 4287 24070 4302
rect 24018 4253 24027 4287
rect 24027 4253 24061 4287
rect 24061 4253 24070 4287
rect 24018 4250 24070 4253
rect 23080 4017 23132 4069
rect 23256 4017 23308 4069
rect 23584 4002 23636 4014
rect 23584 3968 23592 4002
rect 23592 3968 23626 4002
rect 23626 3968 23636 4002
rect 23584 3962 23636 3968
rect 23082 3926 23134 3936
rect 23082 3892 23092 3926
rect 23092 3892 23126 3926
rect 23126 3892 23134 3926
rect 23082 3884 23134 3892
rect 22252 3669 22304 3672
rect 22252 3635 22285 3669
rect 22285 3635 22304 3669
rect 22252 3620 22304 3635
rect 23106 3661 23158 3678
rect 23106 3627 23127 3661
rect 23127 3627 23158 3661
rect 23106 3626 23158 3627
rect 23456 3809 23508 3820
rect 23456 3775 23464 3809
rect 23464 3775 23498 3809
rect 23498 3775 23508 3809
rect 23456 3768 23508 3775
rect 22014 3543 22066 3584
rect 22014 3532 22020 3543
rect 22020 3532 22054 3543
rect 22054 3532 22066 3543
rect 20709 3354 20761 3368
rect 20709 3320 20715 3354
rect 20715 3320 20749 3354
rect 20749 3320 20761 3354
rect 20709 3316 20761 3320
rect 21013 3320 21065 3372
rect 21676 3383 21728 3430
rect 21676 3378 21686 3383
rect 21686 3378 21720 3383
rect 21720 3378 21728 3383
rect 20126 3140 20178 3152
rect 20126 3106 20134 3140
rect 20134 3106 20168 3140
rect 20168 3106 20178 3140
rect 20126 3100 20178 3106
rect 21149 3117 21201 3130
rect 21149 3083 21181 3117
rect 21181 3083 21201 3117
rect 21149 3078 21201 3083
rect 21381 3112 21433 3120
rect 21381 3078 21390 3112
rect 21390 3078 21424 3112
rect 21424 3078 21433 3112
rect 21381 3068 21433 3078
rect 21694 2946 21746 2958
rect 21694 2912 21702 2946
rect 21702 2912 21736 2946
rect 21736 2912 21746 2946
rect 21694 2906 21746 2912
rect 23352 3543 23404 3564
rect 23352 3512 23384 3543
rect 23384 3512 23404 3543
rect 25182 4408 25234 4416
rect 25182 4374 25188 4408
rect 25188 4374 25222 4408
rect 25222 4374 25234 4408
rect 25182 4364 25234 4374
rect 25454 4439 25506 4486
rect 25454 4434 25464 4439
rect 25464 4434 25498 4439
rect 25498 4434 25506 4439
rect 25090 4292 25142 4304
rect 25090 4258 25097 4292
rect 25097 4258 25131 4292
rect 25131 4258 25142 4292
rect 25090 4252 25142 4258
rect 25994 4410 26046 4418
rect 25994 4376 26001 4410
rect 26001 4376 26035 4410
rect 26035 4376 26046 4410
rect 25994 4366 26046 4376
rect 25906 4287 25958 4302
rect 25906 4253 25915 4287
rect 25915 4253 25949 4287
rect 25949 4253 25958 4287
rect 25906 4250 25958 4253
rect 24968 4017 25020 4069
rect 25144 4017 25196 4069
rect 25472 4002 25524 4014
rect 25472 3968 25480 4002
rect 25480 3968 25514 4002
rect 25514 3968 25524 4002
rect 25472 3962 25524 3968
rect 24970 3926 25022 3936
rect 24970 3892 24980 3926
rect 24980 3892 25014 3926
rect 25014 3892 25022 3926
rect 24970 3884 25022 3892
rect 24140 3669 24192 3672
rect 24140 3635 24173 3669
rect 24173 3635 24192 3669
rect 24140 3620 24192 3635
rect 24994 3661 25046 3678
rect 24994 3627 25015 3661
rect 25015 3627 25046 3661
rect 24994 3626 25046 3627
rect 25344 3809 25396 3820
rect 25344 3775 25352 3809
rect 25352 3775 25386 3809
rect 25386 3775 25396 3809
rect 25344 3768 25396 3775
rect 23902 3543 23954 3584
rect 23902 3532 23908 3543
rect 23908 3532 23942 3543
rect 23942 3532 23954 3543
rect 22597 3354 22649 3368
rect 22597 3320 22603 3354
rect 22603 3320 22637 3354
rect 22637 3320 22649 3354
rect 22597 3316 22649 3320
rect 22901 3320 22953 3372
rect 23564 3383 23616 3430
rect 23564 3378 23574 3383
rect 23574 3378 23608 3383
rect 23608 3378 23616 3383
rect 22014 3140 22066 3152
rect 22014 3106 22022 3140
rect 22022 3106 22056 3140
rect 22056 3106 22066 3140
rect 22014 3100 22066 3106
rect 23037 3117 23089 3130
rect 23037 3083 23069 3117
rect 23069 3083 23089 3117
rect 23037 3078 23089 3083
rect 23269 3112 23321 3120
rect 23269 3078 23278 3112
rect 23278 3078 23312 3112
rect 23312 3078 23321 3112
rect 23269 3068 23321 3078
rect 23582 2946 23634 2958
rect 23582 2912 23590 2946
rect 23590 2912 23624 2946
rect 23624 2912 23634 2946
rect 23582 2906 23634 2912
rect 25240 3543 25292 3564
rect 25240 3512 25272 3543
rect 25272 3512 25292 3543
rect 26028 3669 26080 3672
rect 26028 3635 26061 3669
rect 26061 3635 26080 3669
rect 26028 3620 26080 3635
rect 25790 3543 25842 3584
rect 25790 3532 25796 3543
rect 25796 3532 25830 3543
rect 25830 3532 25842 3543
rect 24485 3354 24537 3368
rect 24485 3320 24491 3354
rect 24491 3320 24525 3354
rect 24525 3320 24537 3354
rect 24485 3316 24537 3320
rect 24789 3320 24841 3372
rect 25452 3383 25504 3430
rect 25452 3378 25462 3383
rect 25462 3378 25496 3383
rect 25496 3378 25504 3383
rect 23902 3140 23954 3152
rect 23902 3106 23910 3140
rect 23910 3106 23944 3140
rect 23944 3106 23954 3140
rect 23902 3100 23954 3106
rect 24925 3117 24977 3130
rect 24925 3083 24957 3117
rect 24957 3083 24977 3117
rect 24925 3078 24977 3083
rect 25157 3112 25209 3120
rect 25157 3078 25166 3112
rect 25166 3078 25200 3112
rect 25200 3078 25209 3112
rect 25157 3068 25209 3078
rect 25470 2946 25522 2958
rect 25470 2912 25478 2946
rect 25478 2912 25512 2946
rect 25512 2912 25522 2946
rect 25470 2906 25522 2912
rect 26373 3354 26425 3368
rect 26373 3320 26379 3354
rect 26379 3320 26413 3354
rect 26413 3320 26425 3354
rect 26373 3316 26425 3320
rect 25790 3140 25842 3152
rect 25790 3106 25798 3140
rect 25798 3106 25832 3140
rect 25832 3106 25842 3140
rect 25790 3100 25842 3106
rect -2017 2592 -1709 2708
rect -129 2592 179 2708
rect 1759 2592 2067 2708
rect 3647 2592 3955 2708
rect 5535 2592 5843 2708
rect 7423 2592 7731 2708
rect 9311 2592 9619 2708
rect 11199 2592 11507 2708
rect 13081 2592 13389 2708
rect 14969 2592 15277 2708
rect 16857 2592 17165 2708
rect 18745 2592 19053 2708
rect 20633 2592 20941 2708
rect 22521 2592 22829 2708
rect 24409 2592 24717 2708
rect 26297 2592 26605 2708
<< metal2 >>
rect 4475 5343 4844 5373
rect 4475 5290 4610 5343
rect 4683 5290 4844 5343
rect 4475 5272 4844 5290
rect 19621 5349 19892 5371
rect 19621 5343 19740 5349
rect 19621 5289 19704 5343
rect 19807 5296 19892 5349
rect 19780 5289 19892 5296
rect 19621 5271 19892 5289
rect -1439 5082 -413 5083
rect 446 5082 1472 5084
rect 13643 5082 14669 5084
rect 15544 5082 16570 5083
rect 21211 5082 22237 5086
rect 23115 5082 24141 5083
rect -3546 5020 11208 5082
rect 11562 5020 26308 5082
rect -3544 5004 11208 5020
rect -3544 5002 2740 5004
rect -3544 4950 2282 5002
rect 2334 4950 2389 5002
rect 2441 4950 2495 5002
rect 2547 4950 2611 5002
rect 2663 4952 2740 5002
rect 2792 5003 11208 5004
rect 2792 4952 2874 5003
rect 2663 4951 2874 4952
rect 2926 4951 2991 5003
rect 3043 4951 3096 5003
rect 3148 4951 3202 5003
rect 3254 4951 3299 5003
rect 3351 4951 3396 5003
rect 3448 5002 11208 5003
rect 3448 4999 4622 5002
rect 4674 5001 11208 5002
rect 3448 4951 4171 4999
rect 2663 4950 4171 4951
rect -3544 4947 4171 4950
rect 4223 4947 4278 4999
rect 4330 4947 4384 4999
rect 4436 4947 4500 4999
rect 4552 4950 4622 4999
rect 4681 5000 11208 5001
rect 4552 4949 4629 4950
rect 4681 4949 4763 5000
rect 4552 4948 4763 4949
rect 4815 4948 4880 5000
rect 4932 4948 4985 5000
rect 5037 4948 5091 5000
rect 5143 4948 5188 5000
rect 5240 4948 5285 5000
rect 5337 4948 11208 5000
rect 11563 5008 26308 5020
rect 11563 4956 17391 5008
rect 17443 5006 26308 5008
rect 17443 4956 17503 5006
rect 4552 4947 11208 4948
rect -3544 4894 11208 4947
rect 11562 4954 17503 4956
rect 17555 4954 17610 5006
rect 17662 4954 17712 5006
rect 17764 5004 26308 5006
rect 17764 4954 17838 5004
rect 11562 4952 17838 4954
rect 17890 4952 17992 5004
rect 18044 4952 18129 5004
rect 18181 4952 18226 5004
rect 18278 4952 18326 5004
rect 18378 5003 26308 5004
rect 18378 4952 18415 5003
rect 11562 4951 18415 4952
rect 18467 4951 18511 5003
rect 18563 5002 26308 5003
rect 18563 4951 19225 5002
rect 11562 4950 19225 4951
rect 19277 4950 19319 5002
rect 19371 4950 19418 5002
rect 19470 4950 19526 5002
rect 19578 4950 19622 5002
rect 19674 4950 19720 5002
rect 19772 5001 26308 5002
rect 19772 4950 19839 5001
rect 11562 4949 19839 4950
rect 19891 4949 19953 5001
rect 20005 4949 20070 5001
rect 20122 4949 20197 5001
rect 20249 4949 20312 5001
rect 20364 4949 26308 5001
rect 11562 4894 26308 4949
rect -3326 4637 -2300 4894
rect -2038 4832 -1688 4846
rect -2038 4716 -2017 4832
rect -1709 4716 -1688 4832
rect -2038 4702 -1688 4716
rect -1439 4637 -413 4894
rect -150 4832 200 4846
rect -150 4716 -129 4832
rect 179 4716 200 4832
rect -150 4702 200 4716
rect 446 4637 1472 4894
rect 2150 4886 5358 4894
rect 1738 4832 2088 4846
rect 1738 4716 1759 4832
rect 2067 4716 2088 4832
rect 1738 4702 2088 4716
rect 2150 4637 3470 4886
rect 3626 4832 3976 4846
rect 3626 4716 3647 4832
rect 3955 4716 3976 4832
rect 3626 4702 3976 4716
rect -3544 4590 3470 4637
rect 4034 4633 5358 4886
rect 5514 4832 5864 4846
rect 5514 4716 5535 4832
rect 5843 4716 5864 4832
rect 5514 4702 5864 4716
rect 6115 4633 7141 4894
rect 7402 4832 7752 4846
rect 7402 4716 7423 4832
rect 7731 4716 7752 4832
rect 7402 4702 7752 4716
rect 8010 4633 9036 4894
rect 9290 4832 9640 4846
rect 9290 4716 9311 4832
rect 9619 4716 9640 4832
rect 9290 4702 9640 4716
rect 9879 4633 10905 4894
rect 11178 4832 11528 4846
rect 11178 4716 11199 4832
rect 11507 4716 11528 4832
rect 11178 4702 11528 4716
rect 11756 4637 12782 4894
rect 13060 4832 13410 4846
rect 13060 4716 13081 4832
rect 13389 4716 13410 4832
rect 13060 4702 13410 4716
rect 13643 4637 14669 4894
rect 14948 4832 15298 4846
rect 14948 4716 14969 4832
rect 15277 4716 15298 4832
rect 14948 4702 15298 4716
rect 15544 4637 16570 4894
rect 17248 4886 20456 4894
rect 16836 4832 17186 4846
rect 16836 4716 16857 4832
rect 17165 4716 17186 4832
rect 16836 4702 17186 4716
rect 17248 4637 18568 4886
rect 18724 4832 19074 4846
rect 18724 4716 18745 4832
rect 19053 4716 19074 4832
rect 18724 4702 19074 4716
rect 19132 4637 20456 4886
rect 20612 4832 20962 4846
rect 20612 4716 20633 4832
rect 20941 4716 20962 4832
rect 20612 4702 20962 4716
rect 21211 4637 22237 4894
rect 22500 4832 22850 4846
rect 22500 4716 22521 4832
rect 22829 4716 22850 4832
rect 22500 4702 22850 4716
rect 23115 4637 24141 4894
rect 24388 4832 24738 4846
rect 24388 4716 24409 4832
rect 24717 4716 24738 4832
rect 24388 4702 24738 4716
rect 24991 4637 26017 4894
rect 26276 4832 26626 4846
rect 26276 4716 26297 4832
rect 26605 4716 26626 4832
rect 26276 4702 26626 4716
rect 4034 4590 11208 4633
rect -3544 4528 11208 4590
rect 11562 4590 26307 4637
rect 11562 4556 26306 4590
rect 11554 4528 26306 4556
rect -3102 4422 -3074 4528
rect -2866 4486 -2800 4494
rect -2866 4434 -2860 4486
rect -2808 4434 -2800 4486
rect -2866 4426 -2800 4434
rect -3142 4416 -3074 4422
rect -3142 4364 -3132 4416
rect -3080 4364 -3074 4416
rect -3142 4358 -3074 4364
rect -3232 4304 -3164 4310
rect -3232 4252 -3224 4304
rect -3172 4252 -3164 4304
rect -3232 4242 -3164 4252
rect -3352 4069 -3288 4076
rect -3352 4038 -3346 4069
rect -3544 4017 -3346 4038
rect -3294 4017 -3288 4069
rect -3544 4010 -3288 4017
rect -3544 4008 -3346 4010
rect -3544 4002 -3352 4008
rect -3352 3936 -3286 3942
rect -3352 3884 -3344 3936
rect -3292 3884 -3286 3936
rect -3352 3878 -3286 3884
rect -3352 3756 -3324 3878
rect -3392 3728 -3324 3756
rect -3532 3372 -3464 3378
rect -3532 3320 -3525 3372
rect -3473 3320 -3464 3372
rect -3532 3314 -3464 3320
rect -3532 2698 -3488 3314
rect -3392 3144 -3364 3728
rect -3330 3678 -3268 3684
rect -3330 3626 -3320 3678
rect -3232 3670 -3204 4242
rect -3176 4069 -3112 4076
rect -3176 4017 -3170 4069
rect -3118 4036 -3112 4069
rect -2850 4036 -2800 4426
rect -2328 4424 -2300 4528
rect -2328 4418 -2262 4424
rect -1214 4422 -1186 4528
rect -978 4486 -912 4494
rect -978 4434 -972 4486
rect -920 4434 -912 4486
rect -978 4426 -912 4434
rect -2328 4404 -2320 4418
rect -2326 4366 -2320 4404
rect -2268 4366 -2262 4418
rect -2326 4360 -2262 4366
rect -1254 4416 -1186 4422
rect -1254 4364 -1244 4416
rect -1192 4364 -1186 4416
rect -1254 4358 -1186 4364
rect -2414 4302 -2350 4308
rect -2414 4272 -2408 4302
rect -2624 4250 -2408 4272
rect -2356 4250 -2350 4302
rect -2624 4244 -2350 4250
rect -1344 4304 -1276 4310
rect -1344 4252 -1336 4304
rect -1284 4252 -1276 4304
rect -3118 4020 -2798 4036
rect -3118 4017 -2784 4020
rect -3176 4014 -2784 4017
rect -3176 4008 -2842 4014
rect -2850 3962 -2842 4008
rect -2790 3962 -2784 4014
rect -2850 3956 -2784 3962
rect -2980 3820 -2908 3832
rect -2980 3768 -2970 3820
rect -2918 3768 -2908 3820
rect -2980 3756 -2908 3768
rect -2944 3754 -2908 3756
rect -3232 3642 -2944 3670
rect -3330 3620 -3268 3626
rect -3296 3574 -3268 3620
rect -3296 3570 -3052 3574
rect -3296 3564 -3014 3570
rect -3296 3546 -3074 3564
rect -3080 3512 -3074 3546
rect -3022 3512 -3014 3564
rect -3080 3504 -3014 3512
rect -3392 3130 -3328 3144
rect -2972 3136 -2944 3642
rect -2868 3430 -2802 3438
rect -2868 3378 -2862 3430
rect -2810 3378 -2802 3430
rect -2868 3370 -2802 3378
rect -3392 3078 -3389 3130
rect -3337 3078 -3328 3130
rect -3392 3062 -3328 3078
rect -3158 3120 -2944 3136
rect -3158 3068 -3157 3120
rect -3105 3108 -2944 3120
rect -3105 3068 -3104 3108
rect -3158 3052 -3104 3068
rect -2852 2964 -2802 3370
rect -2624 3126 -2596 4244
rect -1344 4242 -1276 4252
rect -1464 4069 -1400 4076
rect -1464 4038 -1458 4069
rect -2192 4017 -1458 4038
rect -1406 4017 -1400 4069
rect -2192 4010 -1400 4017
rect -2192 4008 -1458 4010
rect -2192 4002 -1464 4008
rect -2292 3672 -2228 3680
rect -2292 3620 -2286 3672
rect -2234 3620 -2228 3672
rect -2292 3612 -2228 3620
rect -2532 3584 -2466 3590
rect -2532 3532 -2524 3584
rect -2472 3554 -2466 3584
rect -2292 3554 -2264 3612
rect -2472 3532 -2264 3554
rect -2532 3526 -2264 3532
rect -2192 3376 -2164 4002
rect -1464 3936 -1398 3942
rect -1464 3884 -1456 3936
rect -1404 3884 -1398 3936
rect -1464 3878 -1398 3884
rect -1464 3756 -1436 3878
rect -1504 3728 -1436 3756
rect -2192 3368 -1880 3376
rect -2192 3340 -1941 3368
rect -2532 3152 -2456 3158
rect -2532 3126 -2524 3152
rect -2624 3100 -2524 3126
rect -2472 3100 -2456 3152
rect -2624 3098 -2456 3100
rect -2532 3094 -2456 3098
rect -2852 2958 -2786 2964
rect -2852 2906 -2844 2958
rect -2792 2936 -2786 2958
rect -2192 2936 -2164 3340
rect -1960 3316 -1941 3340
rect -1889 3316 -1880 3368
rect -1960 3304 -1880 3316
rect -1644 3372 -1576 3378
rect -1644 3320 -1637 3372
rect -1585 3320 -1576 3372
rect -1644 3314 -1576 3320
rect -2792 2908 -2164 2936
rect -2792 2906 -2786 2908
rect -2852 2900 -2786 2906
rect -2038 2708 -1688 2722
rect -2038 2592 -2017 2708
rect -1709 2592 -1688 2708
rect -1644 2698 -1600 3314
rect -1504 3144 -1476 3728
rect -1442 3678 -1380 3684
rect -1442 3626 -1432 3678
rect -1344 3670 -1316 4242
rect -1288 4069 -1224 4076
rect -1288 4017 -1282 4069
rect -1230 4036 -1224 4069
rect -962 4036 -912 4426
rect -440 4424 -412 4528
rect -440 4418 -374 4424
rect 674 4422 702 4528
rect 910 4486 976 4494
rect 910 4434 916 4486
rect 968 4434 976 4486
rect 910 4426 976 4434
rect -440 4404 -432 4418
rect -438 4366 -432 4404
rect -380 4366 -374 4418
rect -438 4360 -374 4366
rect 634 4416 702 4422
rect 634 4364 644 4416
rect 696 4364 702 4416
rect 634 4358 702 4364
rect -526 4302 -462 4308
rect -526 4272 -520 4302
rect -736 4250 -520 4272
rect -468 4250 -462 4302
rect -736 4244 -462 4250
rect 544 4304 612 4310
rect 544 4252 552 4304
rect 604 4252 612 4304
rect -1230 4020 -910 4036
rect -1230 4017 -896 4020
rect -1288 4014 -896 4017
rect -1288 4008 -954 4014
rect -962 3962 -954 4008
rect -902 3962 -896 4014
rect -962 3956 -896 3962
rect -1092 3820 -1020 3832
rect -1092 3768 -1082 3820
rect -1030 3768 -1020 3820
rect -1092 3756 -1020 3768
rect -1056 3754 -1020 3756
rect -1344 3642 -1056 3670
rect -1442 3620 -1380 3626
rect -1408 3574 -1380 3620
rect -1408 3570 -1164 3574
rect -1408 3564 -1126 3570
rect -1408 3546 -1186 3564
rect -1192 3512 -1186 3546
rect -1134 3512 -1126 3564
rect -1192 3504 -1126 3512
rect -1504 3130 -1440 3144
rect -1084 3136 -1056 3642
rect -980 3430 -914 3438
rect -980 3378 -974 3430
rect -922 3378 -914 3430
rect -980 3370 -914 3378
rect -1504 3078 -1501 3130
rect -1449 3078 -1440 3130
rect -1504 3062 -1440 3078
rect -1270 3120 -1056 3136
rect -1270 3068 -1269 3120
rect -1217 3108 -1056 3120
rect -1217 3068 -1216 3108
rect -1270 3052 -1216 3068
rect -964 2964 -914 3370
rect -736 3126 -708 4244
rect 544 4242 612 4252
rect 424 4069 488 4076
rect 424 4038 430 4069
rect -304 4017 430 4038
rect 482 4017 488 4069
rect -304 4010 488 4017
rect -304 4008 430 4010
rect -304 4002 424 4008
rect -404 3672 -340 3680
rect -404 3620 -398 3672
rect -346 3620 -340 3672
rect -404 3612 -340 3620
rect -644 3584 -578 3590
rect -644 3532 -636 3584
rect -584 3554 -578 3584
rect -404 3554 -376 3612
rect -584 3532 -376 3554
rect -644 3526 -376 3532
rect -304 3376 -276 4002
rect 424 3936 490 3942
rect 424 3884 432 3936
rect 484 3884 490 3936
rect 424 3878 490 3884
rect 424 3756 452 3878
rect 384 3728 452 3756
rect -304 3368 8 3376
rect -304 3340 -53 3368
rect -644 3152 -568 3158
rect -644 3126 -636 3152
rect -736 3100 -636 3126
rect -584 3100 -568 3152
rect -736 3098 -568 3100
rect -644 3094 -568 3098
rect -964 2958 -898 2964
rect -964 2906 -956 2958
rect -904 2936 -898 2958
rect -304 2936 -276 3340
rect -72 3316 -53 3340
rect -1 3316 8 3368
rect -72 3304 8 3316
rect 244 3372 312 3378
rect 244 3320 251 3372
rect 303 3320 312 3372
rect 244 3314 312 3320
rect -904 2908 -276 2936
rect -904 2906 -898 2908
rect -964 2900 -898 2906
rect -150 2708 200 2722
rect -2038 2578 -1688 2592
rect -150 2592 -129 2708
rect 179 2592 200 2708
rect 244 2698 288 3314
rect 384 3144 412 3728
rect 446 3678 508 3684
rect 446 3626 456 3678
rect 544 3670 572 4242
rect 600 4069 664 4076
rect 600 4017 606 4069
rect 658 4036 664 4069
rect 926 4036 976 4426
rect 1448 4424 1476 4528
rect 2150 4524 3470 4528
rect 4034 4524 11208 4528
rect 1448 4418 1514 4424
rect 2562 4422 2590 4524
rect 2798 4486 2864 4494
rect 2798 4434 2804 4486
rect 2856 4434 2864 4486
rect 2798 4426 2864 4434
rect 1448 4404 1456 4418
rect 1450 4366 1456 4404
rect 1508 4366 1514 4418
rect 1450 4360 1514 4366
rect 2522 4416 2590 4422
rect 2522 4364 2532 4416
rect 2584 4364 2590 4416
rect 2522 4358 2590 4364
rect 1362 4302 1426 4308
rect 1362 4272 1368 4302
rect 1152 4250 1368 4272
rect 1420 4250 1426 4302
rect 1152 4244 1426 4250
rect 2432 4304 2500 4310
rect 2432 4252 2440 4304
rect 2492 4252 2500 4304
rect 658 4020 978 4036
rect 658 4017 992 4020
rect 600 4014 992 4017
rect 600 4008 934 4014
rect 926 3962 934 4008
rect 986 3962 992 4014
rect 926 3956 992 3962
rect 796 3820 868 3832
rect 796 3768 806 3820
rect 858 3768 868 3820
rect 796 3756 868 3768
rect 832 3754 868 3756
rect 544 3642 832 3670
rect 446 3620 508 3626
rect 480 3574 508 3620
rect 480 3570 724 3574
rect 480 3564 762 3570
rect 480 3546 702 3564
rect 696 3512 702 3546
rect 754 3512 762 3564
rect 696 3504 762 3512
rect 384 3130 448 3144
rect 804 3136 832 3642
rect 908 3430 974 3438
rect 908 3378 914 3430
rect 966 3378 974 3430
rect 908 3370 974 3378
rect 384 3078 387 3130
rect 439 3078 448 3130
rect 384 3062 448 3078
rect 618 3120 832 3136
rect 618 3068 619 3120
rect 671 3108 832 3120
rect 671 3068 672 3108
rect 618 3052 672 3068
rect 924 2964 974 3370
rect 1152 3126 1180 4244
rect 2432 4242 2500 4252
rect 2312 4069 2376 4076
rect 2312 4038 2318 4069
rect 1584 4017 2318 4038
rect 2370 4017 2376 4069
rect 1584 4010 2376 4017
rect 1584 4008 2318 4010
rect 1584 4002 2312 4008
rect 1484 3672 1548 3680
rect 1484 3620 1490 3672
rect 1542 3620 1548 3672
rect 1484 3612 1548 3620
rect 1244 3584 1310 3590
rect 1244 3532 1252 3584
rect 1304 3554 1310 3584
rect 1484 3554 1512 3612
rect 1304 3532 1512 3554
rect 1244 3526 1512 3532
rect 1584 3376 1612 4002
rect 2312 3936 2378 3942
rect 2312 3884 2320 3936
rect 2372 3884 2378 3936
rect 2312 3878 2378 3884
rect 2312 3756 2340 3878
rect 2272 3728 2340 3756
rect 1584 3368 1896 3376
rect 1584 3340 1835 3368
rect 1244 3152 1320 3158
rect 1244 3126 1252 3152
rect 1152 3100 1252 3126
rect 1304 3100 1320 3152
rect 1152 3098 1320 3100
rect 1244 3094 1320 3098
rect 924 2958 990 2964
rect 924 2906 932 2958
rect 984 2936 990 2958
rect 1584 2936 1612 3340
rect 1816 3316 1835 3340
rect 1887 3316 1896 3368
rect 1816 3304 1896 3316
rect 2132 3372 2200 3378
rect 2132 3320 2139 3372
rect 2191 3320 2200 3372
rect 2132 3314 2200 3320
rect 984 2908 1612 2936
rect 984 2906 990 2908
rect 924 2900 990 2906
rect 1738 2708 2088 2722
rect -150 2578 200 2592
rect 1738 2592 1759 2708
rect 2067 2592 2088 2708
rect 2132 2698 2176 3314
rect 2272 3144 2300 3728
rect 2334 3678 2396 3684
rect 2334 3626 2344 3678
rect 2432 3670 2460 4242
rect 2488 4069 2552 4076
rect 2488 4017 2494 4069
rect 2546 4036 2552 4069
rect 2814 4036 2864 4426
rect 3336 4424 3364 4524
rect 3336 4418 3402 4424
rect 4450 4422 4478 4524
rect 4686 4486 4752 4494
rect 4686 4434 4692 4486
rect 4744 4434 4752 4486
rect 4686 4426 4752 4434
rect 3336 4404 3344 4418
rect 3338 4366 3344 4404
rect 3396 4366 3402 4418
rect 3338 4360 3402 4366
rect 4410 4416 4478 4422
rect 4410 4364 4420 4416
rect 4472 4364 4478 4416
rect 4410 4358 4478 4364
rect 3250 4302 3314 4308
rect 3250 4272 3256 4302
rect 3040 4250 3256 4272
rect 3308 4250 3314 4302
rect 3040 4244 3314 4250
rect 4320 4304 4388 4310
rect 4320 4252 4328 4304
rect 4380 4252 4388 4304
rect 2546 4020 2866 4036
rect 2546 4017 2880 4020
rect 2488 4014 2880 4017
rect 2488 4008 2822 4014
rect 2814 3962 2822 4008
rect 2874 3962 2880 4014
rect 2814 3956 2880 3962
rect 2684 3820 2756 3832
rect 2684 3768 2694 3820
rect 2746 3768 2756 3820
rect 2684 3756 2756 3768
rect 2720 3754 2756 3756
rect 2432 3642 2720 3670
rect 2334 3620 2396 3626
rect 2368 3574 2396 3620
rect 2368 3570 2612 3574
rect 2368 3564 2650 3570
rect 2368 3546 2590 3564
rect 2584 3512 2590 3546
rect 2642 3512 2650 3564
rect 2584 3504 2650 3512
rect 2272 3130 2336 3144
rect 2692 3136 2720 3642
rect 2796 3430 2862 3438
rect 2796 3378 2802 3430
rect 2854 3378 2862 3430
rect 2796 3370 2862 3378
rect 2272 3078 2275 3130
rect 2327 3078 2336 3130
rect 2272 3062 2336 3078
rect 2506 3120 2720 3136
rect 2506 3068 2507 3120
rect 2559 3108 2720 3120
rect 2559 3068 2560 3108
rect 2506 3052 2560 3068
rect 2812 2964 2862 3370
rect 3040 3126 3068 4244
rect 4320 4242 4388 4252
rect 4200 4069 4264 4076
rect 4200 4038 4206 4069
rect 3472 4017 4206 4038
rect 4258 4017 4264 4069
rect 3472 4010 4264 4017
rect 3472 4008 4206 4010
rect 3472 4002 4200 4008
rect 3372 3672 3436 3680
rect 3372 3620 3378 3672
rect 3430 3620 3436 3672
rect 3372 3612 3436 3620
rect 3132 3584 3198 3590
rect 3132 3532 3140 3584
rect 3192 3554 3198 3584
rect 3372 3554 3400 3612
rect 3192 3532 3400 3554
rect 3132 3526 3400 3532
rect 3472 3376 3500 4002
rect 4200 3936 4266 3942
rect 4200 3884 4208 3936
rect 4260 3884 4266 3936
rect 4200 3878 4266 3884
rect 4200 3756 4228 3878
rect 4160 3728 4228 3756
rect 3472 3368 3784 3376
rect 3472 3340 3723 3368
rect 3132 3152 3208 3158
rect 3132 3126 3140 3152
rect 3040 3100 3140 3126
rect 3192 3100 3208 3152
rect 3040 3098 3208 3100
rect 3132 3094 3208 3098
rect 2812 2958 2878 2964
rect 2812 2906 2820 2958
rect 2872 2936 2878 2958
rect 3472 2936 3500 3340
rect 3704 3316 3723 3340
rect 3775 3316 3784 3368
rect 3704 3304 3784 3316
rect 4020 3372 4088 3378
rect 4020 3320 4027 3372
rect 4079 3320 4088 3372
rect 4020 3314 4088 3320
rect 2872 2908 3500 2936
rect 2872 2906 2878 2908
rect 2812 2900 2878 2906
rect 3626 2708 3976 2722
rect 1738 2578 2088 2592
rect 3626 2592 3647 2708
rect 3955 2592 3976 2708
rect 4020 2698 4064 3314
rect 4160 3144 4188 3728
rect 4222 3678 4284 3684
rect 4222 3626 4232 3678
rect 4320 3670 4348 4242
rect 4376 4069 4440 4076
rect 4376 4017 4382 4069
rect 4434 4036 4440 4069
rect 4702 4036 4752 4426
rect 5224 4424 5252 4524
rect 5224 4418 5290 4424
rect 6338 4422 6366 4524
rect 6574 4486 6640 4494
rect 6574 4434 6580 4486
rect 6632 4434 6640 4486
rect 6574 4426 6640 4434
rect 5224 4404 5232 4418
rect 5226 4366 5232 4404
rect 5284 4366 5290 4418
rect 5226 4360 5290 4366
rect 6298 4416 6366 4422
rect 6298 4364 6308 4416
rect 6360 4364 6366 4416
rect 6298 4358 6366 4364
rect 5138 4302 5202 4308
rect 5138 4272 5144 4302
rect 4928 4250 5144 4272
rect 5196 4250 5202 4302
rect 4928 4244 5202 4250
rect 6208 4304 6276 4310
rect 6208 4252 6216 4304
rect 6268 4252 6276 4304
rect 4434 4020 4754 4036
rect 4434 4017 4768 4020
rect 4376 4014 4768 4017
rect 4376 4008 4710 4014
rect 4702 3962 4710 4008
rect 4762 3962 4768 4014
rect 4702 3956 4768 3962
rect 4572 3820 4644 3832
rect 4572 3768 4582 3820
rect 4634 3768 4644 3820
rect 4572 3756 4644 3768
rect 4608 3754 4644 3756
rect 4320 3642 4608 3670
rect 4222 3620 4284 3626
rect 4256 3574 4284 3620
rect 4256 3570 4500 3574
rect 4256 3564 4538 3570
rect 4256 3546 4478 3564
rect 4472 3512 4478 3546
rect 4530 3512 4538 3564
rect 4472 3504 4538 3512
rect 4160 3130 4224 3144
rect 4580 3136 4608 3642
rect 4684 3430 4750 3438
rect 4684 3378 4690 3430
rect 4742 3378 4750 3430
rect 4684 3370 4750 3378
rect 4160 3078 4163 3130
rect 4215 3078 4224 3130
rect 4160 3062 4224 3078
rect 4394 3120 4608 3136
rect 4394 3068 4395 3120
rect 4447 3108 4608 3120
rect 4447 3068 4448 3108
rect 4394 3052 4448 3068
rect 4700 2964 4750 3370
rect 4928 3126 4956 4244
rect 6208 4242 6276 4252
rect 6088 4069 6152 4076
rect 6088 4038 6094 4069
rect 5360 4017 6094 4038
rect 6146 4017 6152 4069
rect 5360 4010 6152 4017
rect 5360 4008 6094 4010
rect 5360 4002 6088 4008
rect 5260 3672 5324 3680
rect 5260 3620 5266 3672
rect 5318 3620 5324 3672
rect 5260 3612 5324 3620
rect 5020 3584 5086 3590
rect 5020 3532 5028 3584
rect 5080 3554 5086 3584
rect 5260 3554 5288 3612
rect 5080 3532 5288 3554
rect 5020 3526 5288 3532
rect 5360 3376 5388 4002
rect 6088 3936 6154 3942
rect 6088 3884 6096 3936
rect 6148 3884 6154 3936
rect 6088 3878 6154 3884
rect 6088 3756 6116 3878
rect 6048 3728 6116 3756
rect 5360 3368 5672 3376
rect 5360 3340 5611 3368
rect 5020 3152 5096 3158
rect 5020 3126 5028 3152
rect 4928 3100 5028 3126
rect 5080 3100 5096 3152
rect 4928 3098 5096 3100
rect 5020 3094 5096 3098
rect 4700 2958 4766 2964
rect 4700 2906 4708 2958
rect 4760 2936 4766 2958
rect 5360 2936 5388 3340
rect 5592 3316 5611 3340
rect 5663 3316 5672 3368
rect 5592 3304 5672 3316
rect 5908 3372 5976 3378
rect 5908 3320 5915 3372
rect 5967 3320 5976 3372
rect 5908 3314 5976 3320
rect 4760 2908 5388 2936
rect 4760 2906 4766 2908
rect 4700 2900 4766 2906
rect 5514 2708 5864 2722
rect 3626 2578 3976 2592
rect 5514 2592 5535 2708
rect 5843 2592 5864 2708
rect 5908 2698 5952 3314
rect 6048 3144 6076 3728
rect 6110 3678 6172 3684
rect 6110 3626 6120 3678
rect 6208 3670 6236 4242
rect 6264 4069 6328 4076
rect 6264 4017 6270 4069
rect 6322 4036 6328 4069
rect 6590 4036 6640 4426
rect 7112 4424 7140 4524
rect 7112 4418 7178 4424
rect 8226 4422 8254 4524
rect 8462 4486 8528 4494
rect 8462 4434 8468 4486
rect 8520 4434 8528 4486
rect 8462 4426 8528 4434
rect 7112 4404 7120 4418
rect 7114 4366 7120 4404
rect 7172 4366 7178 4418
rect 7114 4360 7178 4366
rect 8186 4416 8254 4422
rect 8186 4364 8196 4416
rect 8248 4364 8254 4416
rect 8186 4358 8254 4364
rect 7026 4302 7090 4308
rect 7026 4272 7032 4302
rect 6816 4250 7032 4272
rect 7084 4250 7090 4302
rect 6816 4244 7090 4250
rect 8096 4304 8164 4310
rect 8096 4252 8104 4304
rect 8156 4252 8164 4304
rect 6322 4020 6642 4036
rect 6322 4017 6656 4020
rect 6264 4014 6656 4017
rect 6264 4008 6598 4014
rect 6590 3962 6598 4008
rect 6650 3962 6656 4014
rect 6590 3956 6656 3962
rect 6460 3820 6532 3832
rect 6460 3768 6470 3820
rect 6522 3768 6532 3820
rect 6460 3756 6532 3768
rect 6496 3754 6532 3756
rect 6208 3642 6496 3670
rect 6110 3620 6172 3626
rect 6144 3574 6172 3620
rect 6144 3570 6388 3574
rect 6144 3564 6426 3570
rect 6144 3546 6366 3564
rect 6360 3512 6366 3546
rect 6418 3512 6426 3564
rect 6360 3504 6426 3512
rect 6048 3130 6112 3144
rect 6468 3136 6496 3642
rect 6572 3430 6638 3438
rect 6572 3378 6578 3430
rect 6630 3378 6638 3430
rect 6572 3370 6638 3378
rect 6048 3078 6051 3130
rect 6103 3078 6112 3130
rect 6048 3062 6112 3078
rect 6282 3120 6496 3136
rect 6282 3068 6283 3120
rect 6335 3108 6496 3120
rect 6335 3068 6336 3108
rect 6282 3052 6336 3068
rect 6588 2964 6638 3370
rect 6816 3126 6844 4244
rect 8096 4242 8164 4252
rect 7976 4069 8040 4076
rect 7976 4038 7982 4069
rect 7248 4017 7982 4038
rect 8034 4017 8040 4069
rect 7248 4010 8040 4017
rect 7248 4008 7982 4010
rect 7248 4002 7976 4008
rect 7148 3672 7212 3680
rect 7148 3620 7154 3672
rect 7206 3620 7212 3672
rect 7148 3612 7212 3620
rect 6908 3584 6974 3590
rect 6908 3532 6916 3584
rect 6968 3554 6974 3584
rect 7148 3554 7176 3612
rect 6968 3532 7176 3554
rect 6908 3526 7176 3532
rect 7248 3376 7276 4002
rect 7976 3936 8042 3942
rect 7976 3884 7984 3936
rect 8036 3884 8042 3936
rect 7976 3878 8042 3884
rect 7976 3756 8004 3878
rect 7936 3728 8004 3756
rect 7248 3368 7560 3376
rect 7248 3340 7499 3368
rect 6908 3152 6984 3158
rect 6908 3126 6916 3152
rect 6816 3100 6916 3126
rect 6968 3100 6984 3152
rect 6816 3098 6984 3100
rect 6908 3094 6984 3098
rect 6588 2958 6654 2964
rect 6588 2906 6596 2958
rect 6648 2936 6654 2958
rect 7248 2936 7276 3340
rect 7480 3316 7499 3340
rect 7551 3316 7560 3368
rect 7480 3304 7560 3316
rect 7796 3372 7864 3378
rect 7796 3320 7803 3372
rect 7855 3320 7864 3372
rect 7796 3314 7864 3320
rect 6648 2908 7276 2936
rect 6648 2906 6654 2908
rect 6588 2900 6654 2906
rect 7402 2708 7752 2722
rect 5514 2578 5864 2592
rect 7402 2592 7423 2708
rect 7731 2592 7752 2708
rect 7796 2698 7840 3314
rect 7936 3144 7964 3728
rect 7998 3678 8060 3684
rect 7998 3626 8008 3678
rect 8096 3670 8124 4242
rect 8152 4069 8216 4076
rect 8152 4017 8158 4069
rect 8210 4036 8216 4069
rect 8478 4036 8528 4426
rect 9000 4424 9028 4524
rect 9000 4418 9066 4424
rect 10114 4422 10142 4524
rect 10350 4486 10416 4494
rect 10350 4434 10356 4486
rect 10408 4434 10416 4486
rect 10350 4426 10416 4434
rect 9000 4404 9008 4418
rect 9002 4366 9008 4404
rect 9060 4366 9066 4418
rect 9002 4360 9066 4366
rect 10074 4416 10142 4422
rect 10074 4364 10084 4416
rect 10136 4364 10142 4416
rect 10074 4358 10142 4364
rect 8914 4302 8978 4308
rect 8914 4272 8920 4302
rect 8704 4250 8920 4272
rect 8972 4250 8978 4302
rect 8704 4244 8978 4250
rect 9984 4304 10052 4310
rect 9984 4252 9992 4304
rect 10044 4252 10052 4304
rect 8210 4020 8530 4036
rect 8210 4017 8544 4020
rect 8152 4014 8544 4017
rect 8152 4008 8486 4014
rect 8478 3962 8486 4008
rect 8538 3962 8544 4014
rect 8478 3956 8544 3962
rect 8348 3820 8420 3832
rect 8348 3768 8358 3820
rect 8410 3768 8420 3820
rect 8348 3756 8420 3768
rect 8384 3754 8420 3756
rect 8096 3642 8384 3670
rect 7998 3620 8060 3626
rect 8032 3574 8060 3620
rect 8032 3570 8276 3574
rect 8032 3564 8314 3570
rect 8032 3546 8254 3564
rect 8248 3512 8254 3546
rect 8306 3512 8314 3564
rect 8248 3504 8314 3512
rect 7936 3130 8000 3144
rect 8356 3136 8384 3642
rect 8460 3430 8526 3438
rect 8460 3378 8466 3430
rect 8518 3378 8526 3430
rect 8460 3370 8526 3378
rect 7936 3078 7939 3130
rect 7991 3078 8000 3130
rect 7936 3062 8000 3078
rect 8170 3120 8384 3136
rect 8170 3068 8171 3120
rect 8223 3108 8384 3120
rect 8223 3068 8224 3108
rect 8170 3052 8224 3068
rect 8476 2964 8526 3370
rect 8704 3126 8732 4244
rect 9984 4242 10052 4252
rect 9864 4069 9928 4076
rect 9864 4038 9870 4069
rect 9136 4017 9870 4038
rect 9922 4017 9928 4069
rect 9136 4010 9928 4017
rect 9136 4008 9870 4010
rect 9136 4002 9864 4008
rect 9036 3672 9100 3680
rect 9036 3620 9042 3672
rect 9094 3620 9100 3672
rect 9036 3612 9100 3620
rect 8796 3584 8862 3590
rect 8796 3532 8804 3584
rect 8856 3554 8862 3584
rect 9036 3554 9064 3612
rect 8856 3532 9064 3554
rect 8796 3526 9064 3532
rect 9136 3376 9164 4002
rect 9864 3936 9930 3942
rect 9864 3884 9872 3936
rect 9924 3884 9930 3936
rect 9864 3878 9930 3884
rect 9864 3756 9892 3878
rect 9824 3728 9892 3756
rect 9136 3368 9448 3376
rect 9136 3340 9387 3368
rect 8796 3152 8872 3158
rect 8796 3126 8804 3152
rect 8704 3100 8804 3126
rect 8856 3100 8872 3152
rect 8704 3098 8872 3100
rect 8796 3094 8872 3098
rect 8476 2958 8542 2964
rect 8476 2906 8484 2958
rect 8536 2936 8542 2958
rect 9136 2936 9164 3340
rect 9368 3316 9387 3340
rect 9439 3316 9448 3368
rect 9368 3304 9448 3316
rect 9684 3372 9752 3378
rect 9684 3320 9691 3372
rect 9743 3320 9752 3372
rect 9684 3314 9752 3320
rect 8536 2908 9164 2936
rect 8536 2906 8542 2908
rect 8476 2900 8542 2906
rect 9290 2708 9640 2722
rect 7402 2578 7752 2592
rect 9290 2592 9311 2708
rect 9619 2592 9640 2708
rect 9684 2698 9728 3314
rect 9824 3144 9852 3728
rect 9886 3678 9948 3684
rect 9886 3626 9896 3678
rect 9984 3670 10012 4242
rect 10040 4069 10104 4076
rect 10040 4017 10046 4069
rect 10098 4036 10104 4069
rect 10366 4036 10416 4426
rect 10888 4424 10916 4524
rect 10888 4418 10954 4424
rect 11996 4422 12024 4528
rect 12232 4486 12298 4494
rect 12232 4434 12238 4486
rect 12290 4434 12298 4486
rect 12232 4426 12298 4434
rect 10888 4404 10896 4418
rect 10890 4366 10896 4404
rect 10948 4366 10954 4418
rect 10890 4360 10954 4366
rect 11956 4416 12024 4422
rect 11956 4364 11966 4416
rect 12018 4364 12024 4416
rect 11956 4358 12024 4364
rect 10802 4302 10866 4308
rect 10802 4272 10808 4302
rect 10592 4250 10808 4272
rect 10860 4250 10866 4302
rect 10592 4244 10866 4250
rect 11866 4304 11934 4310
rect 11866 4252 11874 4304
rect 11926 4252 11934 4304
rect 10098 4020 10418 4036
rect 10098 4017 10432 4020
rect 10040 4014 10432 4017
rect 10040 4008 10374 4014
rect 10366 3962 10374 4008
rect 10426 3962 10432 4014
rect 10366 3956 10432 3962
rect 10236 3820 10308 3832
rect 10236 3768 10246 3820
rect 10298 3768 10308 3820
rect 10236 3756 10308 3768
rect 10272 3754 10308 3756
rect 9984 3642 10272 3670
rect 9886 3620 9948 3626
rect 9920 3574 9948 3620
rect 9920 3570 10164 3574
rect 9920 3564 10202 3570
rect 9920 3546 10142 3564
rect 10136 3512 10142 3546
rect 10194 3512 10202 3564
rect 10136 3504 10202 3512
rect 9824 3130 9888 3144
rect 10244 3136 10272 3642
rect 10348 3430 10414 3438
rect 10348 3378 10354 3430
rect 10406 3378 10414 3430
rect 10348 3370 10414 3378
rect 9824 3078 9827 3130
rect 9879 3078 9888 3130
rect 9824 3062 9888 3078
rect 10058 3120 10272 3136
rect 10058 3068 10059 3120
rect 10111 3108 10272 3120
rect 10111 3068 10112 3108
rect 10058 3052 10112 3068
rect 10364 2964 10414 3370
rect 10592 3126 10620 4244
rect 11866 4242 11934 4252
rect 11746 4069 11810 4076
rect 11746 4038 11752 4069
rect 11024 4017 11752 4038
rect 11804 4017 11810 4069
rect 11024 4010 11810 4017
rect 11024 4008 11752 4010
rect 11024 4002 11746 4008
rect 10924 3672 10988 3680
rect 10924 3620 10930 3672
rect 10982 3620 10988 3672
rect 10924 3612 10988 3620
rect 10684 3584 10750 3590
rect 10684 3532 10692 3584
rect 10744 3554 10750 3584
rect 10924 3554 10952 3612
rect 10744 3532 10952 3554
rect 10684 3526 10952 3532
rect 11024 3376 11052 4002
rect 11746 3936 11812 3942
rect 11746 3884 11754 3936
rect 11806 3884 11812 3936
rect 11746 3878 11812 3884
rect 11746 3756 11774 3878
rect 11706 3728 11774 3756
rect 11024 3368 11336 3376
rect 11024 3340 11275 3368
rect 10684 3152 10760 3158
rect 10684 3126 10692 3152
rect 10592 3100 10692 3126
rect 10744 3100 10760 3152
rect 10592 3098 10760 3100
rect 10684 3094 10760 3098
rect 10364 2958 10430 2964
rect 10364 2906 10372 2958
rect 10424 2936 10430 2958
rect 11024 2936 11052 3340
rect 11256 3316 11275 3340
rect 11327 3316 11336 3368
rect 11256 3304 11336 3316
rect 11566 3372 11634 3378
rect 11566 3320 11573 3372
rect 11625 3320 11634 3372
rect 11566 3314 11634 3320
rect 10424 2908 11052 2936
rect 10424 2906 10430 2908
rect 10364 2900 10430 2906
rect 11178 2708 11528 2722
rect 9290 2578 9640 2592
rect 11178 2592 11199 2708
rect 11507 2592 11528 2708
rect 11566 2698 11610 3314
rect 11706 3144 11734 3728
rect 11768 3678 11830 3684
rect 11768 3626 11778 3678
rect 11866 3670 11894 4242
rect 11922 4069 11986 4076
rect 11922 4017 11928 4069
rect 11980 4036 11986 4069
rect 12248 4036 12298 4426
rect 12770 4424 12798 4528
rect 12770 4418 12836 4424
rect 13884 4422 13912 4528
rect 14120 4486 14186 4494
rect 14120 4434 14126 4486
rect 14178 4434 14186 4486
rect 14120 4426 14186 4434
rect 12770 4404 12778 4418
rect 12772 4366 12778 4404
rect 12830 4366 12836 4418
rect 12772 4360 12836 4366
rect 13844 4416 13912 4422
rect 13844 4364 13854 4416
rect 13906 4364 13912 4416
rect 13844 4358 13912 4364
rect 12684 4302 12748 4308
rect 12684 4272 12690 4302
rect 12474 4250 12690 4272
rect 12742 4250 12748 4302
rect 12474 4244 12748 4250
rect 13754 4304 13822 4310
rect 13754 4252 13762 4304
rect 13814 4252 13822 4304
rect 11980 4020 12300 4036
rect 11980 4017 12314 4020
rect 11922 4014 12314 4017
rect 11922 4008 12256 4014
rect 12248 3962 12256 4008
rect 12308 3962 12314 4014
rect 12248 3956 12314 3962
rect 12118 3820 12190 3832
rect 12118 3768 12128 3820
rect 12180 3768 12190 3820
rect 12118 3756 12190 3768
rect 12154 3754 12190 3756
rect 11866 3642 12154 3670
rect 11768 3620 11830 3626
rect 11802 3574 11830 3620
rect 11802 3570 12046 3574
rect 11802 3564 12084 3570
rect 11802 3546 12024 3564
rect 12018 3512 12024 3546
rect 12076 3512 12084 3564
rect 12018 3504 12084 3512
rect 11706 3130 11770 3144
rect 12126 3136 12154 3642
rect 12230 3430 12296 3438
rect 12230 3378 12236 3430
rect 12288 3378 12296 3430
rect 12230 3370 12296 3378
rect 11706 3078 11709 3130
rect 11761 3078 11770 3130
rect 11706 3062 11770 3078
rect 11940 3120 12154 3136
rect 11940 3068 11941 3120
rect 11993 3108 12154 3120
rect 11993 3068 11994 3108
rect 11940 3052 11994 3068
rect 12246 2964 12296 3370
rect 12474 3126 12502 4244
rect 13754 4242 13822 4252
rect 13634 4069 13698 4076
rect 13634 4038 13640 4069
rect 12906 4017 13640 4038
rect 13692 4017 13698 4069
rect 12906 4010 13698 4017
rect 12906 4008 13640 4010
rect 12906 4002 13634 4008
rect 12806 3672 12870 3680
rect 12806 3620 12812 3672
rect 12864 3620 12870 3672
rect 12806 3612 12870 3620
rect 12566 3584 12632 3590
rect 12566 3532 12574 3584
rect 12626 3554 12632 3584
rect 12806 3554 12834 3612
rect 12626 3532 12834 3554
rect 12566 3526 12834 3532
rect 12906 3376 12934 4002
rect 13634 3936 13700 3942
rect 13634 3884 13642 3936
rect 13694 3884 13700 3936
rect 13634 3878 13700 3884
rect 13634 3756 13662 3878
rect 13594 3728 13662 3756
rect 12906 3368 13218 3376
rect 12906 3340 13157 3368
rect 12566 3152 12642 3158
rect 12566 3126 12574 3152
rect 12474 3100 12574 3126
rect 12626 3100 12642 3152
rect 12474 3098 12642 3100
rect 12566 3094 12642 3098
rect 12246 2958 12312 2964
rect 12246 2906 12254 2958
rect 12306 2936 12312 2958
rect 12906 2936 12934 3340
rect 13138 3316 13157 3340
rect 13209 3316 13218 3368
rect 13138 3304 13218 3316
rect 13454 3372 13522 3378
rect 13454 3320 13461 3372
rect 13513 3320 13522 3372
rect 13454 3314 13522 3320
rect 12306 2908 12934 2936
rect 12306 2906 12312 2908
rect 12246 2900 12312 2906
rect 13060 2708 13410 2722
rect 11178 2578 11528 2592
rect 13060 2592 13081 2708
rect 13389 2592 13410 2708
rect 13454 2698 13498 3314
rect 13594 3144 13622 3728
rect 13656 3678 13718 3684
rect 13656 3626 13666 3678
rect 13754 3670 13782 4242
rect 13810 4069 13874 4076
rect 13810 4017 13816 4069
rect 13868 4036 13874 4069
rect 14136 4036 14186 4426
rect 14658 4424 14686 4528
rect 14658 4418 14724 4424
rect 15772 4422 15800 4528
rect 16008 4486 16074 4494
rect 16008 4434 16014 4486
rect 16066 4434 16074 4486
rect 16008 4426 16074 4434
rect 14658 4404 14666 4418
rect 14660 4366 14666 4404
rect 14718 4366 14724 4418
rect 14660 4360 14724 4366
rect 15732 4416 15800 4422
rect 15732 4364 15742 4416
rect 15794 4364 15800 4416
rect 15732 4358 15800 4364
rect 14572 4302 14636 4308
rect 14572 4272 14578 4302
rect 14362 4250 14578 4272
rect 14630 4250 14636 4302
rect 14362 4244 14636 4250
rect 15642 4304 15710 4310
rect 15642 4252 15650 4304
rect 15702 4252 15710 4304
rect 13868 4020 14188 4036
rect 13868 4017 14202 4020
rect 13810 4014 14202 4017
rect 13810 4008 14144 4014
rect 14136 3962 14144 4008
rect 14196 3962 14202 4014
rect 14136 3956 14202 3962
rect 14006 3820 14078 3832
rect 14006 3768 14016 3820
rect 14068 3768 14078 3820
rect 14006 3756 14078 3768
rect 14042 3754 14078 3756
rect 13754 3642 14042 3670
rect 13656 3620 13718 3626
rect 13690 3574 13718 3620
rect 13690 3570 13934 3574
rect 13690 3564 13972 3570
rect 13690 3546 13912 3564
rect 13906 3512 13912 3546
rect 13964 3512 13972 3564
rect 13906 3504 13972 3512
rect 13594 3130 13658 3144
rect 14014 3136 14042 3642
rect 14118 3430 14184 3438
rect 14118 3378 14124 3430
rect 14176 3378 14184 3430
rect 14118 3370 14184 3378
rect 13594 3078 13597 3130
rect 13649 3078 13658 3130
rect 13594 3062 13658 3078
rect 13828 3120 14042 3136
rect 13828 3068 13829 3120
rect 13881 3108 14042 3120
rect 13881 3068 13882 3108
rect 13828 3052 13882 3068
rect 14134 2964 14184 3370
rect 14362 3126 14390 4244
rect 15642 4242 15710 4252
rect 15522 4069 15586 4076
rect 15522 4038 15528 4069
rect 14794 4017 15528 4038
rect 15580 4017 15586 4069
rect 14794 4010 15586 4017
rect 14794 4008 15528 4010
rect 14794 4002 15522 4008
rect 14694 3672 14758 3680
rect 14694 3620 14700 3672
rect 14752 3620 14758 3672
rect 14694 3612 14758 3620
rect 14454 3584 14520 3590
rect 14454 3532 14462 3584
rect 14514 3554 14520 3584
rect 14694 3554 14722 3612
rect 14514 3532 14722 3554
rect 14454 3526 14722 3532
rect 14794 3376 14822 4002
rect 15522 3936 15588 3942
rect 15522 3884 15530 3936
rect 15582 3884 15588 3936
rect 15522 3878 15588 3884
rect 15522 3756 15550 3878
rect 15482 3728 15550 3756
rect 14794 3368 15106 3376
rect 14794 3340 15045 3368
rect 14454 3152 14530 3158
rect 14454 3126 14462 3152
rect 14362 3100 14462 3126
rect 14514 3100 14530 3152
rect 14362 3098 14530 3100
rect 14454 3094 14530 3098
rect 14134 2958 14200 2964
rect 14134 2906 14142 2958
rect 14194 2936 14200 2958
rect 14794 2936 14822 3340
rect 15026 3316 15045 3340
rect 15097 3316 15106 3368
rect 15026 3304 15106 3316
rect 15342 3372 15410 3378
rect 15342 3320 15349 3372
rect 15401 3320 15410 3372
rect 15342 3314 15410 3320
rect 14194 2908 14822 2936
rect 14194 2906 14200 2908
rect 14134 2900 14200 2906
rect 14948 2708 15298 2722
rect 13060 2578 13410 2592
rect 14948 2592 14969 2708
rect 15277 2592 15298 2708
rect 15342 2698 15386 3314
rect 15482 3144 15510 3728
rect 15544 3678 15606 3684
rect 15544 3626 15554 3678
rect 15642 3670 15670 4242
rect 15698 4069 15762 4076
rect 15698 4017 15704 4069
rect 15756 4036 15762 4069
rect 16024 4036 16074 4426
rect 16546 4424 16574 4528
rect 17248 4524 18568 4528
rect 19132 4524 20456 4528
rect 16546 4418 16612 4424
rect 17660 4422 17688 4524
rect 17896 4486 17962 4494
rect 17896 4434 17902 4486
rect 17954 4434 17962 4486
rect 17896 4426 17962 4434
rect 16546 4404 16554 4418
rect 16548 4366 16554 4404
rect 16606 4366 16612 4418
rect 16548 4360 16612 4366
rect 17620 4416 17688 4422
rect 17620 4364 17630 4416
rect 17682 4364 17688 4416
rect 17620 4358 17688 4364
rect 16460 4302 16524 4308
rect 16460 4272 16466 4302
rect 16250 4250 16466 4272
rect 16518 4250 16524 4302
rect 16250 4244 16524 4250
rect 17530 4304 17598 4310
rect 17530 4252 17538 4304
rect 17590 4252 17598 4304
rect 15756 4020 16076 4036
rect 15756 4017 16090 4020
rect 15698 4014 16090 4017
rect 15698 4008 16032 4014
rect 16024 3962 16032 4008
rect 16084 3962 16090 4014
rect 16024 3956 16090 3962
rect 15894 3820 15966 3832
rect 15894 3768 15904 3820
rect 15956 3768 15966 3820
rect 15894 3756 15966 3768
rect 15930 3754 15966 3756
rect 15642 3642 15930 3670
rect 15544 3620 15606 3626
rect 15578 3574 15606 3620
rect 15578 3570 15822 3574
rect 15578 3564 15860 3570
rect 15578 3546 15800 3564
rect 15794 3512 15800 3546
rect 15852 3512 15860 3564
rect 15794 3504 15860 3512
rect 15482 3130 15546 3144
rect 15902 3136 15930 3642
rect 16006 3430 16072 3438
rect 16006 3378 16012 3430
rect 16064 3378 16072 3430
rect 16006 3370 16072 3378
rect 15482 3078 15485 3130
rect 15537 3078 15546 3130
rect 15482 3062 15546 3078
rect 15716 3120 15930 3136
rect 15716 3068 15717 3120
rect 15769 3108 15930 3120
rect 15769 3068 15770 3108
rect 15716 3052 15770 3068
rect 16022 2964 16072 3370
rect 16250 3126 16278 4244
rect 17530 4242 17598 4252
rect 17410 4069 17474 4076
rect 17410 4038 17416 4069
rect 16682 4017 17416 4038
rect 17468 4017 17474 4069
rect 16682 4010 17474 4017
rect 16682 4008 17416 4010
rect 16682 4002 17410 4008
rect 16582 3672 16646 3680
rect 16582 3620 16588 3672
rect 16640 3620 16646 3672
rect 16582 3612 16646 3620
rect 16342 3584 16408 3590
rect 16342 3532 16350 3584
rect 16402 3554 16408 3584
rect 16582 3554 16610 3612
rect 16402 3532 16610 3554
rect 16342 3526 16610 3532
rect 16682 3376 16710 4002
rect 17410 3936 17476 3942
rect 17410 3884 17418 3936
rect 17470 3884 17476 3936
rect 17410 3878 17476 3884
rect 17410 3756 17438 3878
rect 17370 3728 17438 3756
rect 16682 3368 16994 3376
rect 16682 3340 16933 3368
rect 16342 3152 16418 3158
rect 16342 3126 16350 3152
rect 16250 3100 16350 3126
rect 16402 3100 16418 3152
rect 16250 3098 16418 3100
rect 16342 3094 16418 3098
rect 16022 2958 16088 2964
rect 16022 2906 16030 2958
rect 16082 2936 16088 2958
rect 16682 2936 16710 3340
rect 16914 3316 16933 3340
rect 16985 3316 16994 3368
rect 16914 3304 16994 3316
rect 17230 3372 17298 3378
rect 17230 3320 17237 3372
rect 17289 3320 17298 3372
rect 17230 3314 17298 3320
rect 16082 2908 16710 2936
rect 16082 2906 16088 2908
rect 16022 2900 16088 2906
rect 16836 2708 17186 2722
rect 14948 2578 15298 2592
rect 16836 2592 16857 2708
rect 17165 2592 17186 2708
rect 17230 2698 17274 3314
rect 17370 3144 17398 3728
rect 17432 3678 17494 3684
rect 17432 3626 17442 3678
rect 17530 3670 17558 4242
rect 17586 4069 17650 4076
rect 17586 4017 17592 4069
rect 17644 4036 17650 4069
rect 17912 4036 17962 4426
rect 18434 4424 18462 4524
rect 18434 4418 18500 4424
rect 19548 4422 19576 4524
rect 19784 4486 19850 4494
rect 19784 4434 19790 4486
rect 19842 4434 19850 4486
rect 19784 4426 19850 4434
rect 18434 4404 18442 4418
rect 18436 4366 18442 4404
rect 18494 4366 18500 4418
rect 18436 4360 18500 4366
rect 19508 4416 19576 4422
rect 19508 4364 19518 4416
rect 19570 4364 19576 4416
rect 19508 4358 19576 4364
rect 18348 4302 18412 4308
rect 18348 4272 18354 4302
rect 18138 4250 18354 4272
rect 18406 4250 18412 4302
rect 18138 4244 18412 4250
rect 19418 4304 19486 4310
rect 19418 4252 19426 4304
rect 19478 4252 19486 4304
rect 17644 4020 17964 4036
rect 17644 4017 17978 4020
rect 17586 4014 17978 4017
rect 17586 4008 17920 4014
rect 17912 3962 17920 4008
rect 17972 3962 17978 4014
rect 17912 3956 17978 3962
rect 17782 3820 17854 3832
rect 17782 3768 17792 3820
rect 17844 3768 17854 3820
rect 17782 3756 17854 3768
rect 17818 3754 17854 3756
rect 17530 3642 17818 3670
rect 17432 3620 17494 3626
rect 17466 3574 17494 3620
rect 17466 3570 17710 3574
rect 17466 3564 17748 3570
rect 17466 3546 17688 3564
rect 17682 3512 17688 3546
rect 17740 3512 17748 3564
rect 17682 3504 17748 3512
rect 17370 3130 17434 3144
rect 17790 3136 17818 3642
rect 17894 3430 17960 3438
rect 17894 3378 17900 3430
rect 17952 3378 17960 3430
rect 17894 3370 17960 3378
rect 17370 3078 17373 3130
rect 17425 3078 17434 3130
rect 17370 3062 17434 3078
rect 17604 3120 17818 3136
rect 17604 3068 17605 3120
rect 17657 3108 17818 3120
rect 17657 3068 17658 3108
rect 17604 3052 17658 3068
rect 17910 2964 17960 3370
rect 18138 3126 18166 4244
rect 19418 4242 19486 4252
rect 19298 4069 19362 4076
rect 19298 4038 19304 4069
rect 18570 4017 19304 4038
rect 19356 4017 19362 4069
rect 18570 4010 19362 4017
rect 18570 4008 19304 4010
rect 18570 4002 19298 4008
rect 18470 3672 18534 3680
rect 18470 3620 18476 3672
rect 18528 3620 18534 3672
rect 18470 3612 18534 3620
rect 18230 3584 18296 3590
rect 18230 3532 18238 3584
rect 18290 3554 18296 3584
rect 18470 3554 18498 3612
rect 18290 3532 18498 3554
rect 18230 3526 18498 3532
rect 18570 3376 18598 4002
rect 19298 3936 19364 3942
rect 19298 3884 19306 3936
rect 19358 3884 19364 3936
rect 19298 3878 19364 3884
rect 19298 3756 19326 3878
rect 19258 3728 19326 3756
rect 18570 3368 18882 3376
rect 18570 3340 18821 3368
rect 18230 3152 18306 3158
rect 18230 3126 18238 3152
rect 18138 3100 18238 3126
rect 18290 3100 18306 3152
rect 18138 3098 18306 3100
rect 18230 3094 18306 3098
rect 17910 2958 17976 2964
rect 17910 2906 17918 2958
rect 17970 2936 17976 2958
rect 18570 2936 18598 3340
rect 18802 3316 18821 3340
rect 18873 3316 18882 3368
rect 18802 3304 18882 3316
rect 19118 3372 19186 3378
rect 19118 3320 19125 3372
rect 19177 3320 19186 3372
rect 19118 3314 19186 3320
rect 17970 2908 18598 2936
rect 17970 2906 17976 2908
rect 17910 2900 17976 2906
rect 18724 2708 19074 2722
rect 16836 2578 17186 2592
rect 18724 2592 18745 2708
rect 19053 2592 19074 2708
rect 19118 2698 19162 3314
rect 19258 3144 19286 3728
rect 19320 3678 19382 3684
rect 19320 3626 19330 3678
rect 19418 3670 19446 4242
rect 19474 4069 19538 4076
rect 19474 4017 19480 4069
rect 19532 4036 19538 4069
rect 19800 4036 19850 4426
rect 20322 4424 20350 4524
rect 20322 4418 20388 4424
rect 21436 4422 21464 4528
rect 21672 4486 21738 4494
rect 21672 4434 21678 4486
rect 21730 4434 21738 4486
rect 21672 4426 21738 4434
rect 20322 4404 20330 4418
rect 20324 4366 20330 4404
rect 20382 4366 20388 4418
rect 20324 4360 20388 4366
rect 21396 4416 21464 4422
rect 21396 4364 21406 4416
rect 21458 4364 21464 4416
rect 21396 4358 21464 4364
rect 20236 4302 20300 4308
rect 20236 4272 20242 4302
rect 20026 4250 20242 4272
rect 20294 4250 20300 4302
rect 20026 4244 20300 4250
rect 21306 4304 21374 4310
rect 21306 4252 21314 4304
rect 21366 4252 21374 4304
rect 19532 4020 19852 4036
rect 19532 4017 19866 4020
rect 19474 4014 19866 4017
rect 19474 4008 19808 4014
rect 19800 3962 19808 4008
rect 19860 3962 19866 4014
rect 19800 3956 19866 3962
rect 19670 3820 19742 3832
rect 19670 3768 19680 3820
rect 19732 3768 19742 3820
rect 19670 3756 19742 3768
rect 19706 3754 19742 3756
rect 19418 3642 19706 3670
rect 19320 3620 19382 3626
rect 19354 3574 19382 3620
rect 19354 3570 19598 3574
rect 19354 3564 19636 3570
rect 19354 3546 19576 3564
rect 19570 3512 19576 3546
rect 19628 3512 19636 3564
rect 19570 3504 19636 3512
rect 19258 3130 19322 3144
rect 19678 3136 19706 3642
rect 19782 3430 19848 3438
rect 19782 3378 19788 3430
rect 19840 3378 19848 3430
rect 19782 3370 19848 3378
rect 19258 3078 19261 3130
rect 19313 3078 19322 3130
rect 19258 3062 19322 3078
rect 19492 3120 19706 3136
rect 19492 3068 19493 3120
rect 19545 3108 19706 3120
rect 19545 3068 19546 3108
rect 19492 3052 19546 3068
rect 19798 2964 19848 3370
rect 20026 3126 20054 4244
rect 21306 4242 21374 4252
rect 21186 4069 21250 4076
rect 21186 4038 21192 4069
rect 20458 4017 21192 4038
rect 21244 4017 21250 4069
rect 20458 4010 21250 4017
rect 20458 4008 21192 4010
rect 20458 4002 21186 4008
rect 20358 3672 20422 3680
rect 20358 3620 20364 3672
rect 20416 3620 20422 3672
rect 20358 3612 20422 3620
rect 20118 3584 20184 3590
rect 20118 3532 20126 3584
rect 20178 3554 20184 3584
rect 20358 3554 20386 3612
rect 20178 3532 20386 3554
rect 20118 3526 20386 3532
rect 20458 3376 20486 4002
rect 21186 3936 21252 3942
rect 21186 3884 21194 3936
rect 21246 3884 21252 3936
rect 21186 3878 21252 3884
rect 21186 3756 21214 3878
rect 21146 3728 21214 3756
rect 20458 3368 20770 3376
rect 20458 3340 20709 3368
rect 20118 3152 20194 3158
rect 20118 3126 20126 3152
rect 20026 3100 20126 3126
rect 20178 3100 20194 3152
rect 20026 3098 20194 3100
rect 20118 3094 20194 3098
rect 19798 2958 19864 2964
rect 19798 2906 19806 2958
rect 19858 2936 19864 2958
rect 20458 2936 20486 3340
rect 20690 3316 20709 3340
rect 20761 3316 20770 3368
rect 20690 3304 20770 3316
rect 21006 3372 21074 3378
rect 21006 3320 21013 3372
rect 21065 3320 21074 3372
rect 21006 3314 21074 3320
rect 19858 2908 20486 2936
rect 19858 2906 19864 2908
rect 19798 2900 19864 2906
rect 20612 2708 20962 2722
rect 18724 2578 19074 2592
rect 20612 2592 20633 2708
rect 20941 2592 20962 2708
rect 21006 2698 21050 3314
rect 21146 3144 21174 3728
rect 21208 3678 21270 3684
rect 21208 3626 21218 3678
rect 21306 3670 21334 4242
rect 21362 4069 21426 4076
rect 21362 4017 21368 4069
rect 21420 4036 21426 4069
rect 21688 4036 21738 4426
rect 22210 4424 22238 4528
rect 22210 4418 22276 4424
rect 23324 4422 23352 4528
rect 23560 4486 23626 4494
rect 23560 4434 23566 4486
rect 23618 4434 23626 4486
rect 23560 4426 23626 4434
rect 22210 4404 22218 4418
rect 22212 4366 22218 4404
rect 22270 4366 22276 4418
rect 22212 4360 22276 4366
rect 23284 4416 23352 4422
rect 23284 4364 23294 4416
rect 23346 4364 23352 4416
rect 23284 4358 23352 4364
rect 22124 4302 22188 4308
rect 22124 4272 22130 4302
rect 21914 4250 22130 4272
rect 22182 4250 22188 4302
rect 21914 4244 22188 4250
rect 23194 4304 23262 4310
rect 23194 4252 23202 4304
rect 23254 4252 23262 4304
rect 21420 4020 21740 4036
rect 21420 4017 21754 4020
rect 21362 4014 21754 4017
rect 21362 4008 21696 4014
rect 21688 3962 21696 4008
rect 21748 3962 21754 4014
rect 21688 3956 21754 3962
rect 21558 3820 21630 3832
rect 21558 3768 21568 3820
rect 21620 3768 21630 3820
rect 21558 3756 21630 3768
rect 21594 3754 21630 3756
rect 21306 3642 21594 3670
rect 21208 3620 21270 3626
rect 21242 3574 21270 3620
rect 21242 3570 21486 3574
rect 21242 3564 21524 3570
rect 21242 3546 21464 3564
rect 21458 3512 21464 3546
rect 21516 3512 21524 3564
rect 21458 3504 21524 3512
rect 21146 3130 21210 3144
rect 21566 3136 21594 3642
rect 21670 3430 21736 3438
rect 21670 3378 21676 3430
rect 21728 3378 21736 3430
rect 21670 3370 21736 3378
rect 21146 3078 21149 3130
rect 21201 3078 21210 3130
rect 21146 3062 21210 3078
rect 21380 3120 21594 3136
rect 21380 3068 21381 3120
rect 21433 3108 21594 3120
rect 21433 3068 21434 3108
rect 21380 3052 21434 3068
rect 21686 2964 21736 3370
rect 21914 3126 21942 4244
rect 23194 4242 23262 4252
rect 23074 4069 23138 4076
rect 23074 4038 23080 4069
rect 22346 4017 23080 4038
rect 23132 4017 23138 4069
rect 22346 4010 23138 4017
rect 22346 4008 23080 4010
rect 22346 4002 23074 4008
rect 22246 3672 22310 3680
rect 22246 3620 22252 3672
rect 22304 3620 22310 3672
rect 22246 3612 22310 3620
rect 22006 3584 22072 3590
rect 22006 3532 22014 3584
rect 22066 3554 22072 3584
rect 22246 3554 22274 3612
rect 22066 3532 22274 3554
rect 22006 3526 22274 3532
rect 22346 3376 22374 4002
rect 23074 3936 23140 3942
rect 23074 3884 23082 3936
rect 23134 3884 23140 3936
rect 23074 3878 23140 3884
rect 23074 3756 23102 3878
rect 23034 3728 23102 3756
rect 22346 3368 22658 3376
rect 22346 3340 22597 3368
rect 22006 3152 22082 3158
rect 22006 3126 22014 3152
rect 21914 3100 22014 3126
rect 22066 3100 22082 3152
rect 21914 3098 22082 3100
rect 22006 3094 22082 3098
rect 21686 2958 21752 2964
rect 21686 2906 21694 2958
rect 21746 2936 21752 2958
rect 22346 2936 22374 3340
rect 22578 3316 22597 3340
rect 22649 3316 22658 3368
rect 22578 3304 22658 3316
rect 22894 3372 22962 3378
rect 22894 3320 22901 3372
rect 22953 3320 22962 3372
rect 22894 3314 22962 3320
rect 21746 2908 22374 2936
rect 21746 2906 21752 2908
rect 21686 2900 21752 2906
rect 22500 2708 22850 2722
rect 20612 2578 20962 2592
rect 22500 2592 22521 2708
rect 22829 2592 22850 2708
rect 22894 2698 22938 3314
rect 23034 3144 23062 3728
rect 23096 3678 23158 3684
rect 23096 3626 23106 3678
rect 23194 3670 23222 4242
rect 23250 4069 23314 4076
rect 23250 4017 23256 4069
rect 23308 4036 23314 4069
rect 23576 4036 23626 4426
rect 24098 4424 24126 4528
rect 24098 4418 24164 4424
rect 25212 4422 25240 4528
rect 25448 4486 25514 4494
rect 25448 4434 25454 4486
rect 25506 4434 25514 4486
rect 25448 4426 25514 4434
rect 24098 4404 24106 4418
rect 24100 4366 24106 4404
rect 24158 4366 24164 4418
rect 24100 4360 24164 4366
rect 25172 4416 25240 4422
rect 25172 4364 25182 4416
rect 25234 4364 25240 4416
rect 25172 4358 25240 4364
rect 24012 4302 24076 4308
rect 24012 4272 24018 4302
rect 23802 4250 24018 4272
rect 24070 4250 24076 4302
rect 23802 4244 24076 4250
rect 25082 4304 25150 4310
rect 25082 4252 25090 4304
rect 25142 4252 25150 4304
rect 23308 4020 23628 4036
rect 23308 4017 23642 4020
rect 23250 4014 23642 4017
rect 23250 4008 23584 4014
rect 23576 3962 23584 4008
rect 23636 3962 23642 4014
rect 23576 3956 23642 3962
rect 23446 3820 23518 3832
rect 23446 3768 23456 3820
rect 23508 3768 23518 3820
rect 23446 3756 23518 3768
rect 23482 3754 23518 3756
rect 23194 3642 23482 3670
rect 23096 3620 23158 3626
rect 23130 3574 23158 3620
rect 23130 3570 23374 3574
rect 23130 3564 23412 3570
rect 23130 3546 23352 3564
rect 23346 3512 23352 3546
rect 23404 3512 23412 3564
rect 23346 3504 23412 3512
rect 23034 3130 23098 3144
rect 23454 3136 23482 3642
rect 23558 3430 23624 3438
rect 23558 3378 23564 3430
rect 23616 3378 23624 3430
rect 23558 3370 23624 3378
rect 23034 3078 23037 3130
rect 23089 3078 23098 3130
rect 23034 3062 23098 3078
rect 23268 3120 23482 3136
rect 23268 3068 23269 3120
rect 23321 3108 23482 3120
rect 23321 3068 23322 3108
rect 23268 3052 23322 3068
rect 23574 2964 23624 3370
rect 23802 3126 23830 4244
rect 25082 4242 25150 4252
rect 24962 4069 25026 4076
rect 24962 4038 24968 4069
rect 24234 4017 24968 4038
rect 25020 4017 25026 4069
rect 24234 4010 25026 4017
rect 24234 4008 24968 4010
rect 24234 4002 24962 4008
rect 24134 3672 24198 3680
rect 24134 3620 24140 3672
rect 24192 3620 24198 3672
rect 24134 3612 24198 3620
rect 23894 3584 23960 3590
rect 23894 3532 23902 3584
rect 23954 3554 23960 3584
rect 24134 3554 24162 3612
rect 23954 3532 24162 3554
rect 23894 3526 24162 3532
rect 24234 3376 24262 4002
rect 24962 3936 25028 3942
rect 24962 3884 24970 3936
rect 25022 3884 25028 3936
rect 24962 3878 25028 3884
rect 24962 3756 24990 3878
rect 24922 3728 24990 3756
rect 24234 3368 24546 3376
rect 24234 3340 24485 3368
rect 23894 3152 23970 3158
rect 23894 3126 23902 3152
rect 23802 3100 23902 3126
rect 23954 3100 23970 3152
rect 23802 3098 23970 3100
rect 23894 3094 23970 3098
rect 23574 2958 23640 2964
rect 23574 2906 23582 2958
rect 23634 2936 23640 2958
rect 24234 2936 24262 3340
rect 24466 3316 24485 3340
rect 24537 3316 24546 3368
rect 24466 3304 24546 3316
rect 24782 3372 24850 3378
rect 24782 3320 24789 3372
rect 24841 3320 24850 3372
rect 24782 3314 24850 3320
rect 23634 2908 24262 2936
rect 23634 2906 23640 2908
rect 23574 2900 23640 2906
rect 24388 2708 24738 2722
rect 22500 2578 22850 2592
rect 24388 2592 24409 2708
rect 24717 2592 24738 2708
rect 24782 2698 24826 3314
rect 24922 3144 24950 3728
rect 24984 3678 25046 3684
rect 24984 3626 24994 3678
rect 25082 3670 25110 4242
rect 25138 4069 25202 4076
rect 25138 4017 25144 4069
rect 25196 4036 25202 4069
rect 25464 4036 25514 4426
rect 25986 4424 26014 4528
rect 25986 4418 26052 4424
rect 25986 4404 25994 4418
rect 25988 4366 25994 4404
rect 26046 4366 26052 4418
rect 25988 4360 26052 4366
rect 25900 4302 25964 4308
rect 25900 4272 25906 4302
rect 25690 4250 25906 4272
rect 25958 4250 25964 4302
rect 25690 4244 25964 4250
rect 25196 4020 25516 4036
rect 25196 4017 25530 4020
rect 25138 4014 25530 4017
rect 25138 4008 25472 4014
rect 25464 3962 25472 4008
rect 25524 3962 25530 4014
rect 25464 3956 25530 3962
rect 25334 3820 25406 3832
rect 25334 3768 25344 3820
rect 25396 3768 25406 3820
rect 25334 3756 25406 3768
rect 25370 3754 25406 3756
rect 25082 3642 25370 3670
rect 24984 3620 25046 3626
rect 25018 3574 25046 3620
rect 25018 3570 25262 3574
rect 25018 3564 25300 3570
rect 25018 3546 25240 3564
rect 25234 3512 25240 3546
rect 25292 3512 25300 3564
rect 25234 3504 25300 3512
rect 24922 3130 24986 3144
rect 25342 3136 25370 3642
rect 25446 3430 25512 3438
rect 25446 3378 25452 3430
rect 25504 3378 25512 3430
rect 25446 3370 25512 3378
rect 24922 3078 24925 3130
rect 24977 3078 24986 3130
rect 24922 3062 24986 3078
rect 25156 3120 25370 3136
rect 25156 3068 25157 3120
rect 25209 3108 25370 3120
rect 25209 3068 25210 3108
rect 25156 3052 25210 3068
rect 25462 2964 25512 3370
rect 25690 3126 25718 4244
rect 26122 4002 26658 4038
rect 26022 3672 26086 3680
rect 26022 3620 26028 3672
rect 26080 3620 26086 3672
rect 26022 3612 26086 3620
rect 25782 3584 25848 3590
rect 25782 3532 25790 3584
rect 25842 3554 25848 3584
rect 26022 3554 26050 3612
rect 25842 3532 26050 3554
rect 25782 3526 26050 3532
rect 26122 3376 26150 4002
rect 26122 3368 26434 3376
rect 26122 3340 26373 3368
rect 25782 3152 25858 3158
rect 25782 3126 25790 3152
rect 25690 3100 25790 3126
rect 25842 3100 25858 3152
rect 25690 3098 25858 3100
rect 25782 3094 25858 3098
rect 25462 2958 25528 2964
rect 25462 2906 25470 2958
rect 25522 2936 25528 2958
rect 26122 2936 26150 3340
rect 26354 3316 26373 3340
rect 26425 3316 26434 3368
rect 26354 3304 26434 3316
rect 25522 2908 26150 2936
rect 25522 2906 25528 2908
rect 25462 2900 25528 2906
rect 26276 2708 26626 2722
rect 24388 2578 24738 2592
rect 26276 2592 26297 2708
rect 26605 2592 26626 2708
rect 26276 2578 26626 2592
<< via2 >>
rect 4610 5290 4683 5343
rect 19740 5343 19807 5349
rect 19740 5296 19780 5343
rect 19780 5296 19807 5343
rect -2011 4746 -1955 4802
rect -1931 4746 -1875 4802
rect -1851 4746 -1795 4802
rect -1771 4746 -1715 4802
rect -123 4746 -67 4802
rect -43 4746 13 4802
rect 37 4746 93 4802
rect 117 4746 173 4802
rect 1765 4746 1821 4802
rect 1845 4746 1901 4802
rect 1925 4746 1981 4802
rect 2005 4746 2061 4802
rect 3653 4746 3709 4802
rect 3733 4746 3789 4802
rect 3813 4746 3869 4802
rect 3893 4746 3949 4802
rect 5541 4746 5597 4802
rect 5621 4746 5677 4802
rect 5701 4746 5757 4802
rect 5781 4746 5837 4802
rect 7429 4746 7485 4802
rect 7509 4746 7565 4802
rect 7589 4746 7645 4802
rect 7669 4746 7725 4802
rect 9317 4746 9373 4802
rect 9397 4746 9453 4802
rect 9477 4746 9533 4802
rect 9557 4746 9613 4802
rect 11205 4746 11261 4802
rect 11285 4746 11341 4802
rect 11365 4746 11421 4802
rect 11445 4746 11501 4802
rect 13087 4746 13143 4802
rect 13167 4746 13223 4802
rect 13247 4746 13303 4802
rect 13327 4746 13383 4802
rect 14975 4746 15031 4802
rect 15055 4746 15111 4802
rect 15135 4746 15191 4802
rect 15215 4746 15271 4802
rect 16863 4746 16919 4802
rect 16943 4746 16999 4802
rect 17023 4746 17079 4802
rect 17103 4746 17159 4802
rect 18751 4746 18807 4802
rect 18831 4746 18887 4802
rect 18911 4746 18967 4802
rect 18991 4746 19047 4802
rect 20639 4746 20695 4802
rect 20719 4746 20775 4802
rect 20799 4746 20855 4802
rect 20879 4746 20935 4802
rect 22527 4746 22583 4802
rect 22607 4746 22663 4802
rect 22687 4746 22743 4802
rect 22767 4746 22823 4802
rect 24415 4746 24471 4802
rect 24495 4746 24551 4802
rect 24575 4746 24631 4802
rect 24655 4746 24711 4802
rect 26303 4746 26359 4802
rect 26383 4746 26439 4802
rect 26463 4746 26519 4802
rect 26543 4746 26599 4802
rect -2011 2622 -1955 2678
rect -1931 2622 -1875 2678
rect -1851 2622 -1795 2678
rect -1771 2622 -1715 2678
rect -123 2622 -67 2678
rect -43 2622 13 2678
rect 37 2622 93 2678
rect 117 2622 173 2678
rect 1765 2622 1821 2678
rect 1845 2622 1901 2678
rect 1925 2622 1981 2678
rect 2005 2622 2061 2678
rect 3653 2622 3709 2678
rect 3733 2622 3789 2678
rect 3813 2622 3869 2678
rect 3893 2622 3949 2678
rect 5541 2622 5597 2678
rect 5621 2622 5677 2678
rect 5701 2622 5757 2678
rect 5781 2622 5837 2678
rect 7429 2622 7485 2678
rect 7509 2622 7565 2678
rect 7589 2622 7645 2678
rect 7669 2622 7725 2678
rect 9317 2622 9373 2678
rect 9397 2622 9453 2678
rect 9477 2622 9533 2678
rect 9557 2622 9613 2678
rect 11205 2622 11261 2678
rect 11285 2622 11341 2678
rect 11365 2622 11421 2678
rect 11445 2622 11501 2678
rect 13087 2622 13143 2678
rect 13167 2622 13223 2678
rect 13247 2622 13303 2678
rect 13327 2622 13383 2678
rect 14975 2622 15031 2678
rect 15055 2622 15111 2678
rect 15135 2622 15191 2678
rect 15215 2622 15271 2678
rect 16863 2622 16919 2678
rect 16943 2622 16999 2678
rect 17023 2622 17079 2678
rect 17103 2622 17159 2678
rect 18751 2622 18807 2678
rect 18831 2622 18887 2678
rect 18911 2622 18967 2678
rect 18991 2622 19047 2678
rect 20639 2622 20695 2678
rect 20719 2622 20775 2678
rect 20799 2622 20855 2678
rect 20879 2622 20935 2678
rect 22527 2622 22583 2678
rect 22607 2622 22663 2678
rect 22687 2622 22743 2678
rect 22767 2622 22823 2678
rect 24415 2622 24471 2678
rect 24495 2622 24551 2678
rect 24575 2622 24631 2678
rect 24655 2622 24711 2678
rect 26303 2622 26359 2678
rect 26383 2622 26439 2678
rect 26463 2622 26519 2678
rect 26543 2622 26599 2678
<< metal3 >>
rect 4475 5343 4844 5373
rect 4475 5290 4610 5343
rect 4683 5290 4844 5343
rect 4475 5272 4844 5290
rect 19618 5349 19894 5374
rect 19618 5347 19740 5349
rect 19618 5291 19739 5347
rect 19807 5296 19894 5349
rect 19799 5291 19894 5296
rect 19618 5270 19894 5291
rect -3552 4802 26658 4904
rect -3552 4746 -2011 4802
rect -1955 4746 -1931 4802
rect -1875 4746 -1851 4802
rect -1795 4746 -1771 4802
rect -1715 4746 -123 4802
rect -67 4746 -43 4802
rect 13 4746 37 4802
rect 93 4746 117 4802
rect 173 4746 1765 4802
rect 1821 4746 1845 4802
rect 1901 4746 1925 4802
rect 1981 4746 2005 4802
rect 2061 4746 3653 4802
rect 3709 4746 3733 4802
rect 3789 4746 3813 4802
rect 3869 4746 3893 4802
rect 3949 4746 5541 4802
rect 5597 4746 5621 4802
rect 5677 4746 5701 4802
rect 5757 4746 5781 4802
rect 5837 4746 7429 4802
rect 7485 4746 7509 4802
rect 7565 4746 7589 4802
rect 7645 4746 7669 4802
rect 7725 4746 9317 4802
rect 9373 4746 9397 4802
rect 9453 4746 9477 4802
rect 9533 4746 9557 4802
rect 9613 4746 11205 4802
rect 11261 4746 11285 4802
rect 11341 4746 11365 4802
rect 11421 4746 11445 4802
rect 11501 4746 13087 4802
rect 13143 4746 13167 4802
rect 13223 4746 13247 4802
rect 13303 4746 13327 4802
rect 13383 4746 14975 4802
rect 15031 4746 15055 4802
rect 15111 4746 15135 4802
rect 15191 4746 15215 4802
rect 15271 4746 16863 4802
rect 16919 4746 16943 4802
rect 16999 4746 17023 4802
rect 17079 4746 17103 4802
rect 17159 4746 18751 4802
rect 18807 4746 18831 4802
rect 18887 4746 18911 4802
rect 18967 4746 18991 4802
rect 19047 4746 20639 4802
rect 20695 4746 20719 4802
rect 20775 4746 20799 4802
rect 20855 4746 20879 4802
rect 20935 4746 22527 4802
rect 22583 4746 22607 4802
rect 22663 4746 22687 4802
rect 22743 4746 22767 4802
rect 22823 4746 24415 4802
rect 24471 4746 24495 4802
rect 24551 4746 24575 4802
rect 24631 4746 24655 4802
rect 24711 4746 26303 4802
rect 26359 4746 26383 4802
rect 26439 4746 26463 4802
rect 26519 4746 26543 4802
rect 26599 4746 26658 4802
rect -3552 4650 26658 4746
rect -3544 2678 26658 2782
rect -3544 2622 -2011 2678
rect -1955 2622 -1931 2678
rect -1875 2622 -1851 2678
rect -1795 2622 -1771 2678
rect -1715 2622 -123 2678
rect -67 2622 -43 2678
rect 13 2622 37 2678
rect 93 2622 117 2678
rect 173 2622 1765 2678
rect 1821 2622 1845 2678
rect 1901 2622 1925 2678
rect 1981 2622 2005 2678
rect 2061 2622 3653 2678
rect 3709 2622 3733 2678
rect 3789 2622 3813 2678
rect 3869 2622 3893 2678
rect 3949 2653 5541 2678
rect 3949 2622 4606 2653
rect -3544 2570 4606 2622
rect 4673 2622 5541 2653
rect 5597 2622 5621 2678
rect 5677 2622 5701 2678
rect 5757 2622 5781 2678
rect 5837 2622 7429 2678
rect 7485 2622 7509 2678
rect 7565 2622 7589 2678
rect 7645 2622 7669 2678
rect 7725 2622 9317 2678
rect 9373 2622 9397 2678
rect 9453 2622 9477 2678
rect 9533 2622 9557 2678
rect 9613 2622 11205 2678
rect 11261 2622 11285 2678
rect 11341 2622 11365 2678
rect 11421 2622 11445 2678
rect 11501 2622 13087 2678
rect 13143 2622 13167 2678
rect 13223 2622 13247 2678
rect 13303 2622 13327 2678
rect 13383 2622 14975 2678
rect 15031 2622 15055 2678
rect 15111 2622 15135 2678
rect 15191 2622 15215 2678
rect 15271 2622 16863 2678
rect 16919 2622 16943 2678
rect 16999 2622 17023 2678
rect 17079 2622 17103 2678
rect 17159 2622 18751 2678
rect 18807 2622 18831 2678
rect 18887 2622 18911 2678
rect 18967 2622 18991 2678
rect 19047 2656 20639 2678
rect 19047 2622 19699 2656
rect 4673 2572 19699 2622
rect 19780 2622 20639 2656
rect 20695 2622 20719 2678
rect 20775 2622 20799 2678
rect 20855 2622 20879 2678
rect 20935 2622 22527 2678
rect 22583 2622 22607 2678
rect 22663 2622 22687 2678
rect 22743 2622 22767 2678
rect 22823 2622 24415 2678
rect 24471 2622 24495 2678
rect 24551 2622 24575 2678
rect 24631 2622 24655 2678
rect 24711 2622 26303 2678
rect 26359 2622 26383 2678
rect 26439 2622 26463 2678
rect 26519 2622 26543 2678
rect 26599 2622 26658 2678
rect 19780 2572 26658 2622
rect 4673 2570 26658 2572
rect -3544 2528 26658 2570
rect -3544 2527 9672 2528
rect 11554 2527 24770 2528
<< via3 >>
rect 4610 5290 4683 5343
rect 19739 5296 19740 5347
rect 19740 5296 19799 5347
rect 19739 5291 19799 5296
rect 4606 2570 4673 2653
rect 19699 2572 19780 2656
<< metal4 >>
rect 4486 5343 4812 5412
rect 4486 5290 4610 5343
rect 4683 5290 4812 5343
rect 4486 2653 4812 5290
rect 4486 2570 4606 2653
rect 4673 2570 4812 2653
rect 4486 2535 4812 2570
rect 19628 5347 19893 5374
rect 19628 5291 19739 5347
rect 19799 5291 19893 5347
rect 19628 2656 19893 5291
rect 19628 2572 19699 2656
rect 19780 2572 19893 2656
rect 19628 2507 19893 2572
<< labels >>
flabel metal1 3688 5062 3894 5220 1 FreeSans 400 0 0 0 RESET1
port 4 n
flabel metal1 18800 5062 18998 5222 1 FreeSans 800 0 0 0 RESET2
port 5 n
flabel metal3 -3552 4650 -2011 4904 1 FreeSans 800 0 0 0 VDD
port 1 n
flabel metal2 -3544 4002 -3352 4038 1 FreeSans 800 0 0 0 IN
port 6 n
flabel metal1 26631 3308 26744 3386 1 FreeSans 400 0 0 0 OUT
port 3 n
flabel metal3 -3544 2527 -2011 2782 1 FreeSans 800 0 0 0 VSS
port 2 n
<< end >>
