magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< pwell >>
rect 10 10 806 146
<< nmoslvt >>
rect 92 36 122 120
rect 178 36 208 120
rect 264 36 294 120
rect 350 36 380 120
rect 436 36 466 120
rect 522 36 552 120
rect 608 36 638 120
rect 694 36 724 120
<< ndiff >>
rect 36 101 92 120
rect 36 67 47 101
rect 81 67 92 101
rect 36 36 92 67
rect 122 101 178 120
rect 122 67 133 101
rect 167 67 178 101
rect 122 36 178 67
rect 208 101 264 120
rect 208 67 219 101
rect 253 67 264 101
rect 208 36 264 67
rect 294 101 350 120
rect 294 67 305 101
rect 339 67 350 101
rect 294 36 350 67
rect 380 101 436 120
rect 380 67 391 101
rect 425 67 436 101
rect 380 36 436 67
rect 466 101 522 120
rect 466 67 477 101
rect 511 67 522 101
rect 466 36 522 67
rect 552 101 608 120
rect 552 67 563 101
rect 597 67 608 101
rect 552 36 608 67
rect 638 101 694 120
rect 638 67 649 101
rect 683 67 694 101
rect 638 36 694 67
rect 724 101 780 120
rect 724 67 735 101
rect 769 67 780 101
rect 724 36 780 67
<< ndiffc >>
rect 47 67 81 101
rect 133 67 167 101
rect 219 67 253 101
rect 305 67 339 101
rect 391 67 425 101
rect 477 67 511 101
rect 563 67 597 101
rect 649 67 683 101
rect 735 67 769 101
<< poly >>
rect 92 201 724 217
rect 92 167 153 201
rect 187 167 221 201
rect 255 167 289 201
rect 323 167 357 201
rect 391 167 425 201
rect 459 167 493 201
rect 527 167 561 201
rect 595 167 629 201
rect 663 167 724 201
rect 92 146 724 167
rect 92 120 122 146
rect 178 120 208 146
rect 264 120 294 146
rect 350 120 380 146
rect 436 120 466 146
rect 522 120 552 146
rect 608 120 638 146
rect 694 120 724 146
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
rect 436 10 466 36
rect 522 10 552 36
rect 608 10 638 36
rect 694 10 724 36
<< polycont >>
rect 153 167 187 201
rect 221 167 255 201
rect 289 167 323 201
rect 357 167 391 201
rect 425 167 459 201
rect 493 167 527 201
rect 561 167 595 201
rect 629 167 663 201
<< locali >>
rect 137 201 679 217
rect 137 167 139 201
rect 187 167 211 201
rect 255 167 283 201
rect 323 167 355 201
rect 391 167 425 201
rect 461 167 493 201
rect 533 167 561 201
rect 605 167 629 201
rect 677 167 679 201
rect 137 151 679 167
rect 47 101 81 117
rect 47 51 81 67
rect 133 101 167 117
rect 133 51 167 67
rect 219 101 253 117
rect 219 51 253 67
rect 305 101 339 117
rect 305 51 339 67
rect 391 101 425 117
rect 391 51 425 67
rect 477 101 511 117
rect 477 51 511 67
rect 563 101 597 117
rect 563 51 597 67
rect 649 101 683 117
rect 649 51 683 67
rect 735 101 769 117
rect 735 51 769 67
<< viali >>
rect 139 167 153 201
rect 153 167 173 201
rect 211 167 221 201
rect 221 167 245 201
rect 283 167 289 201
rect 289 167 317 201
rect 355 167 357 201
rect 357 167 389 201
rect 427 167 459 201
rect 459 167 461 201
rect 499 167 527 201
rect 527 167 533 201
rect 571 167 595 201
rect 595 167 605 201
rect 643 167 663 201
rect 663 167 677 201
rect 47 67 81 101
rect 133 67 167 101
rect 219 67 253 101
rect 305 67 339 101
rect 391 67 425 101
rect 477 67 511 101
rect 563 67 597 101
rect 649 67 683 101
rect 735 67 769 101
<< metal1 >>
rect 127 201 689 213
rect 127 167 139 201
rect 173 167 211 201
rect 245 167 283 201
rect 317 167 355 201
rect 389 167 427 201
rect 461 167 499 201
rect 533 167 571 201
rect 605 167 643 201
rect 677 167 689 201
rect 127 155 689 167
rect 41 101 87 118
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 124 110 176 118
rect 124 51 176 58
rect 213 101 259 118
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 296 110 348 118
rect 296 51 348 58
rect 385 101 431 118
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 468 110 520 118
rect 468 51 520 58
rect 557 101 603 118
rect 557 67 563 101
rect 597 67 603 101
rect 557 -29 603 67
rect 640 110 692 118
rect 640 51 692 58
rect 729 101 775 118
rect 729 67 735 101
rect 769 67 775 101
rect 729 -29 775 67
rect 41 -89 775 -29
<< via1 >>
rect 124 101 176 110
rect 124 67 133 101
rect 133 67 167 101
rect 167 67 176 101
rect 124 58 176 67
rect 296 101 348 110
rect 296 67 305 101
rect 305 67 339 101
rect 339 67 348 101
rect 296 58 348 67
rect 468 101 520 110
rect 468 67 477 101
rect 477 67 511 101
rect 511 67 520 101
rect 468 58 520 67
rect 640 101 692 110
rect 640 67 649 101
rect 649 67 683 101
rect 683 67 692 101
rect 640 58 692 67
<< metal2 >>
rect 117 110 183 118
rect 117 106 124 110
rect 176 106 183 110
rect 117 50 122 106
rect 178 50 183 106
rect 117 34 183 50
rect 289 110 355 118
rect 289 106 296 110
rect 348 106 355 110
rect 289 50 294 106
rect 350 50 355 106
rect 289 34 355 50
rect 461 110 527 118
rect 461 106 468 110
rect 520 106 527 110
rect 461 50 466 106
rect 522 50 527 106
rect 461 34 527 50
rect 633 110 699 118
rect 633 106 640 110
rect 692 106 699 110
rect 633 50 638 106
rect 694 50 699 106
rect 633 34 699 50
<< via2 >>
rect 122 58 124 106
rect 124 58 176 106
rect 176 58 178 106
rect 122 50 178 58
rect 294 58 296 106
rect 296 58 348 106
rect 348 58 350 106
rect 294 50 350 58
rect 466 58 468 106
rect 468 58 520 106
rect 520 58 522 106
rect 466 50 522 58
rect 638 58 640 106
rect 640 58 692 106
rect 692 58 694 106
rect 638 50 694 58
<< metal3 >>
rect 117 106 699 111
rect 117 50 122 106
rect 178 50 294 106
rect 350 50 466 106
rect 522 50 638 106
rect 694 50 699 106
rect 117 45 699 50
<< labels >>
flabel metal3 s 117 45 699 111 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 41 -89 775 -29 0 FreeSans 400 0 0 0 SOURCE
port 2 nsew
flabel metal1 s 127 155 689 213 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel pwell s 80 125 91 139 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 5952358
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5942344
string path 1.600 2.950 1.600 -2.225 
<< end >>
