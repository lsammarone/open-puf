//-----------------------------------------------------------------------------
// BR64 - Bistable Ring PUF 64-bit 
//-----------------------------------------------------------------------------
// dump-vcd: False
// verilator-xinit: zeros
module NBR64 
(
  input wire RESET,
  input wire [63:0] C,
  output wire OUT
);
  supply1 VDD;
  supply0 VSS;
  // empty module
  // see lib file
  
endmodule
