magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< poly >>
rect -3 8942 157 8958
rect -3 8908 26 8942
rect 60 8908 94 8942
rect 128 8908 157 8942
rect -260 8806 -100 8822
rect -260 8772 -231 8806
rect -197 8772 -163 8806
rect -129 8772 -100 8806
rect -3 7674 26 7708
rect 60 7674 94 7708
rect 128 7674 157 7708
rect -3 7658 157 7674
rect -260 6338 -231 6372
rect -197 6338 -163 6372
rect -129 6338 -100 6372
rect -260 6322 -100 6338
rect -3 7600 157 7616
rect -3 7566 26 7600
rect 60 7566 94 7600
rect 128 7566 157 7600
rect -3 6332 26 6366
rect 60 6332 94 6366
rect 128 6332 157 6366
rect -3 6316 157 6332
rect -258 6080 -98 6096
rect -258 6046 -229 6080
rect -195 6046 -161 6080
rect -127 6046 -98 6080
rect -2 6080 158 6096
rect -2 6046 27 6080
rect 61 6046 95 6080
rect 129 6046 158 6080
<< polycont >>
rect 26 8908 60 8942
rect 94 8908 128 8942
rect -231 8772 -197 8806
rect -163 8772 -129 8806
rect 26 7674 60 7708
rect 94 7674 128 7708
rect -231 6338 -197 6372
rect -163 6338 -129 6372
rect 26 7566 60 7600
rect 94 7566 128 7600
rect 26 6332 60 6366
rect 94 6332 128 6366
rect -229 6046 -195 6080
rect -161 6046 -127 6080
rect 27 6046 61 6080
rect 95 6046 129 6080
<< npolyres >>
rect -260 6372 -100 8772
rect -3 7708 157 8908
rect -3 6366 157 7566
rect -258 1174 -98 6046
rect -2 1174 158 6046
rect -258 1014 158 1174
<< locali >>
rect 10 8908 26 8942
rect 60 8908 94 8942
rect 128 8908 144 8942
rect -247 8772 -231 8806
rect -197 8772 -163 8806
rect -129 8772 -113 8806
rect 10 7674 26 7708
rect 60 7674 94 7708
rect 128 7674 144 7708
rect 10 7566 26 7600
rect 60 7566 94 7600
rect 128 7566 144 7600
rect -247 6338 -231 6372
rect -195 6338 -163 6372
rect -123 6338 -113 6372
rect 10 6332 26 6366
rect 60 6332 94 6366
rect 128 6332 144 6366
rect -245 6046 -229 6080
rect -195 6046 -161 6080
rect -123 6046 -111 6080
rect 11 6046 27 6080
rect 61 6046 95 6080
rect 129 6046 145 6080
<< viali >>
rect -229 6338 -197 6372
rect -197 6338 -195 6372
rect -157 6338 -129 6372
rect -129 6338 -123 6372
rect -229 6046 -195 6080
rect -157 6046 -127 6080
rect -127 6046 -123 6080
<< metal1 >>
rect -241 6372 -111 6378
rect -241 6338 -229 6372
rect -195 6338 -157 6372
rect -123 6338 -111 6372
rect -241 6080 -111 6338
rect -241 6046 -229 6080
rect -195 6046 -157 6080
rect -123 6046 -111 6080
rect -241 6040 -111 6046
use sky130_fd_pr__res_bent_po__example_5595914180861  sky130_fd_pr__res_bent_po__example_5595914180861_0
timestamp 1648127584
transform 0 -1 -98 -1 0 6046
box -50 -243 -49 14
use sky130_fd_pr__res_bent_po__example_5595914180862  sky130_fd_pr__res_bent_po__example_5595914180862_0
timestamp 1648127584
transform 0 1 -3 -1 0 8908
box -50 13 1185 14
use sky130_fd_pr__res_bent_po__example_5595914180862  sky130_fd_pr__res_bent_po__example_5595914180862_1
timestamp 1648127584
transform 0 1 -3 -1 0 7566
box -50 13 1185 14
use sky130_fd_pr__res_bent_po__example_5595914180863  sky130_fd_pr__res_bent_po__example_5595914180863_0
timestamp 1648127584
transform 0 1 -260 -1 0 8772
box -50 13 2385 14
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1648127584
transform 1 0 -229 0 1 6338
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1648127584
transform 1 0 -229 0 1 6046
box 0 0 1 1
<< properties >>
string GDS_END 43493888
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43493324
<< end >>
