magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 67 1010 203
rect 29 21 1010 67
rect 29 -17 63 21
<< scnmos >>
rect 79 93 109 177
rect 267 47 297 177
rect 373 47 403 177
rect 457 47 487 177
rect 541 47 571 177
rect 647 47 677 177
rect 731 47 761 177
rect 815 47 845 177
rect 899 47 929 177
<< scpmoshvt >>
rect 79 413 109 497
rect 267 297 297 497
rect 373 297 403 497
rect 457 297 487 497
rect 541 297 571 497
rect 647 297 677 497
rect 731 297 761 497
rect 815 297 845 497
rect 899 297 929 497
<< ndiff >>
rect 27 149 79 177
rect 27 115 35 149
rect 69 115 79 149
rect 27 93 79 115
rect 109 165 161 177
rect 109 131 119 165
rect 153 131 161 165
rect 109 120 161 131
rect 109 93 159 120
rect 217 104 267 177
rect 215 93 267 104
rect 215 59 223 93
rect 257 59 267 93
rect 215 47 267 59
rect 297 115 373 177
rect 297 81 323 115
rect 357 81 373 115
rect 297 47 373 81
rect 403 97 457 177
rect 403 63 413 97
rect 447 63 457 97
rect 403 47 457 63
rect 487 115 541 177
rect 487 81 497 115
rect 531 81 541 115
rect 487 47 541 81
rect 571 97 647 177
rect 571 63 601 97
rect 635 63 647 97
rect 571 47 647 63
rect 677 114 731 177
rect 677 80 687 114
rect 721 80 731 114
rect 677 47 731 80
rect 761 95 815 177
rect 761 61 771 95
rect 805 61 815 95
rect 761 47 815 61
rect 845 163 899 177
rect 845 129 855 163
rect 889 129 899 163
rect 845 95 899 129
rect 845 61 855 95
rect 889 61 899 95
rect 845 47 899 61
rect 929 95 984 177
rect 929 61 939 95
rect 973 61 984 95
rect 929 47 984 61
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 413 79 443
rect 109 472 161 497
rect 109 438 119 472
rect 153 438 161 472
rect 109 413 161 438
rect 215 485 267 497
rect 215 451 223 485
rect 257 451 267 485
rect 215 417 267 451
rect 215 383 223 417
rect 257 383 267 417
rect 215 349 267 383
rect 215 315 223 349
rect 257 315 267 349
rect 215 297 267 315
rect 297 297 373 497
rect 403 297 457 497
rect 487 297 541 497
rect 571 477 647 497
rect 571 443 592 477
rect 626 443 647 477
rect 571 409 647 443
rect 571 375 592 409
rect 626 375 647 409
rect 571 297 647 375
rect 677 477 731 497
rect 677 443 687 477
rect 721 443 731 477
rect 677 409 731 443
rect 677 375 687 409
rect 721 375 731 409
rect 677 341 731 375
rect 677 307 687 341
rect 721 307 731 341
rect 677 297 731 307
rect 761 477 815 497
rect 761 443 771 477
rect 805 443 815 477
rect 761 409 815 443
rect 761 375 771 409
rect 805 375 815 409
rect 761 297 815 375
rect 845 477 899 497
rect 845 443 855 477
rect 889 443 899 477
rect 845 409 899 443
rect 845 375 855 409
rect 889 375 899 409
rect 845 341 899 375
rect 845 307 855 341
rect 889 307 899 341
rect 845 297 899 307
rect 929 477 981 497
rect 929 443 939 477
rect 973 443 981 477
rect 929 409 981 443
rect 929 375 939 409
rect 973 375 981 409
rect 929 297 981 375
<< ndiffc >>
rect 35 115 69 149
rect 119 131 153 165
rect 223 59 257 93
rect 323 81 357 115
rect 413 63 447 97
rect 497 81 531 115
rect 601 63 635 97
rect 687 80 721 114
rect 771 61 805 95
rect 855 129 889 163
rect 855 61 889 95
rect 939 61 973 95
<< pdiffc >>
rect 35 443 69 477
rect 119 438 153 472
rect 223 451 257 485
rect 223 383 257 417
rect 223 315 257 349
rect 592 443 626 477
rect 592 375 626 409
rect 687 443 721 477
rect 687 375 721 409
rect 687 307 721 341
rect 771 443 805 477
rect 771 375 805 409
rect 855 443 889 477
rect 855 375 889 409
rect 855 307 889 341
rect 939 443 973 477
rect 939 375 973 409
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 373 497 403 523
rect 457 497 487 523
rect 541 497 571 523
rect 647 497 677 523
rect 731 497 761 523
rect 815 497 845 523
rect 899 497 929 523
rect 79 265 109 413
rect 267 265 297 297
rect 373 265 403 297
rect 457 265 487 297
rect 541 265 571 297
rect 647 265 677 297
rect 731 265 761 297
rect 815 265 845 297
rect 899 265 929 297
rect 45 249 113 265
rect 45 215 55 249
rect 89 215 113 249
rect 45 199 113 215
rect 199 249 297 265
rect 199 215 209 249
rect 243 215 297 249
rect 199 199 297 215
rect 349 249 403 265
rect 349 215 359 249
rect 393 215 403 249
rect 349 199 403 215
rect 445 249 499 265
rect 445 215 455 249
rect 489 215 499 249
rect 445 199 499 215
rect 541 249 595 265
rect 541 215 551 249
rect 585 215 595 249
rect 541 199 595 215
rect 647 249 929 265
rect 647 215 657 249
rect 691 215 725 249
rect 759 215 793 249
rect 827 215 861 249
rect 895 215 929 249
rect 647 199 929 215
rect 79 177 109 199
rect 267 177 297 199
rect 373 177 403 199
rect 457 177 487 199
rect 541 177 571 199
rect 647 177 677 199
rect 731 177 761 199
rect 815 177 845 199
rect 899 177 929 199
rect 79 67 109 93
rect 267 21 297 47
rect 373 21 403 47
rect 457 21 487 47
rect 541 21 571 47
rect 647 21 677 47
rect 731 21 761 47
rect 815 21 845 47
rect 899 21 929 47
<< polycont >>
rect 55 215 89 249
rect 209 215 243 249
rect 359 215 393 249
rect 455 215 489 249
rect 551 215 585 249
rect 657 215 691 249
rect 725 215 759 249
rect 793 215 827 249
rect 861 215 895 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 17 477 73 527
rect 17 443 35 477
rect 69 443 73 477
rect 17 427 73 443
rect 119 472 157 491
rect 153 438 157 472
rect 119 413 157 438
rect 21 249 89 391
rect 21 215 55 249
rect 21 199 89 215
rect 123 265 157 413
rect 207 485 273 490
rect 207 451 223 485
rect 257 451 273 485
rect 584 477 634 527
rect 207 417 273 451
rect 207 383 223 417
rect 257 383 273 417
rect 207 349 273 383
rect 207 315 223 349
rect 257 315 325 349
rect 123 249 243 265
rect 123 215 209 249
rect 123 199 243 215
rect 123 181 157 199
rect 119 165 157 181
rect 17 149 69 165
rect 17 115 35 149
rect 17 17 69 115
rect 153 131 157 165
rect 291 165 325 315
rect 359 324 431 475
rect 467 357 527 475
rect 584 443 592 477
rect 626 443 634 477
rect 584 409 634 443
rect 584 375 592 409
rect 626 375 634 409
rect 584 359 634 375
rect 679 477 729 493
rect 679 443 687 477
rect 721 443 729 477
rect 679 409 729 443
rect 679 375 687 409
rect 721 375 729 409
rect 359 249 393 324
rect 467 290 505 357
rect 679 341 729 375
rect 763 477 813 527
rect 763 443 771 477
rect 805 443 813 477
rect 763 409 813 443
rect 763 375 771 409
rect 805 375 813 409
rect 763 359 813 375
rect 847 477 897 493
rect 847 443 855 477
rect 889 443 897 477
rect 847 409 897 443
rect 847 375 855 409
rect 889 375 897 409
rect 359 199 393 215
rect 439 249 505 290
rect 439 215 455 249
rect 489 215 505 249
rect 439 199 505 215
rect 551 289 638 323
rect 679 307 687 341
rect 721 325 729 341
rect 847 341 897 375
rect 931 477 981 527
rect 931 443 939 477
rect 973 443 981 477
rect 931 409 981 443
rect 931 375 939 409
rect 973 375 981 409
rect 931 359 981 375
rect 847 325 855 341
rect 721 307 855 325
rect 889 325 897 341
rect 889 307 993 325
rect 679 291 993 307
rect 551 249 585 289
rect 551 199 585 215
rect 619 215 657 249
rect 691 215 725 249
rect 759 215 793 249
rect 827 215 861 249
rect 895 215 911 249
rect 619 165 653 215
rect 945 181 993 291
rect 291 131 653 165
rect 687 163 993 181
rect 687 145 855 163
rect 119 87 157 131
rect 207 93 257 117
rect 207 59 223 93
rect 323 115 357 131
rect 497 115 531 131
rect 323 61 357 81
rect 397 63 413 97
rect 447 63 463 97
rect 207 17 257 59
rect 397 17 463 63
rect 687 114 737 145
rect 497 61 531 81
rect 575 63 601 97
rect 635 63 651 97
rect 575 17 651 63
rect 721 80 737 114
rect 839 129 855 145
rect 889 145 993 163
rect 889 129 905 145
rect 687 51 737 80
rect 771 95 805 111
rect 771 17 805 61
rect 839 95 905 129
rect 839 61 855 95
rect 889 61 905 95
rect 839 51 905 61
rect 939 95 973 111
rect 939 17 973 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
<< metal1 >>
rect 0 561 1012 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 496 1012 527
rect 0 17 1012 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 -48 1012 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 489 425 523 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 489 357 523 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 397 357 431 391 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 397 425 431 459 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 949 153 983 187 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 or4b_4
rlabel metal1 s 0 -48 1012 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_END 1085826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1077394
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.060 0.000 
<< end >>
