magic
tech sky130A
magscale 1 2
timestamp 1654144341
<< nwell >>
rect -396 700 772 1034
rect -16 512 306 700
rect -16 474 210 512
rect -234 -24 976 -22
rect -234 -30 1322 -24
rect -572 -343 1322 -30
rect -572 -351 630 -343
rect 970 -345 1322 -343
rect -234 -422 630 -351
rect -18 -544 304 -422
rect -18 -582 208 -544
<< pwell >>
rect -355 463 -85 645
rect 459 463 729 645
rect 10 218 312 400
rect 54 34 266 134
rect -492 -591 -306 -409
rect 704 -583 890 -401
rect 1009 -585 1283 -429
rect 8 -838 310 -656
rect 52 -1022 264 -922
<< nmos >>
rect 98 244 128 374
rect 194 244 224 374
rect 96 -812 126 -682
rect 192 -812 222 -682
<< scnmos >>
rect -277 489 -247 619
rect -193 489 -163 619
rect 537 489 567 619
rect 621 489 651 619
rect -414 -565 -384 -435
rect 782 -557 812 -427
rect 1087 -559 1117 -455
rect 1175 -559 1205 -455
<< scpmoshvt >>
rect -277 739 -247 939
rect -205 739 -175 939
rect 537 739 567 939
rect 609 739 639 939
rect -414 -315 -384 -115
rect 782 -307 812 -107
rect 1087 -267 1117 -109
rect 1175 -267 1205 -109
<< pmoshvt >>
rect 82 574 112 774
rect 178 574 208 774
rect -140 -322 -110 -122
rect 80 -482 110 -282
rect 176 -482 206 -282
rect 506 -322 536 -122
<< ndiff >>
rect -329 605 -277 619
rect -329 571 -321 605
rect -287 571 -277 605
rect -329 537 -277 571
rect -329 503 -321 537
rect -287 503 -277 537
rect -329 489 -277 503
rect -247 605 -193 619
rect -247 571 -237 605
rect -203 571 -193 605
rect -247 537 -193 571
rect -247 503 -237 537
rect -203 503 -193 537
rect -247 489 -193 503
rect -163 605 -111 619
rect -163 571 -153 605
rect -119 571 -111 605
rect 485 605 537 619
rect -163 537 -111 571
rect 485 571 493 605
rect 527 571 537 605
rect -163 503 -153 537
rect -119 503 -111 537
rect -163 489 -111 503
rect 485 537 537 571
rect 485 503 493 537
rect 527 503 537 537
rect 485 489 537 503
rect 567 605 621 619
rect 567 571 577 605
rect 611 571 621 605
rect 567 537 621 571
rect 567 503 577 537
rect 611 503 621 537
rect 567 489 621 503
rect 651 605 703 619
rect 651 571 661 605
rect 695 571 703 605
rect 651 537 703 571
rect 651 503 661 537
rect 695 503 703 537
rect 651 489 703 503
rect 36 360 98 374
rect 36 326 48 360
rect 82 326 98 360
rect 36 292 98 326
rect 36 258 48 292
rect 82 258 98 292
rect 36 244 98 258
rect 128 360 194 374
rect 128 326 144 360
rect 178 326 194 360
rect 128 292 194 326
rect 128 258 144 292
rect 178 258 194 292
rect 128 244 194 258
rect 224 360 286 374
rect 224 326 240 360
rect 274 326 286 360
rect 224 292 286 326
rect 224 258 240 292
rect 274 258 286 292
rect 224 244 286 258
rect -466 -447 -414 -435
rect -466 -481 -458 -447
rect -424 -481 -414 -447
rect -466 -515 -414 -481
rect -466 -549 -458 -515
rect -424 -549 -414 -515
rect -466 -565 -414 -549
rect -384 -447 -332 -435
rect -384 -481 -374 -447
rect -340 -481 -332 -447
rect -384 -515 -332 -481
rect 730 -439 782 -427
rect 730 -473 738 -439
rect 772 -473 782 -439
rect 730 -507 782 -473
rect -384 -549 -374 -515
rect -340 -549 -332 -515
rect -384 -565 -332 -549
rect 730 -541 738 -507
rect 772 -541 782 -507
rect 730 -557 782 -541
rect 812 -439 864 -427
rect 812 -473 822 -439
rect 856 -473 864 -439
rect 812 -507 864 -473
rect 812 -541 822 -507
rect 856 -541 864 -507
rect 812 -557 864 -541
rect 1035 -500 1087 -455
rect 1035 -534 1043 -500
rect 1077 -534 1087 -500
rect 1035 -559 1087 -534
rect 1117 -513 1175 -455
rect 1117 -547 1129 -513
rect 1163 -547 1175 -513
rect 1117 -559 1175 -547
rect 1205 -483 1257 -455
rect 1205 -517 1215 -483
rect 1249 -517 1257 -483
rect 1205 -559 1257 -517
rect 34 -696 96 -682
rect 34 -730 46 -696
rect 80 -730 96 -696
rect 34 -764 96 -730
rect 34 -798 46 -764
rect 80 -798 96 -764
rect 34 -812 96 -798
rect 126 -696 192 -682
rect 126 -730 142 -696
rect 176 -730 192 -696
rect 126 -764 192 -730
rect 126 -798 142 -764
rect 176 -798 192 -764
rect 126 -812 192 -798
rect 222 -696 284 -682
rect 222 -730 238 -696
rect 272 -730 284 -696
rect 222 -764 284 -730
rect 222 -798 238 -764
rect 272 -798 284 -764
rect 222 -812 284 -798
<< pdiff >>
rect -329 927 -277 939
rect -329 893 -321 927
rect -287 893 -277 927
rect -329 859 -277 893
rect -329 825 -321 859
rect -287 825 -277 859
rect -329 791 -277 825
rect -329 757 -321 791
rect -287 757 -277 791
rect -329 739 -277 757
rect -247 739 -205 939
rect -175 927 -123 939
rect -175 893 -165 927
rect -131 893 -123 927
rect 485 927 537 939
rect -175 859 -123 893
rect 485 893 493 927
rect 527 893 537 927
rect -175 825 -165 859
rect -131 825 -123 859
rect -175 791 -123 825
rect 485 859 537 893
rect 485 825 493 859
rect 527 825 537 859
rect -175 757 -165 791
rect -131 757 -123 791
rect 485 791 537 825
rect -175 739 -123 757
rect 20 759 82 774
rect 20 725 32 759
rect 66 725 82 759
rect 20 691 82 725
rect 20 657 32 691
rect 66 657 82 691
rect 20 623 82 657
rect 20 589 32 623
rect 66 589 82 623
rect 20 574 82 589
rect 112 759 178 774
rect 112 725 128 759
rect 162 725 178 759
rect 112 691 178 725
rect 112 657 128 691
rect 162 657 178 691
rect 112 623 178 657
rect 112 589 128 623
rect 162 589 178 623
rect 112 574 178 589
rect 208 759 270 774
rect 208 725 224 759
rect 258 725 270 759
rect 485 757 493 791
rect 527 757 537 791
rect 485 739 537 757
rect 567 739 609 939
rect 639 927 691 939
rect 639 893 649 927
rect 683 893 691 927
rect 639 859 691 893
rect 639 825 649 859
rect 683 825 691 859
rect 639 791 691 825
rect 639 757 649 791
rect 683 757 691 791
rect 639 739 691 757
rect 208 691 270 725
rect 208 657 224 691
rect 258 657 270 691
rect 208 623 270 657
rect 208 589 224 623
rect 258 589 270 623
rect 208 574 270 589
rect -466 -127 -414 -115
rect -466 -161 -458 -127
rect -424 -161 -414 -127
rect -466 -195 -414 -161
rect -466 -229 -458 -195
rect -424 -229 -414 -195
rect -466 -263 -414 -229
rect -466 -297 -458 -263
rect -424 -297 -414 -263
rect -466 -315 -414 -297
rect -384 -127 -332 -115
rect -384 -161 -374 -127
rect -340 -161 -332 -127
rect -384 -195 -332 -161
rect -384 -229 -374 -195
rect -340 -229 -332 -195
rect -384 -263 -332 -229
rect -384 -297 -374 -263
rect -340 -297 -332 -263
rect -384 -315 -332 -297
rect -198 -137 -140 -122
rect -198 -171 -186 -137
rect -152 -171 -140 -137
rect -198 -205 -140 -171
rect -198 -239 -186 -205
rect -152 -239 -140 -205
rect -198 -273 -140 -239
rect -198 -307 -186 -273
rect -152 -307 -140 -273
rect -198 -322 -140 -307
rect -110 -137 -52 -122
rect -110 -171 -98 -137
rect -64 -171 -52 -137
rect -110 -205 -52 -171
rect 730 -119 782 -107
rect 448 -137 506 -122
rect 448 -171 460 -137
rect 494 -171 506 -137
rect -110 -239 -98 -205
rect -64 -239 -52 -205
rect -110 -273 -52 -239
rect -110 -307 -98 -273
rect -64 -307 -52 -273
rect 448 -205 506 -171
rect 448 -239 460 -205
rect 494 -239 506 -205
rect 448 -273 506 -239
rect -110 -322 -52 -307
rect 18 -297 80 -282
rect 18 -331 30 -297
rect 64 -331 80 -297
rect 18 -365 80 -331
rect 18 -399 30 -365
rect 64 -399 80 -365
rect 18 -433 80 -399
rect 18 -467 30 -433
rect 64 -467 80 -433
rect 18 -482 80 -467
rect 110 -297 176 -282
rect 110 -331 126 -297
rect 160 -331 176 -297
rect 110 -365 176 -331
rect 110 -399 126 -365
rect 160 -399 176 -365
rect 110 -433 176 -399
rect 110 -467 126 -433
rect 160 -467 176 -433
rect 110 -482 176 -467
rect 206 -297 268 -282
rect 206 -331 222 -297
rect 256 -331 268 -297
rect 448 -307 460 -273
rect 494 -307 506 -273
rect 448 -322 506 -307
rect 536 -137 594 -122
rect 536 -171 548 -137
rect 582 -171 594 -137
rect 536 -205 594 -171
rect 536 -239 548 -205
rect 582 -239 594 -205
rect 536 -273 594 -239
rect 536 -307 548 -273
rect 582 -307 594 -273
rect 730 -153 738 -119
rect 772 -153 782 -119
rect 730 -187 782 -153
rect 730 -221 738 -187
rect 772 -221 782 -187
rect 730 -255 782 -221
rect 730 -289 738 -255
rect 772 -289 782 -255
rect 730 -307 782 -289
rect 812 -119 864 -107
rect 812 -153 822 -119
rect 856 -153 864 -119
rect 812 -187 864 -153
rect 812 -221 822 -187
rect 856 -221 864 -187
rect 812 -255 864 -221
rect 812 -289 822 -255
rect 856 -289 864 -255
rect 1035 -129 1087 -109
rect 1035 -163 1043 -129
rect 1077 -163 1087 -129
rect 1035 -197 1087 -163
rect 1035 -231 1043 -197
rect 1077 -231 1087 -197
rect 1035 -267 1087 -231
rect 1117 -129 1175 -109
rect 1117 -163 1129 -129
rect 1163 -163 1175 -129
rect 1117 -197 1175 -163
rect 1117 -231 1129 -197
rect 1163 -231 1175 -197
rect 1117 -267 1175 -231
rect 1205 -129 1257 -109
rect 1205 -163 1215 -129
rect 1249 -163 1257 -129
rect 1205 -210 1257 -163
rect 1205 -244 1215 -210
rect 1249 -244 1257 -210
rect 1205 -267 1257 -244
rect 812 -307 864 -289
rect 536 -322 594 -307
rect 206 -365 268 -331
rect 206 -399 222 -365
rect 256 -399 268 -365
rect 206 -433 268 -399
rect 206 -467 222 -433
rect 256 -467 268 -433
rect 206 -482 268 -467
<< ndiffc >>
rect -321 571 -287 605
rect -321 503 -287 537
rect -237 571 -203 605
rect -237 503 -203 537
rect -153 571 -119 605
rect 493 571 527 605
rect -153 503 -119 537
rect 493 503 527 537
rect 577 571 611 605
rect 577 503 611 537
rect 661 571 695 605
rect 661 503 695 537
rect 48 326 82 360
rect 48 258 82 292
rect 144 326 178 360
rect 144 258 178 292
rect 240 326 274 360
rect 240 258 274 292
rect -458 -481 -424 -447
rect -458 -549 -424 -515
rect -374 -481 -340 -447
rect 738 -473 772 -439
rect -374 -549 -340 -515
rect 738 -541 772 -507
rect 822 -473 856 -439
rect 822 -541 856 -507
rect 1043 -534 1077 -500
rect 1129 -547 1163 -513
rect 1215 -517 1249 -483
rect 46 -730 80 -696
rect 46 -798 80 -764
rect 142 -730 176 -696
rect 142 -798 176 -764
rect 238 -730 272 -696
rect 238 -798 272 -764
<< pdiffc >>
rect -321 893 -287 927
rect -321 825 -287 859
rect -321 757 -287 791
rect -165 893 -131 927
rect 493 893 527 927
rect -165 825 -131 859
rect 493 825 527 859
rect -165 757 -131 791
rect 32 725 66 759
rect 32 657 66 691
rect 32 589 66 623
rect 128 725 162 759
rect 128 657 162 691
rect 128 589 162 623
rect 224 725 258 759
rect 493 757 527 791
rect 649 893 683 927
rect 649 825 683 859
rect 649 757 683 791
rect 224 657 258 691
rect 224 589 258 623
rect -458 -161 -424 -127
rect -458 -229 -424 -195
rect -458 -297 -424 -263
rect -374 -161 -340 -127
rect -374 -229 -340 -195
rect -374 -297 -340 -263
rect -186 -171 -152 -137
rect -186 -239 -152 -205
rect -186 -307 -152 -273
rect -98 -171 -64 -137
rect 460 -171 494 -137
rect -98 -239 -64 -205
rect -98 -307 -64 -273
rect 460 -239 494 -205
rect 30 -331 64 -297
rect 30 -399 64 -365
rect 30 -467 64 -433
rect 126 -331 160 -297
rect 126 -399 160 -365
rect 126 -467 160 -433
rect 222 -331 256 -297
rect 460 -307 494 -273
rect 548 -171 582 -137
rect 548 -239 582 -205
rect 548 -307 582 -273
rect 738 -153 772 -119
rect 738 -221 772 -187
rect 738 -289 772 -255
rect 822 -153 856 -119
rect 822 -221 856 -187
rect 822 -289 856 -255
rect 1043 -163 1077 -129
rect 1043 -231 1077 -197
rect 1129 -163 1163 -129
rect 1129 -231 1163 -197
rect 1215 -163 1249 -129
rect 1215 -244 1249 -210
rect 222 -399 256 -365
rect 222 -467 256 -433
<< psubdiff >>
rect 80 102 240 108
rect 80 68 137 102
rect 171 68 240 102
rect 80 60 240 68
rect 78 -954 238 -948
rect 78 -988 135 -954
rect 169 -988 238 -954
rect 78 -996 238 -988
<< nsubdiff >>
rect 198 961 332 978
rect 198 927 226 961
rect 260 927 332 961
rect 198 908 332 927
rect 196 -95 330 -78
rect 196 -129 224 -95
rect 258 -129 330 -95
rect 196 -148 330 -129
<< psubdiffcont >>
rect 137 68 171 102
rect 135 -988 169 -954
<< nsubdiffcont >>
rect 226 927 260 961
rect 224 -129 258 -95
<< poly >>
rect -277 939 -247 965
rect -205 939 -175 965
rect 537 939 567 965
rect 609 939 639 965
rect 160 855 226 871
rect 160 821 176 855
rect 210 821 226 855
rect 160 805 226 821
rect 82 774 112 800
rect 178 774 208 805
rect -277 707 -247 739
rect -334 691 -247 707
rect -334 657 -319 691
rect -285 657 -247 691
rect -205 707 -175 739
rect -205 691 -101 707
rect -205 677 -151 691
rect -334 641 -247 657
rect -277 619 -247 641
rect -193 657 -151 677
rect -117 657 -101 691
rect -193 641 -101 657
rect -193 619 -163 641
rect 537 707 567 739
rect 480 691 567 707
rect 480 657 495 691
rect 529 657 567 691
rect 609 707 639 739
rect 609 691 713 707
rect 609 677 663 691
rect 480 641 567 657
rect 537 619 567 641
rect 621 657 663 677
rect 697 657 713 691
rect 621 641 713 657
rect 621 619 651 641
rect 82 543 112 574
rect 178 548 208 574
rect 64 527 130 543
rect 64 493 80 527
rect 114 506 130 527
rect 114 493 242 506
rect -277 463 -247 489
rect -193 463 -163 489
rect 64 474 242 493
rect 176 446 242 474
rect 537 463 567 489
rect 621 463 651 489
rect 176 412 192 446
rect 226 412 242 446
rect 98 374 128 400
rect 176 396 242 412
rect 194 374 224 396
rect 98 222 128 244
rect 80 206 146 222
rect 80 172 96 206
rect 130 172 146 206
rect 194 218 224 244
rect 194 188 328 218
rect 80 156 146 172
rect 298 20 328 188
rect 24 -10 506 20
rect -158 -41 -92 -25
rect -158 -75 -142 -41
rect -108 -75 -92 -41
rect -414 -115 -384 -89
rect -158 -91 -92 -75
rect -140 -122 -110 -91
rect -414 -347 -384 -315
rect 24 -168 54 -10
rect 474 -25 506 -10
rect 474 -41 554 -25
rect 474 -75 504 -41
rect 538 -75 554 -41
rect 474 -91 554 -75
rect 474 -92 536 -91
rect 506 -122 536 -92
rect 782 -107 812 -81
rect 24 -198 110 -168
rect 80 -282 110 -198
rect 158 -201 224 -185
rect 158 -235 174 -201
rect 208 -235 224 -201
rect 158 -251 224 -235
rect 176 -282 206 -251
rect -470 -363 -384 -347
rect -140 -353 -110 -322
rect -470 -397 -454 -363
rect -420 -397 -384 -363
rect -470 -413 -384 -397
rect -414 -435 -384 -413
rect -158 -369 -92 -353
rect -158 -403 -142 -369
rect -108 -403 -92 -369
rect -158 -419 -92 -403
rect 1087 -109 1117 -83
rect 1175 -109 1205 -83
rect 1087 -282 1117 -267
rect 1081 -306 1117 -282
rect 506 -353 536 -322
rect 782 -339 812 -307
rect 488 -369 554 -353
rect 488 -403 504 -369
rect 538 -403 554 -369
rect 488 -419 554 -403
rect 726 -355 812 -339
rect 1081 -341 1111 -306
rect 1175 -328 1205 -267
rect 726 -389 742 -355
rect 776 -389 812 -355
rect 726 -405 812 -389
rect 782 -427 812 -405
rect 1035 -357 1111 -341
rect 1035 -391 1045 -357
rect 1079 -391 1111 -357
rect 1035 -407 1111 -391
rect 1153 -344 1207 -328
rect 1153 -378 1163 -344
rect 1197 -378 1207 -344
rect 1153 -394 1207 -378
rect 1081 -416 1111 -407
rect 80 -513 110 -482
rect 176 -508 206 -482
rect 62 -529 128 -513
rect 62 -563 78 -529
rect 112 -550 128 -529
rect 112 -563 240 -550
rect 1081 -440 1117 -416
rect 1087 -455 1117 -440
rect 1175 -455 1205 -394
rect -414 -591 -384 -565
rect 62 -582 240 -563
rect 174 -610 240 -582
rect 782 -583 812 -557
rect 1087 -585 1117 -559
rect 1175 -585 1205 -559
rect 174 -644 190 -610
rect 224 -644 240 -610
rect 96 -682 126 -656
rect 174 -660 240 -644
rect 192 -682 222 -660
rect 96 -834 126 -812
rect 78 -850 144 -834
rect 192 -838 222 -812
rect 78 -884 94 -850
rect 128 -884 144 -850
rect 78 -900 144 -884
<< polycont >>
rect 176 821 210 855
rect -319 657 -285 691
rect -151 657 -117 691
rect 495 657 529 691
rect 663 657 697 691
rect 80 493 114 527
rect 192 412 226 446
rect 96 172 130 206
rect -142 -75 -108 -41
rect 504 -75 538 -41
rect 174 -235 208 -201
rect -454 -397 -420 -363
rect -142 -403 -108 -369
rect 504 -403 538 -369
rect 742 -389 776 -355
rect 1045 -391 1079 -357
rect 1163 -378 1197 -344
rect 78 -563 112 -529
rect 190 -644 224 -610
rect 94 -884 128 -850
<< locali >>
rect -398 1003 -336 1004
rect 68 1003 458 1004
rect -398 970 -327 1003
rect -356 969 -327 970
rect -293 969 -235 1003
rect -201 969 -143 1003
rect -109 969 487 1003
rect 521 969 579 1003
rect 613 969 671 1003
rect 705 969 734 1003
rect -337 927 -271 932
rect -337 893 -321 927
rect -287 893 -271 927
rect -337 859 -271 893
rect -337 825 -321 859
rect -287 825 -271 859
rect -337 791 -271 825
rect -337 757 -321 791
rect -287 775 -271 791
rect -165 927 -99 969
rect -131 893 -99 927
rect 68 963 350 969
rect 68 929 107 963
rect 141 961 350 963
rect 141 929 226 961
rect 68 927 226 929
rect 260 927 350 961
rect 68 894 350 927
rect 477 927 543 932
rect -165 859 -99 893
rect -131 825 -99 859
rect 477 893 493 927
rect 527 893 543 927
rect 477 859 543 893
rect -165 791 -99 825
rect -287 757 -201 775
rect -337 741 -201 757
rect -131 757 -99 791
rect -165 741 -99 757
rect -40 855 226 856
rect -40 821 176 855
rect 210 821 226 855
rect -40 820 226 821
rect -339 700 -269 707
rect -339 666 -321 700
rect -287 691 -269 700
rect -339 657 -319 666
rect -285 657 -269 691
rect -235 621 -201 741
rect -167 696 -97 707
rect -167 691 -148 696
rect -167 657 -151 691
rect -114 662 -97 696
rect -117 657 -97 662
rect -335 605 -287 621
rect -335 571 -321 605
rect -335 537 -287 571
rect -335 503 -321 537
rect -335 459 -287 503
rect -253 605 -187 621
rect -253 580 -237 605
rect -253 546 -239 580
rect -203 571 -187 605
rect -205 546 -187 571
rect -253 537 -187 546
rect -253 503 -237 537
rect -203 503 -187 537
rect -253 493 -187 503
rect -153 605 -99 621
rect -119 571 -99 605
rect -153 537 -99 571
rect -119 503 -99 537
rect -153 459 -99 503
rect -356 425 -327 459
rect -293 425 -235 459
rect -201 425 -143 459
rect -109 425 -80 459
rect -356 214 -322 425
rect -125 122 -91 425
rect -40 206 -6 820
rect 160 818 226 820
rect 477 825 493 859
rect 527 825 543 859
rect 477 791 543 825
rect 32 759 66 778
rect 32 691 66 693
rect 32 655 66 657
rect 32 570 66 589
rect 128 759 162 778
rect 128 691 162 693
rect 128 655 162 657
rect 128 570 162 589
rect 224 759 258 778
rect 477 757 493 791
rect 527 775 543 791
rect 649 927 715 969
rect 683 893 715 927
rect 649 859 715 893
rect 683 825 715 859
rect 649 791 715 825
rect 527 757 613 775
rect 477 741 613 757
rect 683 757 715 791
rect 649 741 715 757
rect 224 691 258 693
rect 475 698 545 707
rect 475 664 491 698
rect 525 691 545 698
rect 475 657 495 664
rect 529 657 545 691
rect 224 655 258 657
rect 579 621 613 741
rect 647 698 717 707
rect 647 691 665 698
rect 647 657 663 691
rect 699 664 717 698
rect 697 657 717 664
rect 224 570 258 589
rect 479 605 527 621
rect 479 571 493 605
rect 479 537 527 571
rect 64 493 80 527
rect 114 493 130 527
rect 479 503 493 537
rect 479 459 527 503
rect 561 605 627 621
rect 561 571 577 605
rect 611 575 627 605
rect 561 541 579 571
rect 613 541 627 575
rect 561 537 627 541
rect 561 503 577 537
rect 611 503 627 537
rect 561 493 627 503
rect 661 605 715 621
rect 695 571 715 605
rect 661 537 715 571
rect 695 503 715 537
rect 661 459 715 503
rect 176 412 192 446
rect 226 412 242 446
rect 458 425 487 459
rect 521 425 579 459
rect 613 425 671 459
rect 705 425 734 459
rect 48 362 82 378
rect 48 292 82 326
rect 48 240 82 256
rect 144 362 178 378
rect 144 292 178 326
rect 144 240 178 256
rect 240 362 274 378
rect 240 292 274 326
rect 274 256 622 280
rect 240 240 622 256
rect -40 172 96 206
rect 130 172 146 206
rect -125 102 270 122
rect -125 97 137 102
rect -125 88 16 97
rect 0 63 16 88
rect 50 68 137 97
rect 171 78 270 102
rect 442 80 488 82
rect 442 78 446 80
rect 171 68 446 78
rect 50 63 446 68
rect 0 46 446 63
rect 480 46 488 80
rect 0 44 488 46
rect 442 38 488 44
rect -459 -51 -425 -44
rect -534 -85 -505 -51
rect -471 -85 -413 -51
rect -379 -85 -321 -51
rect -287 -85 -258 -51
rect -158 -75 -142 -41
rect -108 -75 -92 -41
rect 66 -54 180 -52
rect -466 -127 -424 -85
rect 66 -93 348 -54
rect 488 -75 504 -41
rect 538 -75 554 -41
rect 66 -118 105 -93
rect -466 -161 -458 -127
rect -466 -195 -424 -161
rect -466 -229 -458 -195
rect -466 -263 -424 -229
rect -466 -297 -458 -263
rect -466 -313 -424 -297
rect -390 -127 -324 -119
rect -390 -161 -374 -127
rect -340 -161 -324 -127
rect -390 -195 -324 -161
rect -390 -229 -374 -195
rect -340 -229 -324 -195
rect -390 -263 -324 -229
rect -390 -297 -374 -263
rect -340 -297 -324 -263
rect -390 -315 -324 -297
rect -470 -352 -404 -349
rect -470 -386 -456 -352
rect -422 -363 -404 -352
rect -470 -397 -454 -386
rect -420 -397 -404 -363
rect -470 -447 -424 -431
rect -370 -435 -324 -315
rect -186 -137 -152 -118
rect -100 -127 105 -118
rect 139 -95 348 -93
rect 139 -127 224 -95
rect -100 -129 224 -127
rect 258 -118 348 -95
rect 588 -118 622 240
rect 662 -77 691 -43
rect 725 -77 783 -43
rect 817 -77 875 -43
rect 909 -77 938 -43
rect 258 -129 494 -118
rect -100 -137 494 -129
rect -100 -162 -98 -137
rect -186 -205 -152 -203
rect -186 -241 -152 -239
rect -186 -326 -152 -307
rect -64 -162 460 -137
rect 546 -137 622 -118
rect 546 -158 548 -137
rect -98 -205 -64 -203
rect 158 -235 174 -201
rect 208 -235 224 -201
rect 460 -205 494 -203
rect -98 -241 -64 -239
rect 460 -241 494 -239
rect -98 -326 -64 -307
rect 30 -297 64 -278
rect 30 -365 64 -363
rect -158 -403 -142 -369
rect -108 -403 -92 -369
rect 30 -401 64 -399
rect -470 -481 -458 -447
rect -470 -515 -424 -481
rect -470 -549 -458 -515
rect -470 -595 -424 -549
rect -390 -447 -324 -435
rect -390 -481 -374 -447
rect -340 -481 -324 -447
rect -390 -494 -324 -481
rect 30 -486 64 -467
rect 126 -297 160 -278
rect 126 -365 160 -363
rect 126 -401 160 -399
rect 126 -486 160 -467
rect 222 -297 256 -278
rect 460 -326 494 -307
rect 582 -158 622 -137
rect 730 -119 772 -77
rect 1008 -79 1037 -45
rect 1071 -79 1129 -45
rect 1163 -79 1221 -45
rect 1255 -79 1284 -45
rect 730 -153 738 -119
rect 548 -205 582 -203
rect 548 -241 582 -239
rect 730 -187 772 -153
rect 730 -221 738 -187
rect 730 -255 772 -221
rect 730 -289 738 -255
rect 730 -305 772 -289
rect 806 -119 872 -111
rect 806 -153 822 -119
rect 856 -153 872 -119
rect 806 -187 872 -153
rect 806 -221 822 -187
rect 856 -221 872 -187
rect 806 -255 872 -221
rect 806 -289 822 -255
rect 856 -289 872 -255
rect 806 -307 872 -289
rect 1041 -129 1077 -113
rect 1041 -163 1043 -129
rect 1041 -197 1077 -163
rect 1041 -231 1043 -197
rect 1113 -129 1179 -79
rect 1113 -163 1129 -129
rect 1163 -163 1179 -129
rect 1113 -197 1179 -163
rect 1113 -231 1129 -197
rect 1163 -231 1179 -197
rect 1213 -129 1267 -113
rect 1213 -163 1215 -129
rect 1249 -163 1267 -129
rect 1213 -210 1267 -163
rect 1041 -265 1077 -231
rect 1213 -244 1215 -210
rect 1249 -244 1267 -210
rect 1041 -299 1176 -265
rect 1213 -294 1267 -244
rect 548 -326 582 -307
rect 222 -365 256 -363
rect 634 -341 778 -340
rect 634 -355 792 -341
rect 222 -401 256 -399
rect 488 -368 554 -366
rect 634 -368 742 -355
rect 488 -369 742 -368
rect 488 -403 504 -369
rect 538 -382 742 -369
rect 538 -402 674 -382
rect 726 -389 742 -382
rect 776 -389 792 -355
rect 538 -403 554 -402
rect 726 -439 772 -423
rect 826 -427 872 -307
rect 1142 -328 1176 -299
rect 1029 -357 1097 -335
rect 1029 -358 1045 -357
rect 1029 -392 1043 -358
rect 1079 -391 1097 -357
rect 1077 -392 1097 -391
rect 1029 -409 1097 -392
rect 1142 -344 1197 -328
rect 1142 -378 1163 -344
rect 1142 -394 1197 -378
rect 1231 -344 1267 -294
rect 1231 -346 1272 -344
rect 1231 -380 1236 -346
rect 1270 -380 1272 -346
rect 1231 -382 1272 -380
rect 256 -467 502 -450
rect 222 -484 502 -467
rect 222 -486 256 -484
rect -390 -515 -48 -494
rect -390 -549 -374 -515
rect -340 -526 -48 -515
rect -340 -529 128 -526
rect -340 -530 78 -529
rect -340 -549 -318 -530
rect -390 -554 -318 -549
rect -390 -561 -324 -554
rect -84 -562 78 -530
rect 62 -563 78 -562
rect 112 -563 128 -529
rect 454 -572 502 -484
rect -534 -629 -505 -595
rect -471 -629 -413 -595
rect -379 -629 -321 -595
rect -287 -629 -258 -595
rect -176 -600 -130 -590
rect -176 -634 -170 -600
rect -136 -620 -130 -600
rect 454 -606 462 -572
rect 496 -606 502 -572
rect 726 -473 738 -439
rect 726 -507 772 -473
rect 726 -541 738 -507
rect 726 -587 772 -541
rect 806 -439 872 -427
rect 806 -490 822 -439
rect 856 -490 872 -439
rect 1142 -445 1176 -394
rect 806 -507 872 -490
rect 806 -541 822 -507
rect 856 -541 872 -507
rect 806 -553 872 -541
rect 1043 -479 1176 -445
rect 1231 -454 1267 -382
rect 1043 -500 1077 -479
rect 1215 -483 1267 -454
rect 1043 -555 1077 -534
rect 1113 -547 1129 -513
rect 1163 -547 1179 -513
rect -136 -634 -126 -620
rect -176 -704 -126 -634
rect 174 -644 190 -610
rect 224 -644 240 -610
rect 454 -618 502 -606
rect 662 -621 691 -587
rect 725 -621 783 -587
rect 817 -621 875 -587
rect 909 -621 938 -587
rect 1113 -589 1179 -547
rect 1249 -517 1267 -483
rect 1215 -555 1267 -517
rect 1008 -623 1037 -589
rect 1071 -623 1129 -589
rect 1163 -623 1221 -589
rect 1255 -623 1284 -589
rect -258 -740 -126 -704
rect 46 -694 80 -678
rect 142 -694 176 -678
rect 80 -730 81 -729
rect -258 -788 -222 -740
rect 46 -764 81 -730
rect 80 -766 81 -764
rect 142 -764 176 -730
rect -74 -788 46 -766
rect -258 -800 46 -788
rect 80 -800 82 -766
rect -258 -802 82 -800
rect -258 -824 -38 -802
rect 46 -816 80 -802
rect 142 -816 176 -800
rect 238 -694 272 -678
rect 238 -764 272 -730
rect 238 -816 272 -800
rect 78 -884 94 -850
rect 128 -884 144 -850
rect -2 -954 268 -934
rect -2 -959 135 -954
rect -2 -993 14 -959
rect 48 -988 135 -959
rect 169 -988 268 -954
rect 48 -993 268 -988
rect -2 -1012 268 -993
<< viali >>
rect -327 969 -293 1003
rect -235 969 -201 1003
rect -143 969 -109 1003
rect 487 969 521 1003
rect 579 969 613 1003
rect 671 969 705 1003
rect 107 929 141 963
rect 176 821 210 855
rect -321 691 -287 700
rect -321 666 -319 691
rect -319 666 -287 691
rect -148 691 -114 696
rect -148 662 -117 691
rect -117 662 -114 691
rect -239 571 -237 580
rect -237 571 -205 580
rect -239 546 -205 571
rect -327 425 -293 459
rect -235 425 -201 459
rect -143 425 -109 459
rect -356 180 -322 214
rect 32 725 66 727
rect 32 693 66 725
rect 32 623 66 655
rect 32 621 66 623
rect 128 725 162 727
rect 128 693 162 725
rect 128 623 162 655
rect 128 621 162 623
rect 224 725 258 727
rect 224 693 258 725
rect 491 691 525 698
rect 491 664 495 691
rect 495 664 525 691
rect 224 623 258 655
rect 224 621 258 623
rect 665 691 699 698
rect 665 664 697 691
rect 697 664 699 691
rect 80 493 114 527
rect 579 571 611 575
rect 611 571 613 575
rect 579 541 613 571
rect 192 412 226 446
rect 487 425 521 459
rect 579 425 613 459
rect 671 425 705 459
rect 48 360 82 362
rect 48 328 82 360
rect 48 258 82 290
rect 48 256 82 258
rect 144 360 178 362
rect 144 328 178 360
rect 144 258 178 290
rect 144 256 178 258
rect 240 360 274 362
rect 240 328 274 360
rect 240 258 274 290
rect 240 256 274 258
rect 96 172 130 206
rect 16 63 50 97
rect 446 46 480 80
rect -505 -85 -471 -51
rect -413 -85 -379 -51
rect -321 -85 -287 -51
rect -142 -75 -108 -41
rect 504 -75 538 -41
rect -456 -363 -422 -352
rect -456 -386 -454 -363
rect -454 -386 -422 -363
rect 105 -127 139 -93
rect 691 -77 725 -43
rect 783 -77 817 -43
rect 875 -77 909 -43
rect -186 -171 -152 -169
rect -186 -203 -152 -171
rect -186 -273 -152 -241
rect -186 -275 -152 -273
rect -98 -171 -64 -169
rect -98 -203 -64 -171
rect 460 -171 494 -169
rect 174 -235 208 -201
rect 460 -203 494 -171
rect -98 -273 -64 -241
rect -98 -275 -64 -273
rect 460 -273 494 -241
rect 460 -275 494 -273
rect 30 -331 64 -329
rect 30 -363 64 -331
rect -142 -403 -108 -369
rect 30 -433 64 -401
rect 30 -435 64 -433
rect 126 -331 160 -329
rect 126 -363 160 -331
rect 126 -433 160 -401
rect 126 -435 160 -433
rect 1037 -79 1071 -45
rect 1129 -79 1163 -45
rect 1221 -79 1255 -45
rect 548 -171 582 -169
rect 548 -203 582 -171
rect 548 -273 582 -241
rect 548 -275 582 -273
rect 222 -331 256 -329
rect 222 -363 256 -331
rect 222 -433 256 -401
rect 504 -403 538 -369
rect 222 -435 256 -433
rect 1043 -391 1045 -358
rect 1045 -391 1077 -358
rect 1043 -392 1077 -391
rect 1236 -380 1270 -346
rect 78 -563 112 -529
rect -505 -629 -471 -595
rect -413 -629 -379 -595
rect -321 -629 -287 -595
rect -170 -634 -136 -600
rect 462 -606 496 -572
rect 822 -473 856 -456
rect 822 -490 856 -473
rect 190 -644 224 -610
rect 691 -621 725 -587
rect 783 -621 817 -587
rect 875 -621 909 -587
rect 1037 -623 1071 -589
rect 1129 -623 1163 -589
rect 1221 -623 1255 -589
rect 46 -696 80 -694
rect 46 -728 80 -696
rect 142 -696 176 -694
rect 142 -728 176 -696
rect 46 -798 80 -766
rect 46 -800 80 -798
rect 142 -798 176 -766
rect 142 -800 176 -798
rect 238 -696 272 -694
rect 238 -728 272 -696
rect 238 -798 272 -766
rect 238 -800 272 -798
rect 94 -884 128 -850
rect 14 -993 48 -959
<< metal1 >>
rect -574 1120 1322 1192
rect -574 1004 961 1120
rect 1269 1004 1322 1120
rect -574 1003 1322 1004
rect -574 969 -327 1003
rect -293 969 -235 1003
rect -201 969 -143 1003
rect -109 969 487 1003
rect 521 969 579 1003
rect 613 969 671 1003
rect 705 969 1322 1003
rect -574 963 1322 969
rect -574 938 107 963
rect -514 -20 -436 938
rect 78 929 107 938
rect 141 938 1322 963
rect 141 929 168 938
rect 78 908 168 929
rect 164 872 222 874
rect 164 855 226 872
rect 164 821 176 855
rect 210 821 226 855
rect 164 812 226 821
rect -336 774 30 778
rect 112 774 178 782
rect -336 746 72 774
rect -336 708 -308 746
rect -14 727 72 746
rect -336 700 -270 708
rect -336 666 -321 700
rect -287 666 -270 700
rect -336 654 -270 666
rect -164 704 -96 710
rect -164 652 -154 704
rect -102 652 -96 704
rect -164 646 -96 652
rect -14 693 32 727
rect 66 693 72 727
rect 112 722 118 774
rect 170 722 178 774
rect 112 714 128 722
rect -14 655 72 693
rect -14 621 32 655
rect 66 621 72 655
rect -254 592 -186 598
rect -254 540 -246 592
rect -194 540 -186 592
rect -254 530 -186 540
rect -14 574 72 621
rect 122 693 128 714
rect 162 714 178 722
rect 218 742 546 774
rect 218 727 314 742
rect 162 693 168 714
rect 122 655 168 693
rect 122 621 128 655
rect 162 621 168 655
rect 122 574 168 621
rect 218 693 224 727
rect 258 693 314 727
rect 518 706 546 742
rect 218 655 314 693
rect 218 621 224 655
rect 258 621 314 655
rect 476 698 546 706
rect 476 664 491 698
rect 525 664 546 698
rect 476 646 546 664
rect 652 706 716 712
rect 652 654 658 706
rect 710 654 716 706
rect 652 648 716 654
rect 218 574 314 621
rect -356 459 -80 490
rect -356 425 -327 459
rect -293 425 -235 459
rect -201 425 -143 459
rect -109 425 -80 459
rect -356 394 -80 425
rect -14 374 36 574
rect 68 527 126 542
rect 68 493 80 527
rect 114 493 126 527
rect 68 476 126 493
rect 180 446 238 464
rect 180 412 192 446
rect 226 412 238 446
rect 180 402 238 412
rect 268 374 314 574
rect 564 590 628 596
rect 564 538 570 590
rect 622 538 628 590
rect 564 532 628 538
rect 458 459 734 490
rect 458 425 487 459
rect 521 425 579 459
rect 613 425 671 459
rect 705 425 734 459
rect 458 422 734 425
rect -374 357 -310 364
rect -374 324 -368 357
rect -316 324 -310 357
rect -198 357 -134 364
rect -198 324 -192 357
rect -316 305 -192 324
rect -140 305 -134 357
rect -368 296 -134 305
rect -14 362 88 374
rect -14 328 48 362
rect 82 328 88 362
rect -14 290 88 328
rect 138 362 184 374
rect 138 328 144 362
rect 178 328 184 362
rect 138 308 184 328
rect 234 362 314 374
rect 234 328 240 362
rect 274 328 314 362
rect -14 258 48 290
rect -218 256 48 258
rect 82 256 88 290
rect -218 244 88 256
rect 128 302 194 308
rect 128 250 136 302
rect 188 250 194 302
rect 128 244 194 250
rect 234 290 314 328
rect 234 256 240 290
rect 274 256 314 290
rect 430 394 734 422
rect 234 244 280 256
rect -218 230 36 244
rect -374 224 -308 230
rect -374 172 -366 224
rect -314 172 -308 224
rect -374 166 -308 172
rect -534 -34 -258 -20
rect -534 -51 -342 -34
rect -290 -51 -258 -34
rect -534 -85 -505 -51
rect -471 -85 -413 -51
rect -379 -85 -342 -51
rect -287 -85 -258 -51
rect -534 -86 -342 -85
rect -290 -86 -258 -85
rect -534 -116 -258 -86
rect -218 -120 -190 230
rect 82 206 146 216
rect 82 172 96 206
rect 130 172 402 206
rect 82 154 146 172
rect -2 108 70 120
rect -2 56 8 108
rect 60 56 70 108
rect -2 44 70 56
rect 368 -10 402 172
rect 430 90 458 394
rect 430 80 498 90
rect 430 46 446 80
rect 480 46 498 80
rect 430 32 498 46
rect -158 -38 402 -10
rect -158 -41 -92 -38
rect -158 -75 -142 -41
rect -108 -75 -92 -41
rect -158 -84 -92 -75
rect 76 -93 166 -72
rect -218 -148 -146 -120
rect -192 -169 -146 -148
rect -192 -203 -186 -169
rect -152 -203 -146 -169
rect -192 -241 -146 -203
rect -192 -275 -186 -241
rect -152 -275 -146 -241
rect -192 -322 -146 -275
rect -104 -142 -58 -122
rect 76 -127 105 -93
rect 139 -127 166 -93
rect -104 -148 -36 -142
rect 76 -148 166 -127
rect -104 -169 -96 -148
rect -104 -203 -98 -169
rect -44 -200 -36 -148
rect -64 -203 -36 -200
rect -104 -208 -36 -203
rect 162 -184 220 -182
rect 368 -184 402 -38
rect 488 -41 554 -30
rect 488 -75 504 -41
rect 538 -75 554 -41
rect 488 -86 554 -75
rect 662 -40 1286 -8
rect 662 -43 692 -40
rect 744 -43 1286 -40
rect 662 -77 691 -43
rect 744 -77 783 -43
rect 817 -77 875 -43
rect 909 -45 1286 -43
rect 909 -77 1037 -45
rect 662 -92 692 -77
rect 744 -79 1037 -77
rect 1071 -79 1129 -45
rect 1163 -79 1221 -45
rect 1255 -79 1286 -45
rect 744 -92 1286 -79
rect 662 -110 1286 -92
rect 162 -201 402 -184
rect 446 -128 512 -122
rect 446 -180 454 -128
rect 506 -180 512 -128
rect 446 -186 460 -180
rect -104 -241 -58 -208
rect -104 -275 -98 -241
rect -64 -275 -58 -241
rect 162 -235 174 -201
rect 208 -212 402 -201
rect 454 -203 460 -186
rect 494 -186 512 -180
rect 542 -169 588 -122
rect 494 -203 500 -186
rect 208 -235 400 -212
rect 162 -244 400 -235
rect -104 -322 -58 -275
rect 110 -282 176 -274
rect 24 -286 70 -282
rect -16 -329 70 -286
rect -554 -340 -486 -334
rect -554 -392 -547 -340
rect -495 -346 -486 -340
rect -495 -352 -402 -346
rect -495 -386 -456 -352
rect -422 -386 -402 -352
rect -495 -392 -402 -386
rect -554 -396 -402 -392
rect -158 -369 -92 -358
rect -554 -398 -486 -396
rect -158 -403 -142 -369
rect -108 -403 -92 -369
rect -158 -416 -92 -403
rect -16 -363 30 -329
rect 64 -363 70 -329
rect 110 -334 116 -282
rect 168 -334 176 -282
rect 110 -342 126 -334
rect -16 -401 70 -363
rect -16 -435 30 -401
rect 64 -435 70 -401
rect -16 -482 70 -435
rect 120 -363 126 -342
rect 160 -342 176 -334
rect 216 -329 312 -282
rect 160 -363 166 -342
rect 120 -401 166 -363
rect 120 -435 126 -401
rect 160 -435 166 -401
rect 120 -482 166 -435
rect 216 -363 222 -329
rect 256 -363 312 -329
rect 216 -401 312 -363
rect 216 -435 222 -401
rect 256 -435 312 -401
rect 216 -482 312 -435
rect -16 -536 34 -482
rect -534 -582 -258 -564
rect -534 -595 -411 -582
rect -359 -595 -258 -582
rect -182 -586 -124 -578
rect -534 -629 -505 -595
rect -471 -629 -413 -595
rect -359 -629 -321 -595
rect -287 -629 -258 -595
rect -534 -634 -411 -629
rect -359 -634 -258 -629
rect -534 -660 -258 -634
rect -190 -592 -116 -586
rect -190 -644 -179 -592
rect -127 -644 -116 -592
rect -36 -602 34 -536
rect 66 -529 124 -514
rect 66 -563 78 -529
rect 112 -563 124 -529
rect 66 -580 124 -563
rect -190 -650 -116 -644
rect -182 -656 -124 -650
rect -466 -930 -382 -660
rect -16 -682 34 -602
rect 178 -610 236 -592
rect 178 -644 190 -610
rect 224 -644 236 -610
rect 178 -654 236 -644
rect 266 -682 312 -482
rect -16 -694 86 -682
rect -16 -728 46 -694
rect 80 -728 86 -694
rect -16 -766 86 -728
rect 136 -694 182 -682
rect 136 -728 142 -694
rect 176 -728 182 -694
rect 136 -748 182 -728
rect 232 -694 312 -682
rect 232 -728 238 -694
rect 272 -728 312 -694
rect -16 -800 46 -766
rect 80 -800 86 -766
rect -16 -812 86 -800
rect 126 -754 192 -748
rect 126 -806 134 -754
rect 186 -806 192 -754
rect 126 -812 192 -806
rect 232 -766 312 -728
rect 232 -800 238 -766
rect 272 -800 312 -766
rect 340 -476 400 -244
rect 454 -241 500 -203
rect 454 -275 460 -241
rect 494 -275 500 -241
rect 454 -322 500 -275
rect 542 -203 548 -169
rect 582 -203 588 -169
rect 542 -241 588 -203
rect 542 -275 548 -241
rect 582 -275 588 -241
rect 542 -322 588 -275
rect 1028 -344 1100 -340
rect 488 -369 554 -356
rect 488 -403 504 -369
rect 538 -403 554 -369
rect 488 -412 554 -403
rect 1028 -396 1037 -344
rect 1089 -396 1100 -344
rect 1028 -408 1100 -396
rect 1224 -346 1298 -326
rect 1224 -380 1236 -346
rect 1270 -380 1298 -346
rect 1224 -404 1298 -380
rect 810 -456 868 -442
rect 810 -476 822 -456
rect 340 -490 822 -476
rect 856 -490 868 -456
rect 340 -510 868 -490
rect 232 -812 278 -800
rect 340 -840 400 -510
rect 446 -560 522 -554
rect 446 -612 454 -560
rect 506 -612 522 -560
rect 446 -618 522 -612
rect 662 -587 1284 -556
rect 80 -850 400 -840
rect 80 -884 94 -850
rect 128 -884 400 -850
rect 80 -902 400 -884
rect 662 -621 691 -587
rect 725 -621 783 -587
rect 817 -621 875 -587
rect 909 -589 1284 -587
rect 909 -621 1037 -589
rect 662 -623 1037 -621
rect 1071 -623 1129 -589
rect 1163 -623 1221 -589
rect 1255 -623 1284 -589
rect 662 -654 1284 -623
rect 662 -930 760 -654
rect -566 -959 1322 -930
rect -566 -993 14 -959
rect 48 -993 1322 -959
rect -566 -1004 1322 -993
rect -566 -1120 961 -1004
rect 1269 -1120 1322 -1004
rect -566 -1184 1322 -1120
<< via1 >>
rect 961 1004 1269 1120
rect -154 696 -102 704
rect -154 662 -148 696
rect -148 662 -114 696
rect -114 662 -102 696
rect -154 652 -102 662
rect 118 727 170 774
rect 118 722 128 727
rect 128 722 162 727
rect 162 722 170 727
rect -246 580 -194 592
rect -246 546 -239 580
rect -239 546 -205 580
rect -205 546 -194 580
rect -246 540 -194 546
rect 658 698 710 706
rect 658 664 665 698
rect 665 664 699 698
rect 699 664 710 698
rect 658 654 710 664
rect 570 575 622 590
rect 570 541 579 575
rect 579 541 613 575
rect 613 541 622 575
rect 570 538 622 541
rect -368 305 -316 357
rect -192 305 -140 357
rect 136 290 188 302
rect 136 256 144 290
rect 144 256 178 290
rect 178 256 188 290
rect 136 250 188 256
rect -366 214 -314 224
rect -366 180 -356 214
rect -356 180 -322 214
rect -322 180 -314 214
rect -366 172 -314 180
rect -342 -51 -290 -34
rect -342 -85 -321 -51
rect -321 -85 -290 -51
rect -342 -86 -290 -85
rect 8 97 60 108
rect 8 63 16 97
rect 16 63 50 97
rect 50 63 60 97
rect 8 56 60 63
rect -96 -169 -44 -148
rect -96 -200 -64 -169
rect -64 -200 -44 -169
rect 692 -43 744 -40
rect 692 -77 725 -43
rect 725 -77 744 -43
rect 692 -92 744 -77
rect 454 -169 506 -128
rect 454 -180 460 -169
rect 460 -180 494 -169
rect 494 -180 506 -169
rect -547 -392 -495 -340
rect 116 -329 168 -282
rect 116 -334 126 -329
rect 126 -334 160 -329
rect 160 -334 168 -329
rect -411 -595 -359 -582
rect -411 -629 -379 -595
rect -379 -629 -359 -595
rect -411 -634 -359 -629
rect -179 -600 -127 -592
rect -179 -634 -170 -600
rect -170 -634 -136 -600
rect -136 -634 -127 -600
rect -179 -644 -127 -634
rect 134 -766 186 -754
rect 134 -800 142 -766
rect 142 -800 176 -766
rect 176 -800 186 -766
rect 134 -806 186 -800
rect 1037 -358 1089 -344
rect 1037 -392 1043 -358
rect 1043 -392 1077 -358
rect 1077 -392 1089 -358
rect 1037 -396 1089 -392
rect 454 -572 506 -560
rect 454 -606 462 -572
rect 462 -606 496 -572
rect 496 -606 506 -572
rect 454 -612 506 -606
rect 961 -1120 1269 -1004
<< metal2 >>
rect 940 1120 1290 1134
rect 940 1004 961 1120
rect 1269 1004 1290 1120
rect 940 990 1290 1004
rect -566 816 1322 844
rect -124 710 -96 816
rect 112 774 178 782
rect 112 722 118 774
rect 170 722 178 774
rect 112 714 178 722
rect -164 704 -96 710
rect -164 652 -154 704
rect -102 652 -96 704
rect -164 646 -96 652
rect -254 592 -186 598
rect -254 540 -246 592
rect -194 540 -186 592
rect -254 530 -186 540
rect -374 357 -310 364
rect -374 326 -368 357
rect -566 305 -368 326
rect -316 305 -310 357
rect -566 298 -310 305
rect -566 296 -368 298
rect -566 290 -374 296
rect -374 224 -308 230
rect -374 172 -366 224
rect -314 172 -308 224
rect -374 166 -308 172
rect -374 44 -346 166
rect -414 16 -346 44
rect -554 -340 -486 -334
rect -554 -392 -547 -340
rect -495 -392 -486 -340
rect -554 -398 -486 -392
rect -554 -1014 -510 -398
rect -414 -568 -386 16
rect -352 -34 -290 -28
rect -352 -86 -342 -34
rect -254 -42 -226 530
rect -198 357 -134 364
rect -198 305 -192 357
rect -140 324 -134 357
rect 128 324 178 714
rect 650 712 678 816
rect 650 706 716 712
rect 650 692 658 706
rect 652 654 658 692
rect 710 654 716 706
rect 652 648 716 654
rect 564 590 628 596
rect 564 560 570 590
rect 354 538 570 560
rect 622 538 628 590
rect 354 532 628 538
rect -140 308 180 324
rect -140 305 194 308
rect -198 302 194 305
rect -198 296 136 302
rect 128 250 136 296
rect 188 250 194 302
rect 128 244 194 250
rect -2 108 70 120
rect -2 56 8 108
rect 60 56 70 108
rect -2 44 70 56
rect 34 42 70 44
rect -254 -70 34 -42
rect -352 -92 -290 -86
rect -318 -138 -290 -92
rect -318 -142 -74 -138
rect -318 -148 -36 -142
rect -318 -166 -96 -148
rect -102 -200 -96 -166
rect -44 -200 -36 -148
rect -102 -208 -36 -200
rect -414 -582 -350 -568
rect 6 -576 34 -70
rect 110 -282 176 -274
rect 110 -334 116 -282
rect 168 -334 176 -282
rect 110 -342 176 -334
rect -414 -634 -411 -582
rect -359 -634 -350 -582
rect -414 -650 -350 -634
rect -180 -592 34 -576
rect -180 -644 -179 -592
rect -127 -604 34 -592
rect -127 -644 -126 -604
rect -180 -660 -126 -644
rect 126 -748 176 -342
rect 354 -586 382 532
rect 786 290 1322 326
rect 686 -40 750 -32
rect 686 -92 692 -40
rect 744 -92 750 -40
rect 686 -100 750 -92
rect 446 -128 512 -122
rect 446 -180 454 -128
rect 506 -158 512 -128
rect 686 -158 714 -100
rect 506 -180 714 -158
rect 446 -186 714 -180
rect 786 -336 814 290
rect 786 -344 1098 -336
rect 786 -372 1037 -344
rect 446 -560 522 -554
rect 446 -586 454 -560
rect 354 -612 454 -586
rect 506 -612 522 -560
rect 354 -614 522 -612
rect 446 -618 522 -614
rect 126 -754 192 -748
rect 126 -806 134 -754
rect 186 -776 192 -754
rect 786 -776 814 -372
rect 1018 -396 1037 -372
rect 1089 -396 1098 -344
rect 1018 -408 1098 -396
rect 186 -804 814 -776
rect 186 -806 192 -804
rect 126 -812 192 -806
rect 940 -1004 1290 -990
rect 940 -1120 961 -1004
rect 1269 -1120 1290 -1004
rect 940 -1134 1290 -1120
<< via2 >>
rect 967 1034 1023 1090
rect 1047 1034 1103 1090
rect 1127 1034 1183 1090
rect 1207 1034 1263 1090
rect 967 -1090 1023 -1034
rect 1047 -1090 1103 -1034
rect 1127 -1090 1183 -1034
rect 1207 -1090 1263 -1034
<< metal3 >>
rect -574 1090 1322 1192
rect -574 1034 967 1090
rect 1023 1034 1047 1090
rect 1103 1034 1127 1090
rect 1183 1034 1207 1090
rect 1263 1034 1322 1090
rect -574 938 1322 1034
rect -566 -1034 1322 -930
rect -566 -1090 967 -1034
rect 1023 -1090 1047 -1034
rect 1103 -1090 1127 -1034
rect 1183 -1090 1207 -1034
rect 1263 -1090 1322 -1034
rect -566 -1185 1322 -1090
<< labels >>
flabel metal2 -566 290 -374 326 1 FreeSans 800 0 0 0 IN
port 1 n
flabel metal2 786 290 1322 326 1 FreeSans 800 0 0 0 OUT
port 6 n
flabel metal3 -574 938 967 1192 1 FreeSans 800 0 0 0 VDD
port 5 n
flabel metal3 -566 -1184 961 -930 1 FreeSans 800 0 0 0 VSS
port 4 n
flabel metal2 -554 -1014 -510 -392 1 FreeSans 800 0 0 0 C
port 2 n
flabel metal2 -566 816 1322 844 1 FreeSans 800 0 0 0 RESET
port 3 n
flabel metal1 1270 -404 1298 -326 1 FreeSans 800 0 0 0 buf_out
port 7 n
<< end >>
