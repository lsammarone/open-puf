magic
tech sky130B
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__hvdfm1sd2__example_55959141808449  sky130_fd_pr__hvdfm1sd2__example_55959141808449_0
timestamp 1648127584
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808449  sky130_fd_pr__hvdfm1sd2__example_55959141808449_1
timestamp 1648127584
transform 1 0 160 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 188 85 188 85 0 FreeSans 300 0 0 0 D
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 27731252
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27730194
<< end >>
