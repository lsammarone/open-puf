magic
tech sky130A
magscale 1 2
timestamp 1654298126
<< nwell >>
rect 30250 -2656 30362 -2335
rect 30529 -2656 30618 -2335
<< viali >>
rect 27523 -2576 27557 -2542
rect 29040 -2563 29074 -2529
rect 29208 -2563 29242 -2529
rect 29376 -2563 29410 -2529
rect 29544 -2563 29578 -2529
rect 29712 -2563 29746 -2529
rect 29880 -2563 29914 -2529
rect 30048 -2563 30082 -2529
rect 30788 -2564 30822 -2530
rect 30956 -2564 30990 -2530
rect 31124 -2564 31158 -2530
rect 31292 -2564 31326 -2530
rect 31460 -2564 31494 -2530
rect 31628 -2564 31662 -2530
rect 31796 -2564 31830 -2530
rect 27337 -2702 27371 -2668
rect 27871 -2694 27905 -2660
rect 28599 -2703 28633 -2669
rect 28800 -2698 28834 -2664
rect 28919 -2698 28953 -2664
rect 29038 -2698 29072 -2664
rect 29157 -2698 29191 -2664
rect 29276 -2698 29310 -2664
rect 29395 -2698 29429 -2664
rect 29514 -2698 29548 -2664
rect 30724 -2696 30758 -2662
rect 30843 -2696 30877 -2662
rect 30962 -2696 30996 -2662
rect 31081 -2696 31115 -2662
rect 31200 -2696 31234 -2662
rect 31319 -2696 31353 -2662
rect 31438 -2696 31472 -2662
<< metal1 >>
rect 86 1593 444 1613
rect 86 1592 386 1593
rect 86 1540 110 1592
rect 162 1541 386 1592
rect 438 1541 444 1593
rect 162 1540 444 1541
rect 86 1516 444 1540
rect 27760 -2421 27836 -2325
rect 28664 -2421 28740 -2325
rect 30212 -2421 30399 -2325
rect 30491 -2421 30678 -2325
rect 27513 -2542 27566 -2525
rect 27513 -2576 27523 -2542
rect 27557 -2576 27566 -2542
rect -317 -2668 27389 -2646
rect -317 -2702 27337 -2668
rect 27371 -2702 27389 -2668
rect -317 -2720 27389 -2702
rect 27513 -2647 27566 -2576
rect 29028 -2529 31845 -2504
rect 29028 -2563 29040 -2529
rect 29074 -2563 29208 -2529
rect 29242 -2563 29376 -2529
rect 29410 -2563 29544 -2529
rect 29578 -2563 29712 -2529
rect 29746 -2563 29880 -2529
rect 29914 -2563 30048 -2529
rect 30082 -2530 31845 -2529
rect 30082 -2538 30788 -2530
rect 30082 -2563 30260 -2538
rect 29028 -2590 30260 -2563
rect 30312 -2590 30363 -2538
rect 30415 -2590 30466 -2538
rect 30518 -2590 30569 -2538
rect 30621 -2564 30788 -2538
rect 30822 -2564 30956 -2530
rect 30990 -2564 31124 -2530
rect 31158 -2564 31292 -2530
rect 31326 -2564 31460 -2530
rect 31494 -2564 31628 -2530
rect 31662 -2564 31796 -2530
rect 31830 -2564 31845 -2530
rect 30621 -2590 31845 -2564
rect 29028 -2612 31845 -2590
rect 27513 -2660 27923 -2647
rect 27513 -2694 27871 -2660
rect 27905 -2694 27923 -2660
rect 27513 -2708 27923 -2694
rect 28577 -2662 31768 -2653
rect 28577 -2664 30724 -2662
rect 28577 -2669 28800 -2664
rect 28577 -2703 28599 -2669
rect 28633 -2698 28800 -2669
rect 28834 -2698 28919 -2664
rect 28953 -2698 29038 -2664
rect 29072 -2698 29157 -2664
rect 29191 -2698 29276 -2664
rect 29310 -2698 29395 -2664
rect 29429 -2698 29514 -2664
rect 29548 -2696 30724 -2664
rect 30758 -2696 30843 -2662
rect 30877 -2696 30962 -2662
rect 30996 -2696 31081 -2662
rect 31115 -2696 31200 -2662
rect 31234 -2696 31319 -2662
rect 31353 -2696 31438 -2662
rect 31472 -2696 31768 -2662
rect 29548 -2698 31768 -2696
rect 28633 -2703 31768 -2698
rect 28577 -2710 31768 -2703
rect 27760 -2965 27836 -2869
rect 28664 -2966 28740 -2870
rect 30212 -2965 30399 -2869
rect 30491 -2965 30678 -2869
rect -167 -6186 614 -6171
rect -167 -6194 555 -6186
rect -167 -6246 -150 -6194
rect -98 -6238 555 -6194
rect 607 -6238 614 -6186
rect -98 -6246 614 -6238
rect -167 -6264 614 -6246
<< via1 >>
rect 30296 3154 30348 3206
rect 30413 3154 30465 3206
rect 30530 3154 30582 3206
rect 110 1540 162 1592
rect 386 1541 438 1593
rect 31363 -2407 31415 -2355
rect 31493 -2407 31545 -2355
rect 31623 -2407 31675 -2355
rect 30260 -2590 30312 -2538
rect 30363 -2590 30415 -2538
rect 30466 -2590 30518 -2538
rect 30569 -2590 30621 -2538
rect 31353 -2937 31405 -2885
rect 31466 -2937 31518 -2885
rect 31579 -2937 31631 -2885
rect 31692 -2937 31744 -2885
rect 31805 -2937 31857 -2885
rect 31353 -4826 31405 -4774
rect 31466 -4826 31518 -4774
rect 31579 -4826 31631 -4774
rect 31692 -4826 31744 -4774
rect 31805 -4826 31857 -4774
rect 31353 -4931 31405 -4879
rect 31466 -4931 31518 -4879
rect 31579 -4931 31631 -4879
rect 31692 -4931 31744 -4879
rect 31805 -4931 31857 -4879
rect -150 -6246 -98 -6194
rect 555 -6238 607 -6186
rect 30285 -9075 30337 -9023
rect 30368 -9075 30420 -9023
rect 30451 -9075 30503 -9023
rect 30534 -9075 30586 -9023
<< metal2 >>
rect 60942 6037 60978 6070
rect -159 6001 555 6037
rect 60231 6001 60978 6037
rect -159 -6171 -123 6001
rect 30232 3261 30628 3290
rect 30232 3205 30263 3261
rect 30319 3206 30372 3261
rect 30428 3206 30481 3261
rect 30537 3206 30628 3261
rect 30348 3205 30372 3206
rect 30465 3205 30481 3206
rect 30232 3159 30296 3205
rect 30348 3159 30413 3205
rect 30465 3159 30530 3205
rect 30232 3103 30263 3159
rect 30348 3154 30372 3159
rect 30465 3154 30481 3159
rect 30582 3154 30628 3206
rect 30319 3103 30372 3154
rect 30428 3103 30481 3154
rect 30537 3103 30628 3154
rect 30232 3082 30628 3103
rect 75 1592 173 1619
rect 75 1540 110 1592
rect 162 1540 173 1592
rect 75 1500 173 1540
rect 373 1593 477 1616
rect 373 1541 386 1593
rect 438 1581 477 1593
rect 60942 1581 60978 6001
rect 438 1545 649 1581
rect 60325 1545 60978 1581
rect 438 1541 477 1545
rect 373 1516 477 1541
rect -160 -6194 -49 -6171
rect -160 -6246 -150 -6194
rect -98 -6246 -49 -6194
rect -160 -6286 -49 -6246
rect 107 -10650 143 1500
rect 30233 -1921 30630 -1882
rect 30233 -1977 30256 -1921
rect 30312 -1977 30360 -1921
rect 30416 -1977 30464 -1921
rect 30520 -1977 30568 -1921
rect 30624 -1977 30630 -1921
rect 30233 -2020 30630 -1977
rect 30233 -2076 30256 -2020
rect 30312 -2076 30360 -2020
rect 30416 -2076 30464 -2020
rect 30520 -2076 30568 -2020
rect 30624 -2076 30630 -2020
rect 30233 -2538 30630 -2076
rect 31324 -2351 31725 -2326
rect 31324 -2407 31363 -2351
rect 31419 -2407 31492 -2351
rect 31548 -2407 31621 -2351
rect 31677 -2407 31725 -2351
rect 31324 -2420 31725 -2407
rect 30233 -2590 30260 -2538
rect 30312 -2590 30363 -2538
rect 30415 -2590 30466 -2538
rect 30518 -2590 30569 -2538
rect 30621 -2590 30630 -2538
rect 30233 -3250 30630 -2590
rect 30233 -3306 30269 -3250
rect 30325 -3306 30357 -3250
rect 30413 -3306 30445 -3250
rect 30501 -3306 30533 -3250
rect 30589 -3306 30630 -3250
rect 30233 -3345 30630 -3306
rect 30233 -3401 30269 -3345
rect 30325 -3401 30357 -3345
rect 30413 -3401 30445 -3345
rect 30501 -3401 30533 -3345
rect 30589 -3401 30630 -3345
rect 30233 -3432 30630 -3401
rect 31298 -2885 31965 -2868
rect 31298 -2937 31353 -2885
rect 31405 -2937 31466 -2885
rect 31518 -2937 31579 -2885
rect 31631 -2937 31692 -2885
rect 31744 -2937 31805 -2885
rect 31857 -2937 31965 -2885
rect 31298 -4774 31965 -2937
rect 31298 -4826 31353 -4774
rect 31405 -4826 31466 -4774
rect 31518 -4826 31579 -4774
rect 31631 -4826 31692 -4774
rect 31744 -4826 31805 -4774
rect 31857 -4826 31965 -4774
rect 31298 -4879 31965 -4826
rect 31298 -4931 31353 -4879
rect 31405 -4931 31466 -4879
rect 31518 -4931 31579 -4879
rect 31631 -4931 31692 -4879
rect 31744 -4931 31805 -4879
rect 31857 -4931 31965 -4879
rect 31298 -4979 31965 -4931
rect 548 -6186 618 -6165
rect 548 -6238 555 -6186
rect 607 -6194 618 -6186
rect 607 -6230 878 -6194
rect 60554 -6230 61279 -6194
rect 607 -6238 618 -6230
rect 548 -6269 618 -6238
rect 30233 -8974 30630 -8941
rect 30233 -9030 30274 -8974
rect 30330 -9023 30366 -8974
rect 30422 -9023 30458 -8974
rect 30514 -9023 30550 -8974
rect 30337 -9030 30366 -9023
rect 30422 -9030 30451 -9023
rect 30514 -9030 30534 -9023
rect 30606 -9030 30630 -8974
rect 30233 -9065 30285 -9030
rect 30337 -9065 30368 -9030
rect 30420 -9065 30451 -9030
rect 30503 -9065 30534 -9030
rect 30586 -9065 30630 -9030
rect 30233 -9121 30274 -9065
rect 30337 -9075 30366 -9065
rect 30422 -9075 30451 -9065
rect 30514 -9075 30534 -9065
rect 30330 -9121 30366 -9075
rect 30422 -9121 30458 -9075
rect 30514 -9121 30550 -9075
rect 30606 -9121 30630 -9065
rect 30233 -9147 30630 -9121
rect 61243 -10650 61279 -6230
rect 107 -10686 784 -10650
rect 60460 -10686 61279 -10650
rect 61243 -10697 61279 -10686
<< via2 >>
rect 30263 3206 30319 3261
rect 30372 3206 30428 3261
rect 30481 3206 30537 3261
rect 30263 3205 30296 3206
rect 30296 3205 30319 3206
rect 30372 3205 30413 3206
rect 30413 3205 30428 3206
rect 30481 3205 30530 3206
rect 30530 3205 30537 3206
rect 30263 3154 30296 3159
rect 30296 3154 30319 3159
rect 30372 3154 30413 3159
rect 30413 3154 30428 3159
rect 30481 3154 30530 3159
rect 30530 3154 30537 3159
rect 30263 3103 30319 3154
rect 30372 3103 30428 3154
rect 30481 3103 30537 3154
rect 30256 -1977 30312 -1921
rect 30360 -1977 30416 -1921
rect 30464 -1977 30520 -1921
rect 30568 -1977 30624 -1921
rect 30256 -2076 30312 -2020
rect 30360 -2076 30416 -2020
rect 30464 -2076 30520 -2020
rect 30568 -2076 30624 -2020
rect 31363 -2355 31419 -2351
rect 31363 -2407 31415 -2355
rect 31415 -2407 31419 -2355
rect 31492 -2355 31548 -2351
rect 31492 -2407 31493 -2355
rect 31493 -2407 31545 -2355
rect 31545 -2407 31548 -2355
rect 31621 -2355 31677 -2351
rect 31621 -2407 31623 -2355
rect 31623 -2407 31675 -2355
rect 31675 -2407 31677 -2355
rect 30269 -3306 30325 -3250
rect 30357 -3306 30413 -3250
rect 30445 -3306 30501 -3250
rect 30533 -3306 30589 -3250
rect 30269 -3401 30325 -3345
rect 30357 -3401 30413 -3345
rect 30445 -3401 30501 -3345
rect 30533 -3401 30589 -3345
rect 30274 -9023 30330 -8974
rect 30366 -9023 30422 -8974
rect 30458 -9023 30514 -8974
rect 30550 -9023 30606 -8974
rect 30274 -9030 30285 -9023
rect 30285 -9030 30330 -9023
rect 30366 -9030 30368 -9023
rect 30368 -9030 30420 -9023
rect 30420 -9030 30422 -9023
rect 30458 -9030 30503 -9023
rect 30503 -9030 30514 -9023
rect 30550 -9030 30586 -9023
rect 30586 -9030 30606 -9023
rect 30274 -9075 30285 -9065
rect 30285 -9075 30330 -9065
rect 30366 -9075 30368 -9065
rect 30368 -9075 30420 -9065
rect 30420 -9075 30422 -9065
rect 30458 -9075 30503 -9065
rect 30503 -9075 30514 -9065
rect 30550 -9075 30586 -9065
rect 30586 -9075 30606 -9065
rect 30274 -9121 30330 -9075
rect 30366 -9121 30422 -9075
rect 30458 -9121 30514 -9075
rect 30550 -9121 30606 -9075
<< metal3 >>
rect 30232 3261 30627 3290
rect 30232 3205 30263 3261
rect 30319 3238 30372 3261
rect 30428 3205 30481 3261
rect 30537 3205 30627 3261
rect 30232 3159 30306 3205
rect 30402 3159 30627 3205
rect 30232 3103 30263 3159
rect 30319 3103 30372 3130
rect 30428 3103 30481 3159
rect 30537 3103 30627 3159
rect 30232 3082 30627 3103
rect 30 -135 530 -75
rect 30 -277 530 -217
rect 30 -419 530 -359
rect 30 -561 530 -501
rect 30 -703 530 -643
rect 30 -845 530 -785
rect 30 -987 530 -927
rect 30 -1129 530 -1069
rect 30 -1271 530 -1211
rect 30 -1413 530 -1353
rect 30 -1555 530 -1495
rect 30 -1697 530 -1637
rect 30 -1839 530 -1779
rect 30232 -1921 30629 -1879
rect 30 -1981 530 -1921
rect 30232 -1977 30256 -1921
rect 30312 -1946 30360 -1921
rect 30416 -1977 30464 -1921
rect 30520 -1946 30568 -1921
rect 30624 -1977 30629 -1921
rect 30232 -2020 30297 -1977
rect 30393 -2020 30479 -1977
rect 30575 -2020 30629 -1977
rect 30 -2123 530 -2063
rect 30232 -2076 30256 -2020
rect 30312 -2076 30360 -2054
rect 30416 -2076 30464 -2020
rect 30520 -2076 30568 -2054
rect 30624 -2076 30629 -2020
rect 30232 -2103 30629 -2076
rect 30 -2265 530 -2205
rect 31324 -2337 31725 -2326
rect 30 -2407 530 -2347
rect 31324 -2351 31445 -2337
rect 31619 -2351 31725 -2337
rect 31324 -2407 31363 -2351
rect 31419 -2401 31445 -2351
rect 31619 -2401 31621 -2351
rect 31419 -2407 31492 -2401
rect 31548 -2407 31621 -2401
rect 31677 -2407 31725 -2351
rect 31324 -2420 31725 -2407
rect 30 -2549 530 -2489
rect 30 -2691 530 -2631
rect 30 -2833 530 -2773
rect 30 -2975 530 -2915
rect 30 -3117 530 -3057
rect 30 -3259 530 -3199
rect 30233 -3250 30630 -3192
rect 30233 -3306 30269 -3250
rect 30325 -3269 30357 -3250
rect 30413 -3306 30445 -3250
rect 30501 -3269 30533 -3250
rect 30589 -3306 30630 -3250
rect 30 -3401 530 -3341
rect 30233 -3345 30289 -3306
rect 30385 -3345 30479 -3306
rect 30575 -3345 30630 -3306
rect 30233 -3401 30269 -3345
rect 30325 -3401 30357 -3377
rect 30413 -3401 30445 -3345
rect 30501 -3401 30533 -3377
rect 30589 -3401 30630 -3345
rect 30233 -3432 30630 -3401
rect 30 -3543 530 -3483
rect 30 -3685 530 -3625
rect 30 -3827 530 -3767
rect 30 -3969 530 -3909
rect 30 -4111 530 -4051
rect 30 -4253 530 -4193
rect 30 -4395 530 -4335
rect 30 -4537 530 -4477
rect 30233 -8974 30630 -8941
rect 30233 -9030 30274 -8974
rect 30330 -8998 30366 -8974
rect 30422 -9030 30458 -8974
rect 30514 -8997 30550 -8974
rect 30606 -9030 30630 -8974
rect 30233 -9065 30301 -9030
rect 30397 -9065 30475 -9030
rect 30571 -9065 30630 -9030
rect 30233 -9121 30274 -9065
rect 30330 -9121 30366 -9106
rect 30422 -9121 30458 -9065
rect 30514 -9121 30550 -9105
rect 30606 -9121 30630 -9065
rect 30233 -9147 30630 -9121
<< via3 >>
rect 30306 3205 30319 3238
rect 30319 3205 30372 3238
rect 30372 3205 30402 3238
rect 30306 3159 30402 3205
rect 30306 3130 30319 3159
rect 30319 3130 30372 3159
rect 30372 3130 30402 3159
rect 31369 2236 31493 2402
rect 31568 2236 31692 2402
rect 30297 -1977 30312 -1946
rect 30312 -1977 30360 -1946
rect 30360 -1977 30393 -1946
rect 30479 -1977 30520 -1946
rect 30520 -1977 30568 -1946
rect 30568 -1977 30575 -1946
rect 30297 -2020 30393 -1977
rect 30479 -2020 30575 -1977
rect 30297 -2054 30312 -2020
rect 30312 -2054 30360 -2020
rect 30360 -2054 30393 -2020
rect 30479 -2054 30520 -2020
rect 30520 -2054 30568 -2020
rect 30568 -2054 30575 -2020
rect 31445 -2351 31619 -2337
rect 31445 -2401 31492 -2351
rect 31492 -2401 31548 -2351
rect 31548 -2401 31619 -2351
rect 30289 -3306 30325 -3269
rect 30325 -3306 30357 -3269
rect 30357 -3306 30385 -3269
rect 30479 -3306 30501 -3269
rect 30501 -3306 30533 -3269
rect 30533 -3306 30575 -3269
rect 30289 -3345 30385 -3306
rect 30479 -3345 30575 -3306
rect 30289 -3377 30325 -3345
rect 30325 -3377 30357 -3345
rect 30357 -3377 30385 -3345
rect 30479 -3377 30501 -3345
rect 30501 -3377 30533 -3345
rect 30533 -3377 30575 -3345
rect 30301 -9030 30330 -8998
rect 30330 -9030 30366 -8998
rect 30366 -9030 30397 -8998
rect 30475 -9030 30514 -8997
rect 30514 -9030 30550 -8997
rect 30550 -9030 30571 -8997
rect 30301 -9065 30397 -9030
rect 30475 -9065 30571 -9030
rect 30301 -9106 30330 -9065
rect 30330 -9106 30366 -9065
rect 30366 -9106 30397 -9065
rect 30475 -9105 30514 -9065
rect 30514 -9105 30550 -9065
rect 30550 -9105 30571 -9065
<< metal4 >>
rect 30232 3238 30629 3350
rect 30232 3130 30306 3238
rect 30402 3130 30629 3238
rect 30232 -1442 30629 3130
rect 30231 -1803 30629 -1442
rect 30232 -1946 30629 -1803
rect 30232 -2054 30297 -1946
rect 30393 -2054 30479 -1946
rect 30575 -2054 30629 -1946
rect 30232 -2103 30629 -2054
rect 31317 2402 31721 2521
rect 31317 2236 31369 2402
rect 31493 2236 31568 2402
rect 31692 2236 31721 2402
rect 31317 -2017 31721 2236
rect 31317 -2148 31725 -2017
rect 31324 -2337 31725 -2148
rect 31324 -2401 31445 -2337
rect 31619 -2401 31725 -2337
rect 31324 -2420 31725 -2401
rect 30234 -3269 30630 -3193
rect 30234 -3377 30289 -3269
rect 30385 -3377 30479 -3269
rect 30575 -3377 30630 -3269
rect 30234 -8997 30630 -3377
rect 30234 -8998 30475 -8997
rect 30234 -9106 30301 -8998
rect 30397 -9105 30475 -8998
rect 30571 -9105 30630 -8997
rect 30397 -9106 30630 -9105
rect 30234 -9209 30630 -9106
use BR128half  BR128half_0
timestamp 1654224521
transform 1 0 449 0 1 71
box -430 -58 60604 7443
use BR128half  BR128half_1
timestamp 1654224521
transform -1 0 60660 0 1 -12160
box -430 -58 60604 7443
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 27300 0 1 -2917
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1650294714
transform 1 0 27836 0 1 -2917
box -38 -48 866 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654066915
transform 1 0 28740 0 1 -2917
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654066915
transform 1 0 30656 0 1 -2917
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 30399 0 1 -2917
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1650294714
transform 1 0 27668 0 1 -2917
box -38 -48 130 592
<< end >>
