magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 1 21 355 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
<< ndiff >>
rect 27 127 79 177
rect 27 93 35 127
rect 69 93 79 127
rect 27 47 79 93
rect 109 95 163 177
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 127 247 177
rect 193 93 203 127
rect 237 93 247 127
rect 193 47 247 93
rect 277 95 329 177
rect 277 61 287 95
rect 321 61 329 95
rect 277 47 329 61
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 163 497
rect 193 297 247 497
rect 277 485 329 497
rect 277 451 287 485
rect 321 451 329 485
rect 277 417 329 451
rect 277 383 287 417
rect 321 383 329 417
rect 277 297 329 383
<< ndiffc >>
rect 35 93 69 127
rect 119 61 153 95
rect 203 93 237 127
rect 287 61 321 95
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 287 451 321 485
rect 287 383 321 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 25 249 109 265
rect 25 215 35 249
rect 69 215 109 249
rect 25 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 249 341 265
rect 247 215 297 249
rect 331 215 341 249
rect 247 199 341 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
<< polycont >>
rect 35 215 69 249
rect 161 215 195 249
rect 297 215 331 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 18 485 234 490
rect 18 451 35 485
rect 69 456 234 485
rect 69 451 85 456
rect 18 417 85 451
rect 18 383 35 417
rect 69 383 85 417
rect 18 349 85 383
rect 18 315 35 349
rect 69 315 85 349
rect 18 299 85 315
rect 119 265 166 401
rect 200 333 234 456
rect 287 485 350 527
rect 321 451 350 485
rect 287 417 350 451
rect 321 383 350 417
rect 287 367 350 383
rect 200 299 263 333
rect 18 249 85 265
rect 18 215 35 249
rect 69 215 85 249
rect 18 199 85 215
rect 119 249 195 265
rect 119 215 161 249
rect 119 199 195 215
rect 229 165 263 299
rect 18 131 263 165
rect 297 249 351 333
rect 331 215 351 249
rect 297 131 351 215
rect 18 127 69 131
rect 18 93 35 127
rect 203 127 237 131
rect 18 77 69 93
rect 103 95 169 97
rect 103 61 119 95
rect 153 61 169 95
rect 203 77 237 93
rect 271 95 337 97
rect 103 17 169 61
rect 271 61 287 95
rect 321 61 337 95
rect 271 17 337 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 30 425 64 459 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 306 153 340 187 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor3_1
rlabel metal1 s 0 -48 368 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 2013464
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2009284
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.200 0.000 
<< end >>
