/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/sonos/end_of_life/typical/tt.spice