* NGSPICE file created from BR64_flat.ext - technology: sky130A

.subckt BR64_flat OUT C[63] C[62] C[61] C[60] C[59] C[58] C[57] C[56] C[55] C[54]
+ C[53] C[52] C[51] C[50] C[49] C[48] C[47] C[46] C[45] C[44] C[43] C[42] C[41] C[40]
+ C[39] C[38] C[37] C[36] C[35] C[34] C[33] C[32] C[31] C[30] C[29] C[28] C[27] C[26]
+ C[25] C[24] C[23] C[22] C[21] C[20] C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12]
+ C[11] C[10] C[9] C[8] C[7] C[6] C[5] C[4] C[3] C[2] C[1] C[0] RESET VDD VSS
X0 VSS a_10234_5882# a_10236_6938# VSS sky130_fd_pr__nfet_01v8 ad=1.07957e+14p pd=1.15496e+09u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X2 a_2668_702# a_2078_619# a_2572_702# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X3 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=1.69742e+14p ps=1.6004e+09u w=1e+06u l=150000u
X4 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X5 a_14313_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_2668_702# a_2304_765# a_2572_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X7 a_27110_702# a_28504_619# a_28554_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X8 VDD a_684_702# a_1609_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X9 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X10 a_26753_1923# a_26666_1825# a_26671_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X11 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VSS a_45669_1861# a_59296_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X13 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X14 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_59310_5882# a_58544_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X17 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X18 VSS a_5349_6584# a_5299_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X19 a_10537_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X20 a_43689_5637# a_43716_6378# a_43701_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X21 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X22 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.32e+12p ps=4.064e+07u w=1e+06u l=150000u
X24 a_10222_1758# a_9630_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X25 VDD a_45669_1861# a_53993_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X26 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X27 VSS a_20842_6337# a_20790_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X28 a_42310_702# a_42312_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X29 a_n225_6339# a_190_619# a_240_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X30 VSS a_39722_6337# a_39670_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X31 VDD a_38438_702# a_39363_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X32 a_57769_1923# a_57410_1758# a_57408_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X33 a_19558_702# a_21178_765# a_21002_1825# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X34 a_45583_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X35 a_15343_1923# a_15338_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X36 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X37 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X38 VDD a_24223_6584# a_24173_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X39 a_2572_702# a_2304_765# a_2133_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X40 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X41 a_43689_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X42 a_32872_1758# a_32280_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X43 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X44 VDD a_30571_1861# a_39969_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X45 a_21558_6938# a_20790_6363# a_19572_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X46 a_29110_6938# a_28394_6337# a_27124_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X47 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_15288_619# C[40] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X49 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X51 a_43745_1923# a_43658_1825# a_43663_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X52 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.808e+12p ps=2.944e+07u w=650000u l=150000u
X53 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X54 a_19572_5882# a_18954_6337# a_19172_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X55 VSS RESET sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X56 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=4.32e+12p pd=4.064e+07u as=0p ps=0u w=1e+06u l=150000u
X57 a_2586_5882# a_3856_6337# a_4047_5637# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X58 a_3966_619# C[34] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X59 a_18083_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X60 VDD a_40058_765# a_39882_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X61 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X62 VSS a_45669_1861# a_49321_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X63 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X64 a_18765_625# a_18595_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X65 VDD a_14783_6584# a_14733_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X66 a_34760_1758# a_34394_765# a_32774_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X67 a_6362_5882# a_7580_6363# a_7823_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X68 a_42326_6938# a_41558_6363# a_40340_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X69 a_47459_5637# a_47486_6378# a_47471_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X70 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 a_n315_6584# a_n225_6339# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X73 a_58932_765# a_58706_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X74 a_32335_1923# a_32330_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X75 VDD a_30571_1861# a_30529_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X76 a_46080_702# a_46082_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X77 VDD a_41215_6584# a_41165_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X78 VSS a_54425_6584# a_54375_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X79 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X80 VDD a_13900_702# a_14825_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X81 VDD a_43498_6337# a_43446_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X82 a_19656_1758# a_19064_619# a_17670_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X83 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X84 a_42214_702# a_41946_765# a_41775_1923# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X85 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X86 VSS C[25] a_11408_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X87 a_47459_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X88 a_11219_625# a_11049_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X89 a_36564_5882# a_35946_6337# a_36164_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X90 a_47872_702# a_49266_619# a_49316_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X91 a_35075_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X92 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X93 a_55438_5882# a_56708_6337# a_56899_5637# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X94 VSS a_45380_6337# a_45328_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X95 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X96 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X97 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X98 a_21460_5882# a_20790_6363# a_21060_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X99 VSS a_49760_702# a_50685_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X100 VDD a_31775_6584# a_31725_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X101 VSS a_44985_6584# a_44935_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X102 a_4021_1923# a_4016_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X103 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X104 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X105 a_5991_1923# a_5904_1825# a_5909_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X106 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 a_25332_5882# a_24566_6363# a_25236_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X108 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X109 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X110 a_13406_619# C[39] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X111 a_37439_6584# a_36564_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X112 a_46096_6938# a_45328_6363# a_44116_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X113 VSS a_2682_5882# a_2684_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X114 a_36648_1758# a_36056_619# a_34662_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X115 VSS a_15467_1861# a_19654_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X116 a_8250_5882# a_7632_6337# a_7850_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X117 a_40422_702# a_40058_765# a_40326_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X118 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X119 a_36662_6938# a_36660_5882# a_36963_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X120 VDD a_47268_6337# a_47216_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X121 a_21859_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X122 VDD a_32506_765# a_32330_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X123 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.16e+12p pd=2.032e+07u as=0p ps=0u w=1e+06u l=150000u
X124 VDD a_3461_6584# a_3411_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X125 VSS a_21556_5882# a_21558_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X126 a_53632_702# a_53634_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X127 a_15892_5882# a_15126_6363# a_15796_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X128 a_11611_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X129 a_2078_619# C[33] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X130 a_34394_765# a_34168_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X131 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X132 a_9685_1923# a_9680_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X133 VDD a_369_1861# a_7879_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X134 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_9125_6584# a_8250_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X136 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X137 a_36282_765# a_36056_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X138 VDD a_40326_702# a_41251_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X139 VDD a_55156_765# a_54980_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X140 a_8334_1758# a_7742_619# a_6348_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X141 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X142 a_40326_702# a_39832_619# a_39887_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X143 a_19668_5882# a_18954_6337# a_19572_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X144 a_4572_6938# a_3856_6337# a_2586_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X145 VDD a_1968_6337# a_1916_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X146 a_53097_1923# a_53092_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X147 a_27222_6938# a_27220_5882# a_27523_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X148 VDD a_45669_1861# a_51291_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X149 a_42627_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X150 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X151 VSS C[12] a_35946_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X152 a_54631_625# a_54461_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X153 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X154 a_29094_702# a_28504_619# a_28998_702# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X155 a_5555_625# a_5385_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X156 a_29094_702# a_28730_765# a_28998_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X157 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=1.404e+12p pd=1.472e+07u as=0p ps=0u w=650000u l=150000u
X159 a_41720_619# C[54] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X160 VDD a_28998_702# a_29923_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X161 a_29108_5882# a_28342_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X162 a_13487_5637# a_13514_6378# a_13499_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X163 a_32884_5882# a_32118_6363# a_32788_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X164 a_26317_625# a_26147_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X165 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X166 VSS a_369_1861# a_11573_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X167 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X168 a_27567_1923# a_27208_1758# a_27206_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X169 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X170 VDD a_52537_6584# a_52487_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X171 a_20653_625# a_20483_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X172 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X173 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 a_15381_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X175 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X176 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X177 a_36660_5882# a_35946_6337# a_36564_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X178 a_18559_6584# a_17684_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X179 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X180 a_44214_6938# a_44212_5882# a_44515_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X181 a_13487_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X182 VSS a_684_702# a_1609_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X183 a_9856_765# a_9630_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X184 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X185 a_32870_702# a_32506_765# a_32774_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X186 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X187 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X188 VSS C[19] a_22730_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X189 a_11744_765# a_11518_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X190 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X191 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 a_19668_5882# a_18902_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X193 a_47886_5882# a_47268_6337# a_47486_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X194 a_28504_619# C[47] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X195 a_13543_1923# a_13456_1825# a_13461_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X196 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X197 a_46397_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X198 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X199 a_4570_5882# a_3804_6363# a_4474_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X200 a_25320_1758# a_24728_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X201 a_55520_702# a_55156_765# a_55424_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X202 a_57424_6938# a_56708_6337# a_55438_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X203 VSS a_38438_702# a_39363_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X204 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X205 VDD a_54820_6337# a_54768_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X206 VSS a_15467_1861# a_19119_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X207 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X208 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X209 a_8346_5882# a_7632_6337# a_8250_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X210 a_44559_1923# a_44200_1758# a_44198_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X211 a_12124_6938# a_11356_6363# a_10138_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X212 a_17257_5637# a_17284_6378# a_17269_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X213 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X214 a_32373_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X215 VDD a_47604_765# a_47428_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X216 VSS C[8] a_43498_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X217 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X218 a_47970_1758# a_47378_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X219 a_32774_702# a_32506_765# a_32335_1923# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=0p ps=0u w=650000u l=150000u
X220 a_32774_702# a_32280_619# a_32335_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X221 VDD a_11013_6584# a_10963_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X222 VSS a_24223_6584# a_24173_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X223 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 a_47970_1758# a_47378_619# a_45984_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X225 VDD a_13296_6337# a_13244_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X226 VSS C[10] a_39722_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X227 a_36660_5882# a_35894_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X228 a_47984_6938# a_47982_5882# a_48285_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X229 VDD a_55424_702# a_56349_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X230 a_17257_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X231 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X232 a_55424_702# a_54930_619# a_54985_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X233 a_47984_6938# a_47268_6337# a_45998_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X234 VDD a_30571_1861# a_31343_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X235 a_17670_702# a_19064_619# a_19114_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X236 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X237 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X238 a_25236_5882# a_26506_6337# a_26697_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X239 a_57422_5882# a_56656_6363# a_57326_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X240 VDD a_7968_765# a_7792_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X241 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X242 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X243 a_18765_625# a_18595_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X244 VSS a_30571_1861# a_36111_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X245 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X246 VSS RESET sky130_fd_sc_hd__inv_4_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X247 VSS a_14783_6584# a_14733_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X248 VDD a_27110_702# a_28035_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X249 a_7237_6584# a_6362_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X250 a_34249_5637# a_34276_6378# a_34261_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X251 a_n315_6584# a_n225_6339# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X252 VDD a_58596_6337# a_58814_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X253 a_53646_5882# a_52880_6363# a_53550_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X254 a_32870_702# a_32872_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X255 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X256 VSS a_41215_6584# a_41165_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X257 VSS a_13900_702# a_14825_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X258 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X259 a_8346_5882# a_7580_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X260 VSS C[6] a_47268_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X261 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=2.808e+12p pd=2.944e+07u as=0p ps=0u w=650000u l=150000u
X262 a_57422_5882# a_56708_6337# a_57326_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X263 VSS a_53646_5882# a_53648_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X264 a_12026_5882# a_13244_6363# a_13487_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X265 a_38081_1923# a_37994_1825# a_37999_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X266 VDD a_369_1861# a_3029_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X267 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X268 a_34249_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X269 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X270 VSS a_9738_6378# a_9711_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X271 a_6805_1923# a_6446_1758# a_6444_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X272 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X273 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X274 a_34662_702# a_36056_619# a_36106_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X275 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X276 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 VDD a_17066_6337# a_17014_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X278 a_42228_5882# a_43498_6337# a_43689_5637# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=0p ps=0u w=650000u l=150000u
X279 a_24954_765# a_24728_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X280 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X281 VSS a_32170_6337# a_32118_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X282 a_24809_5637# a_24836_6378# a_24821_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X283 a_26842_765# a_26616_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X284 a_32870_702# a_32280_619# a_32774_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X285 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X286 VSS a_53150_6378# a_53123_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X287 VDD a_30886_702# a_31811_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X288 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X289 a_50217_1923# a_49858_1758# a_49856_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X290 a_23430_702# a_23432_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X291 VSS a_31775_6584# a_31725_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X292 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X293 a_47982_5882# a_47268_6337# a_47886_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X294 a_49872_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X295 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X296 a_55536_6938# a_55534_5882# a_55837_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X297 a_24809_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X298 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X299 a_53135_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X300 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X301 a_13914_5882# a_13296_6337# a_13514_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X302 VDD a_15467_1861# a_21089_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X303 a_12425_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X304 a_24865_1923# a_24778_1825# a_24783_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X305 a_47872_702# a_47378_619# a_47433_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X306 VDD a_369_1861# a_8693_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X307 VSS a_45669_1861# a_57408_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X308 VSS a_30571_1861# a_43663_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X309 VDD a_34058_6337# a_34006_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X310 a_327_1923# a_240_1825# a_245_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X311 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X312 VSS a_3461_6584# a_3411_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X313 a_41801_5637# a_41828_6378# a_41813_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X314 a_30392_619# C[48] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X315 VDD a_45669_1861# a_52105_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X316 a_40422_702# a_40424_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X317 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X318 VSS a_37834_6337# a_37782_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X319 a_32280_619# C[49] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X320 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X321 a_271_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X322 a_8332_702# a_7968_765# a_8236_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X323 a_15880_1758# a_15514_765# a_13900_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X324 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X325 a_59312_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X326 VSS a_40326_702# a_41251_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X327 a_36550_702# a_38170_765# a_37994_1825# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X328 VSS a_45669_1861# a_56873_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X329 VDD a_6080_765# a_5904_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X330 a_13998_1758# a_13406_619# a_12012_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X331 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X332 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X333 VDD a_22335_6584# a_22285_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X334 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X335 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X336 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X337 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X338 VDD C[4] a_51044_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X339 a_49858_1758# a_49266_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X340 a_36564_5882# a_37782_6363# a_38025_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X341 a_14012_6938# a_14010_5882# a_14313_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X342 a_5555_625# a_5385_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X343 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X344 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X345 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X346 a_56818_619# C[62] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X347 a_41857_1923# a_41770_1825# a_41775_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X348 a_51380_765# a_51154_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X349 VSS a_28998_702# a_29923_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X350 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 a_698_5882# a_1968_6337# a_2159_5637# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X352 a_17684_5882# a_17066_6337# a_17284_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X353 a_23430_702# a_23066_765# a_23334_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X354 a_16195_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X355 VSS a_9520_6337# a_9468_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X356 a_8236_702# a_7968_765# a_7797_1923# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X357 VDD a_21178_765# a_21002_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X358 a_8236_702# a_7742_619# a_7797_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X359 a_19064_619# C[42] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X360 a_27110_702# a_28730_765# a_28554_1825# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X361 VSS a_45669_1861# a_47433_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X362 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X363 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X364 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X365 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X366 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X367 a_43309_625# a_43139_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X368 a_32872_1758# a_32506_765# a_30886_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X369 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X370 a_45571_5637# a_45598_6378# a_45583_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X371 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X372 a_20653_625# a_20483_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X373 a_46080_702# a_45716_765# a_45984_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X374 a_7742_619# C[36] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X375 a_30447_1923# a_30442_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X376 a_14357_1923# a_13998_1758# a_13996_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X377 VSS a_52537_6584# a_52487_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X378 VSS C[24] a_13296_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X379 a_9630_619# C[37] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X380 a_47968_702# a_47378_619# a_47872_702# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X381 a_47968_702# a_47604_765# a_47872_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X382 a_18559_6584# a_17684_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X383 VDD a_45984_702# a_46909_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X384 VDD a_37834_6337# a_38052_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X385 a_17768_1758# a_17176_619# a_15782_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X386 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X387 a_23334_702# a_22840_619# a_22895_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X388 a_23334_702# a_23066_765# a_22895_1923# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X389 a_49403_1923# a_49316_1825# a_49321_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X390 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X391 VDD C[1] a_56708_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X392 VSS C[26] a_9520_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X393 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X394 a_n225_6339# a_28_6363# a_271_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X395 a_34676_5882# a_34058_6337# a_34276_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X396 a_17782_6938# a_17780_5882# a_18083_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X397 a_45984_702# a_47378_619# a_47428_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 a_33187_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X399 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X400 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X401 a_22840_619# C[44] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X402 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X403 a_27220_5882# a_26454_6363# a_27124_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X404 a_44214_6938# a_43498_6337# a_42228_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X405 VDD a_41610_6337# a_41558_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X406 a_38452_5882# a_37782_6363# a_38052_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X407 a_2133_1923# a_2128_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X408 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X409 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X410 a_14010_5882# a_13296_6337# a_13914_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X411 a_47872_702# a_47604_765# a_47433_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X412 VDD a_28394_6337# a_28612_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X413 a_23444_5882# a_22678_6363# a_23348_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X414 a_45490_619# C[56] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X415 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 a_53550_5882# a_54820_6337# a_55011_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X417 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X418 VSS a_11013_6584# a_10963_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X419 VSS a_794_5882# a_796_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X420 a_34760_1758# a_34168_619# a_32774_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X421 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X422 VSS C[22] a_17066_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X423 a_6362_5882# a_5744_6337# a_5962_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X424 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X425 a_8332_702# a_7742_619# a_8236_702# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X426 VSS a_55424_702# a_56349_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X427 a_27220_5882# a_26506_6337# a_27124_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X428 VDD a_6348_702# a_7273_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X429 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X430 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X431 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X432 a_57326_5882# a_58544_6363# a_58787_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X433 a_34774_6938# a_34772_5882# a_35075_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X434 VDD a_80_6337# a_298_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X435 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X436 a_34774_6938# a_34058_6337# a_32788_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X437 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X438 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X440 a_29012_5882# a_28342_6363# a_28612_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X441 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X442 VDD a_1573_6584# a_1523_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X443 a_44212_5882# a_43446_6363# a_44116_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X444 a_782_1758# a_190_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X445 a_57410_1758# a_57044_765# a_55424_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X446 VSS a_27110_702# a_28035_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X447 a_35757_625# a_35587_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X448 a_44116_5882# a_45380_6337# a_45571_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X449 a_15514_765# a_15288_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X450 a_2670_1758# a_2078_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X451 a_47872_702# a_49492_765# a_49316_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X452 a_7797_1923# a_7792_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X453 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X454 a_7237_6584# a_6362_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X455 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X456 a_40436_5882# a_39670_6363# a_40340_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X457 a_23430_702# a_22840_619# a_23334_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X458 a_17402_765# a_17176_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X459 a_53634_1758# a_53268_765# a_51648_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X460 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X461 VDD a_21446_702# a_22371_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X462 a_6446_1758# a_5854_619# a_4460_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X463 a_53268_765# a_53042_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X464 a_17780_5882# a_17066_6337# a_17684_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X465 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X466 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X467 a_47886_5882# a_49104_6363# a_49347_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X468 a_25334_6938# a_25332_5882# a_25635_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X469 a_58407_625# a_58237_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X470 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X471 VSS C[13] a_34058_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X472 a_59200_702# a_58596_6337# a_58814_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X473 VSS a_40436_5882# a_40438_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X474 a_46080_702# a_45490_619# a_45984_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X475 VSS a_15467_1861# a_27206_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X476 VSS a_369_1861# a_13461_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X477 a_27220_5882# a_26454_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X478 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X479 a_55438_5882# a_54820_6337# a_55038_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X480 VSS a_30886_702# a_31811_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X481 a_11599_5637# a_11626_6378# a_11611_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X482 a_30996_5882# a_30230_6363# a_30900_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X483 a_10220_702# a_10222_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X484 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X485 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X486 VSS a_28612_6378# a_28585_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X487 a_25679_1923# a_25320_1758# a_25318_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X488 VDD a_45669_1861# a_58843_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X489 a_34772_5882# a_34058_6337# a_34676_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X490 a_42312_1758# a_41720_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X491 a_59298_1758# a_58706_619# a_57312_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X492 a_42326_6938# a_42324_5882# a_42627_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X493 a_11599_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X494 VDD a_49156_6337# a_49374_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X495 a_12012_702# a_13406_619# a_13456_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X496 a_51760_6938# a_50992_6363# a_49774_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X497 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X498 a_17780_5882# a_17014_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X499 a_55522_1758# a_54930_619# a_53536_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X500 a_45998_5882# a_45380_6337# a_45598_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X501 a_11655_1923# a_11568_1825# a_11573_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X502 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X503 VDD a_13632_765# a_13456_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X504 VSS a_30571_1861# a_44198_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X505 a_13998_1758# a_13406_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X506 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X507 a_2682_5882# a_1916_6363# a_2586_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X508 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X509 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X510 a_47378_619# C[57] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X511 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X512 a_55536_6938# a_54820_6337# a_53550_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X513 VDD a_52932_6337# a_52880_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X514 VSS a_15467_1861# a_17231_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X515 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X516 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X517 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X518 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X519 VDD a_15467_1861# a_27567_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X520 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X521 a_6458_5882# a_5744_6337# a_6362_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X522 a_15369_5637# a_15396_6378# a_15381_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X523 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X524 a_30485_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X525 VSS a_22335_6584# a_22285_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X526 sky130_fd_sc_hd__inv_4_0/Y RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X527 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X528 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X529 a_19201_1923# a_19114_1825# a_19119_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X530 VDD C[17] a_26506_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X531 a_2304_765# a_2078_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X532 a_46096_6938# a_46094_5882# a_46397_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X533 VSS C[2] a_54820_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X534 a_15369_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X535 a_794_5882# a_80_6337# a_698_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X536 a_4192_765# a_3966_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X537 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X538 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X539 a_15782_702# a_17176_619# a_17226_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X540 a_36137_5637# a_36164_6378# a_36149_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X541 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X542 a_43309_625# a_43139_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X543 VSS a_30571_1861# a_34223_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X544 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X545 a_39925_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X546 a_2171_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X547 a_5349_6584# a_4474_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X548 a_32361_5637# a_32388_6378# a_32373_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X549 a_51758_5882# a_50992_6363# a_51662_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X550 VDD a_56708_6337# a_56926_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X551 a_59310_5882# a_58596_6337# a_59200_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X552 VSS a_45984_702# a_46909_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X553 a_30982_702# a_30984_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X554 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X555 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X556 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X557 a_6458_5882# a_5692_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X558 VSS C[7] a_45380_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X559 a_19290_765# a_19064_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X560 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X561 a_36193_1923# a_36106_1825# a_36111_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X562 VDD a_369_1861# a_1141_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X563 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X564 VSS a_45669_1861# a_49856_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X565 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X566 OUT a_60125_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X567 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X568 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X569 a_27124_5882# a_28342_6363# a_28585_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X570 a_49870_5882# a_49104_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X571 VSS a_7850_6378# a_7823_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X572 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X573 a_32774_702# a_34168_619# a_34218_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X574 a_4917_1923# a_4558_1758# a_4556_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X575 VDD a_15178_6337# a_15126_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X576 VSS a_369_1861# a_5909_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X577 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X578 VSS a_30282_6337# a_30230_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X579 a_22921_5637# a_22948_6378# a_22933_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X580 a_4047_5637# a_4074_6378# a_4059_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X581 a_4572_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X582 VSS a_51262_6378# a_51235_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X583 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X584 a_21542_702# a_21544_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X585 VSS a_18954_6337# a_18902_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X586 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X587 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X588 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X589 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X590 a_7835_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X591 a_29096_1758# a_28504_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X592 a_17670_702# a_19290_765# a_19114_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X593 a_13900_702# a_13406_619# a_13461_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X594 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X595 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X596 a_10234_5882# a_9468_6363# a_10138_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X597 a_23432_1758# a_23066_765# a_21446_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X598 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X599 a_40340_5882# a_41610_6337# a_41801_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X600 VSS a_369_1861# a_245_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X601 a_51247_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X602 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X603 a_4047_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X604 a_17684_5882# a_18902_6363# a_19145_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X605 a_12026_5882# a_11408_6337# a_11626_6378# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X606 VSS a_6348_702# a_7273_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X607 a_21007_1923# a_21002_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X608 a_38534_702# a_38170_765# a_38438_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X609 a_38534_702# a_37944_619# a_38438_702# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X610 VDD a_30571_1861# a_38081_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X611 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X612 a_4460_702# a_5854_619# a_5904_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=0p ps=0u w=1e+06u l=150000u
X613 a_22977_1923# a_22890_1825# a_22895_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X614 VDD a_369_1861# a_6805_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X615 VSS a_45669_1861# a_55520_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X616 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X617 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X618 VSS a_1573_6584# a_1523_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X619 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X620 a_35757_625# a_35587_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X621 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X622 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X623 VDD a_45669_1861# a_50217_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X624 a_44200_1758# a_43834_765# a_42214_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X625 a_25236_5882# a_24618_6337# a_24836_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X626 VSS a_35946_6337# a_35894_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X627 VDD a_44102_702# a_45027_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X628 a_57424_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X629 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X630 a_30900_5882# a_32170_6337# a_32361_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X631 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X632 VDD C[28] a_5744_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X633 VSS a_21446_702# a_22371_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X634 a_34662_702# a_36282_765# a_36106_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X635 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X636 VSS a_30571_1861# a_41775_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X637 VDD a_15467_1861# a_28641_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X638 VDD a_20447_6584# a_20397_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X639 VDD a_39327_6584# a_39277_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X640 a_38438_702# a_38170_765# a_37999_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X641 a_38438_702# a_37944_619# a_37999_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X642 a_58407_625# a_58237_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X643 a_53648_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X644 a_29096_1758# a_28504_619# a_27110_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X645 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X646 a_34676_5882# a_35894_6363# a_36137_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X647 VDD C[5] a_49156_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X648 a_12124_6938# a_12122_5882# a_12425_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X649 a_48761_6584# a_47886_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X650 VDD a_18954_6337# a_19172_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X651 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X652 a_52743_625# a_52573_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X653 VDD a_15467_1861# a_24865_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X654 a_37944_619# C[52] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X655 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X656 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X657 a_57312_702# a_58706_619# a_58756_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X658 a_25320_1758# a_24728_619# a_23334_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X659 VDD a_369_1861# a_327_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X660 a_15796_5882# a_15178_6337# a_15396_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X661 VDD a_45669_1861# a_59657_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X662 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X663 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X664 a_39832_619# C[53] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X665 VSS a_369_1861# a_13996_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X666 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X667 VSS a_7632_6337# a_7580_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X668 a_41946_765# a_41720_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X669 a_13996_702# a_13406_619# a_13900_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X670 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X671 a_13996_702# a_13632_765# a_13900_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X672 a_14010_5882# a_13244_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X673 a_43834_765# a_43608_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X674 a_6348_702# a_7968_765# a_7792_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X675 a_25334_6938# a_24618_6337# a_23348_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X676 VDD a_22730_6337# a_22678_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X677 a_24429_625# a_24259_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X678 a_30984_1758# a_30618_765# a_28998_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X679 VDD a_29887_6584# a_29837_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X680 a_19572_5882# a_18902_6363# a_19172_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X681 VSS a_51044_6337# a_50992_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X682 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X683 a_57410_1758# a_56818_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X684 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X685 VDD C[0] a_58596_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X686 a_12469_1923# a_12110_1758# a_12108_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X687 a_8348_6938# a_7580_6363# a_6362_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X688 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X689 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X690 VDD a_35946_6337# a_36164_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X691 a_15880_1758# a_15288_619# a_13900_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X692 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X693 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X694 a_47515_1923# a_47428_1825# a_47433_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X695 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X696 VDD a_28730_765# a_28554_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X697 a_13900_702# a_13632_765# a_13461_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X698 a_32788_5882# a_32170_6337# a_32388_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X699 a_15894_6938# a_15892_5882# a_16195_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X700 a_31299_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X701 a_44102_702# a_45490_619# a_45540_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X702 a_15894_6938# a_15178_6337# a_13914_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X703 VSS a_30996_5882# a_30998_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X704 a_2670_1758# a_2304_765# a_684_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X705 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X706 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X707 a_42326_6938# a_41610_6337# a_40340_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X708 VDD a_36550_702# a_37475_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X709 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X710 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X711 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X712 VSS a_56708_6337# a_56656_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X713 a_21556_5882# a_20790_6363# a_21460_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X714 VDD a_26506_6337# a_26724_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X715 a_29108_5882# a_28394_6337# a_29012_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X716 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X717 a_51662_5882# a_52932_6337# a_53123_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X718 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X719 a_30984_1758# a_30392_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X720 a_32872_1758# a_32280_619# a_30886_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X721 a_16239_1923# a_15880_1758# a_15878_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X722 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X723 VDD a_45669_1861# a_49403_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X724 VSS C[23] a_15178_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X725 a_4474_5882# a_3856_6337# a_4074_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X726 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X727 a_25332_5882# a_24618_6337# a_25236_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X728 a_55438_5882# a_56656_6363# a_56899_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X729 a_32886_6938# a_32884_5882# a_33187_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X730 a_32886_6938# a_32170_6337# a_30900_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X731 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X732 a_8250_5882# a_7580_6363# a_7850_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X733 a_42324_5882# a_41558_6363# a_42228_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X734 a_36056_619# C[51] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X735 a_55522_1758# a_55156_765# a_53536_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X736 a_16877_625# a_16707_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X737 VSS a_21060_6378# a_21033_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X738 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X739 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X740 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X741 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X742 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X743 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X744 a_5349_6584# a_4474_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X745 a_12108_702# a_11744_765# a_12012_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X746 a_12108_702# a_11518_619# a_12012_702# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X747 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X748 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X749 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X750 VDD a_43498_6337# a_43716_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X751 a_57044_765# a_56818_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X752 a_51746_1758# a_51380_765# a_49760_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X753 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X754 a_27999_6584# a_27124_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X755 a_4558_1758# a_3966_619# a_2572_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X756 a_15892_5882# a_15178_6337# a_15796_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X757 a_58932_765# a_58706_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X758 VDD a_12012_702# a_12937_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X759 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X760 a_45998_5882# a_47216_6363# a_47459_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X761 a_23446_6938# a_23444_5882# a_23747_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X762 VSS C[14] a_32170_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X763 a_21045_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X764 a_40326_702# a_40058_765# a_39887_1923# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X765 a_55011_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X766 OUT a_60125_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X767 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X768 a_57326_5882# a_56708_6337# a_56926_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X769 a_8334_1758# a_7742_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X770 a_8649_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X771 VSS a_15467_1861# a_25318_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X772 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X773 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X774 a_27110_702# a_26616_619# a_26671_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X775 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X776 VDD a_15467_1861# a_20015_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X777 VSS a_51758_5882# a_51760_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X778 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X779 a_28998_702# a_28504_619# a_28559_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X780 a_28998_702# a_28730_765# a_28559_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X781 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X782 a_46094_5882# a_45328_6363# a_45998_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X783 a_27222_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X784 VDD a_45669_1861# a_56955_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X785 a_11518_619# C[38] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X786 VSS C[29] a_3856_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X787 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 a_23432_1758# a_22840_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X789 a_57410_1758# a_56818_619# a_55424_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X790 a_13406_619# C[39] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X791 VDD a_47268_6337# a_47486_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X792 a_23446_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X793 VDD C[21] a_18954_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X794 VDD C[11] a_37834_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X795 a_10124_702# a_11518_619# a_11568_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X796 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X797 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X798 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X799 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X800 a_46082_1758# a_45490_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X801 a_58761_1923# a_58756_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X802 VSS a_30571_1861# a_42310_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X803 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X804 VDD a_30618_765# a_30442_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X805 VDD a_15467_1861# a_29455_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X806 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X807 a_53648_6938# a_52932_6337# a_51662_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X808 VSS a_44102_702# a_45027_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X809 VSS a_15467_1861# a_15343_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X810 a_32506_765# a_32280_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X811 a_44214_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X812 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X813 a_4570_5882# a_3856_6337# a_4474_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X814 a_40422_702# a_39832_619# a_40326_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X815 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 a_34394_765# a_34168_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X817 VDD a_53268_765# a_53092_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X818 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X819 VDD C[16] a_28394_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X820 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X821 VSS a_20447_6584# a_20397_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X822 VSS a_39327_6584# a_39277_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X823 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X824 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X825 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X826 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X827 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X828 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X829 a_52743_625# a_52573_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X830 a_55156_765# a_54930_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X831 a_35551_6584# a_34676_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X832 a_48761_6584# a_47886_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X833 a_3667_625# a_3497_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X834 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X835 a_27206_702# a_26842_765# a_27110_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X836 a_27206_702# a_26616_619# a_27110_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X837 a_17313_1923# a_17226_1825# a_17231_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X838 VDD C[18] a_24618_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X839 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X840 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X841 VSS C[3] a_52932_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X842 a_13900_702# a_15288_619# a_15338_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X843 VDD a_19290_765# a_19114_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X844 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X845 a_55424_702# a_55156_765# a_54985_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X846 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X847 a_24429_625# a_24259_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X848 a_12012_702# a_13632_765# a_13456_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X849 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X850 a_12124_6938# a_11408_6337# a_10138_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X851 a_48329_1923# a_47970_1758# a_47968_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X852 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X853 VSS a_29887_6584# a_29837_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X854 a_30473_5637# a_30500_6378# a_30485_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X855 a_54930_619# C[61] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X856 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X857 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X858 VSS a_26506_6337# a_26454_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X859 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X860 VSS a_369_1861# a_4556_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X861 a_47984_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X862 a_27110_702# a_26842_765# a_26671_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X863 a_21460_5882# a_22730_6337# a_22921_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X864 a_4570_5882# a_3804_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X865 a_30982_702# a_30618_765# a_30886_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X866 VDD a_15467_1861# a_19201_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X867 a_9856_765# a_9630_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X868 a_34305_1923# a_34218_1825# a_34223_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X869 VDD C[9] a_41610_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X870 a_26616_619# C[46] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X871 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X872 a_25236_5882# a_26454_6363# a_26697_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X873 VSS a_5962_6378# a_5935_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X874 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X875 a_30886_702# a_32280_619# a_32330_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X876 a_3029_1923# a_2670_1758# a_2668_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X877 VSS a_369_1861# a_4021_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X878 a_9723_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X879 a_28504_619# C[47] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X880 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X881 a_39913_5637# a_39940_6378# a_39925_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X882 VSS a_36550_702# a_37475_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X883 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X884 a_12122_5882# a_11356_6363# a_12026_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X885 a_2159_5637# a_2186_6378# a_2171_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X886 a_25320_1758# a_24954_765# a_23334_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X887 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X888 a_2684_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X889 a_38534_702# a_38536_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X890 a_780_702# a_782_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X891 a_5947_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X892 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X893 VDD a_45716_765# a_45540_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X894 a_15782_702# a_17402_765# a_17226_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X895 a_30886_702# a_30618_765# a_30447_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X896 VDD a_13296_6337# a_13514_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X897 a_30886_702# a_30392_619# a_30447_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X898 a_21544_1758# a_21178_765# a_19558_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X899 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 a_38452_5882# a_39722_6337# a_39913_5637# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X901 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X902 a_2159_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X903 a_47604_765# a_47378_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X904 a_15796_5882# a_17014_6363# a_17257_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X905 a_19654_702# a_19064_619# a_19558_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X906 VDD a_30571_1861# a_36193_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X907 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X908 a_19654_702# a_19290_765# a_19558_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X909 a_55520_702# a_54930_619# a_55424_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X910 a_2572_702# a_3966_619# a_4016_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X911 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X912 a_12122_5882# a_11408_6337# a_12026_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X913 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X914 a_27124_5882# a_26506_6337# a_26724_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X915 VDD a_53536_702# a_54461_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X916 a_39969_1923# a_39882_1825# a_39887_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X917 VDD a_369_1861# a_4917_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X918 a_42228_5882# a_43446_6363# a_43689_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X919 a_56313_6584# a_55438_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X920 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X921 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X922 a_16877_625# a_16707_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X923 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X924 a_23348_5882# a_22730_6337# a_22948_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X925 a_42312_1758# a_41946_765# a_40326_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X926 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X927 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X928 a_57422_5882# a_56656_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X929 a_55011_5637# a_55038_6378# a_55023_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X930 VDD a_25222_702# a_26147_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X931 a_55536_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X932 a_29012_5882# a_30282_6337# a_30473_5637# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X933 a_58799_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X934 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X935 VDD a_15467_1861# a_26753_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X936 a_27999_6584# a_27124_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X937 VSS a_12012_702# a_12937_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X938 a_19558_702# a_19290_765# a_19119_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X939 VSS a_58814_6378# a_58787_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X940 a_13914_5882# a_13244_6363# a_13514_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X941 a_19558_702# a_19064_619# a_19119_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X942 a_55881_1923# a_55522_1758# a_55520_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X943 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X944 sky130_fd_sc_hd__inv_4_0/Y RESET VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X945 a_27208_1758# a_26616_619# a_25222_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X946 a_32788_5882# a_34006_6363# a_34249_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X947 a_10236_6938# a_10234_5882# a_10537_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X948 a_46873_6584# a_45998_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X949 a_53042_619# C[60] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X950 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X951 VDD a_17066_6337# a_17284_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X952 a_41421_625# a_41251_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X953 a_41801_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X954 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X955 a_44116_5882# a_43498_6337# a_43716_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X956 a_55424_702# a_56818_619# a_56868_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X957 a_38550_6938# a_37782_6363# a_36564_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X958 a_23432_1758# a_22840_619# a_21446_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X959 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X960 a_55067_1923# a_54980_1825# a_54985_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X961 a_28559_1923# a_28554_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X962 VSS a_369_1861# a_12108_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X963 VSS a_5744_6337# a_5692_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X964 a_24954_765# a_24728_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X965 a_30982_702# a_30392_619# a_30886_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X966 a_4460_702# a_6080_765# a_5904_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X967 a_51648_702# a_53042_619# a_53092_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X968 a_23446_6938# a_22730_6337# a_21460_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X969 VDD a_20842_6337# a_20790_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X970 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X971 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X972 VDD a_39722_6337# a_39670_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X973 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X974 VDD a_9125_6584# a_9075_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X975 a_14012_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X976 a_46082_1758# a_45716_765# a_44102_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X977 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X978 a_59296_702# a_59298_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X979 VDD a_45669_1861# a_57769_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X980 VDD a_30571_1861# a_43745_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X981 a_4474_5882# a_5692_6363# a_5935_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X982 a_23066_765# a_22840_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X983 a_44200_1758# a_43608_619# a_42214_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X984 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X985 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X986 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X987 VDD a_34058_6337# a_34276_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X988 a_45627_1923# a_45540_1825# a_45545_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X989 a_n225_6339# a_416_765# a_240_1825# VSS sky130_fd_pr__nfet_01v8 ad=4.29e+11p pd=3.92e+06u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X990 VSS a_80_6337# a_28_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X991 a_45984_702# a_45716_765# a_45545_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X992 a_45984_702# a_45490_619# a_45545_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X993 a_45571_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X994 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X995 a_796_6938# a_28_6363# a_n225_6339# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X996 VSS a_58596_6337# a_58544_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X997 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X998 a_40438_6938# a_39722_6337# a_38452_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X999 a_30392_619# C[48] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1000 VDD a_17670_702# a_18595_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1001 a_6444_702# a_5854_619# a_6348_702# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1002 a_6444_702# a_6080_765# a_6348_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1003 a_57312_702# a_58932_765# a_58756_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1004 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1005 a_18127_1923# a_17768_1758# a_17766_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1006 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1007 VDD a_24618_6337# a_24836_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1008 a_38548_5882# a_37782_6363# a_38452_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1009 VDD a_5744_6337# a_5962_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1010 a_49774_5882# a_51044_6337# a_51235_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1011 a_17782_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1012 a_3667_625# a_3497_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1013 VDD a_45669_1861# a_47515_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1014 a_35551_6584# a_34676_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1015 a_2586_5882# a_1968_6337# a_2186_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1016 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1017 a_1097_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1018 VSS a_38548_5882# a_38550_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1019 VDD C[25] a_11408_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1020 a_53550_5882# a_54768_6363# a_55011_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1021 a_49492_765# a_49266_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1022 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1023 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1024 VSS a_30571_1861# a_36646_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1025 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1026 a_21542_702# a_21178_765# a_21446_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1027 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1028 a_30998_6938# a_30282_6337# a_29012_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1029 a_51380_765# a_51154_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1030 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1031 a_6362_5882# a_5692_6363# a_5962_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1032 a_6348_702# a_6080_765# a_5909_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1033 a_6348_702# a_5854_619# a_5909_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1034 VDD a_45380_6337# a_45328_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1035 a_17176_619# C[41] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1036 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1037 a_38851_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1038 a_19064_619# C[42] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1039 VSS a_38052_6378# a_38025_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1040 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1041 a_38536_1758# a_37944_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1042 a_35119_1923# a_34760_1758# a_34758_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1043 a_5854_619# C[35] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1044 VDD a_41610_6337# a_41828_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1045 a_44212_5882# a_43498_6337# a_44116_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1046 a_2670_1758# a_2078_619# a_684_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1047 a_7742_619# C[36] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1048 a_12901_6584# a_12026_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1049 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1050 a_34774_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1051 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1052 a_8250_5882# a_9520_6337# a_9711_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1053 a_44116_5882# a_45328_6363# a_45571_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 a_698_5882# a_28_6363# a_298_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1055 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1056 a_2684_6938# a_2682_5882# a_2985_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1057 VSS C[15] a_30282_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1058 a_38037_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1059 a_21446_702# a_21178_765# a_21007_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1060 a_21446_702# a_20952_619# a_21007_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1061 a_2684_6938# a_1968_6337# a_698_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1062 a_51209_1923# a_51204_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1063 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1064 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1065 a_49872_6938# a_49104_6363# a_47886_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1066 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1067 VSS a_6458_5882# a_6460_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1068 a_26111_6584# a_25236_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1069 VSS a_15467_1861# a_23430_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1070 a_20952_619# C[43] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1071 a_21558_6938# a_21556_5882# a_21859_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1072 a_22840_619# C[44] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1073 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1074 VSS a_49870_5882# a_49872_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1075 VDD a_30571_1861# a_37007_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1076 a_12110_1758# a_11744_765# a_10124_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1077 a_25334_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1078 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1079 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1080 a_28597_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1081 VSS C[30] a_1968_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1082 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1083 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1084 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1085 a_45490_619# C[56] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1086 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1087 a_59200_702# a_58544_6363# a_58814_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1088 VDD a_45380_6337# a_45598_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1089 VDD a_50649_6584# a_50599_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1090 a_21558_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1091 VSS a_53536_702# a_54461_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1092 a_16671_6584# a_15796_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1093 VDD C[12] a_35946_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1094 VDD a_4460_702# a_5385_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1095 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1096 a_25222_702# a_26616_619# a_26666_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=6.6e+11p pd=5.32e+06u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1097 a_56873_1923# a_56868_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1098 VSS a_30571_1861# a_40422_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1099 a_56313_6584# a_55438_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1100 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1101 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1102 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1103 VSS a_298_6378# a_271_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1104 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1105 VSS a_59310_5882# a_59312_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1106 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1107 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1108 a_51760_6938# a_51044_6337# a_49774_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1109 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1110 VSS a_25222_702# a_26147_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1111 a_10138_5882# a_9520_6337# a_9738_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1112 a_33869_625# a_33699_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1113 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1114 a_21446_702# a_22840_619# a_22890_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1115 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1116 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1117 a_44212_5882# a_43446_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1118 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1119 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1120 a_42326_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1121 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1122 a_2682_5882# a_1968_6337# a_2586_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1123 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1124 a_21542_702# a_20952_619# a_21446_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1125 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1126 a_49774_5882# a_49104_6363# a_49374_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1127 a_15514_765# a_15288_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1128 VDD a_19558_702# a_20483_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1129 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1130 a_29094_702# a_29096_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1131 VDD a_369_1861# a_13543_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1132 VDD a_36282_765# a_36106_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1133 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1134 a_42671_1923# a_42312_1758# a_42310_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1135 a_56519_625# a_56349_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1136 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1137 VSS C[27] a_7632_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1138 a_41421_625# a_41251_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1139 a_33663_6584# a_32788_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1140 a_46873_6584# a_45998_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1141 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1142 VDD C[19] a_22730_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1143 a_38170_765# a_37944_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1144 a_15425_1923# a_15338_1825# a_15343_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1145 VSS a_45669_1861# a_47968_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1146 a_42214_702# a_43608_619# a_43658_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1147 a_10222_1758# a_9630_619# a_8236_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1148 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1149 a_34772_5882# a_34006_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1150 a_44102_702# a_43608_619# a_43663_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1151 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1152 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1153 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1154 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1155 VSS a_28394_6337# a_28342_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1156 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1157 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1158 a_10236_6938# a_9520_6337# a_8250_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 a_19654_702# a_19656_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1160 a_9331_625# a_9161_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1161 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1162 VSS a_9125_6584# a_9075_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1163 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1164 VSS a_24618_6337# a_24566_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1165 VDD C[8] a_43498_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1166 VDD a_30571_1861# a_44559_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1167 a_40424_1758# a_39832_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1168 a_46096_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1169 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1170 a_19572_5882# a_20842_6337# a_21033_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1171 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1172 a_49359_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1173 VDD a_15467_1861# a_17313_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1174 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1175 VSS a_49374_6378# a_49347_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1176 VDD C[10] a_39722_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1177 a_46441_1923# a_46082_1758# a_46080_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1178 a_32417_1923# a_32330_1825# a_32335_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1179 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1180 a_23348_5882# a_24566_6363# a_24809_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 a_55534_5882# a_54820_6337# a_55438_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1182 VDD a_11744_765# a_11568_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1183 a_28998_702# a_30392_619# a_30442_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1184 VSS a_369_1861# a_2133_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1185 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1186 a_32361_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1187 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1188 VSS a_17670_702# a_18595_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1189 a_13632_765# a_13406_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1190 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1191 a_36646_702# a_36648_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1192 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1193 VDD a_11408_6337# a_11626_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1194 a_38536_1758# a_38170_765# a_36550_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.6e+11p ps=5.32e+06u w=1e+06u l=150000u
X1195 a_48967_625# a_48797_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1196 a_4103_1923# a_4016_1825# a_4021_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1197 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1198 a_58201_6584# a_57326_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1199 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1200 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1201 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1202 a_13914_5882# a_15126_6363# a_15369_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1203 VDD C[6] a_47268_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1204 VDD a_30571_1861# a_34305_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1205 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1206 a_44198_702# a_43834_765# a_44102_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1207 a_44198_702# a_43608_619# a_44102_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1208 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1209 a_53648_6938# a_53646_5882# a_53949_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1210 VDD a_42214_702# a_43139_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1211 sky130_fd_sc_hd__inv_4_0/Y RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1212 a_22921_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1213 a_416_765# a_190_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1214 a_684_702# a_2078_619# a_2128_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1215 a_40340_5882# a_41558_6363# a_41801_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1216 a_19670_6938# a_18902_6363# a_17684_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1217 a_54425_6584# a_53550_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1218 a_9711_5637# a_9738_6378# a_9723_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1219 a_2304_765# a_2078_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1220 a_36550_702# a_36056_619# a_36111_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1221 a_8332_702# a_8334_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1222 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1223 VDD a_32170_6337# a_32118_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1224 a_40424_1758# a_40058_765# a_38438_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1225 a_55534_5882# a_54768_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1226 a_53123_5637# a_53150_6378# a_53135_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1227 VSS a_19668_5882# a_19670_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1228 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1229 a_51744_702# a_51746_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1230 VSS a_49156_6337# a_49104_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1231 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1232 a_59200_702# a_58706_619# a_58761_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1233 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1234 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1235 VSS a_56926_6378# a_56899_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1236 a_12901_6584# a_12026_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1237 a_44102_702# a_43834_765# a_43663_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1238 a_53993_1923# a_53634_1758# a_53632_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1239 VDD a_369_1861# a_5991_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1240 VSS a_45669_1861# a_54985_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1241 a_30900_5882# a_32118_6363# a_32361_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1242 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1243 VDD a_15178_6337# a_15396_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1244 a_9767_1923# a_9680_1825# a_9685_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1245 a_42228_5882# a_41610_6337# a_41828_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1246 a_43608_619# C[55] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1247 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1248 a_53536_702# a_54930_619# a_54980_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1249 a_36662_6938# a_35894_6363# a_34676_5882# VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1250 a_55522_1758# a_54930_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1251 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 a_53179_1923# a_53092_1825# a_53097_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1253 a_26671_1923# a_26666_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1254 VSS a_369_1861# a_10220_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1255 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1256 a_26111_6584# a_25236_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1257 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1258 VSS a_3856_6337# a_3804_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1259 VSS a_29108_5882# a_29110_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1260 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1261 a_21558_6938# a_20842_6337# a_19572_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1262 a_2572_702# a_4192_765# a_4016_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1263 VDD a_37834_6337# a_37782_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1264 VDD a_26842_765# a_26666_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1265 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1266 VSS a_45669_1861# a_45545_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1267 VDD a_7237_6584# a_7187_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1268 a_12124_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1269 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1270 a_12012_702# a_11518_619# a_11573_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 a_57408_702# a_57410_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1272 VDD a_45669_1861# a_55881_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1273 VDD a_30571_1861# a_41857_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1274 a_2586_5882# a_3804_6363# a_4047_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 a_19668_5882# a_18902_6363# a_19572_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1276 a_28730_765# a_28504_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1277 a_42312_1758# a_41720_619# a_40326_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1278 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1279 VSS a_50649_6584# a_50599_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1280 VSS a_4460_702# a_5385_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1281 VDD a_32170_6337# a_32388_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1282 a_36646_702# a_36056_619# a_36550_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1283 a_36646_702# a_36282_765# a_36550_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1284 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1285 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 a_16671_6584# a_15796_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1287 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1288 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1289 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1290 a_47079_625# a_46909_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1291 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1292 VDD a_45669_1861# a_55067_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1293 VSS a_15467_1861# a_17766_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1294 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1295 VSS C[20] a_20842_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1296 a_43663_1923# a_43658_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1297 VDD a_369_1861# a_14357_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1298 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1299 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1300 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1301 VDD a_9520_6337# a_9468_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1302 a_33869_625# a_33699_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1303 a_59296_702# a_58706_619# a_59200_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1304 a_59296_702# a_58932_765# a_59200_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1305 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1306 a_19971_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1307 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1308 VSS a_19172_6378# a_19145_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1309 VSS a_19558_702# a_20483_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1310 a_36564_5882# a_35894_6363# a_36164_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1311 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1312 a_36550_702# a_36282_765# a_36111_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1313 a_49858_1758# a_49492_765# a_47872_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1314 VDD a_3856_6337# a_4074_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1315 a_56519_625# a_56349_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1316 VDD C[24] a_13296_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1317 a_15894_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1318 VDD a_45669_1861# a_45627_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1319 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1320 a_19157_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1321 a_33663_6584# a_32788_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1322 a_50855_625# a_50685_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1323 a_55424_702# a_57044_765# a_56868_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1324 a_46082_1758# a_45490_619# a_44102_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1325 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1326 VDD C[26] a_9520_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1327 a_51662_5882# a_52880_6363# a_53123_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1328 a_10220_702# a_9856_765# a_10124_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1329 VSS a_30571_1861# a_34758_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1330 a_59200_702# a_58932_765# a_58761_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1331 a_37944_619# C[52] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1332 a_40058_765# a_39832_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1333 a_46096_6938# a_45380_6337# a_44116_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1334 a_41946_765# a_41720_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1335 a_9331_625# a_9161_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1336 a_58706_619# C[63] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1337 a_36963_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1338 VDD a_15467_1861# a_18127_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1339 a_8346_5882# a_7580_6363# a_8250_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1340 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1341 a_19656_1758# a_19064_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1342 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1343 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1344 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1345 VSS a_11408_6337# a_11356_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1346 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1347 a_45984_702# a_47604_765# a_47428_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1348 a_5909_1923# a_5904_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1349 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1350 a_32886_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1351 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1352 VDD a_10124_702# a_11049_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1353 VSS a_8346_5882# a_8348_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1354 a_10124_702# a_9630_619# a_9685_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1355 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1356 a_796_6938# a_794_5882# a_1097_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1357 a_36149_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1358 VDD C[22] a_17066_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1359 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1360 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1361 a_33231_1923# a_32872_1758# a_32870_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1362 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1363 a_47984_6938# a_47216_6363# a_45998_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1364 a_12012_702# a_11744_765# a_11573_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1365 VDD a_52932_6337# a_53150_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1366 a_10138_5882# a_11356_6363# a_11599_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1367 VSS a_4570_5882# a_4572_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1368 a_42324_5882# a_41610_6337# a_42228_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1369 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1370 a_24223_6584# a_23348_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1371 VSS a_15467_1861# a_21542_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1372 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1373 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1374 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1375 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1376 VDD a_34662_702# a_35587_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1377 a_10222_1758# a_9856_765# a_8236_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1378 a_25332_5882# a_24566_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1379 a_53550_5882# a_52932_6337# a_53150_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1380 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1381 a_52061_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1382 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1383 a_26709_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1384 a_48967_625# a_48797_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1385 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1386 VSS C[31] a_80_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1387 VSS a_26724_6378# a_26697_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1388 a_23791_1923# a_23432_1758# a_23430_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1389 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1390 a_58201_6584# a_57326_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1391 VDD a_57312_702# a_58237_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1392 a_57326_5882# a_56656_6363# a_56926_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1393 a_38550_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1394 VSS a_42214_702# a_43139_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1395 a_32884_5882# a_32170_6337# a_32788_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1396 a_14783_6584# a_13914_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1397 VDD C[13] a_34058_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1398 a_40438_6938# a_40436_5882# a_40739_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.1e+11p ps=2.42e+06u w=1e+06u l=150000u
X1399 VDD a_n315_6584# a_n365_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1400 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1401 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1402 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1403 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1404 a_23334_702# a_24728_619# a_24778_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1405 a_41215_6584# a_40340_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1406 a_54425_6584# a_53550_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1407 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1408 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1409 VSS a_57422_5882# a_57424_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1410 a_53634_1758# a_53042_619# a_51648_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1411 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1412 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1413 a_34168_619# C[50] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1414 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1415 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1416 a_36056_619# C[51] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1417 a_19558_702# a_20952_619# a_21002_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1418 a_42324_5882# a_41558_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1419 a_40438_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1420 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1421 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1422 a_28585_5637# a_28612_6378# a_28597_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1423 a_47886_5882# a_47216_6363# a_47486_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1424 a_57044_765# a_56818_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1425 a_27206_702# a_27208_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1426 VDD a_15467_1861# a_25679_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1427 VDD a_369_1861# a_11655_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1428 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1429 VSS a_43716_6378# a_43689_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1430 VDD a_17402_765# a_17226_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1431 a_40783_1923# a_40424_1758# a_40422_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1432 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1433 a_17768_1758# a_17176_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1434 a_12110_1758# a_11518_619# a_10124_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1435 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1436 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1437 a_31775_6584# a_30900_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1438 a_39533_625# a_39363_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1439 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1440 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1441 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1442 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1443 a_6446_1758# a_5854_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1444 VSS a_45669_1861# a_46080_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1445 a_40326_702# a_41720_619# a_41770_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1446 a_13461_1923# a_13456_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1447 a_25222_702# a_24728_619# a_24783_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1448 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1449 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1450 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1451 a_25222_702# a_26842_765# a_26666_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1452 VSS a_7237_6584# a_7187_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1453 VSS a_30571_1861# a_32335_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1454 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1455 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1456 a_46094_5882# a_45328_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1457 a_44198_702# a_44200_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1458 VDD a_30571_1861# a_42671_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1459 a_21544_1758# a_20952_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1460 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1461 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 a_3461_6584# a_2586_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1463 a_19656_1758# a_19290_765# a_17670_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1464 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1465 a_11518_619# C[38] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1466 a_36564_5882# a_37834_6337# a_38025_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1467 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1468 a_14012_6938# a_13244_6363# a_12026_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1469 VDD a_15467_1861# a_15425_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1470 VSS a_47486_6378# a_47459_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1471 a_47079_625# a_46909_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1472 a_30529_1923# a_30442_1825# a_30447_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1473 VDD a_12901_6584# a_12851_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1474 a_53646_5882# a_52932_6337# a_53550_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1475 a_21460_5882# a_22678_6363# a_22921_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1476 VDD C[2] a_54820_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1477 a_30473_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1478 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1479 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1480 a_14995_625# a_14825_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1481 VSS a_43498_6337# a_43446_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1482 a_30618_765# a_30392_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1483 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1484 a_53632_702# a_53268_765# a_53536_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1485 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1486 a_27124_5882# a_28394_6337# a_28585_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1487 a_32506_765# a_32280_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1488 VDD a_51380_765# a_51204_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1489 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1490 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1491 a_49266_619# C[58] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1492 a_36648_1758# a_36282_765# a_34662_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1493 a_2215_1923# a_2128_1825# a_2133_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1494 a_50855_625# a_50685_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1495 VDD C[7] a_45380_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1496 VDD a_30571_1861# a_32417_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1497 a_1779_625# a_1609_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1498 a_25318_702# a_24954_765# a_25222_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1499 a_39913_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1500 a_55156_765# a_54930_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1501 VDD a_59200_702# a_60125_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1502 a_37999_1923# a_37994_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1503 a_17782_6938# a_17014_6363# a_15796_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1504 a_38452_5882# a_39670_6363# a_39913_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1505 VDD a_22730_6337# a_22948_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1506 a_52537_6584# a_51662_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1507 a_7823_5637# a_7850_6378# a_7835_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1508 VDD sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1509 a_17670_702# a_17176_619# a_17231_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1510 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1511 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1512 a_53536_702# a_53268_765# a_53097_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1513 VDD a_4192_765# a_4016_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1514 a_6444_702# a_6446_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1515 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1516 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1517 a_53536_702# a_53042_619# a_53097_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1519 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1520 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1521 VDD a_30282_6337# a_30230_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1522 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1523 a_53646_5882# a_52880_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1524 a_51235_5637# a_51262_6378# a_51247_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1525 VDD a_18954_6337# a_18902_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1526 VSS a_369_1861# a_9685_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1527 VSS a_36660_5882# a_36662_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1528 a_6080_765# a_5854_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1529 a_49856_702# a_49858_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1530 a_8334_1758# a_7968_765# a_6348_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1531 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1532 VSS a_47268_6337# a_47216_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1533 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1534 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1535 VSS a_10124_702# a_11049_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1536 a_54930_619# C[61] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1537 VDD a_369_1861# a_4103_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1538 a_7968_765# a_7742_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1539 VSS a_45669_1861# a_53097_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1540 a_32774_702# a_34394_765# a_34218_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1541 a_29012_5882# a_30230_6363# a_30473_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1542 a_27124_5882# a_26454_6363# a_26724_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1543 a_7879_1923# a_7792_1825# a_7797_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1544 VDD a_37439_6584# a_37389_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1545 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1546 a_24728_619# C[45] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1547 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1548 a_34774_6938# a_34006_6363# a_32788_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1549 a_26616_619# C[46] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1550 a_24783_1923# a_24778_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=3.77e+11p pd=3.76e+06u as=0p ps=0u w=650000u l=150000u
X1551 a_11013_6584# a_10138_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1552 a_24223_6584# a_23348_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1553 VSS a_1968_6337# a_1916_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1554 VSS a_27220_5882# a_27222_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1555 a_245_1923# a_240_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1556 VSS a_34662_702# a_35587_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1557 a_38550_6938# a_37834_6337# a_36564_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1558 a_5690_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1559 VDD a_35946_6337# a_35894_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1560 a_51235_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1561 a_12122_5882# a_11356_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1562 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1563 a_40340_5882# a_39722_6337# a_39940_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1564 a_10236_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1565 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1566 a_13107_625# a_12937_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1567 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1568 a_698_5882# a_1916_6363# a_2159_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 a_17684_5882# a_17014_6363# a_17284_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1570 a_13499_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1571 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1572 VSS a_57312_702# a_58237_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1573 a_47886_5882# a_49156_6337# a_49347_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1574 VSS a_13514_6378# a_13487_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1575 a_10581_1923# a_10222_1758# a_10220_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1576 VDD a_369_1861# a_9767_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1577 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1578 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1579 a_45716_765# a_45490_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1580 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1581 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1582 VDD a_30282_6337# a_30500_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1583 a_44116_5882# a_43446_6363# a_43716_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1584 a_17766_702# a_17176_619# a_17670_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1585 a_6460_6938# a_5692_6363# a_4474_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1586 a_17766_702# a_17402_765# a_17670_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1587 a_53632_702# a_53042_619# a_53536_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1588 a_14783_6584# a_13914_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1589 a_47604_765# a_47378_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1590 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1591 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1592 VDD a_51648_702# a_52573_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1593 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1594 VSS a_n315_6584# a_n365_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1595 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1596 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1597 VSS a_15467_1861# a_15878_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1598 a_41775_1923# a_41770_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1599 a_41215_6584# a_40340_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1600 VSS a_44212_5882# a_44214_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1601 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1602 VDD a_7632_6337# a_7580_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1603 a_40424_1758# a_39832_619# a_38438_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1604 a_30900_5882# a_30282_6337# a_30500_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1605 a_190_619# C[32] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1606 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1607 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1608 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1609 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1610 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1611 VDD a_51044_6337# a_50992_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1612 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1613 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1614 a_34676_5882# a_34006_6363# a_34276_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1615 VDD a_39722_6337# a_39940_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1616 a_17670_702# a_17402_765# a_17231_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1617 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1618 VDD a_1968_6337# a_2186_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1619 a_15892_5882# a_15126_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1620 a_4460_702# a_3966_619# a_4021_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1621 a_13996_702# a_13998_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1622 VDD a_369_1861# a_12469_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1623 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1624 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1625 VSS a_54820_6337# a_54768_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1626 a_39533_625# a_39363_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1627 sky130_fd_sc_hd__inv_4_0/Y RESET VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1628 a_51154_619# C[59] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1629 a_17269_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1630 a_31775_6584# a_30900_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1631 a_59312_6938# a_58544_6363# a_57326_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1632 a_53536_702# a_55156_765# a_54980_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1633 VSS a_17284_6378# a_17257_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1634 a_53042_619# C[60] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1635 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1636 a_30984_1758# a_30392_619# a_28998_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1637 a_49321_1923# a_49316_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1638 VSS a_30571_1861# a_32870_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1639 VDD a_58201_6584# a_58151_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1640 a_23444_5882# a_22730_6337# a_23348_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1641 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1642 a_55536_6938# a_54768_6363# a_53550_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1643 a_30998_6938# a_30996_5882# a_31299_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1644 VSS a_13296_6337# a_13244_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1645 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1646 VDD a_43834_765# a_43658_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1647 a_6458_5882# a_5692_6363# a_6362_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1648 VSS a_47982_5882# a_47984_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1649 a_44200_1758# a_43608_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1650 VDD a_56708_6337# a_56656_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1651 a_21178_765# a_20952_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1652 a_44102_702# a_45716_765# a_45540_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1653 a_3461_6584# a_2586_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1654 VDD a_54820_6337# a_55038_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1655 a_30998_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1656 VDD a_7632_6337# a_7850_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1657 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1658 a_23066_765# a_22840_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1659 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1660 VDD a_48761_6584# a_48711_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1661 a_19670_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1662 VDD C[23] a_15178_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1663 VSS a_34276_6378# a_34249_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1664 a_28205_625# a_28035_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1665 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1666 a_31343_1923# a_30984_1758# a_30982_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1667 VSS a_12901_6584# a_12851_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1668 a_794_5882# a_28_6363# a_698_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1669 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1670 a_40436_5882# a_39722_6337# a_40340_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1671 a_8250_5882# a_9468_6363# a_9711_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1672 a_22335_6584# a_21460_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1673 a_14995_625# a_14825_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1674 VSS a_30571_1861# a_38534_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1675 a_6761_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1676 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1677 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1678 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1679 a_49872_6938# a_49156_6337# a_47886_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1680 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1681 VDD a_15782_702# a_16707_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1682 a_4556_702# a_3966_619# a_4460_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1683 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1684 a_4556_702# a_4192_765# a_4460_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1685 a_23444_5882# a_22678_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1686 a_51662_5882# a_51044_6337# a_51262_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1687 a_21033_5637# a_21060_6378# a_21045_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1688 a_50173_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1689 VSS a_17066_6337# a_17014_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1690 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1691 VSS a_24836_6378# a_24809_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1692 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1693 a_21903_1923# a_21544_1758# a_21542_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1694 a_1779_625# a_1609_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1695 VSS a_15467_1861# a_22895_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1696 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1697 a_43103_6584# a_42228_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1698 a_55438_5882# a_54768_6363# a_55038_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1699 a_30996_5882# a_30282_6337# a_30900_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1700 a_31981_625# a_31811_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1701 VDD C[14] a_32170_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1702 VSS a_59200_702# a_60125_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1703 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1704 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1705 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1706 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1707 a_52537_6584# a_51662_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1708 a_49492_765# a_49266_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1709 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1710 a_4460_702# a_4192_765# a_4021_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1711 a_51746_1758# a_51154_619# a_49760_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=4.29e+11p ps=3.92e+06u w=650000u l=150000u
X1712 a_21089_1923# a_21002_1825# a_21007_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1713 VSS a_55534_5882# a_55536_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1714 a_15288_619# C[40] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1715 VSS a_45669_1861# a_53632_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1716 a_283_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1717 a_59613_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1718 a_40436_5882# a_39670_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1719 a_17176_619# C[41] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1720 a_51760_6938# a_51758_5882# a_52061_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1721 a_36648_1758# a_36056_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1722 VDD RESET sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1723 a_21033_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1724 a_3966_619# C[34] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1725 a_13998_1758# a_13632_765# a_12012_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1726 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1727 VSS a_34058_6337# a_34006_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1728 a_45998_5882# a_45328_6363# a_45598_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1729 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1730 a_5854_619# C[35] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1731 a_55837_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1732 a_8348_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1733 a_25318_702# a_25320_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1734 VSS a_41828_6378# a_41801_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1735 VDD a_15467_1861# a_23791_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1736 VDD C[29] a_3856_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1737 VSS a_30571_1861# a_39887_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1738 a_17684_5882# a_18954_6337# a_19145_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1739 a_49870_5882# a_49104_6363# a_49774_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1740 VDD a_58932_765# a_58756_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1741 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1742 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1743 a_59298_1758# a_58706_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1744 VSS a_37439_6584# a_37389_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1745 a_51760_6938# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1746 a_38438_702# a_39832_619# a_39882_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1747 VDD a_15467_1861# a_22977_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1748 a_11573_1923# a_11568_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1749 a_11013_6584# a_10138_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1750 VSS C[4] a_51044_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1751 VSS a_14010_5882# a_14012_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1752 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1753 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1754 a_20952_619# C[43] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1755 a_47982_5882# a_47216_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1756 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1757 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1758 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1759 a_13107_625# a_12937_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1760 VSS a_30571_1861# a_30447_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1761 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1762 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1763 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1764 VDD a_30571_1861# a_40783_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1765 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1766 a_1573_6584# a_698_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1767 a_17768_1758# a_17402_765# a_15782_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1768 VDD a_13265_3394# a_35892_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1769 a_34676_5882# a_35946_6337# a_36137_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.77e+11p ps=3.76e+06u w=650000u l=150000u
X1770 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1771 VSS a_51648_702# a_52573_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1772 VSS a_45598_6378# a_45571_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1773 VDD a_2572_702# a_3497_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1774 a_29110_6938# a_28342_6363# a_27124_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1775 a_2682_5882# a_1916_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1776 a_23334_702# a_24954_765# a_24778_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1777 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1778 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1779 a_19572_5882# a_20790_6363# a_21033_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1780 VDD C[3] a_52932_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1781 a_51758_5882# a_51044_6337# a_51662_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1782 a_19119_1923# a_19114_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1783 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1784 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1785 VDD a_27999_6584# a_27949_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1786 a_30093_625# a_29923_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1787 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1788 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1789 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1790 a_25334_6938# a_24566_6363# a_23348_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1791 a_12110_1758# a_11518_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1792 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1793 VSS C[1] a_56708_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1794 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1795 a_42310_702# a_41946_765# a_42214_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1796 VSS a_17780_5882# a_17782_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1797 VDD a_45669_1861# a_48329_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1798 a_6362_5882# a_7632_6337# a_7823_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1799 VDD a_26506_6337# a_26454_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1800 VDD a_34394_765# a_34218_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1801 a_34760_1758# a_34168_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1802 a_13900_702# a_15514_765# a_15338_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1803 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1804 a_2078_619# C[33] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1805 VSS a_41610_6337# a_41558_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1806 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1807 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1808 VDD a_18559_6584# a_18509_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1809 a_36282_765# a_36056_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1810 a_40326_702# a_41946_765# a_41770_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1811 a_38025_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1812 a_36111_1923# a_36106_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1813 a_15894_6938# a_15126_6363# a_13914_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1814 VDD a_20842_6337# a_21060_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1815 a_50649_6584# a_49774_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1816 VSS a_58201_6584# a_58151_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1817 a_38170_765# a_37944_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1818 VDD a_57044_765# a_56868_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1819 a_5935_5637# a_5962_6378# a_5947_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1820 a_10234_5882# a_9520_6337# a_10138_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1821 a_42214_702# a_41720_619# a_41775_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1822 a_4556_702# a_4558_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1823 a_19670_6938# a_18954_6337# a_17684_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1824 a_51758_5882# a_50992_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1825 a_7443_625# a_7273_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1826 VSS a_369_1861# a_7797_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1827 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1828 VSS a_34772_5882# a_34774_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1829 a_41720_619# C[54] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1830 a_6446_1758# a_6080_765# a_4460_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1831 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1832 a_21460_5882# a_20842_6337# a_21060_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1833 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1834 a_29108_5882# a_28342_6363# a_29012_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1835 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1836 VDD a_369_1861# a_2215_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1837 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1838 a_30886_702# a_32506_765# a_32330_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1839 VSS a_45669_1861# a_51209_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1840 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1841 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1842 a_56911_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1843 a_9711_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1844 a_28205_625# a_28035_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1845 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1846 a_25236_5882# a_24566_6363# a_24836_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1847 VDD a_35551_6584# a_35501_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1848 VSS a_48761_6584# a_48711_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1849 a_32886_6938# a_32118_6363# a_30900_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1850 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1851 a_53123_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1852 a_22541_625# a_22371_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1853 a_782_1758# a_416_765# a_n225_6339# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1854 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1855 a_5935_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1856 a_22895_1923# a_22890_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1857 a_22335_6584# a_21460_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1858 VSS a_25332_5882# a_25334_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1859 a_21544_1758# a_20952_619# a_19558_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1860 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1861 VSS a_15782_702# a_16707_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1862 a_11744_765# a_11518_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1863 a_29411_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1864 a_36662_6938# a_35946_6337# a_34676_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1865 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1866 a_10234_5882# a_9468_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1867 a_13632_765# a_13406_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1868 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1869 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1870 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1871 a_49760_702# a_51154_619# a_51204_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1872 a_59298_1758# a_58932_765# a_57312_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1873 a_15796_5882# a_15126_6363# a_15396_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1874 a_25635_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1875 a_27208_1758# a_26616_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1876 a_58787_5637# a_58814_6378# a_58799_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1877 a_45998_5882# a_47268_6337# a_47459_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1878 VSS a_11626_6378# a_11599_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1879 a_31981_625# a_31811_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1880 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1881 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1882 a_43103_6584# a_42228_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1883 a_42228_5882# a_41558_6363# a_41828_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1884 a_4572_6938# a_3804_6363# a_2586_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1885 a_42310_702# a_41720_619# a_42214_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1886 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1887 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1888 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1889 VDD a_49492_765# a_49316_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1890 a_416_765# a_190_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1891 a_8236_702# a_9630_619# a_9680_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1892 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1893 a_34662_702# a_34168_619# a_34223_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1894 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1895 a_8348_6938# a_7632_6337# a_6362_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X1896 VSS a_42324_5882# a_42326_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1897 a_58787_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1898 VDD a_5744_6337# a_5692_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1899 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1900 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1901 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1902 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 VSS a_15467_1861# a_29094_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1904 a_58843_1923# a_58756_1825# a_58761_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1905 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1906 a_57312_702# a_56818_619# a_56873_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1907 a_32788_5882# a_32118_6363# a_32388_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1908 a_12108_702# a_12110_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1909 VDD a_369_1861# a_10581_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1910 VDD a_9856_765# a_9680_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1911 VDD RESET sky130_fd_sc_hd__inv_4_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1912 VSS a_52932_6337# a_52880_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1913 a_36660_5882# a_35894_6363# a_36564_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1914 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1915 a_57424_6938# a_56656_6363# a_55438_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1916 a_51648_702# a_53268_765# a_53092_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1917 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1918 VDD a_80_6337# a_28_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1919 VSS a_15396_6378# a_15369_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1920 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1921 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1922 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1923 a_53634_1758# a_53042_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1924 a_47433_1923# a_47428_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1925 VSS a_30571_1861# a_30982_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1926 a_15277_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1927 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1928 VDD a_56313_6584# a_56263_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1929 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1930 a_43608_619# C[55] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1931 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1932 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1933 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1934 a_21556_5882# a_20842_6337# a_21460_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X1935 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1936 a_53648_6938# a_52880_6363# a_51662_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1937 VDD a_58596_6337# a_58544_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1938 VSS C[17] a_26506_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1939 a_4474_5882# a_3804_6363# a_4074_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1940 VDD a_24954_765# a_24778_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1941 VDD a_9520_6337# a_9738_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X1942 VSS a_46094_5882# a_46096_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1943 VSS a_36164_6378# a_36137_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1944 a_30996_5882# a_30230_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1945 a_26842_765# a_26616_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1946 a_1573_6584# a_698_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1947 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1948 VSS a_2572_702# a_3497_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1949 a_34758_702# a_34168_619# a_34662_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1950 VDD a_46873_6584# a_46823_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1951 a_28730_765# a_28504_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1952 a_34758_702# a_34394_765# a_34662_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1953 VDD a_32774_702# a_33699_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1954 VSS a_369_1861# a_2668_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1955 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1956 VSS a_32388_6378# a_32361_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1957 a_15878_702# a_15880_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1958 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1959 a_10124_702# a_9856_765# a_9685_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1960 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1961 a_38550_6938# a_38548_5882# a_38851_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1962 a_30093_625# a_29923_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1963 a_10124_702# a_11744_765# a_11568_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X1964 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1965 a_20447_6584# a_19572_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1966 VSS a_27999_6584# a_27949_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1967 a_39327_6584# a_38452_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1968 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1969 a_4873_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1970 a_57408_702# a_56818_619# a_57312_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1971 a_57408_702# a_57044_765# a_57312_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1972 a_21556_5882# a_20790_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1973 a_38025_5637# a_38052_6378# a_38037_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1974 a_796_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1975 a_49760_702# a_49266_619# a_49321_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1976 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1977 a_12026_5882# a_13296_6337# a_13487_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1978 VSS a_15178_6337# a_15126_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1979 VDD a_30571_1861# a_35119_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1980 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1981 a_34662_702# a_34394_765# a_34223_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1982 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1983 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1984 a_4059_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1985 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1986 VSS a_22948_6378# a_22921_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1987 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1988 VSS a_4074_6378# a_4047_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1989 a_32280_619# C[49] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1990 a_38895_1923# a_38536_1758# a_38534_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X1991 a_53550_5882# a_52880_6363# a_53150_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1992 VSS a_15467_1861# a_21007_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1993 a_1141_1923# a_782_1758# a_780_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X1994 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1995 VDD C[15] a_30282_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1996 a_29887_6584# a_29012_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1997 VSS a_18559_6584# a_18509_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1998 VSS a_369_1861# a_8332_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1999 VSS a_13265_3394# a_5690_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2000 a_46094_5882# a_45380_6337# a_45998_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2001 a_57312_702# a_57044_765# a_56873_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2002 a_50649_6584# a_49774_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2003 a_22933_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2004 a_6460_6938# a_6458_5882# a_6761_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2005 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2006 VSS a_45669_1861# a_51744_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2007 a_40058_765# a_39832_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2008 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2009 a_57725_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.1e+11p pd=2.42e+06u as=0p ps=0u w=1e+06u l=150000u
X2010 a_51746_1758# a_51154_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2011 a_7443_625# a_7273_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2012 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2013 a_56818_619# C[62] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2014 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2015 a_49872_6938# a_49870_5882# a_50173_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2016 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2017 a_58706_619# C[63] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2018 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2019 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2020 a_53949_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2021 a_29096_1758# a_28730_765# a_27110_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2022 a_6460_6938# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2023 VDD a_15467_1861# a_21903_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2024 VDD C[30] a_1968_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2025 a_10220_702# a_9630_619# a_10124_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2026 VDD a_23066_765# a_22890_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2027 a_15796_5882# a_17066_6337# a_17257_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2028 a_47982_5882# a_47216_6363# a_47886_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2029 a_43701_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2030 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2031 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2032 VSS a_35551_6584# a_35501_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2033 a_12026_5882# a_11356_6363# a_11626_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2034 VSS a_15467_1861# a_26671_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2035 a_45197_625# a_45027_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2036 VSS C[28] a_5744_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2037 a_22541_625# a_22371_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2038 a_44985_6584# a_44116_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2039 a_9630_619# C[37] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2040 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2041 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2042 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2043 a_271_5637# a_298_6378# a_283_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2044 a_49856_702# a_49266_619# a_49760_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2045 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2046 a_49856_702# a_49492_765# a_49760_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2047 a_6348_702# a_7742_619# a_7792_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2048 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2049 a_59312_6938# a_59310_5882# a_59613_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2050 VSS C[5] a_49156_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2051 VSS a_12122_5882# a_12124_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2052 a_28585_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2053 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2054 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2055 a_28641_1923# a_28554_1825# a_28559_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2056 a_30381_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2057 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2058 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2059 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2060 a_32788_5882# a_34058_6337# a_34249_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2061 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2062 VDD C[27] a_7632_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2063 VSS a_22730_6337# a_22678_6363# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2064 VSS a_35892_2529# a_45479_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2065 a_59657_1923# a_59298_1758# a_59296_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2066 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2067 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2068 a_27222_6938# a_26454_6363# a_25236_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2069 a_49760_702# a_49492_765# a_49321_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2070 a_21446_702# a_23066_765# a_22890_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2071 a_47471_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 VSS C[0] a_58596_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2073 a_17231_1923# a_17226_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2074 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2075 a_15277_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2076 VDD a_26111_6584# a_26061_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2077 VSS a_5690_2529# a_179_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2078 a_14012_6938# a_13296_6337# a_12026_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2079 VDD a_416_765# a_240_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2080 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2081 a_23446_6938# a_22678_6363# a_21460_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2082 VDD a_28394_6337# a_28342_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2083 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2084 a_34168_619# C[50] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2085 VDD a_8236_702# a_9161_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2086 a_45669_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2087 VSS a_15892_5882# a_15894_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2088 a_47968_702# a_47970_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2089 VDD a_45669_1861# a_46441_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2090 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2091 a_4474_5882# a_5744_6337# a_5935_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2092 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2093 a_42214_702# a_43834_765# a_43658_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2094 a_27222_6938# a_26506_6337# a_25236_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2095 VDD a_24618_6337# a_24566_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2096 VDD a_15514_765# a_15338_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2097 a_15880_1758# a_15288_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2098 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2099 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2100 a_37645_625# a_37475_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2101 VDD a_16671_6584# a_16621_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2102 a_44214_6938# a_43446_6363# a_42228_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2103 a_49347_5637# a_49374_6378# a_49359_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2104 a_17402_765# a_17176_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2105 a_4558_1758# a_3966_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2106 a_38438_702# a_40058_765# a_39882_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2107 a_53268_765# a_53042_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2108 a_34223_1923# a_34218_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2109 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2110 a_25318_702# a_24728_619# a_25222_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2111 VDD a_43103_6584# a_43053_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2112 VSS a_56313_6584# a_56263_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2113 VDD a_23334_702# a_24259_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2114 a_n225_6339# a_80_6337# a_271_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2115 a_2668_702# a_2670_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2116 a_30381_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2117 a_40438_6938# a_39670_6363# a_38452_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2118 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2119 a_17782_6938# a_17066_6337# a_15796_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2120 a_49347_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2121 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2122 VSS a_32884_5882# a_32886_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2123 a_4558_1758# a_4192_765# a_2572_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2124 a_38452_5882# a_37834_6337# a_38052_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2125 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2126 a_14010_5882# a_13244_6363# a_13914_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2127 a_57326_5882# a_58596_6337# a_58787_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2128 VDD a_47872_702# a_48797_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2129 a_28998_702# a_30618_765# a_30442_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2130 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2131 a_55023_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2132 VSS a_32774_702# a_33699_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2133 a_7823_5637# a_179_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2134 a_23348_5882# a_22678_6363# a_22948_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2135 a_780_702# a_416_765# a_684_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2136 VDD a_33663_6584# a_33613_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2137 VSS a_46873_6584# a_46823_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2138 a_25222_702# a_24954_765# a_24783_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2139 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2140 a_30998_6938# a_30230_6363# a_29012_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2141 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2142 a_20447_6584# a_19572_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2143 a_39887_1923# a_39882_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2144 a_39327_6584# a_38452_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2145 VSS a_23444_5882# a_23446_6938# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2146 a_38536_1758# a_37944_619# a_36550_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2147 a_29012_5882# a_28394_6337# a_28612_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2148 a_27523_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2149 a_51291_1923# a_51204_1825# a_51209_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.7e+11p ps=5.14e+06u w=1e+06u l=150000u
X2150 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2151 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2152 a_51744_702# a_51154_619# a_51648_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2153 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2154 a_51744_702# a_51380_765# a_51648_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=5.7e+11p pd=5.14e+06u as=0p ps=0u w=1e+06u l=150000u
X2155 a_19670_6938# a_19668_5882# a_19971_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2156 a_30618_765# a_30392_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2157 VSS a_45669_1861# a_58761_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2158 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2159 a_684_702# a_2304_765# a_2128_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2160 VDD a_49156_6337# a_49104_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2161 a_47378_619# C[57] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2162 a_684_702# a_416_765# a_245_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2163 VDD a_35892_2529# a_30571_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2164 a_684_702# a_190_619# a_245_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2165 a_23747_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2166 VDD a_5349_6584# a_5299_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2167 a_56899_5637# a_56926_6378# a_56911_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2168 a_698_5882# a_80_6337# a_298_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2169 a_49266_619# C[58] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2170 a_55520_702# a_55522_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2171 a_40340_5882# a_39670_6363# a_39940_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2172 a_17780_5882# a_17014_6363# a_17684_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2173 a_2684_6938# a_1916_6363# a_698_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2174 a_369_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2175 a_29887_6584# a_29012_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2176 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2177 a_15782_702# a_15288_619# a_15343_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2178 a_6460_6938# a_5744_6337# a_4474_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2179 a_51648_702# a_51380_765# a_51209_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2180 a_56899_5637# a_45479_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2181 a_51648_702# a_51154_619# a_51209_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2182 VDD a_2304_765# a_2128_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2183 VSS sky130_fd_sc_hd__inv_4_0/Y a_13265_3394# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2184 VDD a_3856_6337# a_3804_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2185 a_54985_1923# a_54980_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2186 VDD a_45669_1861# a_53179_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2187 a_29110_6938# a_29108_5882# a_29411_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2188 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2189 a_35892_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2190 VSS C[21] a_18954_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2191 a_44515_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2192 VSS C[11] a_37834_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2193 a_56955_1923# a_56868_1825# a_56873_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2194 a_4192_765# a_3966_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2195 a_782_1758# a_190_619# a_n225_6339# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2196 VDD a_35892_2529# a_30381_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2197 a_30900_5882# a_30230_6363# a_30500_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2198 VDD a_5690_2529# a_15467_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2199 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2200 a_6080_765# a_5854_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2201 a_40739_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2202 a_30571_1861# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2203 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2204 VSS a_35892_2529# a_45669_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2205 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2206 VSS a_5690_2529# a_15467_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2207 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2208 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2209 a_29110_6938# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2210 a_179_5549# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2211 a_796_6938# a_80_6337# a_n225_6339# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2212 a_45197_625# a_45027_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2213 a_7968_765# a_7742_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2214 a_34772_5882# a_34006_6363# a_34676_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2215 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2216 a_47970_1758# a_47604_765# a_45984_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2217 a_49760_702# a_51380_765# a_51204_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2218 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2219 a_45545_1923# a_45540_1825# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2220 a_29455_1923# a_29096_1758# a_29094_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2221 a_44985_6584# a_44116_5882# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2222 VDD a_54425_6584# a_54375_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2223 VSS C[16] a_28394_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2224 a_24728_619# C[45] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2225 a_38548_5882# a_37834_6337# a_38452_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=6e+11p pd=5.2e+06u as=0p ps=0u w=1e+06u l=150000u
X2226 VDD C[20] a_20842_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2227 a_19290_765# a_19064_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2228 a_49774_5882# a_50992_6363# a_51235_5637# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2229 a_59312_6938# a_58596_6337# a_57326_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2230 a_780_702# a_190_619# a_684_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2231 a_32884_5882# a_32118_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2232 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2233 VSS C[18] a_24618_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2234 a_2586_5882# a_1916_6363# a_2186_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2235 VSS a_5690_2529# a_15277_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2236 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2237 a_49774_5882# a_49156_6337# a_49374_6378# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2238 a_19145_5637# a_19172_6378# a_19157_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2239 a_30571_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2240 a_5690_2529# a_13265_3394# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2241 a_11219_625# a_11049_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2242 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2243 a_48285_5317# a_45479_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2244 VSS a_35892_2529# a_30571_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2245 a_17766_702# a_17768_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2246 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2247 VDD a_15467_1861# a_16239_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2248 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2249 a_20015_1923# a_19656_1758# a_19654_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2250 VSS a_5690_2529# a_369_1861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2251 a_15878_702# a_15288_619# a_15782_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2252 VDD a_44985_6584# a_44935_6365# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2253 a_15878_702# a_15514_765# a_15782_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2254 VSS a_369_1861# a_780_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2255 a_45716_765# a_45490_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2256 VDD a_49760_702# a_50685_625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X2257 VSS a_30500_6378# a_30473_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2258 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2259 a_8236_702# a_9856_765# a_9680_1825# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.015e+11p ps=1.92e+06u w=650000u l=150000u
X2260 a_34261_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2261 VSS a_13265_3394# a_35892_2529# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2262 VSS a_26111_6584# a_26061_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2263 a_37439_6584# a_36564_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2264 VDD a_51044_6337# a_51262_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2265 a_2985_5317# a_179_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2266 a_49858_1758# a_49266_619# a_47872_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2267 a_15467_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2268 a_10236_6938# a_9468_6363# a_8250_5882# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2269 VSS a_8236_702# a_9161_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2270 a_190_619# C[32] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2271 VSS C[9] a_41610_6337# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X2272 a_38548_5882# a_37782_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2273 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2274 a_794_5882# a_28_6363# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2275 a_19145_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2276 VDD a_38170_765# a_37994_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6e+11p ps=5.2e+06u w=1e+06u l=150000u
X2277 a_10138_5882# a_11408_6337# a_11599_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2278 a_34758_702# a_34760_1758# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2279 VDD a_30571_1861# a_33231_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2280 a_15782_702# a_15514_765# a_15343_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2281 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2282 a_2572_702# a_2078_619# a_2133_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2283 VDD a_11408_6337# a_11356_6363# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2284 a_59310_5882# a_58544_6363# a_59200_702# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2285 VSS a_39940_6378# a_39913_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2286 VSS a_2186_6378# a_2159_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2287 a_37007_1923# a_36648_1758# a_36646_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2288 a_51662_5882# a_50992_6363# a_51262_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2289 a_37645_625# a_37475_625# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X2290 VSS a_30571_1861# a_37999_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2291 a_24821_5317# a_15277_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2292 a_8348_6938# a_8346_5882# a_8649_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2293 a_13265_3394# sky130_fd_sc_hd__inv_4_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2294 VSS a_16671_6584# a_16621_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2295 a_51154_619# C[59] VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2296 a_9125_6584# a_8250_5882# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2297 VSS a_369_1861# a_6444_702# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2298 VDD a_5690_2529# a_15277_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2299 a_23348_5882# a_24618_6337# a_24809_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2300 a_55534_5882# a_54768_6363# a_55438_5882# VSS sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X2301 a_36662_6938# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2302 VSS a_23334_702# a_24259_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2303 a_15467_1861# a_5690_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2304 a_45669_1861# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2305 VDD a_5690_2529# a_369_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2306 VSS a_43103_6584# a_43053_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2307 a_4572_6938# a_4570_5882# a_4873_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2308 a_35892_2529# a_13265_3394# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2309 VSS a_35892_2529# a_30381_5549# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2310 VDD a_41946_765# a_41770_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2311 a_54631_625# a_54461_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2312 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2313 a_36137_5637# a_30381_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2314 a_39832_619# C[53] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2315 a_179_5549# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2316 VSS a_15467_1861# a_28559_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2317 a_8693_1923# a_8334_1758# a_8332_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2318 a_36550_702# a_37944_619# a_37994_1825# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2319 VSS a_47872_702# a_48797_625# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2320 a_27208_1758# a_26842_765# a_25222_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2321 a_43834_765# a_43608_619# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X2322 VDD C[31] a_80_6337# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2323 VDD a_30571_1861# a_38895_1923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2324 a_26697_5637# a_26724_6378# a_26709_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2325 a_13914_5882# a_15178_6337# a_15369_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2326 a_41813_5317# a_30381_5549# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2327 a_21178_765# a_20952_619# VSS VSS sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X2328 VSS a_55038_6378# a_55011_5637# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2329 a_52105_1923# a_51746_1758# a_51744_702# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2330 a_10138_5882# a_9468_6363# a_9738_6378# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2331 VSS a_15467_1861# a_24783_1923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2332 a_45479_5549# a_35892_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2333 VDD a_35892_2529# a_45479_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2334 VSS a_33663_6584# a_33613_6365# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X2335 a_26317_625# a_26147_625# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X2336 a_45479_5549# a_35892_2529# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2337 VDD a_35892_2529# a_45669_1861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2338 VDD a_5690_2529# a_179_5549# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2339 a_369_1861# a_5690_2529# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2340 a_49870_5882# a_49156_6337# a_49774_5882# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2341 VDD a_13265_3394# a_5690_2529# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2342 a_57424_6938# a_57422_5882# a_57725_5317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2343 a_26697_5637# a_15277_5549# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

