magic
tech sky130A
magscale 1 2
timestamp 1656570806
<< nwell >>
rect 14749 3456 15131 3777
rect 44891 3616 45273 3937
<< nsubdiff >>
rect 45016 3789 45150 3808
rect 45016 3755 45088 3789
rect 45122 3755 45150 3789
rect 45016 3738 45150 3755
rect 14874 3629 15008 3648
rect 14874 3595 14946 3629
rect 14980 3595 15008 3629
rect 14874 3578 15008 3595
<< nsubdiffcont >>
rect 45088 3755 45122 3789
rect 14946 3595 14980 3629
<< locali >>
rect 44813 3789 45356 3809
rect 44813 3755 45088 3789
rect 45122 3755 45356 3789
rect 44813 3737 45356 3755
rect 14671 3629 15214 3649
rect 14671 3595 14946 3629
rect 14980 3595 15214 3629
rect 14671 3577 15214 3595
<< viali >>
rect 43514 3669 43548 3714
rect 43682 3676 43716 3721
rect 43850 3666 43884 3711
rect 44018 3678 44052 3723
rect 44184 3676 44218 3721
rect 44350 3678 44384 3723
rect 44518 3678 44552 3723
rect 44692 3676 44726 3721
rect 45448 3670 45482 3715
rect 45610 3674 45644 3719
rect 45780 3678 45814 3723
rect 45944 3674 45978 3719
rect 46114 3674 46148 3719
rect 46282 3670 46316 3715
rect 46450 3674 46484 3719
rect 46624 3670 46658 3715
rect 43714 3578 43748 3612
rect 43814 3578 43848 3612
rect 43914 3578 43948 3612
rect 44014 3578 44048 3612
rect 44114 3578 44148 3612
rect 44214 3578 44248 3612
rect 44314 3578 44348 3612
rect 44414 3578 44448 3612
rect 45374 3578 45408 3612
rect 45474 3578 45508 3612
rect 45574 3578 45608 3612
rect 45674 3578 45708 3612
rect 45774 3578 45808 3612
rect 45874 3578 45908 3612
rect 45974 3578 46008 3612
rect 46074 3578 46108 3612
rect 13372 3509 13406 3554
rect 13540 3516 13574 3561
rect 13708 3506 13742 3551
rect 13876 3518 13910 3563
rect 14042 3516 14076 3561
rect 14208 3518 14242 3563
rect 14376 3518 14410 3563
rect 14550 3516 14584 3561
rect 15306 3510 15340 3555
rect 15468 3514 15502 3559
rect 15638 3518 15672 3563
rect 15802 3514 15836 3559
rect 15972 3514 16006 3559
rect 16140 3510 16174 3555
rect 16308 3514 16342 3559
rect 16482 3510 16516 3555
rect 13572 3418 13606 3452
rect 13672 3418 13706 3452
rect 13772 3418 13806 3452
rect 13872 3418 13906 3452
rect 13972 3418 14006 3452
rect 14072 3418 14106 3452
rect 14172 3418 14206 3452
rect 14272 3418 14306 3452
rect 15232 3418 15266 3452
rect 15332 3418 15366 3452
rect 15432 3418 15466 3452
rect 15532 3418 15566 3452
rect 15632 3418 15666 3452
rect 15732 3418 15766 3452
rect 15832 3418 15866 3452
rect 15932 3418 15966 3452
<< metal1 >>
rect 14423 4747 14678 5103
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14678 4747
rect 14423 4665 14678 4695
rect 44563 4747 44790 5115
rect 44563 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 44563 4661 44790 4695
rect 7079 4528 7615 4612
rect 22113 4537 22721 4595
rect 37217 4545 37841 4603
rect 52223 4551 52956 4609
rect 44732 3923 45399 3932
rect 44742 3874 45399 3923
rect 14642 3718 15291 3768
rect 14590 3710 15291 3718
rect 37381 3723 52816 3733
rect 37381 3721 44018 3723
rect 37381 3714 43682 3721
rect 37381 3713 37563 3714
rect 37381 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3669 43514 3714
rect 43548 3676 43682 3714
rect 43716 3711 44018 3721
rect 43716 3676 43850 3711
rect 43548 3669 43850 3676
rect 37615 3666 43850 3669
rect 43884 3678 44018 3711
rect 44052 3721 44350 3723
rect 44052 3678 44184 3721
rect 43884 3676 44184 3678
rect 44218 3678 44350 3721
rect 44384 3678 44518 3723
rect 44552 3721 45780 3723
rect 44552 3678 44692 3721
rect 44218 3676 44692 3678
rect 44726 3719 45780 3721
rect 44726 3715 45610 3719
rect 44726 3676 45448 3715
rect 43884 3670 45448 3676
rect 45482 3674 45610 3715
rect 45644 3678 45780 3719
rect 45814 3719 52816 3723
rect 45814 3678 45944 3719
rect 45644 3674 45944 3678
rect 45978 3674 46114 3719
rect 46148 3715 46450 3719
rect 46148 3674 46282 3715
rect 45482 3670 46282 3674
rect 46316 3674 46450 3715
rect 46484 3715 52816 3719
rect 46484 3674 46624 3715
rect 46316 3670 46624 3674
rect 46658 3714 52816 3715
rect 46658 3709 52664 3714
rect 46658 3670 52573 3709
rect 43884 3666 52573 3670
rect 37615 3662 52573 3666
rect 37512 3661 52573 3662
rect 37381 3657 52573 3661
rect 52625 3662 52664 3709
rect 52716 3662 52816 3714
rect 52625 3657 52816 3662
rect 37381 3652 52816 3657
rect 43682 3612 46285 3618
rect 43682 3578 43714 3612
rect 43748 3578 43814 3612
rect 43848 3578 43914 3612
rect 43948 3578 44014 3612
rect 44048 3578 44114 3612
rect 44148 3578 44214 3612
rect 44248 3578 44314 3612
rect 44348 3578 44414 3612
rect 44448 3578 45374 3612
rect 45408 3578 45474 3612
rect 45508 3578 45574 3612
rect 45608 3578 45674 3612
rect 45708 3578 45774 3612
rect 45808 3578 45874 3612
rect 45908 3578 45974 3612
rect 46008 3578 46074 3612
rect 46108 3578 46285 3612
rect 43682 3573 46285 3578
rect 7224 3563 22590 3573
rect 43682 3570 45128 3573
rect 7224 3561 13876 3563
rect 7224 3558 13540 3561
rect 7224 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3554 13540 3558
rect 7413 3509 13372 3554
rect 13406 3516 13540 3554
rect 13574 3551 13876 3561
rect 13574 3516 13708 3551
rect 13406 3509 13708 3516
rect 7413 3506 13708 3509
rect 13742 3518 13876 3551
rect 13910 3561 14208 3563
rect 13910 3518 14042 3561
rect 13742 3516 14042 3518
rect 14076 3518 14208 3561
rect 14242 3518 14376 3563
rect 14410 3561 15638 3563
rect 14410 3518 14550 3561
rect 14076 3516 14550 3518
rect 14584 3559 15638 3561
rect 14584 3555 15468 3559
rect 14584 3516 15306 3555
rect 13742 3510 15306 3516
rect 15340 3514 15468 3555
rect 15502 3518 15638 3559
rect 15672 3559 22590 3563
rect 15672 3518 15802 3559
rect 15502 3514 15802 3518
rect 15836 3514 15972 3559
rect 16006 3555 16308 3559
rect 16006 3514 16140 3555
rect 15340 3510 16140 3514
rect 16174 3514 16308 3555
rect 16342 3556 22590 3559
rect 16342 3555 22475 3556
rect 16342 3514 16482 3555
rect 16174 3510 16482 3514
rect 16516 3549 22475 3555
rect 16516 3510 22376 3549
rect 13742 3506 22376 3510
rect 7224 3497 22376 3506
rect 22428 3504 22475 3549
rect 22527 3504 22590 3556
rect 22428 3497 22590 3504
rect 7224 3492 22590 3497
rect 44978 3569 45128 3570
rect 44978 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3570 46285 3573
rect 45180 3521 45206 3570
rect 45075 3517 45206 3521
rect 44978 3478 45206 3517
rect 13540 3452 16143 3458
rect 13540 3418 13572 3452
rect 13606 3418 13672 3452
rect 13706 3418 13772 3452
rect 13806 3418 13872 3452
rect 13906 3418 13972 3452
rect 14006 3418 14072 3452
rect 14106 3418 14172 3452
rect 14206 3418 14272 3452
rect 14306 3418 15232 3452
rect 15266 3418 15332 3452
rect 15366 3418 15432 3452
rect 15466 3418 15532 3452
rect 15566 3418 15632 3452
rect 15666 3418 15732 3452
rect 15766 3418 15832 3452
rect 15866 3418 15932 3452
rect 15966 3418 16143 3452
rect 13540 3413 16143 3418
rect 13540 3410 14986 3413
rect 14836 3409 14986 3410
rect 14836 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3410 16143 3413
rect 15038 3361 15064 3410
rect 14933 3357 15064 3361
rect 14836 3318 15064 3357
rect 44732 3326 45484 3384
rect 13202 3148 13253 3244
rect 14590 3172 15271 3230
rect 19721 3175 45232 3219
rect 19721 3172 45120 3175
rect 13202 3147 13252 3148
rect 19721 3120 45031 3172
rect 45083 3123 45120 3172
rect 45172 3123 45232 3175
rect 45083 3120 45232 3123
rect 19721 3096 45232 3120
rect 19721 3044 45031 3096
rect 45083 3044 45124 3096
rect 45176 3044 45232 3096
rect 19721 3037 45232 3044
rect 14848 3013 45232 3037
rect 14848 2992 19927 3013
rect 14848 2940 14885 2992
rect 14937 2987 19927 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 19927 2987
rect 14848 2914 19927 2935
rect 14848 2912 14979 2914
rect 7015 2840 7678 2898
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 19927 2914
rect 14937 2860 19927 2862
rect 14848 2831 19927 2860
rect 22113 2852 22741 2910
rect 37125 2852 37888 2910
rect 52315 2843 52966 2901
<< via1 >>
rect 7264 4761 7316 4813
rect 7345 4760 7397 4812
rect 22380 4758 22432 4810
rect 22475 4758 22527 4810
rect 37457 4760 37509 4812
rect 37559 4760 37611 4812
rect 14443 4695 14495 4747
rect 14521 4695 14573 4747
rect 14614 4695 14666 4747
rect 44594 4695 44646 4747
rect 44677 4695 44729 4747
rect 52575 4733 52627 4785
rect 52670 4733 52722 4785
rect 6272 4537 6324 4589
rect 6379 4539 6431 4591
rect 6481 4539 6533 4591
rect 6581 4540 6633 4592
rect 21302 4543 21354 4595
rect 21405 4543 21457 4595
rect 21488 4543 21540 4595
rect 21589 4543 21641 4595
rect 21676 4543 21728 4595
rect 36434 4539 36486 4591
rect 36522 4539 36574 4591
rect 36607 4544 36659 4596
rect 53350 4536 53402 4588
rect 53444 4536 53496 4588
rect 53521 4536 53573 4588
rect 53601 4535 53653 4587
rect 53675 4536 53727 4588
rect 44600 3870 44652 3922
rect 44690 3871 44742 3923
rect 14467 3718 14519 3770
rect 14590 3718 14642 3770
rect 37460 3661 37512 3713
rect 37563 3662 37615 3714
rect 52573 3657 52625 3709
rect 52664 3662 52716 3714
rect 7265 3506 7317 3558
rect 7361 3506 7413 3558
rect 22376 3497 22428 3549
rect 22475 3504 22527 3556
rect 45023 3517 45075 3569
rect 45128 3521 45180 3573
rect 14881 3357 14933 3409
rect 14986 3361 15038 3413
rect 46035 3330 46087 3382
rect 46127 3331 46179 3383
rect 46217 3330 46269 3382
rect 46305 3329 46357 3381
rect 13680 3169 13732 3221
rect 13764 3169 13816 3221
rect 13857 3170 13909 3222
rect 45031 3120 45083 3172
rect 45120 3123 45172 3175
rect 45031 3044 45083 3096
rect 45124 3044 45176 3096
rect 14885 2940 14937 2992
rect 14979 2935 15031 2987
rect 6266 2843 6318 2895
rect 6364 2843 6416 2895
rect 6459 2843 6511 2895
rect 6564 2843 6616 2895
rect 14885 2860 14937 2912
rect 14979 2862 15031 2914
rect 21316 2848 21368 2900
rect 21416 2848 21468 2900
rect 21515 2848 21567 2900
rect 21618 2848 21670 2900
rect 36424 2842 36476 2894
rect 36512 2842 36564 2894
rect 36610 2838 36662 2890
rect 53346 2839 53398 2891
rect 53434 2839 53486 2891
rect 53517 2839 53569 2891
rect 53604 2839 53656 2891
rect 7265 2623 7317 2675
rect 7345 2621 7397 2673
rect 22381 2638 22433 2690
rect 22464 2638 22516 2690
rect 37459 2628 37511 2680
rect 37550 2628 37602 2680
rect 52576 2613 52628 2665
rect 52659 2613 52711 2665
<< metal2 >>
rect 7240 4813 7429 4843
rect 7240 4761 7264 4813
rect 7316 4812 7429 4813
rect 7316 4761 7345 4812
rect 7240 4760 7345 4761
rect 7397 4760 7429 4812
rect 6208 4592 6692 4719
rect 6208 4591 6581 4592
rect 6208 4589 6379 4591
rect 6208 4537 6272 4589
rect 6324 4539 6379 4589
rect 6431 4539 6481 4591
rect 6533 4540 6581 4591
rect 6633 4540 6692 4592
rect 6533 4539 6692 4540
rect 6324 4537 6692 4539
rect 6208 3372 6692 4537
rect 6208 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6692 3372
rect 6208 3257 6692 3316
rect 6208 3201 6275 3257
rect 6331 3201 6389 3257
rect 6445 3201 6503 3257
rect 6559 3201 6692 3257
rect 6208 3142 6692 3201
rect 6208 3086 6275 3142
rect 6331 3086 6389 3142
rect 6445 3086 6503 3142
rect 6559 3086 6692 3142
rect 6208 2895 6692 3086
rect 6208 2843 6266 2895
rect 6318 2843 6364 2895
rect 6416 2843 6459 2895
rect 6511 2843 6564 2895
rect 6616 2843 6692 2895
rect 6208 2729 6692 2843
rect 7240 3558 7429 4760
rect 14423 4747 14683 4818
rect 14423 4695 14443 4747
rect 14495 4695 14521 4747
rect 14573 4695 14614 4747
rect 14666 4695 14683 4747
rect 22351 4810 22540 4833
rect 22351 4758 22380 4810
rect 22432 4758 22475 4810
rect 22527 4758 22540 4810
rect 14423 3770 14683 4695
rect 14423 3718 14467 3770
rect 14519 3718 14590 3770
rect 14642 3718 14683 3770
rect 14423 3674 14683 3718
rect 21264 4595 21731 4697
rect 21264 4543 21302 4595
rect 21354 4543 21405 4595
rect 21457 4543 21488 4595
rect 21540 4543 21589 4595
rect 21641 4543 21676 4595
rect 21728 4543 21731 4595
rect 7240 3506 7265 3558
rect 7317 3506 7361 3558
rect 7413 3506 7429 3558
rect 7240 2675 7429 3506
rect 14848 3413 15054 3458
rect 14848 3409 14986 3413
rect 14848 3357 14881 3409
rect 14933 3361 14986 3409
rect 15038 3361 15054 3413
rect 14933 3357 15054 3361
rect 7240 2623 7265 2675
rect 7317 2673 7429 2675
rect 7317 2623 7345 2673
rect 7240 2621 7345 2623
rect 7397 2621 7429 2673
rect 13629 3222 13982 3268
rect 13629 3221 13857 3222
rect 13629 3169 13680 3221
rect 13732 3169 13764 3221
rect 13816 3170 13857 3221
rect 13909 3170 13982 3222
rect 13816 3169 13982 3170
rect 13629 2811 13982 3169
rect 14848 2992 15054 3357
rect 14848 2940 14885 2992
rect 14937 2987 15054 2992
rect 14937 2940 14979 2987
rect 14848 2935 14979 2940
rect 15031 2935 15054 2987
rect 14848 2914 15054 2935
rect 14848 2912 14979 2914
rect 14848 2860 14885 2912
rect 14937 2862 14979 2912
rect 15031 2862 15054 2914
rect 14937 2860 15054 2862
rect 14848 2831 15054 2860
rect 21264 3282 21731 4543
rect 21264 3226 21314 3282
rect 21370 3226 21418 3282
rect 21474 3226 21522 3282
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21264 3166 21731 3226
rect 21264 3110 21314 3166
rect 21370 3110 21418 3166
rect 21474 3110 21522 3166
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3050 21731 3110
rect 21264 2994 21314 3050
rect 21370 2994 21418 3050
rect 21474 2994 21522 3050
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 21264 2900 21731 2994
rect 21264 2848 21316 2900
rect 21368 2848 21416 2900
rect 21468 2848 21515 2900
rect 21567 2848 21618 2900
rect 21670 2848 21731 2900
rect 13629 2755 13669 2811
rect 13725 2755 13777 2811
rect 13833 2755 13885 2811
rect 13941 2755 13982 2811
rect 13629 2717 13982 2755
rect 21264 2746 21731 2848
rect 22351 3556 22540 4758
rect 37442 4812 37629 4831
rect 37442 4760 37457 4812
rect 37509 4760 37559 4812
rect 37611 4760 37629 4812
rect 22351 3549 22475 3556
rect 22351 3497 22376 3549
rect 22428 3504 22475 3549
rect 22527 3504 22540 3556
rect 22428 3497 22540 3504
rect 13629 2661 13669 2717
rect 13725 2661 13777 2717
rect 13833 2661 13885 2717
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 22351 2690 22540 3497
rect 36380 4596 36680 4695
rect 36380 4591 36607 4596
rect 36380 4539 36434 4591
rect 36486 4539 36522 4591
rect 36574 4544 36607 4591
rect 36659 4544 36680 4596
rect 36574 4539 36680 4544
rect 36380 3631 36680 4539
rect 36380 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36680 3631
rect 36380 3543 36680 3575
rect 36380 3487 36401 3543
rect 36457 3487 36495 3543
rect 36551 3487 36589 3543
rect 36645 3487 36680 3543
rect 36380 3455 36680 3487
rect 36380 3399 36401 3455
rect 36457 3399 36495 3455
rect 36551 3399 36589 3455
rect 36645 3399 36680 3455
rect 36380 2894 36680 3399
rect 36380 2842 36424 2894
rect 36476 2842 36512 2894
rect 36564 2890 36680 2894
rect 36564 2842 36610 2890
rect 36380 2838 36610 2842
rect 36662 2838 36680 2890
rect 36380 2743 36680 2838
rect 37442 3714 37629 4760
rect 44571 4747 44790 4800
rect 44571 4695 44594 4747
rect 44646 4695 44677 4747
rect 44729 4695 44790 4747
rect 44571 3923 44790 4695
rect 44571 3922 44690 3923
rect 44571 3870 44600 3922
rect 44652 3871 44690 3922
rect 44742 3871 44790 3923
rect 44652 3870 44790 3871
rect 44571 3835 44790 3870
rect 52546 4785 52735 4808
rect 52546 4733 52575 4785
rect 52627 4733 52670 4785
rect 52722 4733 52735 4785
rect 37442 3713 37563 3714
rect 37442 3661 37460 3713
rect 37512 3662 37563 3713
rect 37615 3662 37629 3714
rect 37512 3661 37629 3662
rect 22351 2638 22381 2690
rect 22433 2638 22464 2690
rect 22516 2638 22540 2690
rect 22351 2625 22540 2638
rect 37442 2680 37629 3661
rect 52546 3714 52735 4733
rect 52546 3709 52664 3714
rect 52546 3657 52573 3709
rect 52625 3662 52664 3709
rect 52716 3662 52735 3714
rect 52625 3657 52735 3662
rect 44990 3573 45196 3618
rect 44990 3569 45128 3573
rect 44990 3517 45023 3569
rect 45075 3521 45128 3569
rect 45180 3521 45196 3573
rect 45075 3517 45196 3521
rect 44990 3175 45196 3517
rect 44990 3172 45120 3175
rect 44990 3120 45031 3172
rect 45083 3123 45120 3172
rect 45172 3123 45196 3175
rect 45083 3120 45196 3123
rect 44990 3096 45196 3120
rect 44990 3044 45031 3096
rect 45083 3044 45124 3096
rect 45176 3044 45196 3096
rect 44990 3001 45196 3044
rect 45998 3383 46412 3405
rect 45998 3382 46127 3383
rect 45998 3330 46035 3382
rect 46087 3331 46127 3382
rect 46179 3382 46412 3383
rect 46179 3331 46217 3382
rect 46087 3330 46217 3331
rect 46269 3381 46412 3382
rect 46269 3330 46305 3381
rect 45998 3329 46305 3330
rect 46357 3329 46412 3381
rect 37442 2628 37459 2680
rect 37511 2628 37550 2680
rect 37602 2628 37629 2680
rect 7240 2603 7429 2621
rect 37442 2620 37629 2628
rect 45998 2784 46412 3329
rect 45998 2728 46035 2784
rect 46091 2728 46128 2784
rect 46184 2728 46221 2784
rect 46277 2728 46314 2784
rect 46370 2728 46412 2784
rect 45998 2702 46412 2728
rect 45998 2646 46035 2702
rect 46091 2646 46128 2702
rect 46184 2646 46221 2702
rect 46277 2646 46314 2702
rect 46370 2646 46412 2702
rect 45998 2609 46412 2646
rect 52546 2665 52735 3657
rect 53311 4588 53732 4695
rect 53311 4536 53350 4588
rect 53402 4536 53444 4588
rect 53496 4536 53521 4588
rect 53573 4587 53675 4588
rect 53573 4536 53601 4587
rect 53311 4535 53601 4536
rect 53653 4536 53675 4587
rect 53727 4536 53732 4588
rect 53653 4535 53732 4536
rect 53311 3176 53732 4535
rect 53311 3120 53348 3176
rect 53404 3120 53452 3176
rect 53508 3120 53556 3176
rect 53612 3120 53660 3176
rect 53716 3120 53732 3176
rect 53311 3086 53732 3120
rect 53311 3030 53348 3086
rect 53404 3030 53452 3086
rect 53508 3030 53556 3086
rect 53612 3030 53660 3086
rect 53716 3030 53732 3086
rect 53311 2891 53732 3030
rect 53311 2839 53346 2891
rect 53398 2839 53434 2891
rect 53486 2839 53517 2891
rect 53569 2839 53604 2891
rect 53656 2839 53732 2891
rect 53311 2745 53732 2839
rect 52546 2613 52576 2665
rect 52628 2613 52659 2665
rect 52711 2613 52735 2665
rect 52546 2600 52735 2613
<< via2 >>
rect 6275 3316 6331 3372
rect 6389 3316 6445 3372
rect 6503 3316 6559 3372
rect 6275 3201 6331 3257
rect 6389 3201 6445 3257
rect 6503 3201 6559 3257
rect 6275 3086 6331 3142
rect 6389 3086 6445 3142
rect 6503 3086 6559 3142
rect 21314 3226 21370 3282
rect 21418 3226 21474 3282
rect 21522 3226 21578 3282
rect 21626 3226 21682 3282
rect 21314 3110 21370 3166
rect 21418 3110 21474 3166
rect 21522 3110 21578 3166
rect 21626 3110 21682 3166
rect 21314 2994 21370 3050
rect 21418 2994 21474 3050
rect 21522 2994 21578 3050
rect 21626 2994 21682 3050
rect 13669 2755 13725 2811
rect 13777 2755 13833 2811
rect 13885 2755 13941 2811
rect 13669 2661 13725 2717
rect 13777 2661 13833 2717
rect 13885 2661 13941 2717
rect 36401 3575 36457 3631
rect 36495 3575 36551 3631
rect 36589 3575 36645 3631
rect 36401 3487 36457 3543
rect 36495 3487 36551 3543
rect 36589 3487 36645 3543
rect 36401 3399 36457 3455
rect 36495 3399 36551 3455
rect 36589 3399 36645 3455
rect 46035 2728 46091 2784
rect 46128 2728 46184 2784
rect 46221 2728 46277 2784
rect 46314 2728 46370 2784
rect 46035 2646 46091 2702
rect 46128 2646 46184 2702
rect 46221 2646 46277 2702
rect 46314 2646 46370 2702
rect 53348 3120 53404 3176
rect 53452 3120 53508 3176
rect 53556 3120 53612 3176
rect 53660 3120 53716 3176
rect 53348 3030 53404 3086
rect 53452 3030 53508 3086
rect 53556 3030 53612 3086
rect 53660 3030 53716 3086
<< metal3 >>
rect 36378 3631 36682 3645
rect 36378 3575 36401 3631
rect 36457 3575 36495 3631
rect 36551 3575 36589 3631
rect 36645 3575 36682 3631
rect 36378 3543 36682 3575
rect 36378 3487 36401 3543
rect 36457 3532 36495 3543
rect 36551 3533 36589 3543
rect 36645 3533 36682 3543
rect 36551 3487 36568 3533
rect 36378 3455 36414 3487
rect 36501 3455 36568 3487
rect 6274 3398 6616 3431
rect 36378 3399 36401 3455
rect 36551 3421 36568 3455
rect 36655 3421 36682 3533
rect 36457 3399 36495 3420
rect 36551 3399 36589 3421
rect 36645 3399 36682 3421
rect 6206 3372 6695 3398
rect 36378 3379 36682 3399
rect 6206 3316 6275 3372
rect 6331 3316 6389 3372
rect 6445 3316 6503 3372
rect 6559 3316 6695 3372
rect 6206 3257 6695 3316
rect 6206 3229 6275 3257
rect 6331 3229 6389 3257
rect 6445 3235 6503 3257
rect 6559 3235 6695 3257
rect 6206 3138 6272 3229
rect 6358 3201 6389 3229
rect 6559 3201 6568 3235
rect 6358 3144 6423 3201
rect 6509 3144 6568 3201
rect 6654 3144 6695 3235
rect 6358 3142 6695 3144
rect 6358 3138 6389 3142
rect 6206 3086 6275 3138
rect 6331 3086 6389 3138
rect 6445 3086 6503 3142
rect 6559 3086 6695 3142
rect 6206 3031 6695 3086
rect 21264 3282 21731 3336
rect 21264 3239 21314 3282
rect 21370 3239 21418 3282
rect 21264 3155 21312 3239
rect 21405 3226 21418 3239
rect 21474 3239 21522 3282
rect 21474 3226 21479 3239
rect 21578 3226 21626 3282
rect 21682 3226 21731 3282
rect 21405 3166 21479 3226
rect 21572 3166 21731 3226
rect 21405 3155 21418 3166
rect 21264 3110 21314 3155
rect 21370 3110 21418 3155
rect 21474 3155 21479 3166
rect 21474 3110 21522 3155
rect 21578 3110 21626 3166
rect 21682 3110 21731 3166
rect 21264 3078 21731 3110
rect 21264 2994 21312 3078
rect 21405 3050 21479 3078
rect 21572 3050 21731 3078
rect 21405 2994 21418 3050
rect 21474 2994 21479 3050
rect 21578 2994 21626 3050
rect 21682 2994 21731 3050
rect 53311 3183 53733 3204
rect 53311 3176 53355 3183
rect 53439 3176 53476 3183
rect 53560 3176 53614 3183
rect 53698 3176 53733 3183
rect 53311 3120 53348 3176
rect 53439 3120 53452 3176
rect 53612 3120 53614 3176
rect 53716 3120 53733 3176
rect 53311 3086 53355 3120
rect 53439 3086 53476 3120
rect 53560 3086 53614 3120
rect 53698 3086 53733 3120
rect 53311 3030 53348 3086
rect 53439 3030 53452 3086
rect 53612 3030 53614 3086
rect 53716 3030 53733 3086
rect 53311 3025 53355 3030
rect 53439 3025 53476 3030
rect 53560 3025 53614 3030
rect 53698 3025 53733 3030
rect 53311 2996 53733 3025
rect 21264 2950 21731 2994
rect 13629 2811 13982 2834
rect 13629 2763 13669 2811
rect 13725 2763 13777 2811
rect 13833 2763 13885 2811
rect 13629 2694 13653 2763
rect 13730 2694 13756 2763
rect 13833 2694 13859 2763
rect 13941 2755 13982 2811
rect 13936 2717 13982 2755
rect 13629 2661 13669 2694
rect 13725 2661 13777 2694
rect 13833 2661 13885 2694
rect 13941 2661 13982 2717
rect 13629 2635 13982 2661
rect 45998 2808 46413 2851
rect 45998 2807 46176 2808
rect 45998 2784 46036 2807
rect 46120 2784 46176 2807
rect 46260 2784 46304 2808
rect 45998 2728 46035 2784
rect 46120 2728 46128 2784
rect 46277 2728 46304 2784
rect 45998 2702 46036 2728
rect 46120 2702 46176 2728
rect 46260 2702 46304 2728
rect 45998 2646 46035 2702
rect 46120 2649 46128 2702
rect 46277 2650 46304 2702
rect 46388 2650 46413 2808
rect 46091 2646 46128 2649
rect 46184 2646 46221 2650
rect 46277 2646 46314 2650
rect 46370 2646 46413 2650
rect 45998 2610 46413 2646
<< via3 >>
rect 2518 7211 2624 7389
rect 2727 7210 2833 7388
rect 2893 7210 2999 7388
rect 3073 7212 3179 7390
rect 1284 5093 1390 5271
rect 1456 5094 1562 5272
rect 1630 5093 1736 5271
rect 36414 3487 36457 3532
rect 36457 3487 36495 3532
rect 36495 3487 36501 3532
rect 36568 3487 36589 3533
rect 36589 3487 36645 3533
rect 36645 3487 36655 3533
rect 36414 3455 36501 3487
rect 36568 3455 36655 3487
rect 36414 3420 36457 3455
rect 36457 3420 36495 3455
rect 36495 3420 36501 3455
rect 36568 3421 36589 3455
rect 36589 3421 36645 3455
rect 36645 3421 36655 3455
rect 6272 3201 6275 3229
rect 6275 3201 6331 3229
rect 6331 3201 6358 3229
rect 6423 3201 6445 3235
rect 6445 3201 6503 3235
rect 6503 3201 6509 3235
rect 6272 3142 6358 3201
rect 6423 3144 6509 3201
rect 6568 3144 6654 3235
rect 6272 3138 6275 3142
rect 6275 3138 6331 3142
rect 6331 3138 6358 3142
rect 21312 3226 21314 3239
rect 21314 3226 21370 3239
rect 21370 3226 21405 3239
rect 21479 3226 21522 3239
rect 21522 3226 21572 3239
rect 21312 3166 21405 3226
rect 21479 3166 21572 3226
rect 21312 3155 21314 3166
rect 21314 3155 21370 3166
rect 21370 3155 21405 3166
rect 21479 3155 21522 3166
rect 21522 3155 21572 3166
rect 21312 3050 21405 3078
rect 21479 3050 21572 3078
rect 21312 2994 21314 3050
rect 21314 2994 21370 3050
rect 21370 2994 21405 3050
rect 21479 2994 21522 3050
rect 21522 2994 21572 3050
rect 53355 3176 53439 3183
rect 53476 3176 53560 3183
rect 53614 3176 53698 3183
rect 53355 3120 53404 3176
rect 53404 3120 53439 3176
rect 53476 3120 53508 3176
rect 53508 3120 53556 3176
rect 53556 3120 53560 3176
rect 53614 3120 53660 3176
rect 53660 3120 53698 3176
rect 53355 3086 53439 3120
rect 53476 3086 53560 3120
rect 53614 3086 53698 3120
rect 53355 3030 53404 3086
rect 53404 3030 53439 3086
rect 53476 3030 53508 3086
rect 53508 3030 53556 3086
rect 53556 3030 53560 3086
rect 53614 3030 53660 3086
rect 53660 3030 53698 3086
rect 53355 3025 53439 3030
rect 53476 3025 53560 3030
rect 53614 3025 53698 3030
rect 13653 2755 13669 2763
rect 13669 2755 13725 2763
rect 13725 2755 13730 2763
rect 13653 2717 13730 2755
rect 13653 2694 13669 2717
rect 13669 2694 13725 2717
rect 13725 2694 13730 2717
rect 13756 2755 13777 2763
rect 13777 2755 13833 2763
rect 13756 2717 13833 2755
rect 13756 2694 13777 2717
rect 13777 2694 13833 2717
rect 13859 2755 13885 2763
rect 13885 2755 13936 2763
rect 13859 2717 13936 2755
rect 13859 2694 13885 2717
rect 13885 2694 13936 2717
rect 46036 2784 46120 2807
rect 46176 2784 46260 2808
rect 46304 2784 46388 2808
rect 46036 2728 46091 2784
rect 46091 2728 46120 2784
rect 46176 2728 46184 2784
rect 46184 2728 46221 2784
rect 46221 2728 46260 2784
rect 46304 2728 46314 2784
rect 46314 2728 46370 2784
rect 46370 2728 46388 2784
rect 46036 2702 46120 2728
rect 46176 2702 46260 2728
rect 46304 2702 46388 2728
rect 46036 2649 46091 2702
rect 46091 2649 46120 2702
rect 46176 2650 46184 2702
rect 46184 2650 46221 2702
rect 46221 2650 46260 2702
rect 46304 2650 46314 2702
rect 46314 2650 46370 2702
rect 46370 2650 46388 2702
rect 1286 2145 1392 2323
rect 1491 2147 1597 2325
rect 1690 2147 1796 2325
rect 2532 34 2638 212
rect 2753 34 2859 212
rect 2962 34 3068 212
rect 3136 34 3242 212
rect 6260 66 6346 157
rect 6408 66 6494 157
rect 6556 66 6642 157
rect 13779 140 13856 209
rect 13802 21 13879 90
rect 21317 61 21413 169
rect 21450 61 21546 169
rect 21583 61 21679 169
rect 36412 45 36499 157
rect 36581 45 36668 157
rect 46038 32 46122 190
rect 46151 32 46235 190
rect 46266 32 46350 190
rect 53361 42 53445 200
rect 53480 42 53564 200
rect 53609 42 53693 200
<< metal4 >>
rect 2467 7390 3251 7443
rect 2467 7389 3073 7390
rect 2467 7211 2518 7389
rect 2624 7388 3073 7389
rect 2624 7211 2727 7388
rect 2467 7210 2727 7211
rect 2833 7210 2893 7388
rect 2999 7212 3073 7388
rect 3179 7212 3251 7390
rect 2999 7210 3251 7212
rect 1234 5272 1852 5401
rect 1234 5271 1456 5272
rect 1234 5093 1284 5271
rect 1390 5094 1456 5271
rect 1562 5271 1852 5272
rect 1562 5094 1630 5271
rect 1390 5093 1630 5094
rect 1736 5093 1852 5271
rect 1234 2325 1852 5093
rect 1234 2323 1491 2325
rect 1234 2145 1286 2323
rect 1392 2147 1491 2323
rect 1597 2147 1690 2325
rect 1796 2147 1852 2325
rect 1392 2145 1852 2147
rect 1234 2095 1852 2145
rect 2467 212 3251 7210
rect 36378 3533 36683 3690
rect 36378 3532 36568 3533
rect 36378 3420 36414 3532
rect 36501 3421 36568 3532
rect 36655 3421 36683 3533
rect 36501 3420 36683 3421
rect 2467 34 2532 212
rect 2638 34 2753 212
rect 2859 34 2962 212
rect 3068 34 3136 212
rect 3242 34 3251 212
rect 2467 -55 3251 34
rect 6214 3235 6683 3350
rect 6214 3229 6423 3235
rect 6214 3138 6272 3229
rect 6358 3144 6423 3229
rect 6509 3144 6568 3235
rect 6654 3144 6683 3235
rect 6358 3138 6683 3144
rect 6214 157 6683 3138
rect 21264 3239 21731 3364
rect 21264 3155 21312 3239
rect 21405 3155 21479 3239
rect 21572 3155 21731 3239
rect 21264 3078 21731 3155
rect 21264 2994 21312 3078
rect 21405 2994 21479 3078
rect 21572 2994 21731 3078
rect 13629 2763 13983 2835
rect 13629 2694 13653 2763
rect 13730 2694 13756 2763
rect 13833 2694 13859 2763
rect 13936 2694 13983 2763
rect 13629 2634 13983 2694
rect 6214 66 6260 157
rect 6346 66 6408 157
rect 6494 66 6556 157
rect 6642 66 6683 157
rect 6214 -33 6683 66
rect 13705 209 13906 2634
rect 13705 140 13779 209
rect 13856 140 13906 209
rect 13705 90 13906 140
rect 13705 21 13802 90
rect 13879 21 13906 90
rect 13705 -58 13906 21
rect 21264 169 21731 2994
rect 21264 61 21317 169
rect 21413 61 21450 169
rect 21546 61 21583 169
rect 21679 61 21731 169
rect 21264 -8 21731 61
rect 36378 157 36683 3420
rect 53311 3183 53736 3206
rect 53311 3025 53355 3183
rect 53439 3025 53476 3183
rect 53560 3025 53614 3183
rect 53698 3025 53736 3183
rect 36378 45 36412 157
rect 36499 45 36581 157
rect 36668 45 36683 157
rect 36378 -3 36683 45
rect 45998 2808 46412 2897
rect 45998 2807 46176 2808
rect 45998 2649 46036 2807
rect 46120 2650 46176 2807
rect 46260 2650 46304 2808
rect 46388 2650 46412 2808
rect 46120 2649 46412 2650
rect 45998 190 46412 2649
rect 45998 32 46038 190
rect 46122 32 46151 190
rect 46235 32 46266 190
rect 46350 32 46412 190
rect 45998 -56 46412 32
rect 53311 200 53736 3025
rect 53311 42 53361 200
rect 53445 42 53480 200
rect 53564 42 53609 200
rect 53693 42 53736 200
rect 53311 -44 53736 42
use nbrhalf  nbrhalf_0
timestamp 1656566743
transform 1 0 3552 0 1 -2528
box -3552 2527 26658 5446
use nbrhalf  nbrhalf_1
timestamp 1656566743
transform 1 0 33754 0 1 -2528
box -3552 2527 26658 5446
use nbrhalf  nbrhalf_2
timestamp 1656566743
transform -1 0 56430 0 -1 9968
box -3552 2527 26658 5446
use nbrhalf  nbrhalf_3
timestamp 1656566743
transform -1 0 26228 0 -1 9968
box -3552 2527 26658 5446
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654402208
transform 1 0 15169 0 1 3195
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654402208
transform 1 0 13239 0 1 3195
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1654402208
transform 1 0 45311 0 1 3355
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1654402208
transform 1 0 43381 0 1 3355
box -38 -48 1510 592
<< end >>
