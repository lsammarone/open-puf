**.subckt nor_tb
x1 net2 net1 VGND VNB VPB VPWR IN1 sky130_fd_sc_hd__nor2_1
V1 net2 GND PULSE(1.8 0 0ns 10ps 10ps 2ns 5ns)
V2 net1 GND 0
XM1 IN1 net4 out GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 IN1 net3 out out sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 IN2 net3 out GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 IN2 net4 out out sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
V3 out GND 1.8
x2 net4 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__inv_1
V4 net4 GND 1.8
x3 net6 net5 VGND VNB VPB VPWR IN2 sky130_fd_sc_hd__nor2_1
V5 net6 GND PULSE(1.8 0 0ns 10ps 10ps 2ns 5ns)
V6 net5 GND 0
x4 net2 net1 VGND VNB VPB VPWR IN1 sky130_fd_sc_hd__nor2_1
V7 net2 GND PULSE(1.8 0 0ns 10ps 10ps 2ns 5ns)
V8 net1 GND 0
**** begin user architecture code


.lib /farmshare/home/classes/ee/272/PDKs/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /farmshare/home/classes/ee/272/PDKs/open_pdks/sky130/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice






.control
save all
tran 1n 10n
plot out IN1 IN2
.endc


**** end user architecture code
**.ends
.GLOBAL GND
** flattened .save nodes
.end
