* NGSPICE file created from BR128_flat.ext - technology: sky130A

.subckt BR128_flat OUT C[127] C[126] C[125] C[124] C[123] C[122] C[121] C[120] C[119]
+ C[118] C[117] C[116] C[115] C[114] C[113] C[112] C[63] C[62] C[61] C[60] C[59] C[58]
+ C[57] C[56] C[55] C[54] C[53] C[52] C[51] C[50] C[49] C[48] RESET C[111] C[110]
+ C[109] C[108] C[107] C[106] C[105] C[104] C[103] C[102] C[101] C[100] C[99] C[98]
+ C[97] C[96] C[32] C[33] C[34] C[35] C[36] C[37] C[38] C[39] C[40] C[41] C[42] C[43]
+ C[44] C[45] C[46] C[47] C[0] C[1] C[2] C[3] C[4] C[5] C[7] C[8] C[9] C[10] C[11]
+ C[12] C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24] C[25]
+ C[26] C[27] C[28] C[29] C[30] C[6] C[31] C[95] C[94] C[93] C[92] C[91] C[90] C[89]
+ C[88] C[87] C[86] C[85] C[84] C[83] C[82] C[81] C[80] C[79] C[78] C[77] C[76] C[75]
+ C[74] C[73] C[72] C[71] C[70] C[69] C[68] C[67] C[66] C[65] C[64] VSS VDD
X0 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VDD a_18085_739# a_18033_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_4480_928# a_3605_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4 a_13143_510# a_13141_1566# a_13454_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_3701_1566# a_2987_739# a_3605_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VSS a_31072_18706# a_31020_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VSS a_32960_18706# a_32908_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_56214_13071# a_57608_12988# a_57648_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_22197_6419# a_21971_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_48989_5620# a_48397_6509# a_47003_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_22250_18251# a_23520_18706# a_23711_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_58102_13071# a_59496_12988# a_59536_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_26124_19307# a_25408_18706# a_24138_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VDD a_46170_18706# a_46388_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_56228_18251# a_55610_18706# a_55828_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VDD a_19973_739# a_20191_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VDD a_38853_739# a_39071_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_49757_12994# a_49587_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X25 a_58212_18251# a_57498_18706# a_58116_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_10350_6503# a_10180_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X28 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_29802_18251# a_31072_18706# a_31263_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_16078_12988# C[104] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_50330_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VDD a_2758_18706# a_2706_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 VDD a_53722_18706# a_53940_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_17966_12988# C[105] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VSS C[81] a_27525_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_33676_19307# a_32960_18706# a_31690_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 VDD a_42234_928# a_42184_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X42 a_37156_1811# a_37183_1000# a_37168_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_24236_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 a_59725_6509# C[63] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_45217_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X47 VDD a_37301_6419# a_37115_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 VDD C[26] a_10310_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 a_60100_18251# a_59334_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_29900_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X54 VSS a_3591_6676# a_4516_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X55 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X56 a_22250_18251# a_23468_18732# a_23711_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 a_13488_5455# a_13129_5620# a_13127_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_39340_19307# a_39338_18251# a_39651_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X60 a_54569_1566# a_55839_739# a_56030_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X61 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X62 VDD C[31] a_870_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X64 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 a_14651_6419# a_14425_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 VDD C[30] a_2758_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 a_50101_14292# a_50096_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X68 a_16304_13134# a_16078_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X69 a_36846_12988# C[115] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X70 VDD a_56443_6676# a_57368_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X71 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X72 a_475_18953# a_565_18708# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X73 a_29802_18251# a_31020_18732# a_31263_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 VDD a_45775_18953# a_45725_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X75 a_26108_13071# a_25744_13134# a_26012_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 a_27996_13071# a_27632_13134# a_27900_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_30017_6676# a_29749_6419# a_29568_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X78 a_55949_6509# C[61] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 a_10730_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X80 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X81 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_56671_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 VSS a_29018_928# a_28968_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X83 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 a_12912_18251# a_12146_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X85 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X86 a_23856_13134# a_23630_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X87 a_41359_1566# a_40741_739# a_40959_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X88 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X89 VDD a_29413_739# a_29631_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X90 a_41130_18251# a_42348_18732# a_42591_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X91 VDD a_57103_18953# a_57053_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X92 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X93 a_10875_6419# a_10649_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_13031_6676# a_14651_6419# a_14465_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X95 a_13143_510# a_12427_739# a_11157_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X96 VDD a_35077_739# a_35025_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X97 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 VDD C[65] a_57727_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 a_39189_6419# a_38963_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X100 a_18572_19307# a_17804_18732# a_16586_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X101 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X102 a_35184_13134# a_34958_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X103 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X104 VDD a_32794_928# a_32744_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X105 a_46361_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X106 a_27716_1811# a_27743_1000# a_27728_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_10547_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X108 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X109 VSS a_1088_18747# a_1061_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X110 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X111 a_59496_12988# C[127] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 VDD a_27861_6419# a_27675_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 a_32017_510# a_31249_765# a_30031_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X114 VSS a_37679_1566# a_37681_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X115 a_42736_13134# a_42510_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X116 a_16913_510# a_16911_1566# a_17224_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X117 a_47663_18953# a_46788_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X118 VDD a_8987_6419# a_8801_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X119 a_32328_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X120 VSS a_17856_18706# a_17804_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X121 a_53913_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X122 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X123 a_3472_18251# a_2706_18732# a_3376_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X124 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X125 VSS a_42629_739# a_42577_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X126 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X127 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X128 a_58525_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X129 a_9026_13071# a_10646_13134# a_10460_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X130 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_8659_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 VDD a_47003_6676# a_47928_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X132 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X133 a_14704_18251# a_15968_18706# a_16159_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X134 a_37452_19307# a_36684_18732# a_35466_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X135 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X136 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X137 a_20577_6676# a_20309_6419# a_20128_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X138 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_15376_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 a_18572_19307# a_17856_18706# a_16586_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X141 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X142 a_39457_6676# a_39189_6419# a_39008_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X143 a_794_737# a_1206_13134# a_1020_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X144 VDD a_46004_928# a_45954_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X145 a_43116_19307# a_42348_18732# a_41130_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X146 a_9124_14127# a_8532_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X147 a_45004_19307# a_44236_18732# a_43018_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X148 a_31919_1566# a_31301_739# a_31519_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X149 a_26255_1566# a_27473_765# a_27716_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X150 a_56042_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X151 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_48987_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X152 VSS C[23] a_15968_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X153 VSS a_36736_18706# a_36684_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X154 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 a_1474_13071# a_2868_12988# a_2908_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 a_16307_6509# C[40] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X157 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 a_27762_5455# a_27675_5687# a_27680_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 a_1488_18251# a_870_18706# a_1088_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X160 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X161 a_21672_6503# a_21502_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X162 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X163 a_3472_18251# a_2758_18706# a_3376_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X164 a_55994_5455# a_55989_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X165 a_29749_6419# a_29523_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X166 a_17258_5455# a_16899_5620# a_16897_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X167 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X168 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X169 a_23757_14292# a_23670_14194# a_23675_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 VDD a_58102_13071# a_59027_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X171 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X172 a_33578_18251# a_34848_18706# a_35039_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X173 a_18421_6419# a_18195_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 a_37452_19307# a_36736_18706# a_35466_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X175 a_49757_12994# a_49587_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X176 a_32001_6676# a_32003_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 VDD a_4480_928# a_4430_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X178 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X179 VSS a_28239_1566# a_28241_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X180 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_11010_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X181 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X182 a_28225_6676# a_27635_6509# a_28129_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X183 a_28129_6676# a_29749_6419# a_29563_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X184 VSS C[13] a_34848_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X185 VSS C[12] a_36736_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X186 VSS a_56443_6676# a_57368_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X187 a_44708_1811# a_44735_1000# a_44720_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X188 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X189 a_20687_1566# a_19921_765# a_20591_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X190 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_3458_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X191 a_39567_1566# a_38801_765# a_39471_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X192 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X193 VSS a_40346_928# a_40296_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X194 a_33905_510# a_33903_1566# a_34216_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X195 VSS C[9] a_42400_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X196 a_54438_19307# a_54436_18251# a_54749_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X197 a_42637_14292# a_42550_14194# a_42555_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X198 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X199 VDD a_29184_18706# a_29132_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X200 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X201 VSS a_24463_1566# a_24465_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X202 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X203 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X204 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_50875_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X205 a_55765_14292# a_55760_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X206 a_50056_12988# C[122] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X207 a_51944_12988# C[123] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X208 a_18474_18251# a_17804_18732# a_18074_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X209 a_46602_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X210 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X211 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_14470_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X212 a_3605_1566# a_2987_739# a_3205_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X213 a_11253_1566# a_10539_739# a_11157_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X214 a_11012_14127# a_10420_12988# a_9026_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X215 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_40978_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X216 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X217 VSS a_12912_18251# a_12914_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X218 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X219 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X220 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X221 a_9136_18251# a_8370_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X222 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X223 a_1435_6419# a_1209_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X224 a_5479_6676# a_4985_6509# a_5030_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X225 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X226 a_42211_12994# a_42041_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X227 a_33299_6509# C[49] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X228 a_29018_928# a_28143_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X229 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X230 VDD a_18192_13134# a_18006_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X231 a_22561_6676# a_22563_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X232 a_44754_5455# a_44667_5687# a_44672_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 a_14277_18006# a_14304_18747# a_14289_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X234 a_50282_13134# a_50056_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X235 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X236 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X237 a_14241_14292# a_14236_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X238 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_33115_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X239 a_11337_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X240 a_7236_14127# a_6644_12988# a_5250_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X241 a_10420_12988# C[101] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X242 a_60086_13071# a_59722_13134# a_59990_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X243 a_37354_18251# a_36684_18732# a_36954_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X244 a_4756_12988# C[98] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X245 a_18689_6676# a_20309_6419# a_20123_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X246 a_37569_6676# a_39189_6419# a_39003_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X247 a_20446_14127# a_19854_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X248 VDD a_25744_13134# a_25558_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X249 a_18785_6676# a_18195_6509# a_18689_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X250 a_35413_6419# a_35187_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X251 VSS a_47003_6676# a_47928_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X252 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X253 VSS a_58991_18953# a_58941_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X254 a_7248_18251# a_6482_18732# a_7152_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X255 a_57689_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X256 VSS a_45231_1566# a_45233_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X257 a_3785_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X258 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X259 a_25013_18953# a_24138_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X260 a_44906_18251# a_44236_18732# a_44506_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X261 a_45217_6676# a_44627_6509# a_45121_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X262 a_43329_6676# a_42965_6419# a_43233_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X263 a_52438_13071# a_51944_12988# a_51989_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X264 a_5493_1566# a_6763_739# a_6954_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X265 a_52550_19307# a_51782_18732# a_50564_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X266 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X267 a_32565_18953# a_31690_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X268 a_3362_13071# a_4982_13134# a_4796_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X269 a_3094_13134# a_2868_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X270 a_21672_6503# a_21502_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X271 a_9678_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_4982_13134# a_4756_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X273 VDD a_44624_13134# a_44438_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X274 a_3178_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X275 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X276 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X278 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_31538_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X279 VSS a_50393_1000# a_50366_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X280 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X281 VDD a_53556_928# a_53506_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X282 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X283 VSS a_51834_18706# a_51782_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X284 a_35681_6676# a_37075_6509# a_37115_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X285 a_48478_1811# a_48505_1000# a_48490_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X286 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X287 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X288 VSS a_35066_18747# a_35039_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X289 VSS a_36954_18747# a_36927_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X290 a_28227_5620# a_27635_6509# a_26241_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X291 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_21034_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X292 a_28241_510# a_27525_739# a_26255_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X293 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X294 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_56539_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X295 VDD a_3362_13071# a_4287_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X296 a_19578_928# a_18703_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X297 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X298 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X299 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X300 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X301 a_30129_510# a_29361_765# a_28143_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X302 a_33163_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X303 a_12802_13071# a_12308_12988# a_12353_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X304 a_48676_18251# a_49946_18706# a_50137_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X305 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X306 a_52550_19307# a_51834_18706# a_50564_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X307 VSS a_58102_13071# a_59027_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X308 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X309 VDD RESET a_27668_9428# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X310 a_39685_14292# a_39326_14127# a_39324_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X311 a_12898_13071# a_12308_12988# a_12802_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X312 a_20083_6509# C[42] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X313 VDD a_17856_18706# a_18074_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X314 a_40715_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X315 a_30127_1566# a_29361_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 VSS a_57727_739# a_57675_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X317 VSS C[5] a_49946_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X318 a_44122_928# a_43247_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X319 a_29802_18251# a_29184_18706# a_29402_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X320 a_20591_1566# a_21861_739# a_22052_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X321 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X322 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X323 a_35777_6676# a_35187_6509# a_35681_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X324 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_7234_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X325 a_20458_18251# a_19692_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X326 a_58214_19307# a_58212_18251# a_58525_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X327 VDD a_25408_18706# a_25626_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X328 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X329 a_27107_12994# a_26937_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X330 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X331 a_28995_12994# a_28825_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X332 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X333 VDD a_46399_739# a_46347_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X334 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18011_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X335 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X336 VSS a_59833_1000# a_59806_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X337 VDD a_36736_18706# a_36954_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X338 VDD a_38624_18706# a_38842_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X339 VSS a_22346_18251# a_22348_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X340 a_20446_14127# a_20080_13134# a_18460_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X341 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_25563_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X342 a_18787_5620# a_18195_6509# a_16801_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X343 VSS a_49001_1566# a_49003_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X344 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X345 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X346 a_29802_18251# a_29132_18732# a_29402_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X347 a_58331_6676# a_57837_6509# a_57882_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X348 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X349 a_47099_6676# a_46735_6419# a_47003_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X350 a_7000_5455# a_6913_5687# a_6918_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 VDD a_44288_18706# a_44506_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X352 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X353 VDD a_17461_18953# a_17411_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X354 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X355 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_20128_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X356 VSS a_11803_18953# a_11753_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X357 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X358 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X359 a_7138_13071# a_6870_13134# a_6689_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X360 a_45219_5620# a_44627_6509# a_43233_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X361 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_39008_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X362 a_42820_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X363 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_36891_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X364 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_38779_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X365 a_45135_1566# a_46399_739# a_46590_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X366 a_14196_12988# C[103] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X367 VDD a_12032_928# a_11982_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X368 a_42211_12994# a_42041_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X369 a_29523_6509# C[47] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X370 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_15015_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X371 a_20687_1566# a_19921_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X372 a_41457_510# a_41455_1566# a_41768_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X373 a_32017_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X374 a_16815_1566# a_16145_765# a_16415_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X375 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X376 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_34021_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X377 VDD a_29520_13134# a_29334_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X378 a_39567_1566# a_38801_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X379 VSS a_2363_18953# a_2313_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X380 a_2949_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X381 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35909_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X382 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_44443_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X383 VSS a_19578_928# a_19528_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X384 a_1813_1566# a_1047_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X386 a_50412_5455# a_50325_5687# a_50330_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X387 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X388 VSS a_55444_928# a_55394_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X389 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X390 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X391 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X392 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X393 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X394 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X395 a_54667_510# a_53951_739# a_52681_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X396 VDD a_36341_18953# a_36291_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X397 a_5264_18251# a_6482_18732# a_6725_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X399 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X400 a_18059_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X401 a_19947_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X402 a_37667_5620# a_37075_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X403 a_7479_510# a_6711_765# a_5493_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X404 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X405 a_14422_13134# a_14196_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X406 a_25747_6509# C[45] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X407 a_43331_5620# a_42965_6419# a_41345_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X408 a_56030_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X409 VDD a_43893_18953# a_43843_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X410 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X411 a_9122_13071# a_8758_13134# a_9026_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X412 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X413 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X414 a_1799_6676# a_1435_6419# a_1703_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X415 a_40851_6509# C[53] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X416 a_11157_1566# a_10539_739# a_10757_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X417 a_48891_6676# a_48397_6509# a_48442_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X418 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X419 a_26901_18953# a_26026_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X420 VSS a_50164_18747# a_50137_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X421 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X422 a_56175_6419# a_55949_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 VDD C[81] a_27525_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X424 a_30031_1566# a_31249_765# a_31492_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X425 a_35779_5620# a_35187_6509# a_33793_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X426 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X427 a_47231_14292# a_46872_14127# a_46870_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X428 a_20444_13071# a_19854_12988# a_20348_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X429 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X430 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X431 VSS a_3362_13071# a_4287_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X432 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_8888_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X433 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X434 a_8256_928# a_7381_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X435 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X436 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X437 a_54783_14292# a_54424_14127# a_54422_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X438 a_9026_13071# a_8532_12988# a_8577_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X440 VSS C[2] a_55610_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X441 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X442 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X443 VSS a_14086_18706# a_14034_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X444 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_25792_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X445 a_16815_1566# a_18033_765# a_18276_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X446 a_3474_19307# a_3472_18251# a_3785_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X447 a_22577_510# a_21809_765# a_20591_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X448 a_46884_18251# a_46170_18706# a_46788_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X449 a_52681_1566# a_53899_765# a_54142_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X450 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_52300_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X451 a_3458_13071# a_3460_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X452 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X453 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X454 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X455 VDD a_48058_18706# a_48006_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X456 a_56443_6676# a_57837_6509# a_57877_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X457 VDD a_49946_18706# a_49894_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X458 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X459 a_9353_5620# a_8761_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X460 a_33891_5620# a_33525_6419# a_31905_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X461 a_46590_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X462 a_12816_18251# a_14086_18706# a_14277_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X463 a_27107_12994# a_26937_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X464 a_28995_12994# a_28825_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X465 VDD a_43233_6676# a_44158_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X466 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_18785_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X467 a_42739_6509# C[54] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X468 a_60642_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X469 a_5493_1566# a_4823_765# a_5093_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X470 VDD a_51834_18706# a_52052_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X471 a_21823_18006# a_21850_18747# a_21835_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X472 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X473 VSS C[24] a_14086_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X474 a_46735_6419# a_46509_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X475 a_60315_6676# a_60317_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X476 a_27451_14292# a_27446_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X477 a_52765_5620# a_52173_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X478 a_980_12988# C[96] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X479 a_23630_12988# C[108] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X480 OUT a_60915_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X481 a_7465_5620# a_6873_6509# a_5479_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X482 VDD C[6] a_48058_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X483 VSS C[80] a_29413_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X484 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X485 a_33151_18006# a_33178_18747# a_33163_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X486 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X487 a_6771_14292# a_6684_14194# a_6689_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X488 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_51989_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X489 a_56539_6676# a_55949_6509# a_56443_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X490 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X491 a_33115_14292# a_33110_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X492 VDD C[72] a_44517_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X493 a_56228_18251# a_55558_18732# a_55828_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X494 a_59220_928# a_58345_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X495 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_39685_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X496 VSS a_8651_739# a_8599_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X497 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X498 a_40703_18006# a_40730_18747# a_40715_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X499 a_14506_1811# a_14533_1000# a_14518_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X500 a_58331_6676# a_59725_6509# a_59765_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X501 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X502 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X503 VDD a_53951_739# a_53899_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X504 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X505 VDD a_14651_6419# a_14465_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X506 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X507 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X508 a_47003_6676# a_48397_6509# a_48437_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X509 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X510 VSS C[87] a_16197_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X511 VDD a_51439_18953# a_51389_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X512 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X513 a_33660_13071# a_33296_13134# a_33564_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X514 VSS C[68] a_52063_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X515 a_9367_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X516 a_51439_18953# a_50564_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X517 a_46280_12988# C[120] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X518 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X519 a_29520_13134# a_29294_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X520 VDD a_33793_6676# a_34718_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X521 a_16400_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X522 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X523 a_29375_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X524 VSS a_48276_18747# a_48249_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X525 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X526 a_54651_6676# a_54287_6419# a_54555_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X527 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X528 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X529 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X530 a_30129_510# a_29413_739# a_28143_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X531 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X532 a_36927_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X533 VSS a_55828_18747# a_55801_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X534 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X535 a_52779_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X536 a_58200_14127# a_57834_13134# a_56214_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X537 a_56324_18251# a_55558_18732# a_56228_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X538 a_14552_5455# a_14465_5687# a_14470_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X539 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X540 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X541 a_31676_13071# a_31182_12988# a_31227_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X542 a_24220_13071# a_23630_12988# a_24124_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X543 a_52037_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X544 a_11012_14127# a_10420_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X545 VSS a_39071_1000# a_39044_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X546 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X547 a_46774_13071# a_48394_13134# a_48208_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X548 a_11803_18953# a_10928_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X549 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X550 VSS a_23520_18706# a_23468_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X551 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X552 a_58559_14292# a_58200_14127# a_58198_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X553 a_31772_13071# a_31182_12988# a_31676_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X554 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X555 a_58429_5620# a_57837_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X556 VSS a_15029_1566# a_15031_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X557 a_48676_18251# a_48058_18706# a_48276_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X558 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_5936_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X559 VSS a_6368_928# a_6318_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X560 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X561 VDD a_46774_13071# a_47699_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X562 a_15015_6676# a_14425_6509# a_14919_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X563 a_13127_6676# a_12763_6419# a_13031_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X564 a_18801_510# a_18085_739# a_16815_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X565 a_20362_18251# a_21632_18706# a_21823_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X566 a_54326_13071# a_55720_12988# a_55760_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X567 VSS a_43233_6676# a_44158_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X568 a_24236_19307# a_23520_18706# a_22250_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X569 a_47869_12994# a_47699_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X570 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X571 a_12401_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X572 a_56541_5620# a_55949_6509# a_54555_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X573 VSS a_11253_1566# a_11255_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_31788_19307# a_31072_18706# a_29802_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X575 VSS a_42400_18706# a_42348_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X576 a_4985_6509# C[34] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X577 a_58345_1566# a_57675_765# a_57945_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X578 VDD a_23354_928# a_23304_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X579 a_28143_1566# a_29361_765# a_29604_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X580 a_47113_1566# a_46399_739# a_47017_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X581 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X582 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X583 a_18276_1811# a_18303_1000# a_18288_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X584 a_22348_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X585 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X586 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_48758_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X587 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_26337_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X588 a_33392_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X589 VSS C[16] a_29184_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X590 VDD a_18421_6419# a_18235_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X591 a_34682_928# a_33807_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X592 a_39242_18251# a_40512_18706# a_40703_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X593 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X594 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X595 a_20362_18251# a_21580_18732# a_21823_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X596 a_43116_19307# a_42400_18706# a_41130_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X597 a_33344_5455# a_33339_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X598 a_18556_13071# a_18192_13134# a_18460_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X600 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X601 a_56900_5455# a_56541_5620# a_56539_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X602 a_34958_12988# C[114] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X603 OUT a_60915_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X604 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X605 a_28129_6676# a_27635_6509# a_27680_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X606 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X607 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X608 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X609 a_11024_18251# a_10258_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X610 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_54783_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X611 a_54653_5620# a_54287_6419# a_52667_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X612 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X613 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X614 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X615 a_22479_1566# a_21861_739# a_22079_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X616 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X617 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X618 VSS a_33793_6676# a_34718_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X619 VDD C[69] a_50175_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X620 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_60447_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X621 a_3605_1566# a_4823_765# a_5066_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X622 a_39242_18251# a_40460_18732# a_40703_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X623 VSS a_6981_1000# a_6954_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X624 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X625 VDD a_55215_18953# a_55165_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X626 a_37436_13071# a_37072_13134# a_37340_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X627 VDD a_16197_739# a_16145_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X628 a_3472_18251# a_2706_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X629 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X630 a_1813_1566# a_1099_739# a_1717_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X631 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X632 a_20309_6419# a_20083_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X633 a_16684_19307# a_15916_18732# a_14704_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X634 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X635 a_33296_13134# a_33070_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X636 a_48905_1566# a_48235_765# a_48505_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X637 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X638 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X639 a_44988_13071# a_44624_13134# a_44892_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X640 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X641 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X642 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X643 VSS a_18799_1566# a_18801_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X644 a_49085_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X645 a_40848_13134# a_40622_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X646 a_57608_12988# C[126] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X647 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X648 a_45775_18953# a_44906_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X649 a_3460_14127# a_3094_13134# a_1474_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X650 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X651 VSS a_15968_18706# a_15916_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X652 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X653 a_1584_18251# a_818_18732# a_1488_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X654 a_52025_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X655 VSS a_27668_9428# sky130_fd_sc_hd__buf_2_0/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X656 VDD a_40346_928# a_40296_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X657 a_13129_5620# a_12763_6419# a_11143_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X658 a_35268_1811# a_35295_1000# a_35280_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X659 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X660 a_15017_5620# a_14425_6509# a_13031_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X661 a_5030_5455# a_5025_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X662 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X663 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_43329_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X664 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X665 a_35564_19307# a_34796_18732# a_33578_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X666 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_6771_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X667 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X668 a_20210_5455# a_20123_5687# a_20128_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X669 a_39090_5455# a_39003_5687# a_39008_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X670 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_58788_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X671 a_41228_19307# a_40460_18732# a_39242_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X672 a_58102_13071# a_59722_13134# a_59536_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X673 a_7236_14127# a_6644_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X674 a_57834_13134# a_57608_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X675 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X676 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X677 VDD a_54555_6676# a_55480_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X678 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X679 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X680 VSS a_34848_18706# a_34796_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X681 a_794_737# a_980_12988# a_1020_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X682 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X683 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X684 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X685 a_1254_5455# a_1249_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X686 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X687 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X688 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X689 VSS C[94] a_2987_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X690 a_21869_14292# a_21782_14194# a_21787_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X691 VSS a_46774_13071# a_47699_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X692 VSS a_46004_928# a_45954_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X693 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X694 a_60331_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X695 a_47869_12994# a_47699_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X696 VDD a_33189_739# a_33137_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X697 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X698 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X699 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X700 a_34021_14292# a_33662_14127# a_33660_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 VSS C[14] a_32960_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X702 a_8625_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X703 a_13031_6676# a_14425_6509# a_14465_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X704 a_25828_1811# a_25855_1000# a_25840_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X705 VSS a_35791_1566# a_35793_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X706 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1570_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X707 a_40749_14292# a_40662_14194# a_40667_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X708 VDD a_7099_6419# a_6913_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X709 VDD a_27296_18706# a_27244_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X710 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X711 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X712 VSS a_23749_739# a_23697_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X713 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X714 a_53877_14292# a_53872_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X715 a_10144_928# a_9269_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X716 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X717 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X718 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X719 VDD a_27525_739# a_27743_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X720 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X721 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X722 a_14800_18251# a_14034_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X723 a_16586_18251# a_15916_18732# a_16186_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X724 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X726 a_37569_6676# a_37301_6419# a_37120_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X727 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_22098_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X728 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X729 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X730 a_10914_13071# a_10646_13134# a_10465_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X731 a_26241_6676# a_27635_6509# a_27675_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X732 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X733 a_5591_510# a_4875_739# a_3605_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X734 a_54665_1566# a_53951_739# a_54569_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X735 a_7248_18251# a_6482_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X736 VSS a_11024_18251# a_11026_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X737 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X738 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_47099_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X739 a_54154_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X740 a_40323_12994# a_40153_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X741 a_52534_13071# a_52170_13134# a_52438_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X742 VDD C[17] a_27296_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X743 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X744 VDD a_16304_13134# a_16118_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X745 a_25874_5455# a_25787_5687# a_25792_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X746 VSS a_46399_739# a_46347_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X747 a_12389_18006# a_12416_18747# a_12401_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X748 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X749 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X750 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X751 a_1474_13071# a_1206_13134# a_1025_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X752 a_37681_510# a_36913_765# a_35695_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X753 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X754 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_31227_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X755 a_38664_6503# a_38494_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X756 a_48249_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X757 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X758 a_5348_14127# a_4756_12988# a_3362_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X759 a_30440_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X760 a_54106_5455# a_54101_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X761 VSS a_49551_18953# a_49501_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X762 a_2868_12988# C[97] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X763 a_12537_6509# C[38] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X764 a_35466_18251# a_34796_18732# a_35066_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X765 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X766 a_16533_6419# a_16307_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 a_49780_928# a_48905_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X768 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X769 VDD a_23856_13134# a_23670_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X770 a_7236_14127# a_6870_13134# a_5250_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X771 a_30113_6676# a_30115_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X772 VDD a_2592_928# a_2542_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X773 a_4837_18006# a_4864_18747# a_4849_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X774 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X775 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X776 a_1897_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X777 a_35681_6676# a_35187_6509# a_35232_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X778 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_5575_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X779 a_23125_18953# a_22250_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X780 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X781 a_26337_6676# a_25747_6509# a_26241_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X782 VDD a_35184_13134# a_34998_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X783 VSS a_54555_6676# a_55480_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X784 VDD C[88] a_14315_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X785 a_13045_1566# a_14315_739# a_14506_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X786 a_42820_1811# a_42847_1000# a_42832_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X787 a_2126_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X789 a_50662_19307# a_49894_18732# a_48676_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X790 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X791 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X792 a_37679_1566# a_36913_765# a_37583_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X793 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X794 a_30677_18953# a_29802_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X795 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X796 VSS a_21466_928# a_21416_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X797 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X798 VSS a_27514_18747# a_27487_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X799 a_1206_13134# a_980_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X800 VSS C[72] a_44517_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X801 a_18917_14292# a_18558_14127# a_18556_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X802 VDD a_42736_13134# a_42550_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X803 a_20689_510# a_19973_739# a_18703_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X804 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X805 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X806 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X807 a_9255_6676# a_8987_6419# a_8806_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X808 a_16801_6676# a_18195_6509# a_18235_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X809 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X810 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X811 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X812 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_12582_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X813 a_1717_1566# a_1099_739# a_1317_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X814 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X815 a_10914_13071# a_10420_12988# a_10465_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 a_35695_1566# a_36965_739# a_37156_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X817 a_31275_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X818 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X819 a_39880_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X820 a_21000_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X821 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X822 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X823 a_50662_19307# a_49946_18706# a_48676_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X824 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_27762_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X825 a_33380_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X826 a_37797_14292# a_37438_14127# a_37436_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X827 a_11010_13071# a_10420_12988# a_10914_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X828 a_42866_5455# a_42779_5687# a_42784_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X829 a_48774_19307# a_48772_18251# a_49085_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X830 a_27900_13071# a_29294_12988# a_29334_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X831 a_39553_6676# a_39555_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X832 VDD a_15968_18706# a_16186_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X833 a_48758_13071# a_48760_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X834 a_1799_6676# a_1801_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X835 a_27914_18251# a_27296_18706# a_27514_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X836 a_19555_12994# a_19385_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X837 a_29898_18251# a_29184_18706# a_29802_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X838 a_16897_6676# a_16307_6509# a_16801_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X839 a_33525_6419# a_33299_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X840 a_35681_6676# a_37301_6419# a_37115_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X841 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X842 VDD a_23520_18706# a_23738_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X843 a_56326_19307# a_56324_18251# a_56637_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X844 a_25219_12994# a_25049_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X845 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X846 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X847 VSS a_43343_1566# a_43345_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X848 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X849 a_7234_13071# a_6644_12988# a_7138_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X850 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X851 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X852 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_16123_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X853 a_9365_1566# a_8599_765# a_9269_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X854 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X855 a_39242_18251# a_38624_18706# a_38842_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X856 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X857 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X858 a_3703_510# a_3701_1566# a_4014_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X859 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X860 a_43329_6676# a_42739_6509# a_43233_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X861 a_28227_5620# a_27635_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X862 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X863 a_18703_1566# a_19921_765# a_20164_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X864 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X865 a_29898_18251# a_29132_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X866 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X867 VDD a_34848_18706# a_35066_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X868 VSS a_20458_18251# a_20460_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X869 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X870 a_38435_12994# a_38265_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X871 a_38664_6503# a_38494_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X872 VDD a_55610_18706# a_55558_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X873 VDD a_40741_739# a_40689_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X874 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X875 VDD a_42400_18706# a_42618_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X876 a_44099_12994# a_43929_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X877 VDD a_15573_18953# a_15523_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X878 a_45987_12994# a_45817_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X879 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X880 a_33793_6676# a_35187_6509# a_35227_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X881 a_46590_1811# a_46617_1000# a_46602_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X882 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X883 a_26339_5620# a_25747_6509# a_24353_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X884 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X885 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X886 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_26469_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X887 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35003_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X888 a_5250_13071# a_4982_13134# a_4801_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X889 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_38026_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X890 a_12308_12988# C[102] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X891 a_59623_14292# a_59536_14194# a_59541_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X892 a_40323_12994# a_40153_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X893 a_39242_18251# a_38572_18732# a_38842_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X894 a_3097_6509# C[33] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X895 a_22577_510# a_22575_1566# a_22888_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X896 a_50564_18251# a_49894_18732# a_50164_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X897 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_32133_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X898 a_41441_6676# a_41077_6419# a_41345_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X899 a_8613_18006# a_8640_18747# a_8625_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 a_5362_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X901 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X902 a_4048_5455# a_3689_5620# a_3687_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X903 a_13143_510# a_12375_765# a_11157_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X904 VSS a_19962_18747# a_19935_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X905 a_7367_6676# a_8987_6419# a_8801_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X906 a_43247_1566# a_44465_765# a_44708_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X907 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X908 a_5211_6419# a_4985_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X909 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X910 a_37075_6509# C[51] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X911 VDD a_34453_18953# a_34403_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X912 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X913 a_58331_6676# a_58063_6419# a_57882_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X914 a_25242_928# a_24367_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X915 a_3376_18251# a_4594_18732# a_4837_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X916 a_54438_19307# a_53670_18732# a_52452_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X917 VDD a_50282_13134# a_50096_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X918 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X919 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X920 a_29294_12988# C[111] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X921 a_33889_6676# a_33299_6509# a_33793_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X922 a_12534_13134# a_12308_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X923 a_17461_18953# a_16586_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X924 a_24451_5620# a_24085_6419# a_22465_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X925 a_23711_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X926 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X927 a_46636_5455# a_46549_5687# a_46554_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X928 a_21971_6509# C[43] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X929 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X930 a_28323_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X931 VSS a_38842_18747# a_38815_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X932 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X933 a_45219_5620# a_44627_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X934 VSS a_57945_1000# a_57918_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X935 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X936 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X937 a_16899_5620# a_16307_6509# a_14919_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X938 VSS a_47113_1566# a_47115_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X939 a_50875_6676# a_50877_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X940 a_36939_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X941 a_14802_19307# a_14034_18732# a_12816_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X942 a_56443_6676# a_55949_6509# a_55994_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X943 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X944 a_36341_18953# a_35466_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X945 VDD a_50175_739# a_50393_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X946 a_42591_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X947 a_32001_6676# a_31637_6419# a_31905_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X948 a_43331_5620# a_42739_6509# a_41345_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X949 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_37120_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X950 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X951 a_52895_14292# a_52536_14127# a_52534_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X952 a_45135_1566# a_44465_765# a_44735_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X953 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X954 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X955 a_42005_18953# a_41130_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X956 VSS C[3] a_53722_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X957 VDD a_10144_928# a_10094_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X958 VSS a_12198_18706# a_12146_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X959 a_43893_18953# a_43018_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X960 a_11157_1566# a_12427_739# a_12618_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X961 a_30129_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X962 a_1586_19307# a_1584_18251# a_1897_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X963 a_48891_6676# a_48623_6419# a_48442_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X964 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_13127_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X965 a_37679_1566# a_36913_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X966 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X967 a_19555_12994# a_19385_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X968 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X969 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X970 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X971 a_61314_6503# a_61144_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X972 a_10928_18251# a_12198_18706# a_12389_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X973 a_5575_6676# a_4985_6509# a_5479_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X974 a_54340_18251# a_53722_18706# a_53940_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X975 a_25219_12994# a_25049_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X976 a_14802_19307# a_14086_18706# a_12816_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X977 a_43690_5455# a_43331_5620# a_43329_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X978 a_56324_18251# a_55610_18706# a_56228_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X979 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X980 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X981 VDD a_24353_6676# a_25278_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X982 a_49986_6503# a_49816_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X983 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X984 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X985 VDD a_49946_18706# a_50164_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X986 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18917_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X987 a_23859_6509# C[44] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X988 a_53533_12994# a_53363_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X989 a_54142_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X990 VSS C[25] a_12198_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X991 a_12435_14292# a_12348_14194# a_12353_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X992 a_41443_5620# a_41077_6419# a_39457_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X993 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X994 a_7152_18251# a_8422_18706# a_8613_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X995 a_25563_14292# a_25558_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X996 a_21742_12988# C[107] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X997 a_38435_12994# a_38265_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X998 VDD C[7] a_46170_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X999 a_47003_6676# a_46509_6509# a_46554_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1000 a_60329_1566# a_59563_765# a_60219_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1001 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1002 a_31263_18006# a_31290_18747# a_31275_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1003 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1004 a_4883_14292# a_4796_14194# a_4801_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1005 a_54287_6419# a_54061_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1006 a_56443_6676# a_58063_6419# a_57877_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1007 VDD a_59615_739# a_59833_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1008 a_31227_14292# a_31222_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1009 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_50101_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1010 a_44099_12994# a_43929_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1011 VDD C[82] a_25637_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1012 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1013 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1014 a_45987_12994# a_45817_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1015 a_33891_5620# a_33299_6509# a_31905_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1016 a_54340_18251# a_53670_18732# a_53940_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1017 a_35695_1566# a_35025_765# a_35295_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1018 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1019 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1020 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_37797_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1021 a_9138_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1022 a_6368_928# a_5493_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1023 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1024 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1025 a_1815_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1026 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1027 a_9365_1566# a_8599_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1028 a_20080_13134# a_19854_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1029 a_45233_510# a_44517_739# a_43247_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1030 a_7152_18251# a_8370_18732# a_8613_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1031 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1032 a_31772_13071# a_31408_13134# a_31676_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1034 a_44627_6509# C[55] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1035 a_31919_1566# a_31249_765# a_31519_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1036 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1037 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1038 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_50412_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1039 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1040 VSS a_46388_18747# a_46361_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1041 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1042 a_54555_6676# a_55949_6509# a_55989_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1043 VSS a_28789_18953# a_28739_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1044 a_27487_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1045 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1046 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1047 a_14704_18251# a_14034_18732# a_14304_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1048 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1049 VSS a_38853_739# a_38801_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1050 a_7465_5620# a_6873_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1051 a_32003_5620# a_31637_6419# a_30017_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1052 a_28789_18953# a_27914_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1053 a_48772_18251# a_48006_18732# a_48676_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1054 a_8758_13134# a_8532_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1055 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1056 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_45578_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1057 VSS a_52052_18747# a_52025_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1058 VSS a_53940_18747# a_53913_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1059 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1060 a_22236_13071# a_21742_12988# a_21787_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1061 VDD a_41345_6676# a_42270_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1062 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_16897_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1063 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1064 a_56312_14127# a_55946_13134# a_54326_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1065 a_47003_6676# a_48623_6419# a_48437_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1066 a_704_928# a_794_737# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1067 a_50149_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1068 a_22332_13071# a_21742_12988# a_22236_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1069 VDD a_14422_13134# a_14236_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1070 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1071 a_44892_13071# a_46506_13134# a_46320_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1072 a_50877_5620# a_50285_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1073 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1074 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_59623_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1075 a_5577_5620# a_4985_6509# a_3591_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1076 VSS a_21632_18706# a_21580_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1077 a_59951_6419# a_59725_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1078 a_47460_5455# a_47101_5620# a_47099_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1079 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1080 a_28241_510# a_27473_765# a_26255_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1081 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1082 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1083 a_46774_13071# a_48168_12988# a_48208_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1084 a_54651_6676# a_54061_6509# a_54555_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1085 a_61314_6503# a_61144_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1086 a_1572_14127# a_980_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1087 VDD C[73] a_42629_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1088 a_46788_18251# a_46170_18706# a_46388_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1089 VSS a_13920_928# a_13870_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1090 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1091 a_48772_18251# a_48058_18706# a_48676_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1092 a_52438_13071# a_53832_12988# a_53872_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1093 a_18474_18251# a_19744_18706# a_19935_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1094 VSS a_24353_6676# a_25278_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1095 a_49986_6503# a_49816_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1096 a_12618_1811# a_12645_1000# a_12630_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1097 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1098 a_22348_19307# a_21632_18706# a_20362_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1099 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1100 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1101 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1102 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_59852_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1103 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1104 a_45121_6676# a_46509_6509# a_46549_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1105 a_10513_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1106 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1107 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1108 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1109 VSS a_40512_18706# a_40460_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1110 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_37665_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1111 a_7479_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1112 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1113 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1114 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1115 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1116 a_20460_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1117 a_28012_19307# a_28010_18251# a_28323_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1118 VDD a_31905_6676# a_32830_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1119 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_46870_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1120 a_52763_6676# a_52399_6419# a_52667_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1121 VSS a_36570_928# a_36520_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1122 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_57882_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1123 a_41228_19307# a_40512_18706# a_39242_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1124 a_53533_12994# a_53363_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1125 a_16668_13071# a_16304_13134# a_16572_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1126 a_41455_1566# a_40741_739# a_41359_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1127 a_8659_14292# a_8572_14194# a_8577_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1128 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1129 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1130 a_48397_6509# C[57] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1131 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_33889_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1132 a_58441_1566# a_57675_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1133 a_12664_5455# a_12577_5687# a_12582_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1134 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_51007_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1135 a_26255_1566# a_27525_739# a_27716_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1136 a_59220_928# a_58345_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1137 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1138 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_52895_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1139 VDD a_14086_18706# a_14304_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1141 a_704_928# a_794_737# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1142 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1143 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1144 a_56541_5620# a_55949_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1145 VSS a_13141_1566# a_13143_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1146 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1147 VDD a_53327_18953# a_53277_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1148 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1149 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1150 a_1584_18251# a_818_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1151 a_35548_13071# a_35184_13134# a_35452_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1152 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1153 a_31408_13134# a_31182_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1154 a_48168_12988# C[121] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1155 a_13127_6676# a_12537_6509# a_13031_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1156 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_14241_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1157 VSS a_41345_6676# a_42270_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1158 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 a_58200_14127# a_57608_12988# a_56214_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1160 a_47197_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1161 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1162 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_48442_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1163 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1164 a_1572_14127# a_1206_13134# a_794_737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1165 a_54653_5620# a_54061_6509# a_52667_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1166 a_56457_1566# a_55787_765# a_56057_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1167 VDD a_21466_928# a_21416_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1168 VSS a_37183_1000# a_37156_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1169 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1170 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1171 a_33807_1566# a_35025_765# a_35268_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1172 a_16388_1811# a_16415_1000# a_16400_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1173 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1174 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_24449_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1175 a_31504_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1176 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1177 VDD a_13691_18953# a_13641_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1178 VSS a_14315_739# a_14263_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1179 a_15802_928# a_14933_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1180 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1181 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1182 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_2995_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1183 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_4883_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1184 a_48394_13134# a_48168_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1185 a_33676_19307# a_32908_18732# a_31690_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1186 a_55215_18953# a_54340_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1187 a_51668_928# a_50793_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1188 VSS a_25408_18706# a_25356_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1189 a_16014_6503# a_15844_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1190 a_49780_928# a_48905_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1191 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1192 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1193 a_5348_14127# a_4756_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1194 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1195 a_55946_13134# a_55720_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1196 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1197 a_55012_5455# a_54653_5620# a_54651_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1198 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1199 VDD a_48662_13071# a_49587_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1200 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1201 a_28129_6676# a_27861_6419# a_27680_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1202 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1203 a_52765_5620# a_52399_6419# a_50779_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1204 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1205 VSS C[90] a_10539_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1206 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1207 VSS a_31905_6676# a_32830_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1208 a_14289_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1209 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1210 a_24581_14292# a_24222_14127# a_24220_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1211 a_16434_5455# a_16347_5687# a_16352_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1212 a_15029_1566# a_14263_765# a_14933_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1213 VSS C[18] a_25408_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1214 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1215 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1216 a_15017_5620# a_14425_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1217 VSS C[15] a_31072_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1218 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1219 a_52681_1566# a_53951_739# a_54142_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1220 VSS a_27743_1000# a_27716_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1221 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1222 VDD a_19744_18706# a_19692_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1223 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 a_20673_6676# a_20675_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1225 VSS a_16911_1566# a_16913_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1226 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1227 a_3190_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1228 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1229 sky130_fd_sc_hd__buf_2_0/X a_27668_9428# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1230 a_26241_6676# a_25747_6509# a_25792_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1231 VSS C[78] a_33189_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1232 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1233 VSS a_475_18953# a_425_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1234 a_43461_14292# a_43102_14127# a_43100_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1235 a_33380_1811# a_33407_1000# a_33392_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1236 a_13129_5620# a_12537_6509# a_11143_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1237 a_3142_5455# a_3137_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1238 VSS a_12032_928# a_11982_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1239 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1240 a_56310_13071# a_56312_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1241 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_41441_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1242 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1243 a_11255_510# a_10539_739# a_9269_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1244 a_28239_1566# a_27473_765# a_28143_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1245 a_18689_6676# a_18421_6419# a_18240_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1246 VDD C[22] a_17856_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1247 VDD a_38624_18706# a_38572_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1248 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1249 a_32771_12994# a_32601_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1250 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1251 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_56900_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 a_37202_5455# a_37115_5687# a_37120_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 a_5360_18251# a_4594_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1254 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_23675_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1255 a_31112_6503# a_30942_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1256 VDD a_52667_6676# a_53592_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1257 a_50646_13071# a_50282_13134# a_50550_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1258 VDD a_44288_18706# a_44236_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1259 a_26026_18251# a_25356_18732# a_25626_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1260 a_27914_18251# a_27244_18732# a_27514_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1261 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1262 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1263 a_45121_6676# a_44853_6419# a_44672_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1264 a_10501_18006# a_10528_18747# a_10513_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1265 a_19784_6503# a_19614_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1266 VSS a_40741_739# a_40689_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1267 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1268 a_58102_13071# a_57834_13134# a_57653_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1269 a_59990_13071# a_59722_13134# a_59541_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1270 VSS a_47663_18953# a_47613_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1271 a_3460_14127# a_2868_12988# a_1474_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1272 a_33578_18251# a_32908_18732# a_33178_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1273 VDD a_20080_13134# a_19894_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1274 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_15147_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 VDD a_21968_13134# a_21782_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1276 a_11241_5620# a_10875_6419# a_9255_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1277 VSS a_7248_18251# a_7250_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1278 a_5348_14127# a_4982_13134# a_3362_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1279 VDD C[11] a_38624_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1280 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1281 a_16014_6503# a_15844_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1282 VDD a_6763_739# a_6981_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1283 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1284 a_58214_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1285 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 a_21237_18953# a_20362_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1287 a_16801_6676# a_16307_6509# a_16352_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1288 a_35793_510# a_35077_739# a_33807_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1289 a_30127_1566# a_29361_765# a_30031_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1290 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1291 a_24085_6419# a_23859_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1292 a_26241_6676# a_27861_6419# a_27675_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1293 VSS a_44735_1000# a_44708_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1294 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1295 VDD C[8] a_44288_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1296 VSS a_18074_18747# a_18047_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1297 a_23940_1811# a_23967_1000# a_23952_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1298 a_11010_13071# a_10646_13134# a_10914_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1299 VDD a_33296_13134# a_33110_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1300 VSS a_33903_1566# a_33905_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1301 a_5066_1811# a_5093_1000# a_5078_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1302 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1303 a_58116_18251# a_59334_18732# a_59577_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1304 a_18799_1566# a_18033_765# a_18703_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1305 a_43233_6676# a_42739_6509# a_42784_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1306 VSS a_25626_18747# a_25599_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1307 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1308 VDD a_5211_6419# a_5025_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1309 a_9269_1566# a_10487_765# a_10730_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1310 VDD a_40848_13134# a_40662_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1311 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1312 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1313 a_17029_14292# a_16670_14127# a_16668_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1314 a_26122_18251# a_25356_18732# a_26026_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1315 a_27861_6419# a_27635_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1316 a_8854_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1317 a_28010_18251# a_27244_18732# a_27914_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1318 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1319 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1320 VDD a_25637_739# a_25855_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1321 a_40117_18953# a_39242_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1322 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1323 a_14425_6509# C[39] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1324 VDD a_31301_739# a_31249_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 VSS a_48662_13071# a_49587_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1326 a_35681_6676# a_35413_6419# a_35232_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1327 a_8806_5455# a_8801_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1328 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_20210_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1329 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_39090_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1330 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1331 a_28357_14292# a_27998_14127# a_27996_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1332 a_24353_6676# a_25747_6509# a_25787_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1333 a_42510_12988# C[118] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1334 a_52777_1566# a_52063_739# a_52681_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1335 a_18474_18251# a_17856_18706# a_18074_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1336 a_52266_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1337 VSS a_44506_18747# a_44479_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1338 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1339 a_23986_5455# a_23899_5687# a_23904_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1340 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1341 a_26012_13071# a_27406_12988# a_27446_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1342 a_35909_14292# a_35550_14127# a_35548_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1343 a_18801_510# a_18033_765# a_16815_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1344 a_46886_19307# a_46884_18251# a_47197_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1345 VDD a_11143_6676# a_12068_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1346 a_36776_6503# a_36606_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1347 a_26026_18251# a_25408_18706# a_25626_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1348 a_17667_12994# a_17497_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1349 a_54667_510# a_53899_765# a_52681_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1350 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1351 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1352 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1353 a_5250_13071# a_4756_12988# a_4801_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1354 a_10649_6509# C[37] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1355 a_28010_18251# a_27296_18706# a_27914_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1356 a_16801_6676# a_18421_6419# a_18235_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1357 VSS a_29413_739# a_29361_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1358 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1359 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1360 a_37340_13071# a_38734_12988# a_38774_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1361 a_5346_13071# a_4756_12988# a_5250_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1362 a_1570_13071# a_1572_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1363 a_33793_6676# a_33299_6509# a_33344_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1364 a_28143_1566# a_29413_739# a_29604_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1365 a_2592_928# a_1717_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1366 a_37354_18251# a_36736_18706# a_36954_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1367 a_43004_13071# a_44624_13134# a_44438_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1368 a_24449_6676# a_23859_6509# a_24353_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1369 a_31112_6503# a_30942_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1370 a_41077_6419# a_40851_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1371 a_43233_6676# a_44853_6419# a_44667_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1372 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1373 a_39338_18251# a_38624_18706# a_39242_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1374 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1375 VSS a_52667_6676# a_53592_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1376 VDD C[89] a_12427_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1377 a_40932_1811# a_40959_1000# a_40944_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1378 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1379 VDD a_32960_18706# a_33178_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1380 a_44906_18251# a_44288_18706# a_44506_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1381 a_36547_12994# a_36377_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1382 VDD a_53722_18706# a_53670_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1383 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1384 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1385 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1386 a_19784_6503# a_19614_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1387 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1388 VDD a_41116_13071# a_42041_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1389 VDD a_43004_13071# a_43929_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1390 VDD a_21861_739# a_21809_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1391 VSS C[82] a_25637_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1392 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1393 VDD a_40512_18706# a_40730_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1394 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_29650_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1395 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1396 a_32771_12994# a_32601_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1397 a_7367_6676# a_7099_6419# a_6918_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1398 a_14919_6676# a_16307_6509# a_16347_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1399 VSS a_48505_1000# a_48478_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1400 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1401 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1402 VDD a_44853_6419# a_44667_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1403 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1404 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_24581_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1405 a_3362_13071# a_3094_13134# a_2913_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1406 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_19146_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1407 VDD a_42629_739# a_42847_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1408 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1409 a_16815_1566# a_18085_739# a_18276_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1410 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1411 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_30245_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1412 a_22561_6676# a_22197_6419# a_22465_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1413 a_41345_6676# a_42739_6509# a_42779_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1414 VDD a_25013_18953# a_24963_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1415 a_6725_18006# a_6752_18747# a_6737_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1416 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1417 a_8462_6503# a_8292_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1418 a_37992_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1419 a_10928_18251# a_12146_18732# a_12389_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1420 VDD a_26901_18953# a_26851_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1421 VDD C[4] a_51834_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1422 a_3474_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1423 a_31492_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1424 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_25874_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1425 a_40978_5455# a_40891_5687# a_40896_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1426 VSS C[70] a_48287_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1427 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1428 a_37665_6676# a_37667_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1429 a_8532_12988# C[100] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1430 a_18195_6509# C[41] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1431 VSS a_27130_928# a_27080_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1432 a_28239_1566# a_27473_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1433 VDD a_32565_18953# a_32515_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1434 VDD C[0] a_59386_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1435 a_14786_13071# a_14422_13134# a_14690_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1436 a_1488_18251# a_2706_18732# a_2949_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1437 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_43461_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1438 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1439 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1440 a_31637_6419# a_31411_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1441 a_33793_6676# a_35413_6419# a_35227_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1442 a_10646_13134# a_10420_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1443 a_27406_12988# C[110] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1444 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1445 a_15573_18953# a_14704_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1446 VSS a_29402_18747# a_29375_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1447 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1448 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1449 a_21823_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1450 a_34250_5455# a_33891_5620# a_33889_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1451 a_7477_1566# a_6711_765# a_7381_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1452 a_1815_510# a_1813_1566# a_2126_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1453 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1454 a_41441_6676# a_40851_6509# a_41345_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1455 a_26339_5620# a_25747_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1456 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1457 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1458 a_39326_14127# a_38960_13134# a_37340_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1459 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1460 a_33151_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1461 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 VSS a_11143_6676# a_12068_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1463 a_36776_6503# a_36606_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1464 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1465 a_12914_19307# a_12146_18732# a_10928_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1466 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1467 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1468 a_27900_13071# a_29520_13134# a_29334_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1469 a_27632_13134# a_27406_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1470 a_34453_18953# a_33578_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1471 a_39651_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1472 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1473 a_46872_14127# a_46280_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1474 a_31905_6676# a_33299_6509# a_33339_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1475 a_40703_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1476 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_18240_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1477 a_51007_14292# a_50648_14127# a_50646_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1478 a_24451_5620# a_23859_6509# a_22465_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1479 a_26255_1566# a_25585_765# a_25855_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1480 a_60100_18251# a_59334_18732# a_59990_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1481 a_45315_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1482 VSS a_41455_1566# a_41457_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1483 a_1209_6509# C[32] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1484 VDD a_27900_13071# a_28825_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1485 a_39569_510# a_39567_1566# a_39880_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1486 a_9351_6676# a_9353_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1487 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1488 a_17667_12994# a_17497_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1489 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1490 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_42866_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1491 a_48524_5455# a_48437_5687# a_48442_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1492 a_58991_18953# a_58116_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1493 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1494 a_9122_13071# a_8532_12988# a_9026_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1495 VDD a_48623_6419# a_48437_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1496 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1497 a_3323_6419# a_3097_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1498 a_5479_6676# a_7099_6419# a_6913_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1499 a_24367_1566# a_25585_765# a_25828_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1500 a_52452_18251# a_51834_18706# a_52052_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1501 a_53090_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1502 a_56443_6676# a_56175_6419# a_55994_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1503 a_35187_6509# C[50] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1504 a_45231_1566# a_44465_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1505 VSS a_8422_18706# a_8370_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1506 a_54436_18251# a_53722_18706# a_54340_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1507 a_24810_5455# a_24451_5620# a_24449_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1508 a_32001_6676# a_31411_6509# a_31905_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1509 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1510 a_52763_6676# a_52765_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1511 a_51645_12994# a_51475_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1512 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1513 a_10547_14292# a_10460_14194# a_10465_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1514 a_5575_6676# a_5577_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1515 a_22563_5620# a_22197_6419# a_20577_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1516 a_60100_18251# a_59386_18706# a_59990_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1517 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1519 a_5264_18251# a_6534_18706# a_6725_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1520 a_23675_14292# a_23670_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1521 a_36547_12994# a_36377_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1522 a_38963_6509# C[52] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1523 a_57538_6503# a_57368_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1524 a_9138_19307# a_8422_18706# a_7152_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1525 a_8462_6503# a_8292_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1526 VDD C[76] a_36965_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 VSS a_41116_13071# a_42041_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1528 a_43331_5620# a_42739_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1529 a_52681_1566# a_52063_739# a_52281_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1530 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1531 a_1107_14292# a_1020_14194# a_1025_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1532 a_2995_14292# a_2908_14194# a_2913_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1533 VSS a_43004_13071# a_43929_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1534 a_3591_6676# a_4985_6509# a_5025_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1535 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1536 a_52452_18251# a_51782_18732# a_52052_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1537 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1538 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1539 a_50511_6419# a_50285_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1540 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1541 a_54555_6676# a_54061_6509# a_54106_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1542 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1543 a_7250_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1544 a_41228_19307# a_41226_18251# a_41539_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1545 a_22332_13071# a_21968_13134# a_22236_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1546 a_5591_510# a_4823_765# a_3605_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1547 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1548 a_10121_12994# a_9951_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1549 a_46884_18251# a_46118_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1550 a_41443_5620# a_40851_6509# a_39457_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1551 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_35232_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1552 a_48772_18251# a_48006_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1553 a_42555_14292# a_42550_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1554 a_43247_1566# a_42577_765# a_42847_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1555 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1556 VSS a_19349_18953# a_19299_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1557 a_18047_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1558 a_19935_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1559 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1560 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1561 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_11239_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1562 a_35791_1566# a_35025_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1563 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1564 a_19349_18953# a_18474_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1565 a_47003_6676# a_46735_6419# a_46554_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1566 a_8842_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1567 a_25599_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1568 a_48760_14127# a_48394_13134# a_46774_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 a_36570_928# a_35695_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1570 a_54667_510# a_54665_1566# a_54978_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1571 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1572 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1573 a_3687_6676# a_3097_6509# a_3591_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1574 a_46884_18251# a_46118_18732# a_46788_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1575 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1576 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_26698_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1577 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1578 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1579 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1580 a_20348_13071# a_19854_12988# a_19899_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1581 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1582 VDD a_22465_6676# a_23390_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1583 a_41802_5455# a_41443_5620# a_41441_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1584 a_20460_19307# a_19692_18732# a_18474_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1585 a_54424_14127# a_54058_13134# a_52438_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1586 a_8987_6419# a_8761_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1587 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1588 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1589 a_58754_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1590 VSS a_38229_18953# a_38179_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1591 a_52254_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1592 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1593 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1594 VDD a_12534_13134# a_12348_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1595 a_38229_18953# a_37354_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1596 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1597 a_32015_1566# a_31301_739# a_31919_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1598 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_57735_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1599 a_49001_1566# a_48235_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1600 a_58427_6676# a_58429_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1601 a_44479_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1602 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1603 a_44892_13071# a_46280_12988# a_46320_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 a_54061_6509# C[60] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1605 a_52399_6419# a_52173_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1606 VSS a_31301_739# a_31249_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1607 a_3605_1566# a_4875_739# a_5066_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1608 a_60413_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 a_58200_14127# a_57608_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1610 VDD C[83] a_23749_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1611 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1612 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1613 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1614 a_32003_5620# a_31411_6509# a_30017_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1615 a_33807_1566# a_33137_765# a_33407_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1616 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1617 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1618 a_54326_13071# a_55946_13134# a_55760_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1619 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_6918_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1620 VSS a_14533_1000# a_14506_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1621 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1622 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1623 a_4251_18953# a_3376_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1624 a_20460_19307# a_19744_18706# a_18474_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1625 VSS a_27900_13071# a_28825_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1626 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1627 a_13031_6676# a_12537_6509# a_12582_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1628 a_7477_1566# a_6711_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1629 a_26353_510# a_25637_739# a_24367_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1630 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1631 VSS C[21] a_19744_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1632 VDD a_54326_13071# a_55251_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1633 a_57538_6503# a_57368_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1634 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1635 a_26124_19307# a_26122_18251# a_26435_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1636 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1637 a_52667_6676# a_54061_6509# a_54101_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1638 a_50889_1566# a_50123_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1639 a_47017_1566# a_46347_765# a_46617_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1640 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1641 a_5577_5620# a_4985_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1642 VSS a_19973_739# a_19921_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1643 a_3701_1566# a_2935_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1644 a_51645_12994# a_51475_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1645 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_43690_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1646 VSS a_55839_739# a_55787_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1647 a_22575_1566# a_21861_739# a_22479_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1648 VDD a_39457_6676# a_40382_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1649 a_42234_928# a_41359_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1650 a_22064_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1651 a_18703_1566# a_19973_739# a_20164_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1652 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_58198_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1653 a_47101_5620# a_46735_6419# a_45121_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1654 a_37681_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1655 a_39324_13071# a_39326_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1656 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1657 a_22016_5455# a_22011_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1658 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1659 a_45004_19307# a_45002_18251# a_45315_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1660 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1661 VSS C[69] a_50175_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1662 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1663 VDD a_12198_18706# a_12416_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1664 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1665 a_3689_5620# a_3097_6509# a_1703_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1666 VDD a_31072_18706# a_31020_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1667 a_15785_12994# a_15615_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1668 VDD a_32960_18706# a_32908_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1669 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1670 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1671 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1672 a_52763_6676# a_52173_6509# a_52667_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1673 VDD C[74] a_40741_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1674 a_29421_14292# a_29334_14194# a_29339_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1675 a_10121_12994# a_9951_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1676 a_46774_13071# a_46506_13134# a_46325_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1677 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1678 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1679 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1680 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1681 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1682 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1683 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_12353_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1684 VSS a_22465_6676# a_23390_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1685 VSS a_30906_928# a_30856_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1686 a_10730_1811# a_10757_1000# a_10742_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1687 a_1717_1566# a_1047_765# a_1317_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1688 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1689 a_56312_14127# a_55720_12988# a_54326_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1690 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1691 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_35777_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1692 a_24236_19307# a_23468_18732# a_22250_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1693 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1694 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1695 VSS a_18303_1000# a_18276_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1696 a_1801_5620# a_1435_6419# a_565_18708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1697 VDD a_30017_6676# a_30942_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1698 VDD a_12427_739# a_12645_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1699 a_50875_6676# a_50511_6419# a_50779_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1700 VSS a_17690_928# a_17640_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1701 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1702 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1107_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1703 a_31788_19307# a_31020_18732# a_29802_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1704 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1705 a_46506_13134# a_46280_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1706 VSS a_53556_928# a_53506_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1707 a_53327_18953# a_52452_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1708 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_42784_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1709 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1710 a_11143_6676# a_12537_6509# a_12577_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1711 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1712 a_52779_510# a_52063_739# a_50793_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1713 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1714 a_3460_14127# a_2868_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1715 a_46509_6509# C[56] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1716 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_32001_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1717 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1718 VDD a_8758_13134# a_8572_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1719 a_54058_13134# a_53832_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1720 a_10776_5455# a_10689_5687# a_10694_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1721 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1722 a_57332_928# a_56457_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1723 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1724 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1725 a_8027_18953# a_7152_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1726 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1727 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_47460_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1728 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1729 VDD C[70] a_48287_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1730 a_22693_14292# a_22334_14127# a_22332_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1731 VSS C[19] a_23520_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1732 a_13691_18953# a_12816_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1733 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1734 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1735 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1736 a_11239_6676# a_10649_6509# a_11143_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1737 VSS a_39457_6676# a_40382_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1738 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1739 VSS a_54326_13071# a_55251_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1740 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1741 VDD a_17856_18706# a_17804_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1742 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1743 a_58102_13071# a_57608_12988# a_57653_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1744 a_46870_13071# a_46872_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1745 a_59990_13071# a_59496_12988# a_59541_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1746 VDD a_1703_6676# a_2628_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1747 a_54569_1566# a_53899_765# a_54169_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1748 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1749 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1750 a_41573_14292# a_41214_14127# a_41212_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1751 VSS a_35295_1000# a_35268_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1752 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1753 VDD a_19744_18706# a_19962_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1754 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1755 a_58198_13071# a_57608_12988# a_58102_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1756 a_31690_18251# a_31072_18706# a_31290_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1757 a_54422_13071# a_54424_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1758 a_23331_12994# a_23161_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1759 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_22561_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1760 a_20689_510# a_19921_765# a_18703_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1761 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1762 a_50793_1566# a_52011_765# a_52254_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1763 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1764 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1765 a_33674_18251# a_32960_18706# a_33578_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1766 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1767 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1768 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_3687_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1769 a_60102_19307# a_60100_18251# a_60413_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1770 a_47892_928# a_47017_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1771 VDD C[23] a_15968_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1772 VDD a_36736_18706# a_36684_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1773 a_30883_12994# a_30713_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1774 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_19899_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1775 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_12664_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1776 a_18322_5455# a_18235_5687# a_18240_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1777 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1778 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_21787_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1779 VDD a_8422_18706# a_8640_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1780 a_15785_12994# a_15615_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1781 a_24138_18251# a_23468_18732# a_23738_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1782 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1783 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1784 a_26241_6676# a_25973_6419# a_25792_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1785 a_15029_1566# a_14263_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1786 a_50877_5620# a_50511_6419# a_48891_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1787 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1788 VSS a_45775_18953# a_45725_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1789 a_1572_14127# a_980_12988# a_794_737# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1790 a_31690_18251# a_31020_18732# a_31290_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1791 a_48774_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1792 VSS a_30017_6676# a_30942_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1793 VSS a_18085_739# a_18033_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1794 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1795 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1796 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1797 a_45233_510# a_44465_765# a_43247_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1798 a_58443_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1799 VDD C[13] a_34848_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1800 VSS a_5360_18251# a_5362_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1801 VDD C[12] a_36736_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1802 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1803 a_27336_6503# a_27166_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1804 a_56326_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1805 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1806 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_40667_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1807 a_13129_5620# a_12537_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1808 a_57332_928# a_56457_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1809 VSS a_57103_18953# a_57053_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1810 a_6689_14292# a_6684_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1811 VSS a_6763_739# a_6711_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1812 VDD C[9] a_42400_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1813 VSS a_16186_18747# a_16159_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1814 a_43018_18251# a_42348_18732# a_42618_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1815 VSS a_25855_1000# a_25828_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1816 VDD a_31408_13134# a_31222_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1817 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1818 a_18570_18251# a_17804_18732# a_18474_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1819 a_1302_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1820 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1821 VSS a_23738_18747# a_23711_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1822 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1823 a_24353_6676# a_23859_6509# a_23904_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1824 a_26110_14127# a_25744_13134# a_24124_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1825 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1826 VDD a_36965_739# a_37183_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1827 a_11241_5620# a_10649_6509# a_9255_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1828 a_31492_1811# a_31519_1000# a_31504_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1829 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1830 a_13045_1566# a_12375_765# a_12645_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1831 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1832 a_21835_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1833 a_33070_12988# C[113] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1834 a_14690_13071# a_16304_13134# a_16118_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1835 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_29421_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1836 a_16801_6676# a_16533_6419# a_16352_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1837 a_16572_13071# a_17966_12988# a_18006_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1838 a_26469_14292# a_26110_14127# a_26108_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1839 VDD a_35413_6419# a_35227_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1840 a_35314_5455# a_35227_5687# a_35232_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1841 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1842 a_16586_18251# a_15968_18706# a_16186_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1843 a_37450_18251# a_36684_18732# a_37354_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1844 a_40622_12988# C[117] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1845 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1846 VSS a_42618_18747# a_42591_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1847 VDD a_50779_6676# a_51704_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1848 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1849 a_18570_18251# a_17856_18706# a_18474_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1850 VSS a_1703_6676# a_2628_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1851 a_9269_1566# a_8651_739# a_8869_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1852 a_8613_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1853 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1854 a_22236_13071# a_23630_12988# a_23670_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1855 a_43233_6676# a_42965_6419# a_42784_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1856 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1857 a_43114_18251# a_42348_18732# a_43018_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1858 a_24124_13071# a_25518_12988# a_25558_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1859 a_17896_6503# a_17726_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1860 a_11600_5455# a_11241_5620# a_11239_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1861 a_43247_1566# a_44517_739# a_44708_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1862 a_45002_18251# a_44236_18732# a_44906_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1863 VSS a_21861_739# a_21809_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1864 a_60329_1566# a_59615_739# a_60219_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1865 a_28552_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1866 a_3362_13071# a_2868_12988# a_2913_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1867 a_22052_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1868 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1869 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1870 a_33564_13071# a_35184_13134# a_34998_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1871 a_7099_6419# a_6873_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1872 a_45121_6676# a_44627_6509# a_44672_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1873 a_31538_5455# a_31451_5687# a_31456_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1874 VSS a_10310_18706# a_10258_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1875 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1876 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1877 a_35452_13071# a_36846_12988# a_36886_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1878 a_45349_14292# a_44990_14127# a_44988_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1879 a_28225_6676# a_28227_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1880 a_18799_1566# a_18033_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1881 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1882 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1883 a_3458_13071# a_2868_12988# a_3362_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1884 VSS a_4480_928# a_4430_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1885 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1886 a_35466_18251# a_34848_18706# a_35066_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1887 a_58198_13071# a_58200_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1888 a_41116_13071# a_42736_13134# a_42550_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1889 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_16668_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1890 a_24353_6676# a_25973_6419# a_25787_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1891 a_16913_510# a_16197_739# a_14933_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1892 VSS a_42847_1000# a_42820_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1893 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1894 a_37450_18251# a_36736_18706# a_37354_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1895 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18556_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1896 VDD a_33564_13071# a_34489_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1897 a_22197_6419# a_21971_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1898 VDD a_704_928# a_654_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1899 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1900 a_9040_18251# a_10310_18706# a_10501_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1901 VDD a_31072_18706# a_31290_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1902 a_43004_13071# a_44398_12988# a_44438_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 a_3178_1811# a_3205_1000# a_3190_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1904 a_11026_19307# a_10310_18706# a_9040_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1905 a_23331_12994# a_23161_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1906 a_34659_12994# a_34489_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1907 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1908 a_12914_19307# a_12198_18706# a_10928_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1909 a_43018_18251# a_42400_18706# a_42618_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1910 VDD a_51834_18706# a_51782_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1911 a_45002_18251# a_44288_18706# a_44906_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1912 a_41345_6676# a_40851_6509# a_40896_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1913 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1914 a_48295_14292# a_48208_14194# a_48213_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1915 a_565_18708# a_870_18706# a_1061_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1916 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1917 a_30883_12994# a_30713_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1918 a_25973_6419# a_25747_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1919 a_6966_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1920 a_3474_19307# a_2758_18706# a_1488_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1921 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1922 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1923 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1924 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1925 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1926 VDD a_25973_6419# a_25787_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1927 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1928 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_22693_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1929 a_27336_6503# a_27166_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1930 a_32794_928# a_31919_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1931 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1932 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1933 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_37436_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1934 a_33793_6676# a_33525_6419# a_33344_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1935 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1936 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_37202_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1937 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1938 a_22465_6676# a_23859_6509# a_23899_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1939 a_50889_1566# a_50175_739# a_50793_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1940 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1941 a_9040_18251# a_10258_18732# a_10501_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1942 VDD a_23125_18953# a_23075_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1943 VDD C[5] a_49946_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1944 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1945 a_50378_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1946 a_1586_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1947 a_9138_19307# a_9136_18251# a_9449_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1948 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1949 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_13488_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1950 a_19854_12988# C[106] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1951 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1952 VDD a_9255_6676# a_10180_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1953 a_34888_6503# a_34718_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1954 VDD a_30677_18953# a_30627_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1955 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1956 a_6644_12988# C[99] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1957 VDD a_1099_739# a_1047_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1958 a_565_18708# a_818_18732# a_1061_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1959 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1960 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1961 a_12898_13071# a_12534_13134# a_12802_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1962 a_45544_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1963 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_41573_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1964 a_14919_6676# a_16533_6419# a_16347_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1965 a_29886_14127# a_29294_12988# a_27900_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1966 a_25518_12988# C[109] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1967 a_18883_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1968 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1969 a_1717_1566# a_2935_765# a_3178_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1970 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1971 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1972 a_45217_6676# a_45219_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1973 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1974 VSS a_3701_1566# a_3703_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1975 VDD a_42005_18953# a_41955_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1976 a_29898_18251# a_29132_18732# a_29802_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1977 a_31905_6676# a_31411_6509# a_31456_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1978 a_22561_6676# a_21971_6509# a_22465_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1979 a_39189_6419# a_38963_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1980 VSS a_50779_6676# a_51704_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1981 VDD C[90] a_10539_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1982 VDD a_44517_739# a_44735_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1983 VSS a_39338_18251# a_39340_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1984 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1985 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1986 a_18192_13134# a_17966_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1987 a_38734_12988# C[116] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1988 a_25013_18953# a_24138_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1989 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1990 a_6870_13134# a_6644_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1991 a_31263_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1992 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1993 a_17896_6503# a_17726_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1994 a_43233_6676# a_44627_6509# a_44667_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1995 a_56030_1811# a_56057_1000# a_56042_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1996 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1997 a_26012_13071# a_27632_13134# a_27446_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1998 a_25744_13134# a_25518_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1999 a_44398_12988# C[119] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2000 VDD a_38853_739# a_38801_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2001 a_11026_19307# a_10258_18732# a_9040_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2002 a_32565_18953# a_31690_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2003 a_37763_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2004 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2005 a_5479_6676# a_5211_6419# a_5030_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2006 a_42965_6419# a_42739_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2007 VSS a_46617_1000# a_46590_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2008 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2009 VDD a_18460_13071# a_19385_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2010 VDD a_42965_6419# a_42779_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2011 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2012 a_32017_510# a_32015_1566# a_32328_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2013 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2014 a_59818_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2015 a_43427_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2016 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2017 a_7138_13071# a_6644_12988# a_6689_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2018 VSS a_22575_1566# a_22577_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2019 a_37340_13071# a_38960_13134# a_38774_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2020 VDD a_26012_13071# a_26937_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2021 a_37072_13134# a_36846_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2022 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2023 a_7250_19307# a_6482_18732# a_5264_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2024 a_38960_13134# a_38734_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2025 a_20673_6676# a_20309_6419# a_20577_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2026 a_39457_6676# a_40851_6509# a_40891_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2027 VDD a_57727_739# a_57945_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2028 a_6574_6503# a_6404_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2029 a_39553_6676# a_39189_6419# a_39457_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2030 a_52254_1811# a_52281_1000# a_52266_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2031 a_60447_14292# a_60088_14127# a_60086_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2032 a_57103_18953# a_56228_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2033 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2034 a_50550_13071# a_51944_12988# a_51984_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2035 a_44624_13134# a_44398_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2036 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2037 a_50564_18251# a_49946_18706# a_50164_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2038 a_16307_6509# C[40] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2039 a_26351_1566# a_25585_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2040 a_52548_18251# a_51834_18706# a_52452_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2041 VDD a_37340_13071# a_38265_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2042 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2043 VSS a_6534_18706# a_6482_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2044 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2045 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2046 a_29749_6419# a_29523_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2047 VSS C[95] a_1099_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2048 a_56076_5455# a_55989_5687# a_55994_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2049 a_3591_6676# a_3097_6509# a_3142_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2050 a_31411_6509# C[48] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2051 a_27130_928# a_26255_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2052 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2053 VSS a_33564_13071# a_34489_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2054 VDD a_44892_13071# a_45817_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2055 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_17258_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2056 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2057 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2058 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2059 a_3376_18251# a_4646_18706# a_4837_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2060 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2061 a_21787_14292# a_21782_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2062 a_32362_5455# a_32003_5620# a_32001_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2063 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2064 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2065 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2066 a_34659_12994# a_34489_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2067 VDD C[86] a_18085_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2068 a_5589_1566# a_4823_765# a_5493_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2069 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2070 a_7250_19307# a_6534_18706# a_5264_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2071 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 a_24451_5620# a_23859_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2073 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2074 a_59770_5455# a_59765_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2075 a_31788_19307# a_31786_18251# a_32099_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2076 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_50646_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2077 VSS C[28] a_6534_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2078 a_33660_13071# a_33662_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2079 VSS a_9255_6676# a_10180_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2080 a_34888_6503# a_34718_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2081 a_48987_6676# a_48989_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2082 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2083 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2084 a_60219_6676# a_59615_739# a_59833_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2085 VDD C[2] a_55610_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2086 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_44754_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2087 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2088 VDD a_14086_18706# a_14034_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2089 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2090 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2091 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2092 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2093 a_20444_13071# a_20080_13134# a_20348_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2094 a_30017_6676# a_31411_6509# a_31451_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2095 VDD a_48287_739# a_48505_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2096 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_16352_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2097 a_40667_14292# a_40662_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2098 a_22563_5620# a_21971_6509# a_20577_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2099 a_24367_1566# a_23697_765# a_23967_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2100 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2101 a_7790_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2102 a_16159_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2103 a_29788_13071# a_29520_13134# a_29339_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2104 a_1290_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2105 VSS a_17461_18953# a_17411_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2106 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2107 VDD a_51668_928# a_51618_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2108 a_7463_6676# a_7465_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2109 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2110 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2111 a_3703_510# a_2987_739# a_1717_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2112 a_58212_18251# a_57446_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2113 VDD a_46735_6419# a_46549_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2114 a_17690_928# a_16815_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2115 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2116 a_28012_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2117 a_46872_14127# a_46506_13134# a_44892_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2118 a_1435_6419# a_1209_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2119 a_59426_6503# a_59256_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2120 a_3591_6676# a_5211_6419# a_5025_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2121 a_51202_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2122 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2123 a_33299_6509# C[49] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2124 a_35793_510# a_35025_765# a_33807_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2125 VDD C[24] a_14086_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2126 a_22922_5455# a_22563_5620# a_22561_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2127 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2128 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_57964_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2129 VSS a_54436_18251# a_54438_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2130 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_48295_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2131 a_53832_12988# C[124] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2132 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2133 a_27914_18251# a_29132_18732# a_29375_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2134 a_35039_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2135 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2136 a_44122_928# a_43247_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2137 a_47892_928# a_47017_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2138 VSS a_36341_18953# a_36291_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2139 a_20675_5620# a_20309_6419# a_18689_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2140 a_39555_5620# a_39189_6419# a_37569_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2141 VDD a_10646_13134# a_10460_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2142 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2143 a_52861_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2144 a_48760_14127# a_48168_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2145 a_47099_6676# a_46509_6509# a_47003_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2146 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2147 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2148 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_55847_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2149 VDD C[77] a_35077_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2150 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2151 VSS a_43893_18953# a_43843_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2152 a_6574_6503# a_6404_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2153 a_50793_1566# a_50175_739# a_50393_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2154 a_28241_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2155 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2156 a_9915_18953# a_9040_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2157 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2158 VSS a_18460_13071# a_19385_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2159 a_1703_6676# a_3097_6509# a_3137_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2160 a_52170_13134# a_51944_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2161 a_52438_13071# a_54058_13134# a_53872_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2162 a_52667_6676# a_52173_6509# a_52218_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2163 VSS C[73] a_42629_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2164 a_2363_18953# a_1488_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2165 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2166 VSS a_14304_18747# a_14277_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2167 VSS a_26012_13071# a_26937_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2168 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2169 a_9367_510# a_9365_1566# a_9678_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2170 a_16684_19307# a_16682_18251# a_16995_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2171 a_59722_13134# a_59496_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2172 a_41359_1566# a_40689_765# a_40959_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2173 a_18572_19307# a_18570_18251# a_18883_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2174 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2175 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2176 a_18556_13071# a_18558_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2177 VDD a_52438_13071# a_53363_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2178 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2179 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2180 VDD a_59615_739# a_59563_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2181 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2182 a_33807_1566# a_35077_739# a_35268_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2183 a_24236_19307# a_24234_18251# a_24547_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2184 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2185 VSS a_37340_13071# a_38265_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2186 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2187 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_48524_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2188 a_6954_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2189 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2190 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2191 VDD a_59990_13071# a_60915_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2192 a_34682_928# a_33807_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2193 a_58441_1566# a_57675_765# a_58345_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2194 a_52779_510# a_52777_1566# a_53090_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2195 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2196 a_1799_6676# a_1209_6509# a_1703_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2197 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2198 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2199 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2200 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_24810_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2201 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2202 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2203 VSS a_44892_13071# a_45817_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2204 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2205 VDD a_20577_6676# a_21502_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2206 VSS a_44122_928# a_44072_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2207 a_37452_19307# a_37450_18251# a_37763_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2208 a_9483_14292# a_9124_14127# a_9122_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2209 a_8761_6509# C[36] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2210 a_56866_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2211 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2212 a_14704_18251# a_14086_18706# a_14304_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2213 a_37436_13071# a_37438_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2214 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_56310_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2215 a_13031_6676# a_12763_6419# a_12582_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2216 a_43345_510# a_42629_739# a_41359_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2217 a_50366_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2218 VDD a_23520_18706# a_23468_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2219 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2220 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2221 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2222 a_30127_1566# a_29413_739# a_30031_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2223 VDD a_10310_18706# a_10528_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2224 a_43116_19307# a_43114_18251# a_43427_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2225 a_48989_5620# a_48397_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2226 a_13897_12994# a_13727_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2227 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2228 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2229 a_45233_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2230 a_8256_928# a_7381_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2231 a_21968_13134# a_21742_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2232 a_52173_6509# C[59] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2233 a_59426_6503# a_59256_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2234 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2235 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2236 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2237 a_48760_14127# a_48168_12988# a_46774_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2238 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_5030_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2239 VSS a_12645_1000# a_12618_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2240 VDD a_42400_18706# a_42348_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2241 a_47101_5620# a_46509_6509# a_45121_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2242 a_5589_1566# a_4823_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2243 a_56214_13071# a_55946_13134# a_55765_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2244 a_11143_6676# a_10649_6509# a_10694_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2245 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2246 a_49001_1566# a_48235_765# a_48905_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2247 VDD C[16] a_29184_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2248 a_22348_19307# a_21580_18732# a_20362_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2249 VSS a_58212_18251# a_58214_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2250 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_13259_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2251 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2252 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2253 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2254 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2255 a_50137_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2256 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_8577_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2257 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2258 VSS a_51439_18953# a_51389_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2259 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2260 a_59577_18006# a_59604_18747# a_59589_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2261 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2262 a_50779_6676# a_52173_6509# a_52213_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2263 a_59541_14292# a_59536_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2264 a_55720_12988# C[125] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2265 a_51439_18953# a_50564_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2266 a_56637_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2267 a_3689_5620# a_3097_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2268 a_11255_510# a_10487_765# a_9269_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2269 a_59806_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2270 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2271 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_41802_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2272 a_41359_1566# a_42577_765# a_42820_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2273 a_20687_1566# a_19973_739# a_20591_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2274 a_39567_1566# a_38853_739# a_39471_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2275 a_20176_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2276 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2277 VDD a_6870_13134# a_6684_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2278 a_23354_928# a_22479_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2279 a_39056_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2280 VDD a_6139_18953# a_6089_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2281 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2282 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2283 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2284 a_6139_18953# a_5264_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2285 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2286 a_15342_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2287 a_10501_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2288 a_1801_5620# a_1209_6509# a_565_18708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2289 a_3605_1566# a_2935_765# a_3205_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2290 a_40851_6509# C[53] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2291 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2292 a_20805_14292# a_20446_14127# a_20444_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2293 a_15015_6676# a_15017_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2294 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2295 a_15113_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2296 a_11803_18953# a_10928_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2297 VSS C[20] a_21632_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2298 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2299 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2300 a_11143_6676# a_12763_6419# a_12577_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2301 a_46004_928# a_45135_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2302 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2303 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2304 VSS a_20577_6676# a_21502_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2305 VDD a_14315_739# a_14533_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2306 VSS a_52438_13071# a_53363_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2307 a_57837_6509# C[62] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2308 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2309 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2310 VDD C[66] a_55839_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2311 a_14933_1566# a_14315_739# a_14533_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2312 VDD a_15968_18706# a_15916_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2313 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2314 a_32133_14292# a_31774_14127# a_31772_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2315 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2316 a_22250_18251# a_21632_18706# a_21850_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2317 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2318 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2319 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2320 a_56214_13071# a_55720_12988# a_55765_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2321 a_60331_510# a_60329_1566# a_60642_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2322 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2323 a_24234_18251# a_23520_18706# a_24138_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2324 VSS a_59990_13071# a_60915_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2325 a_12763_6419# a_12537_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2326 a_9269_1566# a_10539_739# a_10730_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2327 VSS a_16415_1000# a_16388_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2328 a_50662_19307# a_50660_18251# a_50973_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2329 VDD a_12763_6419# a_12577_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2330 VSS C[10] a_40512_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2331 a_52550_19307# a_52548_18251# a_52861_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2332 a_21443_12994# a_21273_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2333 a_56310_13071# a_55720_12988# a_56214_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2334 VDD a_10539_739# a_10757_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2335 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2336 a_52534_13071# a_52536_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2337 a_29616_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2338 a_31786_18251# a_31072_18706# a_31690_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2339 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_49348_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2340 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2341 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2342 a_9255_6676# a_10649_6509# a_10689_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2343 VSS C[65] a_57727_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2344 VDD a_34848_18706# a_34796_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2345 a_22052_1811# a_22079_1000# a_22064_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2346 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_30113_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2347 a_41130_18251# a_40512_18706# a_40730_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2348 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2349 a_13897_12994# a_13727_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2350 a_48662_13071# a_48394_13134# a_48213_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2351 a_22250_18251# a_21580_18732# a_21850_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2352 a_43114_18251# a_42400_18706# a_43018_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2353 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2354 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2355 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2356 a_55444_928# a_54569_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2357 a_50891_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2358 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2359 a_46886_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2360 a_60676_5455# a_60317_5620# a_60315_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2361 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2362 a_12353_14292# a_12348_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2363 VDD C[71] a_46399_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2364 VDD C[14] a_32960_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2365 VSS a_3472_18251# a_3474_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2366 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2367 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2368 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2369 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2370 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2371 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2372 a_46788_18251# a_48006_18732# a_48249_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2373 a_2949_18006# a_2976_18747# a_2961_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2374 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2375 VSS a_55215_18953# a_55165_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2376 VSS a_59220_928# a_59170_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2377 a_41130_18251# a_40460_18732# a_40730_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2378 a_4801_14292# a_4796_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2379 a_29568_5455# a_29563_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2380 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2381 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2382 a_59496_12988# C[127] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2383 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_9483_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2384 a_18785_6676# a_18787_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2385 a_16682_18251# a_15916_18732# a_16586_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2386 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2387 a_30031_1566# a_29413_739# a_29631_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2388 a_52681_1566# a_52011_765# a_52281_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2389 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2390 VSS a_21850_18747# a_21823_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2391 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_14552_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2392 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2393 a_24222_14127# a_23856_13134# a_22236_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2394 VDD a_18085_739# a_18303_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2395 VSS a_33407_1000# a_33380_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2396 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2397 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_39553_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2398 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2399 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2400 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_1799_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2401 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2402 a_31182_12988# C[112] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2403 VSS a_33178_18747# a_33151_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2404 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_27533_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2405 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2406 a_14277_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2407 VSS a_36965_739# a_36913_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2408 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2409 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2410 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2411 a_14690_13071# a_16078_12988# a_16118_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2412 a_35562_18251# a_34796_18732# a_35466_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2413 a_30211_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2414 VDD a_16533_6419# a_16347_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2415 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_10776_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2416 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2417 a_27998_14127# a_27406_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2418 a_29224_6503# a_29054_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2419 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2420 a_16682_18251# a_15968_18706# a_16586_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2421 VSS a_40730_18747# a_40703_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2422 a_6725_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2423 a_43102_14127# a_42736_13134# a_41116_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2424 a_44990_14127# a_44624_13134# a_43004_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2425 a_24124_13071# a_25744_13134# a_25558_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2426 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2427 a_13141_1566# a_12375_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2428 a_24353_6676# a_24085_6419# a_23904_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2429 a_41226_18251# a_40460_18732# a_41130_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2430 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2431 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2432 a_1474_13071# a_980_12988# a_1025_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2433 a_13920_928# a_13045_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2434 a_31676_13071# a_33296_13134# a_33110_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2435 a_56555_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2436 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2437 a_26353_510# a_25585_765# a_24367_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2438 VDD a_24124_13071# a_25049_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2439 a_25448_6503# a_25278_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2440 a_56457_1566# a_57675_765# a_57918_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2441 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2442 a_33564_13071# a_34958_12988# a_34998_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2443 a_1570_13071# a_980_12988# a_1474_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2444 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2445 a_11241_5620# a_10649_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2446 a_20591_1566# a_19973_739# a_20191_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2447 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2448 a_33578_18251# a_32960_18706# a_33178_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2449 a_39471_1566# a_38853_739# a_39071_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2450 a_35562_18251# a_34848_18706# a_35466_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2451 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2452 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2453 VSS a_23967_1000# a_23940_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2454 a_39228_13071# a_40622_12988# a_40662_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2455 VDD a_31676_13071# a_32601_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2456 a_41116_13071# a_42510_12988# a_42550_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2457 VDD a_8256_928# a_8206_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2458 VSS a_5093_1000# a_5066_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2459 VSS a_59386_18706# a_59334_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2460 a_21443_12994# a_21273_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2461 a_35777_6676# a_35779_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2462 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2463 a_22465_6676# a_21971_6509# a_22016_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2464 a_37301_6419# a_37075_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2465 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2466 VDD a_35077_739# a_35295_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2467 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2468 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2469 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_27996_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2470 a_46407_14292# a_46320_14194# a_46325_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2471 a_56228_18251# a_57498_18706# a_57689_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2472 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2473 a_11157_1566# a_10487_765# a_10757_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2474 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2475 a_58116_18251# a_59386_18706# a_59577_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2476 a_1586_19307# a_870_18706# a_565_18708# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2477 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2478 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_20805_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2479 VSS a_34682_928# a_34632_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2480 a_14802_19307# a_14800_18251# a_15113_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2481 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2482 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_33660_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2483 VDD a_29413_739# a_29361_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2484 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35548_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2485 a_33905_510# a_33189_739# a_31919_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2486 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_54651_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2487 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_18322_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2488 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2489 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2490 a_33426_5455# a_33339_5687# a_33344_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2491 VDD a_21237_18953# a_21187_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2492 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2493 VDD a_33525_6419# a_33339_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2494 a_46216_6503# a_46046_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2495 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2496 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2497 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2498 a_16078_12988# C[104] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2499 a_8577_14292# a_8572_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2500 a_17966_12988# C[105] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2501 a_24367_1566# a_25637_739# a_25828_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2502 a_4756_12988# C[98] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2503 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2504 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2505 a_26664_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2506 a_26110_14127# a_25518_12988# a_24124_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2507 a_20164_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2508 a_27998_14127# a_27406_12988# a_26012_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2509 VSS C[66] a_55839_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2510 a_39044_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2511 a_16995_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2512 a_18787_5620# a_18195_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2513 a_26337_6676# a_26339_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2514 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2515 a_29886_14127# a_29520_13134# a_27900_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2516 a_16911_1566# a_16145_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2517 VDD a_40117_18953# a_40067_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2518 a_15031_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2519 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2520 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2521 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2522 a_7234_13071# a_6870_13134# a_7138_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2523 a_20309_6419# a_20083_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2524 VSS a_40959_1000# a_40932_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2525 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2526 a_16572_13071# a_18192_13134# a_18006_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2527 a_39326_14127# a_38734_12988# a_37340_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2528 a_16304_13134# a_16078_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2529 a_29224_6503# a_29054_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2530 a_23125_18953# a_22250_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2531 a_36846_12988# C[115] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2532 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2533 a_3094_13134# a_2868_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2534 a_4982_13134# a_4756_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2535 a_1290_1811# a_1317_1000# a_1302_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2536 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2537 a_43004_13071# a_42736_13134# a_42555_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2538 a_39338_18251# a_38572_18732# a_39242_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2539 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2540 a_35875_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2541 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2542 a_23856_13134# a_23630_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2543 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2544 VDD a_19973_739# a_19921_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2545 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2546 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2547 a_30677_18953# a_29802_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2548 a_50660_18251# a_49894_18732# a_50564_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2549 a_31919_1566# a_33137_765# a_33380_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2550 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2551 VDD a_16572_13071# a_17497_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2552 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_53959_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2553 a_25448_6503# a_25278_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2554 a_5112_5455# a_5025_5687# a_5030_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2555 VSS a_12427_739# a_12375_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2556 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2557 a_35184_13134# a_34958_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2558 a_49551_18953# a_48676_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2559 a_35452_13071# a_37072_13134# a_36886_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2560 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_35314_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2561 a_5362_19307# a_4594_18732# a_3376_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2562 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2563 a_20577_6676# a_21971_6509# a_22011_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2564 a_45231_1566# a_44465_765# a_45135_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2565 a_56312_14127# a_55720_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2566 a_29604_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2567 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2568 a_48662_13071# a_50056_12988# a_50096_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2569 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_11600_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2570 a_58443_510# a_57727_739# a_56457_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2571 a_42736_13134# a_42510_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2572 a_1336_5455# a_1249_5687# a_1254_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2573 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2574 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2575 VSS a_24124_13071# a_25049_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2576 VDD a_35452_13071# a_36377_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2577 VSS a_4646_18706# a_4594_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2578 a_50660_18251# a_49946_18706# a_50564_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2579 VSS C[64] a_59615_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2580 a_43656_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2581 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2582 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2583 VSS a_35077_739# a_35025_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2584 VSS a_31676_13071# a_32601_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2585 a_11371_14292# a_11012_14127# a_11010_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2586 a_35779_5620# a_35187_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2587 a_1488_18251# a_2758_18706# a_2949_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2588 a_52218_5455# a_52213_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2589 a_44853_6419# a_44627_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2590 VSS a_1813_1566# a_1815_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2591 a_5362_19307# a_4646_18706# a_3376_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2592 a_24220_13071# a_24222_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2593 a_29884_13071# a_29294_12988# a_29788_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2594 a_20673_6676# a_20083_6509# a_20577_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2595 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2596 a_57701_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2597 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2598 a_39553_6676# a_38963_6509# a_39457_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2599 a_50793_1566# a_52063_739# a_52254_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2600 a_46216_6503# a_46046_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2601 a_29900_19307# a_29898_18251# a_30211_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2602 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_39324_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2603 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2604 VSS C[29] a_4646_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2605 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2606 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2607 a_27635_6509# C[46] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2608 VSS C[79] a_31301_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2609 VDD a_36965_739# a_36913_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2610 a_54142_1811# a_54169_1000# a_54154_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2611 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2612 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2613 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2614 VDD C[3] a_53722_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2615 a_3591_6676# a_3323_6419# a_3142_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2616 VDD a_12198_18706# a_12146_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2617 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_7000_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2618 VSS a_10144_928# a_10094_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2619 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2620 sky130_fd_sc_hd__buf_2_0/X a_27668_9428# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2621 a_35791_1566# a_35025_765# a_35695_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2622 a_30129_510# a_30127_1566# a_30440_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2623 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2624 a_43100_13071# a_43102_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2625 VSS a_15573_18953# a_15523_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2626 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2627 a_27900_13071# a_27632_13134# a_27451_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2628 a_58063_6419# a_57837_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2629 VSS a_39567_1566# a_39569_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2630 VDD a_58063_6419# a_57877_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2631 VDD a_55839_739# a_56057_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2632 a_4686_6503# a_4516_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2633 a_37665_6676# a_37301_6419# a_37569_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2634 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2635 a_56324_18251# a_55558_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2636 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2637 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_10694_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2638 a_26124_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2639 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2640 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_10465_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2641 a_39228_13071# a_38960_13134# a_38779_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2642 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2643 VDD C[25] a_12198_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2644 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2645 a_54424_14127# a_53832_12988# a_52438_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2646 a_50056_12988# C[122] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2647 a_51944_12988# C[123] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2648 a_54188_5455# a_54101_5687# a_54106_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2649 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2650 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1025_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2651 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_46407_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2652 a_1703_6676# a_1209_6509# a_1254_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2653 VDD a_54287_6419# a_54101_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2654 a_25242_928# a_24367_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2655 VSS a_49780_928# a_49730_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2656 VSS a_34453_18953# a_34403_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2657 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2658 a_5264_18251# a_4594_18732# a_4864_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2659 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2660 a_60088_14127# a_59496_12988# a_58102_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2661 a_57930_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2662 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2663 a_54436_18251# a_53670_18732# a_54340_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2664 a_30474_5455# a_30115_5620# a_30113_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2665 a_50973_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2666 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2667 VDD C[87] a_16197_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2668 a_45004_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2669 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2670 a_37354_18251# a_38572_18732# a_38815_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2671 VDD a_8651_739# a_8599_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2672 a_57882_5455# a_57877_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2673 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2674 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2675 VSS a_16572_13071# a_17497_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2676 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2677 a_9138_19307# a_8370_18732# a_7152_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2678 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2679 a_50550_13071# a_52170_13134# a_51984_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2680 VDD a_4982_13134# a_4796_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2681 a_50282_13134# a_50056_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2682 a_58345_1566# a_59563_765# a_59806_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2683 a_48623_6419# a_48397_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2684 a_10420_12988# C[101] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2685 VSS a_12416_18747# a_12389_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2686 VDD a_46399_739# a_46617_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2687 a_22479_1566# a_21809_765# a_22079_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2688 a_9351_6676# a_8987_6419# a_9255_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2689 VDD a_52063_739# a_52011_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2690 a_5902_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2691 a_14800_18251# a_14034_18732# a_14704_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2692 a_16668_13071# a_16670_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2693 VDD a_50550_13071# a_51475_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2694 VSS a_4864_18747# a_4837_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2695 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2696 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2697 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2698 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2699 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2700 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2701 VSS a_35452_13071# a_36377_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2702 VSS C[91] a_8651_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2703 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2704 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_36138_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2705 a_15147_14292# a_14788_14127# a_14786_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2706 a_15802_928# a_14933_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2707 VSS a_54665_1566# a_54667_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2708 a_1073_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2709 a_1703_6676# a_3323_6419# a_3137_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2710 a_2961_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2711 a_27996_13071# a_27998_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2712 a_10914_13071# a_12534_13134# a_12348_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2713 a_39228_13071# a_38734_12988# a_38779_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2714 a_16913_510# a_16145_765# a_14933_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2715 a_47017_1566# a_48235_765# a_48478_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2716 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2717 a_12802_13071# a_14196_12988# a_14236_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2718 a_39914_5455# a_39555_5620# a_39553_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2719 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2720 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2721 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_56076_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2722 a_33676_19307# a_33674_18251# a_33987_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2723 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2724 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2725 a_7595_14292# a_7236_14127# a_7234_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2726 a_2160_5455# a_1801_5620# a_1799_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2727 a_52779_510# a_52011_765# a_50793_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2728 a_12816_18251# a_12198_18706# a_12416_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2729 a_35564_19307# a_35562_18251# a_35875_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2730 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_54422_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2731 VSS a_27525_739# a_27473_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2732 a_42234_928# a_41359_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2733 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2734 VSS C[27] a_8422_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2735 VDD a_21632_18706# a_21580_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2736 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2737 a_35548_13071# a_35550_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2738 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2739 a_14800_18251# a_14086_18706# a_14704_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2740 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_32362_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2741 a_37667_5620# a_37301_6419# a_35681_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2742 a_13920_928# a_13045_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2743 VDD a_10914_13071# a_11839_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2744 a_18093_14292# a_18006_14194# a_18011_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2745 a_980_12988# C[96] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2746 a_19981_14292# a_19894_14194# a_19899_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2747 a_12009_12994# a_11839_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2748 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2749 a_4686_6503# a_4516_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2750 VDD C[78] a_33189_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2751 a_26353_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2752 a_9040_18251# a_8422_18706# a_8640_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2753 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2754 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2755 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2756 a_565_18708# a_1209_6509# a_1249_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2757 a_9367_510# a_8651_739# a_7381_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2758 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2759 a_46872_14127# a_46280_12988# a_44892_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2760 a_50779_6676# a_50285_6509# a_50330_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2761 VSS C[83] a_23749_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2762 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2763 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2764 VDD a_6534_18706# a_6752_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2765 a_8233_12994# a_8063_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2766 VDD a_40512_18706# a_40460_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2767 VSS a_48772_18251# a_48774_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2768 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2769 VDD C[80] a_29413_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2770 a_7479_510# a_7477_1566# a_7790_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2771 a_38861_14292# a_38774_14194# a_38779_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2772 a_54326_13071# a_54058_13134# a_53877_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2773 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2774 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2775 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2776 VSS a_56324_18251# a_56326_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2777 a_46280_12988# C[120] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2778 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2779 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_11371_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2780 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2781 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_6689_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2782 a_44525_14292# a_44438_14194# a_44443_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2783 a_38458_928# a_37583_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2784 VDD a_57727_739# a_57675_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2785 a_3097_6509# C[33] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2786 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_46636_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2787 a_14933_1566# a_16197_739# a_16388_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2788 a_9040_18251# a_8370_18732# a_8640_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2789 a_57689_18006# a_57716_18747# a_57701_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2790 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2791 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2792 a_32794_928# a_31919_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2793 a_56553_1566# a_55787_765# a_56457_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2794 a_54749_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2795 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2796 a_50891_510# a_50889_1566# a_51202_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2797 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_3819_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2798 VSS C[71] a_46399_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2799 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2800 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_22922_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2801 a_9353_5620# a_8987_6419# a_7367_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2802 a_60102_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2803 VSS a_25242_928# a_25192_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2804 VDD a_37569_6676# a_38494_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2805 a_54978_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2806 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2807 a_6873_6509# C[35] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2808 VDD C[93] a_4875_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2809 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2810 VDD a_4251_18953# a_4201_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2811 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2812 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2813 a_11143_6676# a_10875_6419# a_10694_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2814 a_24465_510# a_23749_739# a_22479_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2815 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2816 a_14196_12988# C[103] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2817 a_60331_510# a_59615_739# a_58345_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2818 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2819 a_56310_13071# a_55946_13134# a_56214_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2820 a_47101_5620# a_46509_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2821 VSS a_870_18706# a_818_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2822 a_7381_1566# a_8599_765# a_8842_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2823 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2824 a_21971_6509# C[43] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2825 a_43345_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2826 a_13225_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2827 a_12238_6503# a_12068_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2828 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2829 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2830 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2831 a_50285_6509# C[58] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2832 VSS a_8640_18747# a_8613_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2833 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2834 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_3142_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2835 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2836 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2837 VSS a_53951_739# a_53899_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2838 VSS a_10757_1000# a_10730_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2839 a_51236_5455# a_50877_5620# a_50875_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2840 a_48662_13071# a_48168_12988# a_48213_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2841 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2842 VSS a_50550_13071# a_51475_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2843 a_54555_6676# a_56175_6419# a_55989_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2844 a_30245_14292# a_29886_14127# a_29884_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2845 a_6737_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2846 a_14422_13134# a_14196_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2847 a_54326_13071# a_53832_12988# a_53877_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2848 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2849 a_20362_18251# a_19744_18706# a_19962_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2850 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_40749_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2851 a_48758_13071# a_48168_12988# a_48662_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2852 a_22346_18251# a_21632_18706# a_22250_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2853 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2854 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2855 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2856 a_60315_6676# a_59951_6419# a_60219_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2857 a_4480_928# a_3605_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2858 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2859 VSS a_46170_18706# a_46118_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2860 a_49003_510# a_48287_739# a_47017_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2861 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2862 VDD a_25408_18706# a_25356_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2863 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2864 a_50646_13071# a_50648_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2865 VDD a_14690_13071# a_15615_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2866 a_48987_6676# a_48623_6419# a_48891_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2867 a_57918_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2868 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2869 a_22479_1566# a_23697_765# a_23940_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2870 a_44906_18251# a_46170_18706# a_46361_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2871 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2872 VSS a_10914_13071# a_11839_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2873 VDD a_13920_928# a_13870_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2874 a_37679_1566# a_36965_739# a_37583_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2875 a_48774_19307# a_48058_18706# a_46788_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2876 a_56555_510# a_56553_1566# a_56866_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2877 a_37168_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2878 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2879 a_41226_18251# a_40512_18706# a_41130_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2880 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2881 a_12009_12994# a_11839_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2882 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2883 a_20362_18251# a_19692_18732# a_19962_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2884 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2885 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2886 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2887 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2888 a_59725_6509# C[63] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2889 a_13454_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2890 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2891 VDD C[18] a_25408_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2892 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2893 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2894 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2895 a_16682_18251# a_15916_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2896 a_10465_14292# a_10460_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2897 a_52071_14292# a_51984_14194# a_51989_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2898 a_45121_6676# a_46735_6419# a_46549_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2899 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2900 a_8233_12994# a_8063_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2901 a_13127_6676# a_13129_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2902 VDD C[15] a_31072_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2903 VSS a_1584_18251# a_1586_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2904 VSS a_51668_928# a_51618_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2905 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2906 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2907 a_14651_6419# a_14425_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2908 a_1061_18006# a_1088_18747# a_1073_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2909 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2910 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2911 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2912 a_44906_18251# a_46118_18732# a_46361_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2913 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2914 VSS a_53327_18953# a_53277_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2915 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2916 a_1025_14292# a_1020_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2917 a_2913_14292# a_2908_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2918 VSS a_37569_6676# a_38494_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2919 a_55949_6509# C[61] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2920 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2921 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2922 VDD C[67] a_53951_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2923 a_16670_14127# a_16304_13134# a_14690_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2924 a_57608_12988# C[126] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2925 a_3703_510# a_2935_765# a_1717_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2926 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_7595_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2927 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2928 a_35562_18251# a_34796_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2929 a_56228_18251# a_57446_18732# a_57689_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2930 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2931 a_10875_6419# a_10649_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2932 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18093_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2933 a_23630_12988# C[108] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2934 VDD a_8027_18953# a_7977_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2935 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2936 VDD a_10875_6419# a_10689_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2937 VDD a_9915_18953# a_9865_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2938 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2939 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2940 a_12238_6503# a_12068_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2941 a_27728_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2942 a_1570_13071# a_1206_13134# a_1474_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2943 a_9365_1566# a_8651_739# a_9269_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2944 VSS C[84] a_21861_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2945 a_60219_6676# a_59563_765# a_59833_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2946 a_5591_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2947 a_12389_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2948 VSS a_31290_18747# a_31263_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2949 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_25645_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2950 VSS a_13691_18953# a_13641_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2951 a_35550_14127# a_35184_13134# a_33564_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2952 a_57834_13134# a_57608_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2953 a_20164_1811# a_20191_1000# a_20176_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2954 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2955 a_33674_18251# a_32908_18732# a_33578_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2956 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2957 a_60317_5620# a_59951_6419# a_58331_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2958 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_55994_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2959 a_41214_14127# a_40848_13134# a_39228_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2960 a_22236_13071# a_23856_13134# a_23670_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2961 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2962 a_53556_928# a_52681_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2963 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_36973_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2964 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_38861_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2965 a_48989_5620# a_48623_6419# a_47003_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2966 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2967 a_56553_1566# a_55787_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2968 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2969 VDD a_24085_6419# a_23899_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2970 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2971 a_48905_1566# a_50123_765# a_50366_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2972 a_24138_18251# a_23520_18706# a_23738_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2973 a_29788_13071# a_31408_13134# a_31222_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2974 a_29520_13134# a_29294_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2975 VDD a_58331_6676# a_59256_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2976 a_59951_6419# a_59725_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2977 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2978 a_26122_18251# a_25408_18706# a_26026_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2979 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_44525_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2980 a_39326_14127# a_38734_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2981 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2982 a_58214_19307# a_57446_18732# a_56228_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2983 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2984 VDD a_22236_13071# a_23161_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2985 a_1717_1566# a_2987_739# a_3178_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2986 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2987 a_31676_13071# a_33070_12988# a_33110_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2988 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2989 VDD a_21632_18706# a_21850_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2990 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2991 a_44990_14127# a_44398_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2992 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2993 a_27680_5455# a_27675_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2994 VDD a_29788_13071# a_30713_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2995 a_54653_5620# a_54061_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2996 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2997 VSS a_57498_18706# a_57446_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2998 a_16897_6676# a_16899_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2999 VSS a_14690_13071# a_15615_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3000 a_18421_6419# a_18195_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3001 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3002 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3003 a_50793_1566# a_50123_765# a_50393_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3004 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3005 VDD a_16197_739# a_16415_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3006 VSS a_31519_1000# a_31492_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3007 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3008 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_26108_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3009 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3010 a_29604_1811# a_29631_1000# a_29616_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3011 VSS a_52063_739# a_52011_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3012 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3013 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_46554_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3014 a_52765_5620# a_52173_6509# a_50779_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3015 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3016 a_12914_19307# a_12912_18251# a_13225_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3017 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_31772_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3018 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3019 a_14933_1566# a_16145_765# a_16388_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3020 VDD a_38458_928# a_38408_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3021 VDD a_60219_6676# a_61144_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3022 VSS C[1] a_57498_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3023 a_57735_14292# a_57648_14194# a_57653_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3024 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3025 a_40346_928# a_39471_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3026 VDD a_48891_6676# a_49816_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3027 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3028 a_18558_14127# a_17966_12988# a_16572_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3029 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3030 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_44988_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3031 a_2868_12988# C[97] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3032 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3033 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3034 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3035 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_60676_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3036 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3037 a_12032_928# a_11157_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3038 a_58441_1566# a_57727_739# a_58345_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3039 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3040 a_54667_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3041 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3042 a_39338_18251# a_38572_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3043 VSS a_28010_18251# a_28012_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3044 a_27998_14127# a_27632_13134# a_26012_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3045 a_475_18953# a_565_18708# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3046 a_33564_13071# a_33296_13134# a_33115_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3047 a_37583_1566# a_36965_739# a_37183_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3048 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3049 a_5346_13071# a_4982_13134# a_5250_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3050 a_44672_5455# a_44667_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3051 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3052 a_29339_14292# a_29334_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3053 a_37438_14127# a_36846_12988# a_35452_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3054 a_26435_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3055 a_34958_12988# C[114] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3056 VSS a_3205_1000# a_3178_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3057 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3058 a_21237_18953# a_20362_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3059 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3060 a_1206_13134# a_980_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3061 a_35039_18006# a_35066_18747# a_35051_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3062 a_20577_6676# a_20083_6509# a_20128_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3063 a_35413_6419# a_35187_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3064 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_9351_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3065 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3066 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3067 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3068 a_36927_18006# a_36954_18747# a_36939_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3069 a_43102_14127# a_42510_12988# a_41116_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3070 a_39457_6676# a_38963_6509# a_39008_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3071 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3072 a_32099_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3073 a_44990_14127# a_44398_12988# a_43004_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3074 VDD a_33189_739# a_33407_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3075 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3076 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3077 a_33987_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3078 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3079 a_15015_6676# a_14651_6419# a_14919_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3080 a_59990_13071# a_59334_18732# a_59604_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3081 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3082 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3083 VSS a_58331_6676# a_59256_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3084 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3085 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_52071_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3086 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3087 VDD a_27525_739# a_27473_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3088 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_52763_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3089 a_47663_18953# a_46788_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3090 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3091 a_33296_13134# a_33070_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3092 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_16434_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3093 a_3474_19307# a_2706_18732# a_1488_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3094 a_40117_18953# a_39242_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3095 a_54424_14127# a_53832_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3096 VDD a_31637_6419# a_31451_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3097 a_50891_510# a_50175_739# a_48905_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3098 a_26351_1566# a_25585_765# a_26255_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3099 a_49001_1566# a_48287_739# a_48905_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3100 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3101 VDD a_59722_13134# a_59536_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3102 a_44328_6503# a_44158_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3103 a_20689_510# a_20687_1566# a_21000_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3104 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3105 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3106 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3107 a_40848_13134# a_40622_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3108 a_29018_928# a_28143_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3109 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3110 VSS a_22236_13071# a_23161_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3111 a_60088_14127# a_59496_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3112 VSS a_2758_18706# a_2706_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3113 a_24776_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3114 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3115 a_37156_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3116 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3117 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3118 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3119 a_27900_13071# a_27406_12988# a_27451_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3120 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3121 a_48261_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3122 VSS a_29788_13071# a_30713_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3123 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3124 a_16899_5620# a_16307_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3125 VSS a_60219_6676# a_61144_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3126 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3127 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3128 VSS C[26] a_10310_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3129 a_22348_19307# a_22346_18251# a_22659_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3130 a_13143_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3131 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3132 a_22332_13071# a_22334_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3133 a_26108_13071# a_25518_12988# a_26012_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3134 a_27996_13071# a_27406_12988# a_27900_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3135 a_30017_6676# a_29523_6509# a_29568_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3136 a_55813_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3137 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3138 a_20083_6509# C[42] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3139 VSS a_48891_6676# a_49816_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3140 VDD a_4875_739# a_5093_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3141 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3142 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3143 VSS C[31] a_870_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3144 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3145 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3146 a_21034_5455# a_20675_5620# a_20673_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3147 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3148 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3149 VSS C[30] a_2758_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3150 VSS a_56057_1000# a_56030_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3151 a_39324_13071# a_38734_12988# a_39228_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3152 a_18460_13071# a_18192_13134# a_18011_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3153 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3154 a_16911_1566# a_16145_765# a_16815_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3155 VSS a_32015_1566# a_32017_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3156 a_3224_5455# a_3137_5687# a_3142_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3157 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3158 a_41212_13071# a_41214_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3159 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_60086_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3160 VDD a_3323_6419# a_3137_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3161 a_30113_6676# a_29749_6419# a_30017_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3162 a_26012_13071# a_25744_13134# a_25563_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3163 a_14933_1566# a_14263_765# a_14533_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3164 VDD a_44517_739# a_44465_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3165 a_18572_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3166 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_33426_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3167 VSS a_52281_1000# a_52254_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3168 a_18689_6676# a_20083_6509# a_20123_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3169 a_18785_6676# a_18421_6419# a_18689_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3170 a_37569_6676# a_38963_6509# a_39003_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3171 a_43343_1566# a_42577_765# a_43247_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3172 a_54436_18251# a_53670_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3173 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3174 a_27716_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3175 VDD a_8422_18706# a_8370_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3176 VDD a_59386_18706# a_59604_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3177 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3178 a_15017_5620# a_14651_6419# a_13031_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3179 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3180 a_16586_18251# a_17804_18732# a_18047_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3181 a_6918_5455# a_6913_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3182 VSS a_25013_18953# a_24963_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3183 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3184 a_37340_13071# a_37072_13134# a_36891_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3185 VSS a_26901_18953# a_26851_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3186 a_26353_510# a_26351_1566# a_26664_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3187 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3188 a_12816_18251# a_12146_18732# a_12416_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3189 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3190 a_29294_12988# C[111] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3191 VDD a_59220_928# a_59170_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3192 a_41768_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3193 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3194 a_52536_14127# a_51944_12988# a_50550_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3195 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3196 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3197 VSS a_16197_739# a_16145_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3198 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3199 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3200 a_44892_13071# a_44624_13134# a_44443_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3201 a_48098_6503# a_47928_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3202 VSS a_32565_18953# a_32515_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3203 a_50137_18006# a_50164_18747# a_50149_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3204 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_49119_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3205 a_29523_6509# C[47] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3206 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3207 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3208 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3209 a_37452_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3210 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_59541_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3211 a_33891_5620# a_33299_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3212 a_43345_510# a_42577_765# a_41359_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3213 a_52548_18251# a_51782_18732# a_52452_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3214 a_3376_18251# a_2706_18732# a_2976_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3215 a_8842_1811# a_8869_1000# a_8854_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3216 a_50330_5455# a_50325_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3217 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3218 a_60088_14127# a_59722_13134# a_58102_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3219 a_55444_928# a_54569_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3220 a_35466_18251# a_36684_18732# a_36927_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3221 a_43116_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3222 a_44328_6503# a_44158_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3223 VSS a_4875_739# a_4823_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3224 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3225 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3226 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3227 a_48662_13071# a_50282_13134# a_50096_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3228 VDD a_3094_13134# a_2908_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3229 a_25747_6509# C[45] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3230 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3231 a_41345_6676# a_42965_6419# a_42779_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3232 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3233 a_43018_18251# a_44236_18732# a_44479_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3234 VDD a_58991_18953# a_58941_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3235 a_39324_13071# a_38960_13134# a_39228_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3236 a_58345_1566# a_57727_739# a_57945_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3237 VSS a_10528_18747# a_10501_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3238 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3239 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3240 a_1703_6676# a_1435_6419# a_1254_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3241 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_5112_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3242 a_28129_6676# a_29523_6509# a_29563_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3243 a_33903_1566# a_33137_765# a_33807_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3244 a_27861_6419# a_27635_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3245 VSS C[88] a_14315_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3246 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3247 a_12912_18251# a_12146_18732# a_12816_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3248 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3249 a_56175_6419# a_55949_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3250 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3251 VDD a_14919_6676# a_15844_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3252 VDD a_56175_6419# a_55989_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3253 a_8888_5455# a_8801_5687# a_8806_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3254 VDD a_53951_739# a_54169_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3255 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3256 a_2798_6503# a_2628_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3257 VDD a_49780_928# a_49730_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3258 a_35777_6676# a_35413_6419# a_35681_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3259 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3260 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3261 a_13259_14292# a_12900_14127# a_12898_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3262 a_44708_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3263 a_30031_1566# a_29361_765# a_29631_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3264 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3265 a_59589_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3266 a_26108_13071# a_26110_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3267 a_49314_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3268 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3269 a_41359_1566# a_42629_739# a_42820_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3270 a_58991_18953# a_58116_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3271 a_30115_5620# a_29749_6419# a_28129_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3272 VSS a_29184_18706# a_29132_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3273 a_5707_14292# a_5348_14127# a_5346_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3274 a_10914_13071# a_12308_12988# a_12348_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3275 VSS C[76] a_36965_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3276 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_60315_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3277 VDD a_52399_6419# a_52213_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3278 a_23354_928# a_22479_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3279 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3280 a_10928_18251# a_10310_18706# a_10528_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3281 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3282 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_52534_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3283 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3284 a_9351_6676# a_8761_6509# a_9255_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3285 a_18787_5620# a_18421_6419# a_16801_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3286 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3287 a_12912_18251# a_12198_18706# a_12816_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3288 a_16205_14292# a_16118_14194# a_16123_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3289 VSS a_2592_928# a_2542_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3290 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3291 VDD a_28129_6676# a_29054_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3292 a_31905_6676# a_33525_6419# a_33339_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3293 a_27914_18251# a_29184_18706# a_29375_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3294 a_48905_1566# a_48287_739# a_48505_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3295 a_44988_13071# a_44990_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3296 a_60086_13071# a_59496_12988# a_59990_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3297 VDD a_6763_739# a_6711_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3298 a_7152_18251# a_6534_18706# a_6752_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3299 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3300 a_9136_18251# a_8422_18706# a_9040_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3301 a_42739_6509# C[54] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3302 a_46735_6419# a_46509_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3303 VDD a_2758_18706# a_2976_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3304 VDD a_4646_18706# a_4864_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3305 VDD C[21] a_19744_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3306 VSS a_46884_18251# a_46886_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3307 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3308 a_6345_12994# a_6175_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3309 a_48098_6503# a_47928_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3310 VSS a_9365_1566# a_9367_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3311 a_35085_14292# a_34998_14194# a_35003_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3312 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3313 a_36973_14292# a_36886_14194# a_36891_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3314 a_52438_13071# a_52170_13134# a_51989_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3315 a_7463_6676# a_7099_6419# a_7367_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3316 VDD a_50175_739# a_50123_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3317 a_39471_1566# a_38801_765# a_39071_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3318 a_20591_1566# a_19921_765# a_20191_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3319 a_4014_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3320 a_48249_18006# a_48276_18747# a_48261_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3321 a_30906_928# a_30031_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3322 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3323 a_48213_14292# a_48208_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3324 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3325 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_2913_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3326 a_14518_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3327 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_4801_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3328 a_55801_18006# a_55828_18747# a_55813_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3329 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3330 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_34250_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3331 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3332 a_7152_18251# a_6482_18732# a_6752_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3333 a_39569_510# a_38853_739# a_37583_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3334 VSS a_52777_1566# a_52779_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3335 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1931_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3336 VDD a_11803_18953# a_11753_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3337 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3338 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3339 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3340 a_38026_5455# a_37667_5620# a_37665_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3341 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3342 a_50564_18251# a_51782_18732# a_52025_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3343 VDD a_18689_6676# a_19614_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3344 a_40346_928# a_39471_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3345 VDD a_2363_18953# a_2313_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3346 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3347 a_35779_5620# a_35413_6419# a_33793_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3348 a_48478_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3349 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3350 a_12308_12988# C[102] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3351 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_30474_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3352 a_43343_1566# a_42577_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3353 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3354 a_54422_13071# a_54058_13134# a_54326_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3355 a_54555_6676# a_54287_6419# a_54106_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3356 a_28239_1566# a_27525_739# a_28143_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3357 VSS a_14919_6676# a_15844_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3358 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3359 a_2798_6503# a_2628_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3360 VDD C[79] a_31301_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3361 a_24465_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3362 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3363 VSS a_6752_18747# a_6725_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3364 a_55650_6503# a_55480_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3365 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3366 a_9124_14127# a_8758_13134# a_7138_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3367 a_14470_5455# a_14465_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3368 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_31309_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3369 a_46774_13071# a_46280_12988# a_46325_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3370 a_41443_5620# a_40851_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3371 a_9353_5620# a_8761_6509# a_7367_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3372 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3373 a_18460_13071# a_19854_12988# a_19894_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3374 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3375 a_26901_18953# a_26026_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3376 a_4849_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3377 a_12802_13071# a_14422_13134# a_14236_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3378 a_12534_13134# a_12308_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3379 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3380 a_58443_510# a_57675_765# a_56457_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3381 a_5591_510# a_5589_1566# a_5902_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3382 a_31774_14127# a_31182_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3383 a_46870_13071# a_46280_12988# a_46774_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3384 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3385 a_4251_18953# a_3376_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3386 a_33662_14127# a_33070_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3387 VDD a_37072_13134# a_36886_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3388 a_37583_1566# a_38801_765# a_39044_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3389 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3390 a_20458_18251# a_19744_18706# a_20362_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3391 VSS a_28129_6676# a_29054_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3392 a_19578_928# a_18703_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3393 VDD a_55839_739# a_55787_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3394 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3395 a_1209_6509# C[32] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3396 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_33344_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3397 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3398 VDD a_12802_13071# a_13727_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3399 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3400 a_9712_5455# a_9353_5620# a_9351_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3401 a_30906_928# a_30031_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3402 a_54665_1566# a_53899_765# a_54569_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3403 a_7138_13071# a_8532_12988# a_8572_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3404 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3405 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_39914_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3406 a_7465_5620# a_7099_6419# a_5479_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3407 a_18799_1566# a_18085_739# a_18703_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3408 a_14126_6503# a_13956_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3409 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_2160_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3410 a_46886_19307# a_46170_18706# a_44906_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3411 a_60086_13071# a_60088_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3412 VDD a_35681_6676# a_36606_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3413 a_18288_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3414 a_4985_6509# C[34] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3415 a_56539_6676# a_56175_6419# a_56443_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3416 VDD C[94] a_2987_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3417 a_53124_5455# a_52765_5620# a_52763_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3418 a_5936_5455# a_5577_5620# a_5575_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3419 a_45231_1566# a_44517_739# a_45135_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3420 a_54340_18251# a_55610_18706# a_55801_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3421 VDD C[19] a_23520_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3422 a_58214_19307# a_57498_18706# a_56228_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3423 a_41457_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3424 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3425 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3426 a_38963_6509# C[52] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3427 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3428 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3429 a_50183_14292# a_50096_14194# a_50101_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3430 a_6345_12994# a_6175_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3431 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3432 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3433 a_48168_12988# C[121] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3434 a_56457_1566# a_57727_739# a_57918_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3435 a_56539_6676# a_56541_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3436 a_47113_1566# a_46347_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3437 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3438 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3439 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3440 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3441 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3442 VSS a_18689_6676# a_19614_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3443 a_52667_6676# a_54287_6419# a_54101_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3444 a_26122_18251# a_25356_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3445 a_50511_6419# a_50285_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3446 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3447 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_5707_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3448 VSS a_60329_1566# a_60331_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3449 a_33674_18251# a_32908_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3450 a_54340_18251# a_55558_18732# a_55801_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3451 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3452 a_2592_928# a_1717_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3453 a_58443_510# a_58441_1566# a_58754_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3454 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3455 a_21742_12988# C[107] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3456 a_60315_6676# a_59725_6509# a_60219_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3457 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3458 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_16205_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3459 a_15031_510# a_14315_739# a_13045_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3460 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3461 a_48394_13134# a_48168_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3462 a_31774_14127# a_31182_12988# a_29788_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3463 a_58198_13071# a_57834_13134# a_58102_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3464 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3465 a_24234_18251# a_23468_18732# a_24138_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3466 VDD a_7367_6676# a_8292_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3467 a_55650_6503# a_55480_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3468 VDD a_14315_739# a_14263_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3469 a_20771_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3470 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_23757_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3471 a_18558_14127# a_17966_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3472 VSS a_22079_1000# a_22052_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3473 a_45002_18251# a_44236_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3474 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3475 a_14802_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3476 a_33662_14127# a_33296_13134# a_31676_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3477 a_55946_13134# a_55720_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3478 a_33905_510# a_33137_765# a_31919_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3479 a_13141_1566# a_12375_765# a_13045_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3480 a_35791_1566# a_35077_739# a_35695_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3481 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3482 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3483 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3484 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3485 a_31786_18251# a_31020_18732# a_31690_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3486 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3487 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3488 VSS a_44517_739# a_44465_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3489 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_55012_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3490 VSS a_41226_18251# a_41228_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3491 a_20348_13071# a_21968_13134# a_21782_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3492 a_20080_13134# a_19854_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3493 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3494 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35085_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3495 VDD a_29018_928# a_28968_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3496 a_11566_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3497 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3498 a_49003_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3499 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3500 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3501 VDD C[91] a_8651_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3502 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3503 a_58788_5455# a_58429_5620# a_58427_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3504 a_8027_18953# a_7152_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3505 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_42637_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3506 a_37438_14127# a_36846_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3507 a_56326_19307# a_55558_18732# a_54340_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3508 VDD a_20348_13071# a_21273_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3509 a_20128_5455# a_20123_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3510 a_29788_13071# a_31182_12988# a_31222_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3511 a_39008_5455# a_39003_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3512 VSS a_48058_18706# a_48006_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3513 a_54061_6509# C[60] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3514 VSS a_49946_18706# a_49894_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3515 a_8758_13134# a_8532_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3516 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3517 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3518 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3519 a_14126_6503# a_13956_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3520 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3521 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3522 a_50875_6676# a_50285_6509# a_50779_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3523 VSS a_35681_6676# a_36606_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3524 VSS C[74] a_40741_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3525 VDD C[68] a_52063_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3526 a_39228_13071# a_40848_13134# a_40662_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3527 a_46788_18251# a_48058_18706# a_48249_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3528 VSS a_12802_13071# a_13727_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3529 a_28143_1566# a_27525_739# a_27743_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3530 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3531 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3532 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_24220_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3533 VDD a_39228_13071# a_40153_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3534 a_38827_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3535 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3536 VSS C[6] a_48058_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3537 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3538 a_31919_1566# a_33189_739# a_33380_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3539 a_7477_1566# a_6763_739# a_7381_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3540 a_11026_19307# a_11024_18251# a_11337_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3541 a_3703_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3542 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3543 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_29884_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3544 VDD a_23749_739# a_23967_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3545 a_18570_18251# a_17804_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3546 VDD a_19578_928# a_19528_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3547 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3548 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3549 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3550 a_55847_14292# a_55760_14194# a_55765_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3551 a_14506_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3552 VSS a_42234_928# a_42184_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3553 a_60317_5620# a_59725_6509# a_58331_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3554 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_54106_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3555 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3556 a_19112_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3557 a_16670_14127# a_16078_12988# a_14690_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3558 a_41457_510# a_40741_739# a_39471_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3559 a_51668_928# a_50793_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3560 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_43100_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3561 VDD a_10310_18706# a_10258_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3562 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3563 a_9122_13071# a_9124_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3564 a_54665_1566# a_53899_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3565 a_18558_14127# a_18192_13134# a_16572_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3566 VDD a_22197_6419# a_22011_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3567 a_22098_5455# a_22011_5687# a_22016_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3568 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3569 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3570 VDD a_15802_928# a_15752_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3571 a_24124_13071# a_23856_13134# a_23675_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3572 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3573 VSS a_7367_6676# a_8292_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3574 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3575 a_37450_18251# a_36684_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3576 a_6368_928# a_5493_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3577 a_25840_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3578 VSS a_26122_18251# a_26124_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3579 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3580 a_55421_12994# a_55251_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3581 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3582 a_14323_14292# a_14236_14194# a_14241_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3583 a_18703_1566# a_18085_739# a_18303_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3584 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3585 a_3458_13071# a_3094_13134# a_3362_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3586 a_31676_13071# a_31408_13134# a_31227_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3587 a_25792_5455# a_25787_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3588 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3589 a_27487_18006# a_27514_18747# a_27499_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3590 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3591 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_46325_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3592 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3593 a_35550_14127# a_34958_12988# a_33564_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3594 a_24547_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3595 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3596 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3597 a_12537_6509# C[38] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3598 a_37438_14127# a_37072_13134# a_35452_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3599 a_16533_6419# a_16307_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3600 a_45135_1566# a_44517_739# a_44735_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3601 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3602 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3603 VSS a_45002_18251# a_45004_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3604 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3605 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3606 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_50183_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3607 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3608 a_50877_5620# a_50285_6509# a_48891_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3609 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3610 a_60331_510# a_59563_765# a_58345_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3611 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3612 VDD a_40741_739# a_40959_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3613 a_7381_1566# a_8651_739# a_8842_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3614 a_45775_18953# a_44906_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3615 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3616 a_31408_13134# a_31182_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3617 VDD a_36570_928# a_36520_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3618 a_39471_1566# a_40689_765# a_40932_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3619 a_1586_19307# a_818_18732# a_565_18708# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3620 a_42510_12988# C[118] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3621 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3622 a_52536_14127# a_51944_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3623 VDD a_57834_13134# a_57648_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3624 a_21466_928# a_20591_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3625 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3626 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3627 a_36104_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3628 a_18460_13071# a_17966_12988# a_18011_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3629 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3630 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3631 VSS a_20348_13071# a_21273_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3632 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_23986_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3633 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_59770_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3634 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3635 a_10144_928# a_9269_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3636 a_56553_1566# a_55839_739# a_56457_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3637 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3638 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3639 a_24124_13071# a_23630_12988# a_23675_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3640 a_18556_13071# a_17966_12988# a_18460_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3641 a_18276_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3642 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3643 a_46373_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3644 a_26012_13071# a_25518_12988# a_25563_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3645 a_42832_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3646 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3647 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3648 a_49003_510# a_48235_765# a_47017_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3649 a_20460_19307# a_20458_18251# a_20771_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3650 a_35695_1566# a_35077_739# a_35295_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3651 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3652 a_20444_13071# a_20446_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3653 a_42784_5455# a_42779_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3654 a_53925_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3655 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3656 a_37340_13071# a_36846_12988# a_36891_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3657 VSS a_59615_739# a_59563_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3658 VSS a_1317_1000# a_1290_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3659 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3660 VSS a_39228_13071# a_40153_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3661 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3662 a_33525_6419# a_33299_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3663 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_7463_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3664 a_37569_6676# a_37075_6509# a_37120_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3665 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3666 a_31772_13071# a_31774_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3667 a_37436_13071# a_36846_12988# a_37340_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3668 VSS RESET a_27668_9428# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3669 VDD a_31301_739# a_31519_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3670 a_58345_1566# a_59615_739# a_59806_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3671 a_44892_13071# a_44398_12988# a_44443_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3672 a_16572_13071# a_16304_13134# a_16123_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3673 a_11024_18251# a_10310_18706# a_10928_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3674 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3675 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3676 VDD C[64] a_59615_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3677 a_43100_13071# a_42510_12988# a_43004_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3678 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3679 a_44988_13071# a_44398_12988# a_44892_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3680 VSS C[75] a_38853_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3681 a_19935_18006# a_19962_18747# a_19947_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3682 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3683 VDD a_25637_739# a_25585_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3684 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3685 a_16684_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3686 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3687 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3688 a_24463_1566# a_23697_765# a_24367_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3689 a_37681_510# a_37679_1566# a_37992_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3690 VDD a_6534_18706# a_6482_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3691 a_52548_18251# a_51782_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3692 VDD a_57498_18706# a_57716_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3693 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3694 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3695 a_59197_12994# a_59027_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3696 a_14704_18251# a_15916_18732# a_16159_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3697 a_35452_13071# a_35184_13134# a_35003_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3698 VSS a_23125_18953# a_23075_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3699 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3700 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3701 a_10928_18251# a_10258_18732# a_10528_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3702 a_41130_18251# a_42400_18706# a_42591_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3703 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3704 a_50648_14127# a_50056_12988# a_48662_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3705 a_27406_12988# C[110] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3706 a_26337_6676# a_25973_6419# a_26241_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3707 a_22888_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3708 a_45004_19307# a_44288_18706# a_43018_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3709 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3710 a_55421_12994# a_55251_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3711 a_47017_1566# a_48287_739# a_48478_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3712 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3713 a_7381_1566# a_6763_739# a_6981_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3714 a_35268_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3715 VSS a_30677_18953# a_30627_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3716 a_38815_18006# a_38842_18747# a_38827_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3717 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_47231_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3718 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3719 a_35564_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3720 a_52536_14127# a_52170_13134# a_50550_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3721 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_57653_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3722 a_30113_6676# a_29523_6509# a_30017_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3723 a_41345_6676# a_41077_6419# a_40896_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3724 a_15029_1566# a_14315_739# a_14933_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3725 a_1488_18251# a_818_18732# a_1088_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3726 a_3687_6676# a_3689_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3727 a_11255_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3728 VDD C[28] a_6534_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3729 a_5211_6419# a_4985_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3730 VSS a_57332_928# a_57282_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3731 a_41228_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3732 VSS a_60100_18251# a_60102_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3733 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3734 a_9255_6676# a_8761_6509# a_8806_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3735 a_33578_18251# a_34796_18732# a_35039_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3736 VDD a_49551_18953# a_49501_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3737 a_37075_6509# C[51] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3738 VDD a_2987_739# a_3205_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3739 VSS a_42005_18953# a_41955_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3740 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3741 a_42440_6503# a_42270_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3742 a_56555_510# a_55839_739# a_54569_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3743 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3744 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3745 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3746 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3747 a_27632_13134# a_27406_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3748 VSS a_54169_1000# a_54142_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3749 VDD a_1206_13134# a_1020_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3750 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3751 a_22465_6676# a_24085_6419# a_23899_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3752 a_9367_510# a_8599_765# a_7381_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3753 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3754 a_46554_5455# a_46549_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3755 VSS a_30127_1566# a_30129_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3756 a_12900_14127# a_12534_13134# a_10914_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3757 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3758 VDD a_1435_6419# a_1249_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3759 a_28241_510# a_28239_1566# a_28552_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3760 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3761 a_11024_18251# a_10258_18732# a_10928_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3762 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3763 VDD a_42629_739# a_42577_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3764 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_14323_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3765 a_29788_13071# a_29294_12988# a_29339_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3766 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3767 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3768 a_16897_6676# a_16533_6419# a_16801_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3769 a_41455_1566# a_40689_765# a_41359_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3770 a_29900_19307# a_29132_18732# a_27914_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3771 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3772 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3773 a_25828_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3774 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3775 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3776 a_14788_14127# a_14196_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3777 a_31905_6676# a_31637_6419# a_31456_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3778 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3779 a_24465_510# a_24463_1566# a_24776_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3780 VDD a_57332_928# a_57282_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3781 a_57103_18953# a_56228_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3782 a_9026_13071# a_10420_12988# a_10460_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3783 VSS a_27296_18706# a_27244_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3784 a_3819_14292# a_3460_14127# a_3458_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3785 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3786 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3787 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3788 a_7099_6419# a_6873_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3789 a_33000_6503# a_32830_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3790 a_24465_510# a_23697_765# a_22479_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3791 a_18801_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3792 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3793 a_54569_1566# a_55787_765# a_56030_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3794 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3795 a_52534_13071# a_51944_12988# a_52438_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3796 a_28586_5455# a_28227_5620# a_28225_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3797 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3798 a_26026_18251# a_27296_18706# a_27487_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3799 a_5250_13071# a_6644_12988# a_6684_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3800 a_29900_19307# a_29184_18706# a_27914_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3801 a_26339_5620# a_25973_6419# a_24353_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3802 a_5264_18251# a_4646_18706# a_4864_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3803 VSS sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3804 a_43329_6676# a_43331_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3805 a_33903_1566# a_33137_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3806 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3807 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3808 a_7248_18251# a_6534_18706# a_7152_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3809 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3810 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3811 a_23859_6509# C[44] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3812 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3813 VSS C[17] a_27296_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3814 a_27533_14292# a_27446_14194# a_27451_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3815 a_39457_6676# a_41077_6419# a_40891_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3816 VDD C[84] a_21861_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3817 VDD a_8651_739# a_8869_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3818 VDD a_870_18706# a_1088_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3819 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3820 a_37354_18251# a_38624_18706# a_38815_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3821 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3822 a_4457_12994# a_4287_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3823 a_56457_1566# a_55839_739# a_56057_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3824 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_3224_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3825 a_47115_510# a_46347_765# a_45135_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3826 a_32015_1566# a_31249_765# a_31919_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3827 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_14786_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3828 a_33197_14292# a_33110_14194# a_33115_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3829 a_50550_13071# a_50282_13134# a_50101_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3830 a_25973_6419# a_25747_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3831 a_45233_510# a_45231_1566# a_45544_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3832 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3833 a_46361_18006# a_46388_18747# a_46373_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3834 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3835 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3836 a_7367_6676# a_8761_6509# a_8801_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3837 VSS a_32794_928# a_32744_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3838 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3839 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3840 a_46325_14292# a_46320_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3841 a_32003_5620# a_31411_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3842 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3843 a_59197_12994# a_59027_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3844 a_54287_6419# a_54061_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3845 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3846 VDD a_47892_928# a_47842_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3847 VDD a_52063_739# a_52281_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3848 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3849 a_52025_18006# a_52052_18747# a_52037_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3850 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3851 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3852 a_33889_6676# a_33525_6419# a_33793_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3853 a_39340_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3854 a_53913_18006# a_53940_18747# a_53925_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3855 a_42440_6503# a_42270_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3856 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3857 a_50662_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3858 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3859 a_47426_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3860 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3861 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3862 a_22479_1566# a_23749_739# a_23940_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3863 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3864 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3865 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3866 a_50366_1811# a_50393_1000# a_50378_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3867 a_48676_18251# a_49894_18732# a_50137_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3868 a_30115_5620# a_29523_6509# a_28129_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3869 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_23904_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3870 VSS C[86] a_18085_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3871 a_46870_13071# a_46506_13134# a_46774_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3872 VDD a_50511_6419# a_50325_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3873 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3874 a_21466_928# a_20591_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3875 a_7463_6676# a_6873_6509# a_7367_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3876 a_44627_6509# C[55] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3877 VSS C[67] a_53951_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3878 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3879 a_14788_14127# a_14196_12988# a_12802_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3880 a_16899_5620# a_16533_6419# a_14919_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3881 a_24463_1566# a_23697_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3882 a_35793_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3883 a_45578_5455# a_45219_5620# a_45217_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3884 VDD a_26241_6676# a_27166_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3885 a_30017_6676# a_31637_6419# a_31451_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3886 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3887 a_32017_510# a_31301_739# a_30031_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3888 a_47017_1566# a_46399_739# a_46617_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3889 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3890 VDD a_4875_739# a_4823_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3891 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3892 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3893 a_60219_6676# a_59725_6509# a_59770_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3894 a_17461_18953# a_16586_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3895 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3896 a_3701_1566# a_2935_765# a_3605_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3897 a_9915_18953# a_9040_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3898 VSS a_9136_18251# a_9138_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3899 a_8532_12988# C[100] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3900 a_22563_5620# a_21971_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3901 VDD C[75] a_38853_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3902 a_24222_14127# a_23630_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3903 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3904 a_50891_510# a_50123_765# a_48905_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3905 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3906 a_1061_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3907 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3908 VSS a_7477_1566# a_7479_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3909 a_10646_13134# a_10420_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3910 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3911 a_33000_6503# a_32830_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3912 a_42965_6419# a_42739_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3913 a_47099_6676# a_47101_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3914 a_2363_18953# a_1488_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3915 a_7561_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3916 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3917 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3918 a_29886_14127# a_29294_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3919 a_5575_6676# a_5211_6419# a_5479_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3920 a_37583_1566# a_36913_765# a_37183_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3921 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3922 VSS a_10539_739# a_10487_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3923 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3924 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3925 a_20675_5620# a_20083_6509# a_18689_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3926 a_59806_1811# a_59833_1000# a_59818_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3927 a_36341_18953# a_35466_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3928 a_39555_5620# a_38963_6509# a_37569_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3929 VSS a_50889_1566# a_50891_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3930 a_7138_13071# a_8758_13134# a_8572_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3931 VDD a_59951_6419# a_59765_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3932 a_43102_14127# a_42510_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3933 a_49003_510# a_49001_1566# a_49314_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3934 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3935 a_42005_18953# a_41130_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3936 a_25611_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3937 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3938 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3939 a_43893_18953# a_43018_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3940 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3941 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_40896_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3942 VSS a_55610_18706# a_55558_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3943 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3944 VDD a_16801_6676# a_17726_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3945 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3946 VDD a_7138_13071# a_8063_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3947 VSS a_33189_739# a_33137_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3948 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3949 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3950 a_31411_6509# C[48] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3951 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_29568_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3952 a_41455_1566# a_40689_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3953 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3954 a_52667_6676# a_52399_6419# a_52218_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3955 a_26351_1566# a_25637_739# a_26255_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3956 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3957 a_52452_18251# a_53722_18706# a_53913_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3958 VDD C[20] a_21632_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3959 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3960 a_36570_928# a_35695_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3961 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3962 a_56326_19307# a_55610_18706# a_54340_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3963 a_22577_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3964 a_12630_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3965 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3966 a_48905_1566# a_50175_739# a_50366_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3967 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3968 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3969 a_11010_13071# a_11012_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3970 a_4457_12994# a_4287_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3971 a_44491_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3972 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3973 a_48397_6509# C[57] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3974 a_59852_5455# a_59765_5687# a_59770_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3975 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3976 a_53762_6503# a_53592_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3977 a_12582_5455# a_12577_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3978 a_9269_1566# a_8599_765# a_8869_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3979 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3980 a_49348_5455# a_48989_5620# a_48987_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3981 a_24234_18251# a_23468_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3982 a_54438_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3983 VDD a_29184_18706# a_29402_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3984 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3985 VDD C[10] a_40512_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3986 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3987 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3988 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3989 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_4048_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3990 a_31786_18251# a_31020_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3991 a_52452_18251# a_53670_18732# a_53913_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3992 a_22334_14127# a_21742_12988# a_20348_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3993 VSS a_26241_6676# a_27166_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3994 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3995 a_58427_6676# a_58063_6419# a_58331_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3996 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3997 a_14690_13071# a_14422_13134# a_14241_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3998 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_31456_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3999 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_29339_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4000 a_46506_13134# a_46280_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4001 a_7824_5455# a_7465_5620# a_7463_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4002 a_52777_1566# a_52011_765# a_52681_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4003 a_22346_18251# a_21580_18732# a_22250_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4004 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4005 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4006 a_16670_14127# a_16078_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4007 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_20673_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4008 a_43114_18251# a_42348_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4009 a_12914_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4010 VSS a_31786_18251# a_31788_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4011 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4012 a_31774_14127# a_31408_13134# a_29788_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4013 a_54058_13134# a_53832_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4014 a_5577_5620# a_5211_6419# a_3591_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4015 VSS a_56553_1566# a_56555_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4016 a_16911_1566# a_16197_739# a_16815_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4017 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4018 VDD a_27668_9428# sky130_fd_sc_hd__buf_2_0/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4019 a_46004_928# a_45135_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4020 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4021 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4022 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4023 a_41214_14127# a_40622_12988# a_39228_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4024 VSS a_47892_928# a_47842_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4025 VDD C[95] a_1099_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4026 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4027 a_18460_13071# a_20080_13134# a_19894_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4028 a_12816_18251# a_14034_18732# a_14277_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4029 VDD a_28789_18953# a_28739_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4030 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_33197_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4031 a_43343_1566# a_42629_739# a_43247_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4032 a_48774_19307# a_48006_18732# a_46788_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4033 VSS a_6139_18953# a_6089_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4034 a_28789_18953# a_27914_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4035 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4036 a_20348_13071# a_21742_12988# a_21782_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4037 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4038 a_6139_18953# a_5264_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4039 a_35550_14127# a_34958_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4040 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4041 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4042 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4043 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4044 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_45349_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4045 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4046 a_54651_6676# a_54653_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4047 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4048 VSS a_16801_6676# a_17726_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4049 a_50779_6676# a_52399_6419# a_52213_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4050 a_29387_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4051 VSS C[93] a_4875_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4052 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4053 a_16352_5455# a_16347_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4054 a_47115_510# a_46399_739# a_45135_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4055 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4056 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_22332_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4057 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4058 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_9712_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4059 VSS C[92] a_6763_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4060 VSS C[7] a_46170_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4061 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4062 VDD a_5479_6676# a_6404_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4063 a_53762_6503# a_53592_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4064 VDD a_12427_739# a_12375_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4065 VSS a_7138_13071# a_8063_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4066 VSS a_20191_1000# a_20164_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4067 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4068 a_11253_1566# a_10487_765# a_11157_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4069 a_33903_1566# a_33189_739# a_33807_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4070 a_14786_13071# a_14788_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4071 a_53959_14292# a_53872_14194# a_53877_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4072 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4073 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4074 a_48891_6676# a_50285_6509# a_50325_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4075 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4076 a_58429_5620# a_58063_6419# a_56443_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4077 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_53124_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4078 a_8761_6509# C[36] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4079 VSS a_25637_739# a_25585_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4080 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_41212_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4081 a_12032_928# a_11157_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4082 VDD a_27130_928# a_27080_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4083 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4084 a_28010_18251# a_27244_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4085 a_7250_19307# a_7248_18251# a_7561_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4086 a_47115_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4087 VSS a_16682_18251# a_16684_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4088 a_7234_13071# a_7236_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4089 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4090 VDD C[92] a_6763_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4091 VSS a_18570_18251# a_18572_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4092 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4093 a_22236_13071# a_21968_13134# a_21787_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4094 a_18047_18006# a_18074_18747# a_18059_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4095 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4096 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4097 VSS a_8256_928# a_8206_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4098 a_18011_14292# a_18006_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4099 a_19899_14292# a_19894_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4100 a_37120_5455# a_37115_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4101 VSS a_24234_18251# a_24236_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4102 a_14919_6676# a_14425_6509# a_14470_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4103 a_52173_6509# C[59] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4104 VDD a_59386_18706# a_59334_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4105 a_7479_510# a_6763_739# a_5493_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4106 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4107 a_25599_18006# a_25626_18747# a_25611_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4108 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4109 a_33662_14127# a_33070_12988# a_31676_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4110 VSS a_48287_739# a_48235_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4111 a_22659_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4112 a_45135_1566# a_46347_765# a_46590_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4113 a_48676_18251# a_48006_18732# a_48276_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4114 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4115 a_9255_6676# a_10875_6419# a_10689_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4116 VSS a_37450_18251# a_37452_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4117 a_39044_1811# a_39071_1000# a_39056_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4118 a_26255_1566# a_25637_739# a_25855_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4119 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4120 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4121 a_41116_13071# a_40848_13134# a_40667_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4122 a_60317_5620# a_59725_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4123 VSS a_29631_1000# a_29604_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4124 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_8806_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4125 a_15031_510# a_15029_1566# a_15342_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4126 VSS a_43114_18251# a_43116_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4127 a_38779_14292# a_38774_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4128 a_33070_12988# C[113] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4129 a_5589_1566# a_4875_739# a_5493_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4130 a_24220_13071# a_23856_13134# a_24124_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4131 VDD a_48394_13134# a_48208_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4132 a_24085_6419# a_23859_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4133 a_5078_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4134 a_44479_18006# a_44506_18747# a_44491_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4135 a_44443_14292# a_44438_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4136 VDD a_17690_928# a_17640_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4137 VDD a_21861_739# a_22079_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4138 a_41539_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4139 a_40622_12988# C[117] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4140 a_50648_14127# a_50056_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4141 VDD a_54058_13134# a_53872_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4142 VDD a_55946_13134# a_55760_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4143 VSS a_23354_928# a_23304_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4144 a_12618_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4145 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4146 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4147 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4148 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_52218_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4149 a_17224_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4150 a_22577_510# a_21861_739# a_20591_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4151 a_11255_510# a_11253_1566# a_11566_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4152 a_16572_13071# a_16078_12988# a_16123_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4153 VDD a_44122_928# a_44072_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4154 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4155 a_55215_18953# a_54340_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4156 VDD a_20309_6419# a_20123_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4157 a_52777_1566# a_52011_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4158 VDD a_39189_6419# a_39003_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4159 a_5493_1566# a_6711_765# a_6954_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4160 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4161 a_43100_13071# a_42736_13134# a_43004_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4162 a_14425_6509# C[39] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4163 a_16668_13071# a_16078_12988# a_16572_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4164 VSS a_5479_6676# a_6404_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4165 a_23952_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4166 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4167 a_15376_5455# a_15017_5620# a_15015_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4168 a_37583_1566# a_38853_739# a_39044_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4169 VSS a_59604_18747# a_59577_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4170 a_49119_14292# a_48760_14127# a_48758_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4171 a_23904_5455# a_23899_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4172 a_16815_1566# a_16197_739# a_16415_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4173 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4174 a_57837_6509# C[62] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4175 a_35452_13071# a_34958_12988# a_35003_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4176 a_10649_6509# C[37] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4177 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4178 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4179 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4180 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4181 a_18689_6676# a_18195_6509# a_18240_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4182 a_43247_1566# a_42629_739# a_42847_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4183 a_16684_19307# a_15968_18706# a_14704_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4184 a_41116_13071# a_40622_12988# a_40667_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4185 a_29884_13071# a_29886_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4186 a_43004_13071# a_42510_12988# a_42555_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4187 a_35548_13071# a_34958_12988# a_35452_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4188 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4189 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4190 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4191 a_56214_13071# a_57834_13134# a_57648_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4192 a_12763_6419# a_12537_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4193 a_6954_1811# a_6981_1000# a_6966_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4194 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4195 a_41212_13071# a_40622_12988# a_41116_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4196 a_41077_6419# a_40851_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4197 VDD a_48058_18706# a_48276_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4198 VDD a_41077_6419# a_40891_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4199 a_58116_18251# a_57498_18706# a_57716_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4200 a_20591_1566# a_21809_765# a_22052_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4201 VDD a_34682_928# a_34632_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4202 a_59990_13071# a_59386_18706# a_59604_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4203 a_1584_18251# a_870_18706# a_1488_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4204 VDD a_475_18953# a_425_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4205 VDD a_56214_13071# a_57139_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4206 a_44720_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4207 VSS a_20687_1566# a_20689_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4208 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4209 VDD a_29749_6419# a_29563_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4210 a_31690_18251# a_32960_18706# a_33151_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4211 VDD a_4646_18706# a_4594_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4212 a_50660_18251# a_49894_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4213 a_18801_510# a_18799_1566# a_19112_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4214 a_35564_19307# a_34848_18706# a_33578_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4215 VDD a_55610_18706# a_55828_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4216 a_19854_12988# C[106] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4217 a_57309_12994# a_57139_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4218 a_34216_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4219 VSS a_21237_18953# a_21187_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4220 a_29375_18006# a_29402_18747# a_29387_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4221 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4222 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_48213_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4223 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4224 a_25518_12988# C[109] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4225 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4226 VDD a_30906_928# a_30856_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4227 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4228 a_16388_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4229 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4230 a_11253_1566# a_10487_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4231 a_31788_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4232 VSS a_50660_18251# a_50662_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4233 VSS a_52548_18251# a_52550_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4234 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4235 a_50648_14127# a_50282_13134# a_48662_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4236 a_22465_6676# a_22197_6419# a_22016_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4237 a_40944_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4238 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4239 a_24138_18251# a_25356_18732# a_25599_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4240 a_26026_18251# a_27244_18732# a_27487_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4241 a_33676_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4242 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4243 VDD a_13031_6676# a_13956_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4244 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4245 a_33807_1566# a_33189_739# a_33407_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4246 a_51989_14292# a_51984_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4247 a_18192_13134# a_17966_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4248 a_40896_5455# a_40891_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4249 a_15031_510# a_14263_765# a_13045_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4250 VDD C[29] a_4646_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4251 a_38734_12988# C[116] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4252 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4253 a_31690_18251# a_32908_18732# a_33151_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4254 VDD a_47663_18953# a_47613_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4255 a_18195_6509# C[41] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4256 a_29650_5455# a_29563_5687# a_29568_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4257 VSS a_704_928# a_654_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4258 VSS a_40117_18953# a_40067_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4259 a_29884_13071# a_29520_13134# a_29788_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4260 a_1815_510# a_1047_765# a_794_737# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4261 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_58559_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4262 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4263 a_23560_6503# a_23390_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4264 a_27130_928# a_26255_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4265 a_44398_12988# C[119] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4266 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4267 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4268 a_25744_13134# a_25518_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4269 a_31637_6419# a_31411_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4270 a_19146_5455# a_18787_5620# a_18785_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4271 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4272 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4273 a_33889_6676# a_33891_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4274 VDD a_6368_928# a_6318_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4275 a_11012_14127# a_10646_13134# a_9026_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4276 a_37072_13134# a_36846_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4277 VSS C[85] a_19973_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4278 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4279 a_38960_13134# a_38734_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4280 a_28225_6676# a_27861_6419# a_28129_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4281 VDD a_23749_739# a_23697_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4282 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_12435_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4283 a_22575_1566# a_21809_765# a_22479_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4284 a_26124_19307# a_25356_18732# a_24138_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4285 VSS a_2976_18747# a_2949_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4286 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4287 VSS a_15802_928# a_15752_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4288 a_28012_19307# a_27244_18732# a_26026_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4289 a_49551_18953# a_48676_18251# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4290 a_44624_13134# a_44398_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4291 a_35793_510# a_35791_1566# a_36104_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4292 a_39569_510# a_38801_765# a_37583_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4293 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4294 VSS a_19744_18706# a_19692_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4295 a_55801_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4296 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4297 VSS a_26351_1566# a_26353_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4298 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4299 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4300 a_5360_18251# a_4594_18732# a_5264_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4301 a_12900_14127# a_12308_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4302 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4303 a_24449_6676# a_24085_6419# a_24353_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4304 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4305 a_50550_13071# a_50056_12988# a_50101_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4306 a_39340_19307# a_38572_18732# a_37354_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4307 a_5493_1566# a_4875_739# a_5093_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4308 a_48490_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4309 a_16586_18251# a_17856_18706# a_18047_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4310 a_13141_1566# a_12427_739# a_13045_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4311 VSS a_8869_1000# a_8842_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4312 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4313 a_794_737# a_1099_739# a_1290_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4314 a_1474_13071# a_3094_13134# a_2908_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4315 a_50646_13071# a_50056_12988# a_50550_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4316 a_48442_5455# a_48437_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4317 VDD a_9026_13071# a_9951_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4318 a_24138_18251# a_25408_18706# a_25599_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4319 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4320 a_3323_6419# a_3097_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4321 VSS C[22] a_17856_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4322 a_3362_13071# a_4756_12988# a_4796_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4323 a_7367_6676# a_6873_6509# a_6918_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4324 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4325 a_28012_19307# a_27296_18706# a_26026_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4326 VSS a_38624_18706# a_38572_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4327 a_35187_6509# C[50] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4328 VDD a_1099_739# a_1317_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4329 a_3376_18251# a_2758_18706# a_2976_18747# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4330 a_40552_6503# a_40382_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4331 a_24449_6676# a_24451_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4332 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4333 a_5360_18251# a_4646_18706# a_5264_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4334 VDD a_1474_13071# a_2399_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4335 a_36138_5455# a_35779_5620# a_35777_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4336 VSS a_44288_18706# a_44236_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4337 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4338 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4339 a_25645_14292# a_25558_14194# a_25563_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4340 a_20577_6676# a_22197_6419# a_22011_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4341 a_35466_18251# a_36736_18706# a_36927_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4342 a_2569_12994# a_2399_12994# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4343 a_37301_6419# a_37075_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4344 a_39340_19307# a_38624_18706# a_37354_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4345 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4346 a_31309_14292# a_31222_14194# a_31227_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4347 VSS a_56214_13071# a_57139_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4348 VSS a_50175_739# a_50123_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4349 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_12898_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4350 a_43018_18251# a_44288_18706# a_44479_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4351 VSS a_13031_6676# a_13956_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4352 a_45217_6676# a_44853_6419# a_45121_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4353 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4354 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4355 a_57309_12994# a_57139_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4356 VSS C[11] a_38624_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4357 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4358 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4359 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4360 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4361 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4362 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_5346_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4363 a_23560_6503# a_23390_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4364 a_28143_1566# a_27473_765# a_27743_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4365 VSS C[8] a_44288_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4366 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4367 a_5066_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4368 VDD C[27] a_8422_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4369 a_57653_14292# a_57648_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4370 a_53832_12988# C[124] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4371 VDD a_55444_928# a_55394_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4372 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4373 a_28227_5620# a_27861_6419# a_26241_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4374 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4375 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_58427_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4376 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4377 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4378 a_16913_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4379 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4380 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4381 a_12900_14127# a_12308_12988# a_10914_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4382 a_26698_5455# a_26339_5620# a_26337_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4383 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4384 VSS a_14800_18251# a_14802_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4385 a_14788_14127# a_14422_13134# a_12802_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4386 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4387 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_19981_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4388 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_21869_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4389 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4390 a_41441_6676# a_41443_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4391 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4392 a_52170_13134# a_51944_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4393 a_32015_1566# a_31249_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4394 a_23940_1811# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4395 a_15573_18953# a_14704_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4396 a_9124_14127# a_8532_12988# a_7138_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4397 a_8987_6419# a_8761_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4398 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4399 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4400 a_6644_12988# C[99] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4401 VDD C[85] a_19973_739# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4402 a_39471_1566# a_40741_739# a_40932_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4403 a_22334_14127# a_21742_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4404 a_37665_6676# a_37075_6509# a_37569_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4405 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4406 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4407 VDD a_27632_13134# a_27446_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4408 a_54569_1566# a_53951_739# a_54169_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4409 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4410 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_42555_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4411 a_59722_13134# a_59496_12988# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4412 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4413 a_59577_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4414 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_1336_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4415 a_9136_18251# a_8370_18732# a_9040_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4416 a_5673_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4417 a_5479_6676# a_6873_6509# a_6913_5687# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4418 VDD a_48287_739# a_48235_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4419 a_43345_510# a_43343_1566# a_43656_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4420 a_18703_1566# a_18033_765# a_18303_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4421 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4422 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4423 a_30115_5620# a_29523_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4424 a_52399_6419# a_52173_6509# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4425 a_47113_1566# a_46347_765# a_47017_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4426 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4427 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4428 a_16171_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4429 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4430 a_34453_18953# a_33578_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4431 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4432 a_40552_6503# a_40382_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4433 a_5250_13071# a_6870_13134# a_6684_14194# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4434 a_54422_13071# a_53832_12988# a_54326_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4435 a_6870_13134# a_6644_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4436 a_41214_14127# a_40622_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4437 a_60102_19307# a_59334_18732# a_58116_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4438 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4439 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4440 a_23723_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4441 a_1801_5620# a_1209_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4442 VSS a_53722_18706# a_53670_18732# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4443 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_22016_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4444 a_45219_5620# a_44853_6419# a_43233_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4445 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4446 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4447 VSS a_9026_13071# a_9951_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4448 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4449 VDD a_870_18706# a_818_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4450 a_38458_928# a_37583_1566# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4451 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4452 VDD a_5250_13071# a_6175_12994# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4453 a_33905_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4454 a_14690_13071# a_14196_12988# a_14241_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4455 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_28586_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4456 a_22575_1566# a_21809_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4457 a_50564_18251# a_51834_18706# a_52025_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4458 a_35051_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4459 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4460 VSS a_38458_928# a_38408_763# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4461 a_54438_19307# a_53722_18706# a_52452_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4462 VSS a_1474_13071# a_2399_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4463 BR128half_0/sky130_fd_sc_hd__inv_16_0/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4464 a_52300_5455# a_52213_5687# a_52218_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4465 a_44853_6419# a_44627_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4466 a_2569_12994# a_2399_12994# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4467 a_14786_13071# a_14196_12988# a_14690_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4468 VDD a_2987_739# a_2935_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4469 a_42603_17686# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4470 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4471 a_60219_6676# a_59951_6419# a_59770_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4472 a_40932_1811# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4473 VSS C[4] a_51834_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4474 a_60102_19307# a_59386_18706# a_58116_18251# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4475 a_1813_1566# a_1047_765# a_1717_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4476 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_9122_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4477 a_20675_5620# a_20083_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4478 a_27635_6509# C[46] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4479 a_39555_5620# a_38963_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4480 a_52550_19307# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4481 a_1815_510# a_1099_739# a_794_737# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4482 a_22346_18251# a_21580_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4483 VDD a_27296_18706# a_27514_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4484 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4485 VSS a_5589_1566# a_5591_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4486 VSS C[0] a_59386_18706# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4487 VDD a_46170_18706# a_46118_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4488 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4489 a_13045_1566# a_12427_739# a_12645_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4490 a_3687_6676# a_3323_6419# a_3591_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4491 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4492 VDD BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4493 a_20446_14127# a_19854_12988# a_18460_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4494 a_48758_13071# a_48394_13134# a_48662_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4495 a_13045_1566# a_14263_765# a_14506_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4496 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4497 a_12802_13071# a_12534_13134# a_12353_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4498 a_58063_6419# a_57837_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4499 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4500 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4501 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_17029_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4502 a_22334_14127# a_21968_13134# a_20348_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4503 a_57918_1811# a_57945_1000# a_57930_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4504 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4505 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4506 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_27451_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4507 a_37667_5620# a_37075_6509# a_35681_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4508 a_20458_18251# a_19692_18732# a_20362_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4509 a_47115_510# a_47113_1566# a_47426_2061# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4510 VDD a_45121_6676# a_46046_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4511 a_41226_18251# a_40460_18732# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4512 VSS a_29898_18251# a_29900_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4513 VDD a_19349_18953# a_19299_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4514 a_11026_19307# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4515 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4516 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4517 a_9026_13071# a_8758_13134# a_8577_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4518 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4519 a_19349_18953# a_18474_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4520 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4521 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4522 a_565_18708# a_1435_6419# a_1249_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4523 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4524 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_27680_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4525 a_35695_1566# a_36913_765# a_37156_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4526 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4527 a_26110_14127# a_25518_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4528 a_50779_6676# a_50511_6419# a_50330_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4529 a_41457_510# a_40689_765# a_39471_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4530 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4531 a_46886_19307# a_46118_18732# a_44906_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4532 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4533 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4534 a_24463_1566# a_23749_739# a_24367_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4535 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_54188_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4536 VSS a_4251_18953# a_4201_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4537 a_4837_18006# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4538 a_17690_928# a_16815_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4539 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4540 a_39569_510# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4541 a_20689_510# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4542 a_9449_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4543 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4544 a_53556_928# a_52681_1566# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4545 a_10742_2061# BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4546 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4547 VDD a_38960_13134# a_38774_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4548 VSS a_2987_739# a_2935_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4549 a_794_737# a_1047_765# a_1290_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4550 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4551 a_46509_6509# C[56] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4552 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4553 a_57964_5455# a_57877_5687# a_57882_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4554 VDD a_38229_18953# a_38179_18734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4555 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4556 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4557 a_51874_6503# a_51704_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4558 a_10694_5455# a_10689_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4559 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4560 a_38229_18953# a_37354_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4561 a_7381_1566# a_6711_765# a_6981_1000# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4562 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4563 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4564 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4565 a_48623_6419# a_48397_6509# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4566 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4567 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4568 a_27499_17686# BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4569 VSS C[89] a_12427_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4570 VSS a_58441_1566# a_58443_510# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4571 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4572 a_58427_6676# a_57837_6509# a_58331_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4573 a_58331_6676# a_59951_6419# a_59765_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4574 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4575 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4576 VSS BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_20444_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4577 a_50889_1566# a_50123_765# a_50793_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4578 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4579 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4580 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4581 VSS a_5250_13071# a_6175_12994# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4582 a_3689_5620# a_3323_6419# a_1703_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4583 a_12898_13071# a_12900_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4584 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4585 a_56671_14292# a_56312_14127# a_56310_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4586 VSS C[77] a_35077_739# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4587 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4588 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4589 VSS BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y a_44672_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4590 a_5362_19307# a_5360_18251# a_5673_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4591 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4592 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4593 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4594 a_5346_13071# a_5348_14127# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4595 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4596 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4597 a_20348_13071# a_20080_13134# a_19899_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4598 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4599 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4600 a_16159_18006# a_16186_18747# a_16171_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4601 VSS BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4602 a_16123_14292# a_16118_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4603 a_24222_14127# a_23630_12988# a_22236_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4604 VSS a_45121_6676# a_46046_6503# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4605 a_18240_5455# a_18235_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4606 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4607 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4608 VDD a_57498_18706# a_57446_18732# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4609 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4610 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4611 VDD BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4612 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4613 a_23711_18006# a_23738_18747# a_23723_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4614 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4615 a_10350_6503# a_10180_6503# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4616 a_48891_6676# a_50511_6419# a_50325_5687# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4617 a_48987_6676# a_48397_6509# a_48891_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4618 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4619 a_46788_18251# a_46118_18732# a_46388_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4620 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_28357_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4621 VSS a_33674_18251# a_33676_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4622 VSS a_35562_18251# a_35564_19307# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4623 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_1254_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4624 a_18474_18251# a_19692_18732# a_19935_18006# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4625 VDD BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4626 BR128half_0/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4627 a_35003_14292# a_34998_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4628 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_53877_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4629 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_55765_14292# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4630 a_36891_14292# a_36886_14194# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4631 a_21968_13134# a_21742_12988# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4632 a_31182_12988# C[112] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4633 VDD BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_7824_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4634 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4635 VDD C[1] a_57498_18706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4636 a_58116_18251# a_57446_18732# a_57716_18747# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4637 VDD a_3591_6676# a_4516_6503# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4638 a_37681_510# a_36965_739# a_35695_1566# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4639 VDD a_10539_739# a_10487_765# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4640 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4641 VSS a_8027_18953# a_7977_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4642 a_42591_18006# a_42618_18747# a_42603_17686# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4643 BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4644 VDD a_46506_13134# a_46320_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4645 a_51874_6503# a_51704_6503# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4646 VSS a_9915_18953# a_9865_18734# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4647 VDD sky130_fd_sc_hd__inv_8_0/Y BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4648 VDD a_52170_13134# a_51984_14194# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4649 VDD BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4650 a_11157_1566# a_12375_765# a_12618_1811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4651 a_58429_5620# a_57837_6509# a_56443_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4652 VDD BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_3/Y a_51236_5455# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4653 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4654 a_6873_6509# C[35] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4655 BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4656 VDD a_25242_928# a_25192_763# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4657 BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4658 a_11239_6676# a_10875_6419# a_11143_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4659 a_53327_18953# a_52452_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4660 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4661 VSS BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_28225_6676# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4662 a_35280_2061# BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4663 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4664 BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4665 a_41212_13071# a_40848_13134# a_41116_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4666 a_30031_1566# a_31301_739# a_31492_1811# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4667 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_1/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4668 VSS BR128half_0/sky130_fd_sc_hd__inv_16_0/A BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4669 BR128half_0/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4670 a_55720_12988# C[125] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4671 a_35232_5455# a_35227_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4672 a_50285_6509# C[58] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4673 a_38815_18006# BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4674 VSS a_57716_18747# a_57689_18006# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4675 VDD BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4676 a_14919_6676# a_14651_6419# a_14470_5455# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4677 a_60329_1566# a_59563_765# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4678 VSS BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A BR128half_0/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4679 a_58212_18251# a_57446_18732# a_58116_18251# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4680 a_11239_6676# a_11241_5620# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4681 BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_0/sky130_fd_sc_hd__inv_16_0/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4682 a_33564_13071# a_33070_12988# a_33115_14292# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4683 a_56541_5620# a_56175_6419# a_54555_6676# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4684 a_56555_510# a_55787_765# a_54569_1566# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4685 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4686 BR128half_1/brbufhalf_2/sky130_fd_sc_hd__inv_16_3/Y BR128half_1/brbufhalf_1/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4687 a_13691_18953# a_12816_18251# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4688 a_1931_14292# a_1572_14127# a_1570_13071# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4689 VSS a_1099_739# a_1047_765# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4690 a_24367_1566# a_23749_739# a_23967_1000# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4691 a_33660_13071# a_33070_12988# a_33564_13071# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4692 a_31456_5455# a_31451_5687# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4693 VSS BR128half_1/brbufhalf_0/sky130_fd_sc_hd__inv_16_3/A BR128half_1/brbufhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

