magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 271 1418 582
rect -38 261 199 271
rect 525 261 1418 271
<< pwell >>
rect 279 176 488 229
rect 736 176 931 203
rect 279 157 931 176
rect 1103 157 1379 203
rect 1 40 1379 157
rect 1 21 271 40
rect 517 21 1379 40
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 367 119 397 203
rect 477 66 507 150
rect 622 47 652 125
rect 717 47 747 131
rect 823 47 853 177
rect 1011 47 1041 131
rect 1083 47 1113 131
rect 1179 47 1209 177
rect 1263 47 1293 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 447 413 477 497
rect 571 413 601 497
rect 643 413 673 497
rect 831 297 861 497
rect 927 369 957 497
rect 1083 369 1113 497
rect 1179 297 1209 497
rect 1263 297 1293 497
<< ndiff >>
rect 27 102 79 131
rect 27 68 35 102
rect 69 68 79 102
rect 27 47 79 68
rect 109 89 163 131
rect 109 55 119 89
rect 153 55 163 89
rect 109 47 163 55
rect 193 102 245 131
rect 193 68 203 102
rect 237 68 245 102
rect 193 47 245 68
rect 305 165 367 203
rect 305 131 313 165
rect 347 131 367 165
rect 305 119 367 131
rect 397 150 462 203
rect 397 119 477 150
rect 412 66 477 119
rect 507 125 557 150
rect 762 131 823 177
rect 667 125 717 131
rect 507 112 622 125
rect 507 78 575 112
rect 609 78 622 112
rect 507 66 622 78
rect 543 47 622 66
rect 652 47 717 125
rect 747 106 823 131
rect 747 72 779 106
rect 813 72 823 106
rect 747 47 823 72
rect 853 107 905 177
rect 1129 131 1179 177
rect 853 73 863 107
rect 897 73 905 107
rect 853 47 905 73
rect 959 108 1011 131
rect 959 74 967 108
rect 1001 74 1011 108
rect 959 47 1011 74
rect 1041 47 1083 131
rect 1113 93 1179 131
rect 1113 59 1135 93
rect 1169 59 1179 93
rect 1113 47 1179 59
rect 1209 101 1263 177
rect 1209 67 1219 101
rect 1253 67 1263 101
rect 1209 47 1263 67
rect 1293 161 1353 177
rect 1293 127 1309 161
rect 1343 127 1353 161
rect 1293 93 1353 127
rect 1293 59 1309 93
rect 1343 59 1353 93
rect 1293 47 1353 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 369 351 451
rect 381 413 447 497
rect 477 485 571 497
rect 477 451 512 485
rect 546 451 571 485
rect 477 413 571 451
rect 601 413 643 497
rect 673 477 725 497
rect 673 443 683 477
rect 717 443 725 477
rect 673 413 725 443
rect 779 471 831 497
rect 779 437 787 471
rect 821 437 831 471
rect 381 369 431 413
rect 779 368 831 437
rect 779 334 787 368
rect 821 334 831 368
rect 779 297 831 334
rect 861 471 927 497
rect 861 437 871 471
rect 905 437 927 471
rect 861 369 927 437
rect 957 485 1083 497
rect 957 451 1018 485
rect 1052 451 1083 485
rect 957 417 1083 451
rect 957 383 1018 417
rect 1052 383 1083 417
rect 957 369 1083 383
rect 1113 476 1179 497
rect 1113 442 1135 476
rect 1169 442 1179 476
rect 1113 369 1179 442
rect 861 297 911 369
rect 1129 297 1179 369
rect 1209 475 1263 497
rect 1209 441 1219 475
rect 1253 441 1263 475
rect 1209 349 1263 441
rect 1209 315 1219 349
rect 1253 315 1263 349
rect 1209 297 1263 315
rect 1293 485 1353 497
rect 1293 451 1309 485
rect 1343 451 1353 485
rect 1293 417 1353 451
rect 1293 383 1309 417
rect 1343 383 1353 417
rect 1293 349 1353 383
rect 1293 315 1309 349
rect 1343 315 1353 349
rect 1293 297 1353 315
<< ndiffc >>
rect 35 68 69 102
rect 119 55 153 89
rect 203 68 237 102
rect 313 131 347 165
rect 575 78 609 112
rect 779 72 813 106
rect 863 73 897 107
rect 967 74 1001 108
rect 1135 59 1169 93
rect 1219 67 1253 101
rect 1309 127 1343 161
rect 1309 59 1343 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 451 341 485
rect 512 451 546 485
rect 683 443 717 477
rect 787 437 821 471
rect 787 334 821 368
rect 871 437 905 471
rect 1018 451 1052 485
rect 1018 383 1052 417
rect 1135 442 1169 476
rect 1219 441 1253 475
rect 1219 315 1253 349
rect 1309 451 1343 485
rect 1309 383 1343 417
rect 1309 315 1343 349
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 447 497 477 523
rect 571 497 601 523
rect 643 497 673 523
rect 831 497 861 523
rect 927 497 957 523
rect 1083 497 1113 523
rect 1179 497 1209 523
rect 1263 497 1293 523
rect 447 375 477 413
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 22 264 76 280
rect 163 272 193 363
rect 351 337 381 369
rect 22 230 32 264
rect 66 230 76 264
rect 22 214 76 230
rect 118 262 193 272
rect 327 321 381 337
rect 447 365 529 375
rect 447 331 479 365
rect 513 331 529 365
rect 447 321 529 331
rect 327 287 337 321
rect 371 287 381 321
rect 327 271 381 287
rect 571 279 601 413
rect 643 373 673 413
rect 643 357 747 373
rect 643 323 687 357
rect 721 323 747 357
rect 643 307 747 323
rect 118 228 134 262
rect 168 228 193 262
rect 118 218 193 228
rect 351 248 381 271
rect 477 249 601 279
rect 351 218 397 248
rect 46 176 76 214
rect 163 176 193 218
rect 367 203 397 218
rect 46 146 109 176
rect 79 131 109 146
rect 163 146 290 176
rect 163 131 193 146
rect 260 51 290 146
rect 477 150 507 249
rect 579 197 652 207
rect 579 163 595 197
rect 629 163 652 197
rect 579 153 652 163
rect 367 93 397 119
rect 622 125 652 153
rect 717 131 747 307
rect 831 265 861 297
rect 927 265 957 369
rect 1083 287 1113 369
rect 792 249 861 265
rect 792 215 802 249
rect 836 215 861 249
rect 792 199 861 215
rect 903 249 957 265
rect 903 215 913 249
rect 947 215 957 249
rect 1037 271 1113 287
rect 1037 237 1047 271
rect 1081 237 1113 271
rect 1179 265 1209 297
rect 1263 265 1293 297
rect 1037 221 1113 237
rect 903 199 957 215
rect 823 177 853 199
rect 477 51 507 66
rect 79 21 109 47
rect 163 21 193 47
rect 260 21 507 51
rect 927 176 957 199
rect 927 146 1041 176
rect 1011 131 1041 146
rect 1083 131 1113 221
rect 1155 249 1293 265
rect 1155 215 1165 249
rect 1199 215 1293 249
rect 1155 199 1293 215
rect 1179 177 1209 199
rect 1263 177 1293 199
rect 622 21 652 47
rect 717 21 747 47
rect 823 21 853 47
rect 1011 21 1041 47
rect 1083 21 1113 47
rect 1179 21 1209 47
rect 1263 21 1293 47
<< polycont >>
rect 32 230 66 264
rect 479 331 513 365
rect 337 287 371 321
rect 687 323 721 357
rect 134 228 168 262
rect 595 163 629 197
rect 802 215 836 249
rect 913 215 947 249
rect 1047 237 1081 271
rect 1165 215 1199 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 203 409 248 443
rect 291 485 364 527
rect 291 451 307 485
rect 341 451 364 485
rect 496 451 512 485
rect 546 451 646 485
rect 291 439 364 451
rect 69 375 156 393
rect 35 359 156 375
rect 18 264 66 325
rect 18 255 32 264
rect 18 221 30 255
rect 64 221 66 230
rect 18 197 66 221
rect 122 278 156 359
rect 237 405 248 409
rect 237 375 529 405
rect 203 371 529 375
rect 122 262 168 278
rect 122 228 134 262
rect 122 212 168 228
rect 122 157 156 212
rect 35 123 156 157
rect 35 102 69 123
rect 203 102 256 371
rect 479 365 529 371
rect 306 321 443 337
rect 306 287 337 321
rect 371 287 443 321
rect 35 52 69 68
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 237 68 256 102
rect 203 52 256 68
rect 297 165 363 181
rect 297 131 313 165
rect 347 131 363 165
rect 297 17 363 131
rect 397 57 443 287
rect 513 331 529 365
rect 479 197 529 331
rect 612 265 646 451
rect 680 477 740 527
rect 680 443 683 477
rect 717 443 740 477
rect 680 427 740 443
rect 783 471 827 487
rect 783 437 787 471
rect 821 437 827 471
rect 783 373 827 437
rect 863 471 920 527
rect 863 437 871 471
rect 905 437 920 471
rect 863 402 920 437
rect 1002 485 1068 493
rect 1002 451 1018 485
rect 1052 451 1068 485
rect 1002 417 1068 451
rect 1115 476 1185 527
rect 1115 442 1135 476
rect 1169 442 1185 476
rect 1115 426 1185 442
rect 1219 475 1272 491
rect 1253 441 1272 475
rect 687 368 827 373
rect 1002 383 1018 417
rect 1052 383 1068 417
rect 1002 379 1068 383
rect 687 357 787 368
rect 721 334 787 357
rect 821 334 947 368
rect 1002 345 1185 379
rect 721 323 947 334
rect 687 307 947 323
rect 612 249 836 265
rect 612 231 802 249
rect 711 215 802 231
rect 711 199 836 215
rect 870 249 947 307
rect 870 215 913 249
rect 1042 271 1097 287
rect 1042 255 1047 271
rect 1081 237 1097 271
rect 1076 221 1097 237
rect 1151 265 1185 345
rect 1219 349 1272 441
rect 1253 315 1272 349
rect 1219 299 1272 315
rect 1151 249 1199 265
rect 870 199 947 215
rect 1151 215 1165 249
rect 479 163 595 197
rect 629 163 645 197
rect 711 112 745 199
rect 870 123 917 199
rect 1151 187 1199 215
rect 986 153 1199 187
rect 986 124 1030 153
rect 559 78 575 112
rect 609 78 745 112
rect 779 106 829 122
rect 813 72 829 106
rect 779 17 829 72
rect 863 107 917 123
rect 897 73 917 107
rect 863 51 917 73
rect 967 108 1030 124
rect 1233 119 1272 299
rect 1306 485 1362 527
rect 1306 451 1309 485
rect 1343 451 1362 485
rect 1306 417 1362 451
rect 1306 383 1309 417
rect 1343 383 1362 417
rect 1306 349 1362 383
rect 1306 315 1309 349
rect 1343 315 1362 349
rect 1306 297 1362 315
rect 1001 74 1030 108
rect 967 58 1030 74
rect 1135 93 1169 109
rect 1135 17 1169 59
rect 1212 101 1272 119
rect 1212 67 1219 101
rect 1253 67 1272 101
rect 1212 51 1272 67
rect 1306 161 1362 177
rect 1306 127 1309 161
rect 1343 127 1362 161
rect 1306 93 1362 127
rect 1306 59 1309 93
rect 1343 59 1362 93
rect 1306 17 1362 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 30 230 32 255
rect 32 230 64 255
rect 30 221 64 230
rect 1042 237 1047 255
rect 1047 237 1076 255
rect 1042 221 1076 237
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 18 255 76 261
rect 18 221 30 255
rect 64 252 76 255
rect 1030 255 1088 261
rect 1030 252 1042 255
rect 64 224 1042 252
rect 64 221 76 224
rect 18 215 76 221
rect 1030 221 1042 224
rect 1076 221 1088 255
rect 1030 215 1088 221
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
flabel locali s 306 289 340 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 1226 85 1260 119 0 FreeSans 200 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1226 425 1260 459 0 FreeSans 200 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 1226 357 1260 391 0 FreeSans 200 0 0 0 GCLK
port 7 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 dlclkp_2
rlabel locali s 1042 221 1097 287 1 CLK
port 1 nsew clock input
rlabel metal1 s 1030 252 1088 261 1 CLK
port 1 nsew clock input
rlabel metal1 s 1030 215 1088 224 1 CLK
port 1 nsew clock input
rlabel metal1 s 18 252 76 261 1 CLK
port 1 nsew clock input
rlabel metal1 s 18 224 1088 252 1 CLK
port 1 nsew clock input
rlabel metal1 s 18 215 76 224 1 CLK
port 1 nsew clock input
rlabel metal1 s 0 -48 1380 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_END 2642408
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2632154
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 34.500 13.600 
<< end >>
