magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 6571 2023 7265 2239
rect 14401 1739 14733 2233
<< pwell >>
rect 868 1853 1120 2267
rect 86 1367 738 1376
rect 86 58 850 1367
rect 764 52 850 58
<< mvnmos >>
rect 894 2088 1094 2188
rect 894 1932 1094 2032
rect 112 1197 712 1297
rect 112 1041 712 1141
rect 112 885 712 985
rect 112 729 712 829
rect 112 573 712 673
rect 112 417 712 517
rect 112 137 712 237
<< mvpmos >>
rect 6690 2089 6890 2173
rect 6946 2089 7146 2173
rect 14467 2014 14667 2114
rect 14467 1858 14667 1958
<< mvndiff >>
rect 894 2233 1094 2241
rect 894 2199 906 2233
rect 940 2199 974 2233
rect 1008 2199 1042 2233
rect 1076 2199 1094 2233
rect 894 2188 1094 2199
rect 894 2077 1094 2088
rect 894 2043 906 2077
rect 940 2043 974 2077
rect 1008 2043 1042 2077
rect 1076 2043 1094 2077
rect 894 2032 1094 2043
rect 894 1921 1094 1932
rect 894 1887 906 1921
rect 940 1887 974 1921
rect 1008 1887 1042 1921
rect 1076 1887 1094 1921
rect 894 1879 1094 1887
rect 112 1342 712 1350
rect 112 1308 190 1342
rect 224 1308 258 1342
rect 292 1308 326 1342
rect 360 1308 394 1342
rect 428 1308 462 1342
rect 496 1308 530 1342
rect 564 1308 598 1342
rect 632 1308 666 1342
rect 700 1308 712 1342
rect 112 1297 712 1308
rect 112 1186 712 1197
rect 112 1152 190 1186
rect 224 1152 258 1186
rect 292 1152 326 1186
rect 360 1152 394 1186
rect 428 1152 462 1186
rect 496 1152 530 1186
rect 564 1152 598 1186
rect 632 1152 666 1186
rect 700 1152 712 1186
rect 112 1141 712 1152
rect 112 1030 712 1041
rect 112 996 190 1030
rect 224 996 258 1030
rect 292 996 326 1030
rect 360 996 394 1030
rect 428 996 462 1030
rect 496 996 530 1030
rect 564 996 598 1030
rect 632 996 666 1030
rect 700 996 712 1030
rect 112 985 712 996
rect 112 874 712 885
rect 112 840 190 874
rect 224 840 258 874
rect 292 840 326 874
rect 360 840 394 874
rect 428 840 462 874
rect 496 840 530 874
rect 564 840 598 874
rect 632 840 666 874
rect 700 840 712 874
rect 112 829 712 840
rect 112 718 712 729
rect 112 684 190 718
rect 224 684 258 718
rect 292 684 326 718
rect 360 684 394 718
rect 428 684 462 718
rect 496 684 530 718
rect 564 684 598 718
rect 632 684 666 718
rect 700 684 712 718
rect 112 673 712 684
rect 112 562 712 573
rect 112 528 190 562
rect 224 528 258 562
rect 292 528 326 562
rect 360 528 394 562
rect 428 528 462 562
rect 496 528 530 562
rect 564 528 598 562
rect 632 528 666 562
rect 700 528 712 562
rect 112 517 712 528
rect 112 406 712 417
rect 112 372 190 406
rect 224 372 258 406
rect 292 372 326 406
rect 360 372 394 406
rect 428 372 462 406
rect 496 372 530 406
rect 564 372 598 406
rect 632 372 666 406
rect 700 372 712 406
rect 112 364 712 372
rect 112 282 712 290
rect 112 248 190 282
rect 224 248 258 282
rect 292 248 326 282
rect 360 248 394 282
rect 428 248 462 282
rect 496 248 530 282
rect 564 248 598 282
rect 632 248 666 282
rect 700 248 712 282
rect 112 237 712 248
rect 112 126 712 137
rect 112 92 190 126
rect 224 92 258 126
rect 292 92 326 126
rect 360 92 394 126
rect 428 92 462 126
rect 496 92 530 126
rect 564 92 598 126
rect 632 92 666 126
rect 700 92 712 126
rect 112 84 712 92
<< mvpdiff >>
rect 6637 2161 6690 2173
rect 6637 2127 6645 2161
rect 6679 2127 6690 2161
rect 6637 2089 6690 2127
rect 6890 2161 6946 2173
rect 6890 2127 6901 2161
rect 6935 2127 6946 2161
rect 6890 2089 6946 2127
rect 7146 2161 7199 2173
rect 7146 2127 7157 2161
rect 7191 2127 7199 2161
rect 7146 2089 7199 2127
rect 14467 2159 14667 2167
rect 14467 2125 14479 2159
rect 14513 2125 14547 2159
rect 14581 2125 14615 2159
rect 14649 2125 14667 2159
rect 14467 2114 14667 2125
rect 14467 2003 14667 2014
rect 14467 1969 14479 2003
rect 14513 1969 14547 2003
rect 14581 1969 14615 2003
rect 14649 1969 14667 2003
rect 14467 1958 14667 1969
rect 14467 1847 14667 1858
rect 14467 1813 14479 1847
rect 14513 1813 14547 1847
rect 14581 1813 14615 1847
rect 14649 1813 14667 1847
rect 14467 1805 14667 1813
<< mvndiffc >>
rect 906 2199 940 2233
rect 974 2199 1008 2233
rect 1042 2199 1076 2233
rect 906 2043 940 2077
rect 974 2043 1008 2077
rect 1042 2043 1076 2077
rect 906 1887 940 1921
rect 974 1887 1008 1921
rect 1042 1887 1076 1921
rect 190 1308 224 1342
rect 258 1308 292 1342
rect 326 1308 360 1342
rect 394 1308 428 1342
rect 462 1308 496 1342
rect 530 1308 564 1342
rect 598 1308 632 1342
rect 666 1308 700 1342
rect 190 1152 224 1186
rect 258 1152 292 1186
rect 326 1152 360 1186
rect 394 1152 428 1186
rect 462 1152 496 1186
rect 530 1152 564 1186
rect 598 1152 632 1186
rect 666 1152 700 1186
rect 190 996 224 1030
rect 258 996 292 1030
rect 326 996 360 1030
rect 394 996 428 1030
rect 462 996 496 1030
rect 530 996 564 1030
rect 598 996 632 1030
rect 666 996 700 1030
rect 190 840 224 874
rect 258 840 292 874
rect 326 840 360 874
rect 394 840 428 874
rect 462 840 496 874
rect 530 840 564 874
rect 598 840 632 874
rect 666 840 700 874
rect 190 684 224 718
rect 258 684 292 718
rect 326 684 360 718
rect 394 684 428 718
rect 462 684 496 718
rect 530 684 564 718
rect 598 684 632 718
rect 666 684 700 718
rect 190 528 224 562
rect 258 528 292 562
rect 326 528 360 562
rect 394 528 428 562
rect 462 528 496 562
rect 530 528 564 562
rect 598 528 632 562
rect 666 528 700 562
rect 190 372 224 406
rect 258 372 292 406
rect 326 372 360 406
rect 394 372 428 406
rect 462 372 496 406
rect 530 372 564 406
rect 598 372 632 406
rect 666 372 700 406
rect 190 248 224 282
rect 258 248 292 282
rect 326 248 360 282
rect 394 248 428 282
rect 462 248 496 282
rect 530 248 564 282
rect 598 248 632 282
rect 666 248 700 282
rect 190 92 224 126
rect 258 92 292 126
rect 326 92 360 126
rect 394 92 428 126
rect 462 92 496 126
rect 530 92 564 126
rect 598 92 632 126
rect 666 92 700 126
<< mvpdiffc >>
rect 6645 2127 6679 2161
rect 6901 2127 6935 2161
rect 7157 2127 7191 2161
rect 14479 2125 14513 2159
rect 14547 2125 14581 2159
rect 14615 2125 14649 2159
rect 14479 1969 14513 2003
rect 14547 1969 14581 2003
rect 14615 1969 14649 2003
rect 14479 1813 14513 1847
rect 14547 1813 14581 1847
rect 14615 1813 14649 1847
<< psubdiff >>
rect 790 1317 824 1341
rect 790 1248 824 1283
rect 790 1179 824 1214
rect 790 1110 824 1145
rect 790 1041 824 1076
rect 790 972 824 1007
rect 790 903 824 938
rect 790 834 824 869
rect 790 765 824 800
rect 790 696 824 731
rect 790 626 824 662
rect 790 556 824 592
rect 790 486 824 522
rect 790 416 824 452
rect 790 346 824 382
rect 790 276 824 312
rect 790 206 824 242
rect 790 136 824 172
rect 790 78 824 102
<< psubdiffcont >>
rect 790 1283 824 1317
rect 790 1214 824 1248
rect 790 1145 824 1179
rect 790 1076 824 1110
rect 790 1007 824 1041
rect 790 938 824 972
rect 790 869 824 903
rect 790 800 824 834
rect 790 731 824 765
rect 790 662 824 696
rect 790 592 824 626
rect 790 522 824 556
rect 790 452 824 486
rect 790 382 824 416
rect 790 312 824 346
rect 790 242 824 276
rect 790 172 824 206
rect 790 102 824 136
<< poly >>
rect 6691 2255 6891 2271
rect 1124 2209 1190 2225
rect 1124 2188 1140 2209
rect 862 2088 894 2188
rect 1094 2175 1140 2188
rect 1174 2175 1190 2209
rect 6691 2221 6707 2255
rect 6741 2221 6841 2255
rect 6875 2221 6891 2255
rect 6691 2205 6891 2221
rect 6947 2255 7147 2271
rect 6947 2221 6963 2255
rect 6997 2221 7097 2255
rect 7131 2221 7147 2255
rect 6947 2205 7147 2221
rect 1094 2138 1190 2175
rect 6690 2173 6890 2205
rect 6946 2173 7146 2205
rect 1094 2104 1140 2138
rect 1174 2104 1190 2138
rect 1094 2088 1190 2104
rect 14369 2098 14467 2114
rect 6690 2057 6890 2089
rect 6946 2057 7146 2089
rect 14369 2064 14385 2098
rect 14419 2064 14467 2098
rect 862 1932 894 2032
rect 1094 2016 1190 2032
rect 1094 1982 1140 2016
rect 1174 1982 1190 2016
rect 1094 1945 1190 1982
rect 1094 1932 1140 1945
rect 1124 1911 1140 1932
rect 1174 1911 1190 1945
rect 1124 1895 1190 1911
rect 14369 2014 14467 2064
rect 14667 2014 14699 2114
rect 14369 2003 14435 2014
rect 14369 1969 14385 2003
rect 14419 1969 14435 2003
rect 14369 1958 14435 1969
rect 14369 1908 14467 1958
rect 14369 1874 14385 1908
rect 14419 1874 14467 1908
rect 14369 1858 14467 1874
rect 14667 1858 14699 1958
rect 14 1281 112 1297
rect 14 1247 30 1281
rect 64 1247 112 1281
rect 14 1212 112 1247
rect 14 1178 30 1212
rect 64 1197 112 1212
rect 712 1197 744 1297
rect 64 1178 80 1197
rect 14 1143 80 1178
rect 14 1109 30 1143
rect 64 1141 80 1143
rect 64 1109 112 1141
rect 14 1074 112 1109
rect 14 1040 30 1074
rect 64 1041 112 1074
rect 712 1041 744 1141
rect 64 1040 80 1041
rect 14 1005 80 1040
rect 14 971 30 1005
rect 64 985 80 1005
rect 64 971 112 985
rect 14 935 112 971
rect 14 901 30 935
rect 64 901 112 935
rect 14 885 112 901
rect 712 885 744 985
rect 14 813 112 829
rect 14 779 30 813
rect 64 779 112 813
rect 14 744 112 779
rect 14 710 30 744
rect 64 729 112 744
rect 712 729 744 829
rect 64 710 80 729
rect 14 675 80 710
rect 14 641 30 675
rect 64 673 80 675
rect 64 641 112 673
rect 14 606 112 641
rect 14 572 30 606
rect 64 573 112 606
rect 712 573 744 673
rect 64 572 80 573
rect 14 537 80 572
rect 14 503 30 537
rect 64 517 80 537
rect 64 503 112 517
rect 14 467 112 503
rect 14 433 30 467
rect 64 433 112 467
rect 14 417 112 433
rect 712 417 744 517
rect 14 238 80 254
rect 14 204 30 238
rect 64 237 80 238
rect 64 204 112 237
rect 14 170 112 204
rect 14 136 30 170
rect 64 137 112 170
rect 712 137 744 237
rect 64 136 80 137
rect 14 120 80 136
<< polycont >>
rect 1140 2175 1174 2209
rect 6707 2221 6741 2255
rect 6841 2221 6875 2255
rect 6963 2221 6997 2255
rect 7097 2221 7131 2255
rect 1140 2104 1174 2138
rect 14385 2064 14419 2098
rect 1140 1982 1174 2016
rect 1140 1911 1174 1945
rect 14385 1969 14419 2003
rect 14385 1874 14419 1908
rect 30 1247 64 1281
rect 30 1178 64 1212
rect 30 1109 64 1143
rect 30 1040 64 1074
rect 30 971 64 1005
rect 30 901 64 935
rect 30 779 64 813
rect 30 710 64 744
rect 30 641 64 675
rect 30 572 64 606
rect 30 503 64 537
rect 30 433 64 467
rect 30 204 64 238
rect 30 136 64 170
<< locali >>
rect 890 2199 906 2233
rect 940 2199 974 2233
rect 1014 2199 1042 2233
rect 1086 2199 1092 2233
rect 6691 2221 6703 2255
rect 6741 2221 6841 2255
rect 6879 2221 6891 2255
rect 6947 2221 6959 2255
rect 6997 2221 7097 2255
rect 7135 2221 7147 2255
rect 1140 2163 1174 2175
rect 6645 2174 6679 2177
rect 824 2077 1091 2109
rect 1140 2088 1174 2104
rect 6676 2161 6679 2174
rect 6642 2127 6645 2140
rect 6642 2111 6679 2127
rect 6901 2161 6935 2177
rect 6901 2111 6935 2127
rect 7157 2174 7191 2177
rect 6642 2102 6676 2111
rect 824 2043 906 2077
rect 940 2043 974 2077
rect 1008 2043 1042 2077
rect 1076 2043 1092 2077
rect 7157 2102 7191 2127
rect 14463 2162 14666 2168
rect 14463 2159 14568 2162
rect 14602 2159 14640 2162
rect 14463 2125 14479 2159
rect 14513 2125 14547 2159
rect 14602 2128 14615 2159
rect 14581 2125 14615 2128
rect 14649 2125 14666 2128
rect 14463 2114 14666 2125
rect 14385 2102 14419 2114
rect 14411 2098 14419 2102
rect 14377 2064 14385 2068
rect 824 1990 1091 2043
rect 1140 2020 1174 2032
rect 14377 2030 14419 2064
rect 14411 2003 14419 2030
rect 14509 2003 14604 2009
rect 1140 1945 1174 1982
rect 905 1887 906 1921
rect 940 1887 950 1921
rect 1008 1887 1042 1921
rect 1076 1887 1092 1921
rect 1140 1895 1174 1907
rect 14463 1975 14475 2003
rect 14463 1969 14479 1975
rect 14513 1969 14547 2003
rect 14581 1975 14604 2003
rect 14581 1969 14615 1975
rect 14649 1969 14665 2003
rect 14385 1908 14419 1969
rect 14385 1858 14419 1874
rect 14463 1813 14479 1847
rect 14513 1813 14547 1847
rect 14587 1813 14615 1847
rect 14659 1813 14665 1847
rect 174 1308 190 1342
rect 224 1308 258 1342
rect 292 1308 326 1342
rect 360 1308 394 1342
rect 428 1308 453 1342
rect 496 1308 526 1342
rect 564 1308 598 1342
rect 632 1308 666 1342
rect 704 1308 716 1342
rect 790 1329 824 1341
rect 30 1281 64 1297
rect 30 1212 64 1247
rect 790 1254 824 1283
rect 30 1143 64 1160
rect 174 1152 190 1186
rect 224 1152 258 1186
rect 292 1152 326 1186
rect 360 1152 394 1186
rect 428 1152 462 1186
rect 496 1152 530 1186
rect 564 1152 598 1186
rect 632 1152 635 1186
rect 700 1152 707 1186
rect 790 1179 824 1214
rect 30 1107 64 1109
rect 30 1019 64 1040
rect 790 1110 824 1145
rect 790 1041 824 1070
rect 174 996 190 1030
rect 224 996 258 1030
rect 292 996 326 1030
rect 360 996 394 1030
rect 428 996 453 1030
rect 496 996 525 1030
rect 564 996 598 1030
rect 632 996 666 1030
rect 700 996 716 1030
rect 30 935 64 971
rect 30 885 64 897
rect 790 972 824 995
rect 790 903 824 920
rect 174 840 190 874
rect 224 840 258 874
rect 292 840 326 874
rect 360 840 394 874
rect 428 840 462 874
rect 496 840 530 874
rect 564 840 598 874
rect 632 840 635 874
rect 700 840 707 874
rect 790 834 824 845
rect 30 817 64 829
rect 30 744 64 779
rect 790 765 824 770
rect 790 728 824 731
rect 30 675 64 695
rect 174 684 190 718
rect 224 684 258 718
rect 292 684 326 718
rect 360 684 394 718
rect 428 684 462 718
rect 509 684 530 718
rect 581 684 598 718
rect 632 684 666 718
rect 700 684 716 718
rect 30 606 64 607
rect 30 552 64 572
rect 790 652 824 662
rect 790 576 824 592
rect 174 528 190 562
rect 224 528 258 562
rect 292 528 326 562
rect 360 528 394 562
rect 428 528 462 562
rect 496 528 530 562
rect 564 528 598 562
rect 632 528 635 562
rect 700 528 707 562
rect 30 467 64 503
rect 30 417 64 429
rect 790 500 824 522
rect 790 424 824 452
rect 174 372 190 406
rect 224 372 258 406
rect 292 372 326 406
rect 360 372 394 406
rect 428 372 462 406
rect 509 372 530 406
rect 581 372 598 406
rect 632 372 666 406
rect 700 372 716 406
rect 790 348 824 382
rect 30 242 64 254
rect 174 248 190 282
rect 224 248 258 282
rect 292 248 326 282
rect 360 248 394 282
rect 428 248 462 282
rect 496 248 530 282
rect 564 248 598 282
rect 632 248 635 282
rect 700 248 707 282
rect 790 276 824 312
rect 34 238 64 242
rect 0 204 30 208
rect 0 170 64 204
rect 0 166 30 170
rect 34 132 64 136
rect 30 120 64 132
rect 790 206 824 238
rect 790 136 824 162
rect 174 92 190 126
rect 224 92 258 126
rect 292 92 326 126
rect 360 92 394 126
rect 428 92 462 126
rect 496 92 530 126
rect 564 92 598 126
rect 662 92 666 126
rect 700 92 705 126
rect 790 78 824 86
<< viali >>
rect 980 2199 1008 2233
rect 1008 2199 1014 2233
rect 1052 2199 1076 2233
rect 1076 2199 1086 2233
rect 1140 2209 1174 2242
rect 6703 2221 6707 2255
rect 6707 2221 6737 2255
rect 6845 2221 6875 2255
rect 6875 2221 6879 2255
rect 6959 2221 6963 2255
rect 6963 2221 6993 2255
rect 7101 2221 7131 2255
rect 7131 2221 7135 2255
rect 1140 2208 1174 2209
rect 1140 2138 1174 2163
rect 1140 2129 1174 2138
rect 6642 2161 6676 2174
rect 6642 2140 6645 2161
rect 6645 2140 6676 2161
rect 7157 2161 7191 2174
rect 7157 2140 7191 2161
rect 6642 2068 6676 2102
rect 14568 2159 14602 2162
rect 14640 2159 14674 2162
rect 14568 2128 14581 2159
rect 14581 2128 14602 2159
rect 14640 2128 14649 2159
rect 14649 2128 14674 2159
rect 7157 2068 7191 2102
rect 14377 2098 14411 2102
rect 14377 2068 14385 2098
rect 14385 2068 14411 2098
rect 1140 2016 1174 2020
rect 1140 1986 1174 2016
rect 14377 2003 14411 2030
rect 14475 2003 14509 2009
rect 14604 2003 14638 2009
rect 14377 1996 14385 2003
rect 14385 1996 14411 2003
rect 871 1887 905 1921
rect 950 1887 974 1921
rect 974 1887 984 1921
rect 1140 1911 1174 1941
rect 1140 1907 1174 1911
rect 14475 1975 14479 2003
rect 14479 1975 14509 2003
rect 14604 1975 14615 2003
rect 14615 1975 14638 2003
rect 14553 1813 14581 1847
rect 14581 1813 14587 1847
rect 14625 1813 14649 1847
rect 14649 1813 14659 1847
rect 453 1308 462 1342
rect 462 1308 487 1342
rect 526 1308 530 1342
rect 530 1308 560 1342
rect 598 1308 632 1342
rect 670 1308 700 1342
rect 700 1308 704 1342
rect 790 1317 824 1329
rect 30 1178 64 1194
rect 790 1295 824 1317
rect 790 1248 824 1254
rect 790 1220 824 1248
rect 30 1160 64 1178
rect 635 1152 666 1186
rect 666 1152 669 1186
rect 707 1152 741 1186
rect 30 1074 64 1107
rect 30 1073 64 1074
rect 790 1145 824 1179
rect 790 1076 824 1104
rect 790 1070 824 1076
rect 30 1005 64 1019
rect 30 985 64 1005
rect 453 996 462 1030
rect 462 996 487 1030
rect 525 996 530 1030
rect 530 996 559 1030
rect 790 1007 824 1029
rect 30 901 64 931
rect 30 897 64 901
rect 790 995 824 1007
rect 790 938 824 954
rect 790 920 824 938
rect 635 840 666 874
rect 666 840 669 874
rect 707 840 741 874
rect 790 869 824 879
rect 790 845 824 869
rect 30 813 64 817
rect 30 783 64 813
rect 30 710 64 729
rect 790 800 824 804
rect 790 770 824 800
rect 30 695 64 710
rect 475 684 496 718
rect 496 684 509 718
rect 547 684 564 718
rect 564 684 581 718
rect 790 696 824 728
rect 790 694 824 696
rect 30 607 64 641
rect 790 626 824 652
rect 790 618 824 626
rect 30 537 64 552
rect 30 518 64 537
rect 635 528 666 562
rect 666 528 669 562
rect 707 528 741 562
rect 790 556 824 576
rect 790 542 824 556
rect 30 433 64 463
rect 30 429 64 433
rect 790 486 824 500
rect 790 466 824 486
rect 790 416 824 424
rect 475 372 496 406
rect 496 372 509 406
rect 547 372 564 406
rect 564 372 581 406
rect 790 390 824 416
rect 790 346 824 348
rect 790 314 824 346
rect 635 248 666 282
rect 666 248 669 282
rect 707 248 741 282
rect 0 238 34 242
rect 0 208 30 238
rect 30 208 34 238
rect 0 136 30 166
rect 30 136 34 166
rect 0 132 34 136
rect 790 242 824 272
rect 790 238 824 242
rect 790 172 824 196
rect 790 162 824 172
rect 628 92 632 126
rect 632 92 662 126
rect 705 92 739 126
rect 790 102 824 120
rect 790 86 824 102
<< metal1 >>
rect 155 1381 185 2964
rect 8007 2888 14977 2916
rect 33 1351 185 1381
rect 33 1206 63 1351
rect 24 1194 70 1206
rect 24 1160 30 1194
rect 64 1160 70 1194
rect 24 1107 70 1160
rect 24 1073 30 1107
rect 64 1073 70 1107
rect 24 1019 70 1073
rect 24 985 30 1019
rect 64 985 70 1019
rect 24 931 70 985
rect 24 897 30 931
rect 64 897 70 931
rect 24 885 70 897
tri 181 840 215 874 se
rect 215 841 243 2882
rect 676 2026 728 2425
rect 2730 2299 2736 2351
rect 2788 2299 2800 2351
rect 2852 2299 2858 2351
rect 2730 2291 2858 2299
tri 2772 2257 2806 2291 ne
rect 1134 2242 1180 2254
rect 968 2233 1098 2239
rect 968 2199 980 2233
rect 1014 2199 1052 2233
rect 1086 2199 1098 2233
rect 968 2193 1098 2199
tri 1026 2174 1045 2193 ne
rect 1045 2174 1098 2193
tri 1045 2167 1052 2174 ne
rect 1052 2071 1098 2174
rect 1134 2208 1140 2242
rect 1174 2208 1180 2242
rect 1134 2163 1180 2208
rect 1134 2129 1140 2163
rect 1174 2129 1180 2163
rect 1134 2117 1180 2129
rect 2806 2080 2858 2291
rect 292 1990 366 1996
rect 292 1938 314 1990
rect 292 1917 366 1938
rect 292 1865 314 1917
rect 292 1858 366 1865
rect 292 1847 355 1858
tri 355 1847 366 1858 nw
rect 676 1953 728 1974
rect 292 1392 328 1847
tri 328 1820 355 1847 nw
tri 292 1356 328 1392 ne
tri 328 1382 362 1416 sw
rect 328 1356 362 1382
tri 362 1356 388 1382 sw
tri 650 1356 676 1382 se
rect 676 1356 728 1901
rect 859 2019 865 2071
rect 917 2019 938 2071
rect 990 2019 996 2071
rect 1052 2019 1058 2071
rect 1110 2019 1131 2071
rect 1183 2019 1189 2071
tri 6613 2318 6639 2344 se
rect 6639 2318 7358 2344
rect 6613 2301 7358 2318
rect 6613 2186 6659 2301
tri 6659 2282 6678 2301 nw
tri 6923 2282 6942 2301 ne
rect 6942 2298 7358 2301
rect 6942 2282 7147 2298
tri 6942 2277 6947 2282 ne
rect 6691 2219 6697 2271
rect 6749 2219 6765 2271
rect 6817 2219 6833 2271
rect 6885 2219 6891 2271
rect 6691 2215 6891 2219
rect 6947 2255 7147 2282
tri 7147 2280 7165 2298 nw
tri 7279 2280 7297 2298 ne
rect 7297 2280 7358 2298
tri 7297 2277 7300 2280 ne
rect 7300 2277 7358 2280
tri 7300 2271 7306 2277 ne
rect 7306 2271 7358 2277
tri 7306 2270 7307 2271 ne
rect 6947 2221 6959 2255
rect 6993 2221 7101 2255
rect 7135 2221 7147 2255
rect 6947 2215 7147 2221
tri 6759 2205 6769 2215 ne
rect 6769 2205 6805 2215
tri 6805 2205 6815 2215 nw
rect 6613 2174 6682 2186
rect 6613 2140 6642 2174
rect 6676 2140 6682 2174
rect 6613 2102 6682 2140
rect 6769 2113 6804 2205
tri 6804 2204 6805 2205 nw
rect 7151 2174 7197 2186
rect 7151 2140 7157 2174
rect 7191 2140 7197 2174
tri 6804 2113 6805 2114 sw
tri 6758 2102 6769 2113 se
rect 6769 2102 6805 2113
tri 6805 2102 6816 2113 sw
rect 7151 2102 7197 2140
rect 6613 2068 6642 2102
rect 6676 2068 6682 2102
tri 6753 2097 6758 2102 se
rect 6758 2097 6816 2102
tri 6816 2097 6821 2102 sw
rect 7151 2097 7157 2102
rect 7191 2097 7197 2102
rect 6613 2056 6682 2068
rect 6718 2045 6724 2097
rect 6776 2045 6791 2097
rect 6843 2045 6849 2097
rect 7109 2045 7115 2097
rect 7167 2045 7182 2068
rect 7234 2045 7240 2097
tri 7305 2064 7307 2066 se
rect 7307 2064 7358 2271
rect 8007 2139 8035 2888
rect 14949 2491 14977 2888
rect 14489 2315 14782 2351
tri 7286 2045 7305 2064 se
rect 7305 2045 7358 2064
tri 7358 2045 7377 2064 sw
rect 7832 2057 7838 2109
rect 7890 2057 7902 2109
rect 7954 2057 7960 2109
rect 14371 2102 14417 2114
rect 14371 2068 14377 2102
rect 14411 2068 14417 2102
rect 859 1921 996 2019
rect 1134 1986 1140 2019
rect 1174 1986 1180 2019
rect 1134 1941 1180 1986
rect 2806 2016 2858 2028
tri 7283 2042 7286 2045 se
rect 7286 2042 7377 2045
tri 7377 2042 7380 2045 sw
rect 7283 1990 7289 2042
rect 7341 1990 7356 2042
rect 7408 1990 7414 2042
rect 14371 2030 14417 2068
rect 14371 1996 14377 2030
rect 14411 1996 14417 2030
rect 14489 2015 14525 2315
rect 14556 2162 14882 2168
rect 14556 2128 14568 2162
rect 14602 2128 14640 2162
rect 14674 2130 14882 2162
rect 14674 2128 14758 2130
rect 14556 2122 14758 2128
rect 14752 2078 14758 2122
rect 14810 2078 14824 2130
rect 14876 2078 14882 2130
rect 14371 1984 14417 1996
rect 14463 2009 14650 2015
rect 14463 1975 14475 2009
rect 14509 1975 14604 2009
rect 14638 1975 14650 2009
rect 14463 1969 14650 1975
rect 2806 1958 2858 1964
rect 1134 1927 1140 1941
rect 1174 1927 1180 1941
rect 859 1887 871 1921
rect 905 1887 950 1921
rect 984 1887 996 1921
rect 859 1881 996 1887
rect 1052 1875 1058 1927
rect 1110 1875 1131 1927
rect 1183 1875 1189 1927
rect 14752 1913 14758 1965
rect 14810 1913 14824 1965
rect 14876 1913 14882 1965
tri 14748 1875 14752 1879 se
tri 14726 1853 14748 1875 se
rect 14748 1853 14752 1875
rect 14541 1847 14752 1853
rect 14541 1813 14553 1847
rect 14587 1813 14625 1847
rect 14659 1813 14752 1847
rect 14541 1806 14752 1813
tri 14723 1777 14752 1806 ne
tri 328 1342 342 1356 ne
rect 342 1348 388 1356
tri 388 1348 396 1356 sw
tri 642 1348 650 1356 se
rect 650 1348 728 1356
rect 342 1342 396 1348
tri 396 1342 402 1348 sw
rect 441 1342 728 1348
tri 342 1341 343 1342 ne
rect 343 1341 402 1342
tri 402 1341 403 1342 sw
tri 343 1323 361 1341 ne
rect 361 1323 403 1341
tri 361 1317 367 1323 ne
rect 215 840 242 841
tri 242 840 243 841 nw
tri 170 829 181 840 se
rect 181 829 231 840
tri 231 829 242 840 nw
rect 24 817 206 829
rect 24 783 30 817
rect 64 804 206 817
tri 206 804 231 829 nw
rect 64 786 188 804
tri 188 786 206 804 nw
rect 64 783 89 786
rect 24 770 89 783
tri 89 770 105 786 nw
rect 367 770 403 1323
rect 441 1308 453 1342
rect 487 1308 526 1342
rect 560 1308 598 1342
rect 632 1308 670 1342
rect 704 1308 728 1342
rect 441 1300 728 1308
rect 784 1329 830 1341
rect 441 1295 595 1300
tri 595 1295 600 1300 nw
rect 784 1295 790 1329
rect 824 1295 830 1329
rect 441 1030 571 1295
tri 571 1271 595 1295 nw
rect 784 1254 830 1295
rect 784 1220 790 1254
rect 824 1220 830 1254
rect 441 996 453 1030
rect 487 996 525 1030
rect 559 996 571 1030
rect 441 990 571 996
rect 623 1186 753 1192
rect 623 1152 635 1186
rect 669 1152 707 1186
rect 741 1152 753 1186
rect 623 874 753 1152
rect 623 840 635 874
rect 669 840 707 874
rect 741 840 753 874
tri 403 770 420 787 sw
rect 24 729 70 770
tri 70 751 89 770 nw
rect 24 695 30 729
rect 64 695 70 729
rect 24 641 70 695
rect 367 728 420 770
tri 420 728 462 770 sw
rect 367 727 462 728
tri 462 727 463 728 sw
rect 367 718 593 727
rect 367 686 475 718
tri 367 684 369 686 ne
rect 369 684 475 686
rect 509 684 547 718
rect 581 684 593 718
tri 369 652 401 684 ne
rect 401 652 593 684
rect 24 607 30 641
rect 64 607 70 641
tri 401 618 435 652 ne
rect 435 618 593 652
rect 24 552 70 607
tri 435 590 463 618 ne
rect 24 518 30 552
rect 64 518 70 552
rect 24 463 70 518
rect 24 429 30 463
rect 64 429 70 463
rect 24 417 70 429
rect 463 406 593 618
rect 463 372 475 406
rect 509 372 547 406
rect 581 372 593 406
rect 463 366 593 372
rect 623 562 753 840
rect 623 528 635 562
rect 669 528 707 562
rect 741 528 753 562
rect 623 282 753 528
rect -6 242 40 254
rect 623 248 635 282
rect 669 248 707 282
rect 741 248 753 282
rect 623 242 753 248
rect 784 1179 830 1220
rect 784 1145 790 1179
rect 824 1145 830 1179
rect 784 1104 830 1145
rect 784 1070 790 1104
rect 824 1070 830 1104
rect 784 1029 830 1070
rect 784 995 790 1029
rect 824 995 830 1029
rect 784 954 830 995
rect 784 920 790 954
rect 824 920 830 954
rect 784 879 830 920
rect 784 845 790 879
rect 824 845 830 879
rect 784 804 830 845
rect 784 770 790 804
rect 824 770 830 804
rect 784 728 830 770
rect 784 694 790 728
rect 824 694 830 728
rect 784 652 830 694
rect 784 618 790 652
rect 824 618 830 652
rect 784 576 830 618
rect 784 542 790 576
rect 824 542 830 576
rect 784 500 830 542
rect 784 466 790 500
rect 824 466 830 500
rect 784 424 830 466
rect 784 390 790 424
rect 824 390 830 424
rect 784 348 830 390
rect 784 314 790 348
rect 824 314 830 348
rect 784 272 830 314
rect -6 208 0 242
rect 34 208 40 242
rect -6 166 40 208
rect 784 238 790 272
rect 824 238 830 272
rect 784 196 830 238
rect -6 132 0 166
rect 34 132 40 166
tri 780 162 784 166 se
rect 784 162 790 196
rect 824 162 830 196
tri 750 132 780 162 se
rect 780 132 830 162
rect -6 120 40 132
rect 616 126 830 132
rect 616 92 628 126
rect 662 92 705 126
rect 739 120 830 126
rect 739 92 790 120
rect 616 86 790 92
rect 824 86 830 120
tri 772 74 784 86 ne
rect 784 74 830 86
<< via1 >>
rect 2736 2299 2788 2351
rect 2800 2299 2852 2351
rect 314 1938 366 1990
rect 314 1865 366 1917
rect 676 1974 728 2026
rect 676 1901 728 1953
rect 865 2019 917 2071
rect 938 2019 990 2071
rect 1058 2019 1110 2071
rect 1131 2020 1183 2071
rect 1131 2019 1140 2020
rect 1140 2019 1174 2020
rect 1174 2019 1183 2020
rect 2806 2028 2858 2080
rect 6697 2255 6749 2271
rect 6697 2221 6703 2255
rect 6703 2221 6737 2255
rect 6737 2221 6749 2255
rect 6697 2219 6749 2221
rect 6765 2219 6817 2271
rect 6833 2255 6885 2271
rect 6833 2221 6845 2255
rect 6845 2221 6879 2255
rect 6879 2221 6885 2255
rect 6833 2219 6885 2221
rect 6724 2045 6776 2097
rect 6791 2045 6843 2097
rect 7115 2068 7157 2097
rect 7157 2068 7167 2097
rect 7182 2068 7191 2097
rect 7191 2068 7234 2097
rect 7115 2045 7167 2068
rect 7182 2045 7234 2068
rect 7838 2057 7890 2109
rect 7902 2057 7954 2109
rect 2806 1964 2858 2016
rect 7289 1990 7341 2042
rect 7356 1990 7408 2042
rect 14758 2078 14810 2130
rect 14824 2078 14876 2130
rect 1058 1875 1110 1927
rect 1131 1907 1140 1927
rect 1140 1907 1174 1927
rect 1174 1907 1183 1927
rect 1131 1875 1183 1907
rect 14758 1913 14810 1965
rect 14824 1913 14876 1965
<< metal2 >>
rect 2730 2299 2736 2351
rect 2788 2299 2800 2351
rect 2852 2329 2858 2351
rect 2852 2299 7713 2329
rect 6691 2219 6697 2271
rect 6749 2219 6765 2271
rect 6817 2219 6833 2271
rect 6885 2219 6891 2271
tri 7211 2097 7223 2109 se
rect 7223 2097 7838 2109
rect 6718 2093 6724 2097
tri 3231 2086 3238 2093 se
rect 3238 2086 6724 2093
rect 2806 2080 2858 2086
rect 676 2026 728 2032
rect 314 1990 366 1996
rect 314 1917 366 1938
rect 676 1953 728 1974
rect 859 2019 865 2071
rect 917 2019 938 2071
rect 990 2019 996 2071
rect 1052 2019 1058 2071
rect 1110 2019 1131 2071
rect 1183 2019 1189 2071
tri 3216 2071 3231 2086 se
rect 3231 2071 6724 2086
tri 3190 2045 3216 2071 se
rect 3216 2045 6724 2071
rect 6776 2045 6791 2097
rect 6843 2093 6849 2097
rect 7109 2093 7115 2097
rect 6843 2045 7115 2093
rect 7167 2045 7182 2097
rect 7234 2074 7838 2097
rect 7234 2057 7252 2074
tri 7252 2057 7269 2074 nw
rect 7832 2057 7838 2074
rect 7890 2057 7902 2109
rect 7954 2057 7960 2109
rect 14752 2078 14758 2130
rect 14810 2078 14824 2130
rect 14876 2078 14882 2130
rect 7234 2045 7240 2057
tri 7240 2045 7252 2057 nw
tri 3187 2042 3190 2045 se
rect 3190 2042 3260 2045
tri 3260 2042 3263 2045 nw
rect 859 2016 996 2019
tri 996 2016 999 2019 sw
rect 2806 2016 2858 2028
tri 3165 2020 3187 2042 se
rect 3187 2020 3238 2042
tri 3238 2020 3260 2042 nw
tri 7261 2020 7283 2042 se
rect 7283 2020 7289 2042
tri 3164 2019 3165 2020 se
rect 3165 2019 3233 2020
rect 859 2015 999 2016
tri 999 2015 1000 2016 sw
rect 859 1991 1000 2015
tri 1000 1991 1024 2015 sw
rect 859 1964 2806 1991
tri 3160 2015 3164 2019 se
rect 3164 2015 3233 2019
tri 3233 2015 3238 2020 nw
tri 7256 2015 7261 2020 se
rect 7261 2015 7289 2020
tri 3135 1990 3160 2015 se
rect 3160 1990 3208 2015
tri 3208 1990 3233 2015 nw
tri 3262 1990 3287 2015 se
rect 3287 1990 7289 2015
rect 7341 1990 7356 2042
rect 7408 1990 7414 2042
tri 3110 1965 3135 1990 se
rect 3135 1966 3184 1990
tri 3184 1966 3208 1990 nw
tri 3238 1966 3262 1990 se
rect 3262 1967 7414 1990
rect 3262 1966 3310 1967
rect 3135 1965 3183 1966
tri 3183 1965 3184 1966 nw
tri 3237 1965 3238 1966 se
rect 3238 1965 3310 1966
tri 3310 1965 3312 1967 nw
rect 14752 1965 14882 2078
rect 859 1958 2858 1964
tri 3103 1958 3110 1965 se
rect 3110 1958 3165 1965
tri 3092 1947 3103 1958 se
rect 3103 1947 3165 1958
tri 3165 1947 3183 1965 nw
tri 3219 1947 3237 1965 se
rect 3237 1947 3287 1965
tri 3087 1942 3092 1947 se
rect 3092 1942 3160 1947
tri 3160 1942 3165 1947 nw
tri 3214 1942 3219 1947 se
rect 3219 1942 3287 1947
tri 3287 1942 3310 1965 nw
tri 3072 1927 3087 1942 se
rect 3087 1927 3145 1942
tri 3145 1927 3160 1942 nw
tri 3199 1927 3214 1942 se
rect 3214 1927 3258 1942
rect 728 1901 1058 1927
tri 366 1875 380 1889 sw
rect 676 1879 1058 1901
rect 1052 1875 1058 1879
rect 1110 1875 1131 1927
rect 1183 1913 3131 1927
tri 3131 1913 3145 1927 nw
tri 3185 1913 3199 1927 se
rect 3199 1913 3258 1927
tri 3258 1913 3287 1942 nw
rect 14752 1913 14758 1965
rect 14810 1913 14824 1965
rect 14876 1913 14882 1965
rect 1183 1895 3113 1913
tri 3113 1895 3131 1913 nw
tri 3167 1895 3185 1913 se
rect 3185 1895 3214 1913
rect 1183 1893 3111 1895
tri 3111 1893 3113 1895 nw
tri 3165 1893 3167 1895 se
rect 3167 1893 3214 1895
rect 1183 1889 3107 1893
tri 3107 1889 3111 1893 nw
tri 3161 1889 3165 1893 se
rect 3165 1889 3214 1893
rect 1183 1879 3097 1889
tri 3097 1879 3107 1889 nw
tri 3151 1879 3161 1889 se
rect 3161 1879 3214 1889
rect 1183 1875 1189 1879
tri 3147 1875 3151 1879 se
rect 3151 1875 3214 1879
rect 366 1869 380 1875
tri 380 1869 386 1875 sw
tri 3141 1869 3147 1875 se
rect 3147 1869 3214 1875
tri 3214 1869 3258 1913 nw
rect 14752 1908 14882 1913
rect 366 1865 386 1869
rect 314 1849 386 1865
tri 386 1849 406 1869 sw
tri 3121 1849 3141 1869 se
rect 3141 1849 3194 1869
tri 3194 1849 3214 1869 nw
rect 314 1844 406 1849
tri 406 1844 411 1849 sw
tri 1223 1844 1228 1849 se
rect 1228 1844 3189 1849
tri 3189 1844 3194 1849 nw
rect 314 1801 3146 1844
tri 3146 1801 3189 1844 nw
rect 314 1796 1268 1801
tri 1268 1796 1273 1801 nw
use sky130_fd_pr__nfet_01v8__example_55959141808484  sky130_fd_pr__nfet_01v8__example_55959141808484_0
timestamp 1648127584
transform 0 -1 712 1 0 137
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808485  sky130_fd_pr__nfet_01v8__example_55959141808485_0
timestamp 1648127584
transform 0 1 894 -1 0 2188
box -28 0 284 97
use sky130_fd_pr__nfet_01v8__example_55959141808513  sky130_fd_pr__nfet_01v8__example_55959141808513_0
timestamp 1648127584
transform 0 -1 712 1 0 417
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808513  sky130_fd_pr__nfet_01v8__example_55959141808513_1
timestamp 1648127584
transform 0 -1 712 -1 0 1297
box -28 0 440 267
use sky130_fd_pr__pfet_01v8__example_55959141808482  sky130_fd_pr__pfet_01v8__example_55959141808482_0
timestamp 1648127584
transform 1 0 6946 0 -1 2173
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808482  sky130_fd_pr__pfet_01v8__example_55959141808482_1
timestamp 1648127584
transform 1 0 6690 0 -1 2173
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808512  sky130_fd_pr__pfet_01v8__example_55959141808512_0
timestamp 1648127584
transform 0 1 14467 1 0 1858
box -28 0 284 97
<< labels >>
flabel comment s 7808 2309 7808 2309 0 FreeSans 280 0 0 0 PGB_AMX_VDDA_H_N(I105 DECODER)
<< properties >>
string GDS_END 48423346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48403670
<< end >>
