magic
tech sky130B
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_0
timestamp 1648127584
transform 1 0 160 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_1
timestamp 1648127584
transform 1 0 376 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_2
timestamp 1648127584
transform 1 0 592 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_0
timestamp 1648127584
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_1
timestamp 1648127584
transform 1 0 808 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 836 97 836 97 0 FreeSans 300 0 0 0 S
flabel comment s 620 97 620 97 0 FreeSans 300 0 0 0 D
flabel comment s 404 97 404 97 0 FreeSans 300 0 0 0 S
flabel comment s 188 97 188 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 3278334
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3275870
<< end >>
