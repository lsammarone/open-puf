magic
tech sky130A
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_0
timestamp 1648127584
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808243  sky130_fd_pr__hvdfm1sd2__example_55959141808243_1
timestamp 1648127584
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 85 128 85 0 FreeSans 300 0 0 0 D
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 31287922
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31286992
<< end >>
