* NGSPICE file created from NBR128_flat.ext - technology: sky130A

.subckt NBR128_flat RESET C[0] C[1] C[2] C[3] C[4] C[5] C[7] C[8] C[9] C[10] C[11]
+ C[12] C[13] C[14] C[15] C[16] C[17] C[18] C[19] C[20] C[21] C[22] C[23] C[24] C[25]
+ C[26] C[27] C[28] C[29] C[30] C[6] C[31] C[32] C[33] C[34] C[35] C[36] C[37] C[38]
+ C[39] C[40] C[41] C[42] C[43] C[44] C[45] C[46] C[47] C[48] C[49] C[50] C[51] C[52]
+ C[53] C[54] C[55] C[56] C[57] C[58] C[59] C[60] C[61] C[62] C[95] C[96] C[97] C[98]
+ C[99] C[100] C[101] C[102] C[103] C[104] C[105] C[106] C[107] C[108] C[109] C[110]
+ C[111] C[112] C[113] C[114] C[115] C[116] C[117] C[118] C[119] C[120] C[121] C[122]
+ C[123] C[124] C[125] C[126] C[127] C[63] C[64] C[65] C[66] C[67] C[68] C[69] C[70]
+ C[71] C[72] C[73] C[74] C[75] C[76] C[77] C[78] C[79] C[80] C[81] C[82] C[83] C[84]
+ C[85] C[86] C[87] C[88] C[89] C[90] C[91] C[92] C[93] C[94] OUT VDD VSS
X0 VDD a_57289_5630# a_57816_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 VSS a_1152_508# a_1102_343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_10168_861# a_11173_1079# a_11113_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_38440_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_34901_18776# a_34477_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X6 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_14574_6924# a_14404_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X8 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_12924_12574# C[101] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_43003_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VDD a_49999_19374# a_49949_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X14 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_33645_13118# a_32526_13079# a_33563_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_59960_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_9025_13912# a_7984_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_3361_13118# a_2324_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VSS a_19535_5630# a_20062_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X21 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_28099_518# a_28143_670# a_27154_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_19087_6923# a_18811_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VSS a_31919_671# a_31935_1080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_37018_1105# a_36594_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X26 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_47002_5835# a_47125_6923# a_47849_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_12772_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_21194_14117# a_20470_12574# a_20347_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_13881_6668# a_13429_6923# a_13030_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_8475_19374# a_8051_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X35 a_1677_1557# a_2616_1406# a_2574_1682# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 VDD a_30634_14118# a_31161_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X39 a_54529_1556# a_54585_1079# a_53580_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 VDD a_6816_507# a_6766_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X41 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_3332_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_26410_12574# a_26134_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 a_1555_13912# a_1242_861# a_1473_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 VSS a_37018_1105# a_36968_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X48 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_10363_19374# a_9939_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X50 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X51 VSS a_53288_13079# a_53811_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X52 a_27899_13118# a_28298_12574# a_28750_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_29000_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_6392_1405# a_7397_1079# a_7341_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 VDD a_17422_13079# a_17945_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X56 VSS a_17714_1406# a_16775_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X57 a_923_19373# a_1013_19128# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X58 a_38253_18584# a_39242_19167# a_39198_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X59 a_1444_19298# a_1504_18801# a_1013_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X60 a_40074_14117# a_39350_12574# a_39227_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 a_33242_507# a_32818_862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X62 a_54525_518# a_54585_1079# a_53580_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X63 a_41962_14117# a_41238_12574# a_41115_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 VSS a_28975_5630# a_29502_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X66 a_11993_6668# a_11265_6923# a_11142_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 VDD a_28750_13079# a_29273_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X69 a_8009_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_9107_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 VSS a_40370_861# a_39427_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X73 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X74 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X75 VDD a_51629_6668# a_52152_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X76 a_22435_518# a_23378_861# a_23336_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_45091_518# a_45135_670# a_44146_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 VDD a_36302_13079# a_36825_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X79 a_28251_6923# C[45] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X80 a_36079_6923# a_35803_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X81 a_11989_5630# a_11265_6923# a_11142_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X83 a_19797_18776# a_19373_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X84 a_27874_18261# a_28813_18040# a_28771_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X85 VDD a_21914_507# a_21864_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X86 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X87 VSS a_13715_18040# a_12776_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X88 a_18344_6924# a_18174_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X89 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X90 a_38253_18584# a_39258_18802# a_39198_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X91 a_46744_19298# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X92 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X93 a_52093_13117# a_51923_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X94 a_53981_13117# a_53811_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X95 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X96 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X97 a_53580_861# a_54569_670# a_54525_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X98 a_33538_18261# a_34477_18040# a_34435_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 a_48636_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X100 a_20347_13912# a_19306_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X101 a_50778_6629# a_49741_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X102 VSS a_27578_1105# a_27528_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X103 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X104 VSS a_4275_18040# a_3336_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X105 a_9377_6923# C[35] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 a_42682_507# a_42258_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X107 VDD a_2811_18776# a_2761_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X108 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X109 a_24123_13912# a_24246_12574# a_24970_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X110 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_56295_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X111 a_11113_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X112 a_26011_13912# a_26134_12574# a_26858_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X113 a_20470_12574# C[105] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 a_1242_317# a_1733_1080# a_1673_519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X116 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X117 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X118 a_33563_13912# a_32522_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X119 a_16462_6379# a_16292_6379# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X120 a_38677_18776# a_38253_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X121 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_26240_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X122 a_14918_5834# a_15041_6922# a_15765_5629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X123 VSS a_10928_19167# a_10944_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X124 a_27899_13912# a_28298_12574# a_28746_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X125 a_17651_6668# a_17199_6923# a_16800_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X126 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_24352_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X127 VSS a_23802_1105# a_23752_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X128 a_11117_1556# a_11157_670# a_10168_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X129 a_10884_19299# a_11827_18584# a_11785_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 a_45992_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X132 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X133 VSS a_23149_18584# a_22206_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X134 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_17418_14117# a_16970_12574# a_16571_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X136 a_33563_13912# a_33962_12574# a_34410_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X137 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X138 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X139 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 VDD a_50228_1105# a_50178_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X141 a_13001_518# a_13061_1079# a_12056_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X142 a_15603_18040# a_16602_18801# a_16546_18260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X143 a_39112_6924# a_38942_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X144 a_23082_14117# a_22634_12574# a_22235_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X145 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X146 a_18811_6923# C[40] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X147 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X148 a_25461_18776# a_25037_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X149 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X150 a_24970_14117# a_24522_12574# a_24123_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X151 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X152 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X153 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X154 a_60071_13119# a_58952_13079# a_59989_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X156 a_26858_14117# a_26134_12574# a_26011_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 a_31125_18775# a_30701_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X159 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X160 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X161 VDD C[65] a_56457_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X162 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X163 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X164 a_56098_6380# a_55928_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X165 VSS a_42029_18584# a_41086_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X166 a_53309_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X167 VDD a_14139_19374# a_14089_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X168 VSS a_43917_18584# a_42974_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X169 a_28813_18040# a_29818_18802# a_29762_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X170 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 a_8996_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X172 a_28210_6629# a_27091_6668# a_28128_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X173 a_35336_6924# a_35166_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X174 VSS C[64] a_58345_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X175 a_14139_19374# a_13715_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X176 a_37339_13118# a_36302_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X177 VSS a_57064_13079# a_57587_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X178 a_44341_18776# a_43917_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X179 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X180 a_43850_14117# a_43402_12574# a_43003_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X181 VSS a_15769_6667# a_16292_6923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X182 VSS a_44570_1105# a_44520_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X183 VSS a_3605_670# a_3621_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X184 a_48861_518# a_48905_670# a_47916_1406# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X185 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X186 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X187 a_29991_1556# a_30047_1079# a_29042_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X188 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X189 a_6587_19374# a_6163_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X190 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X191 VSS a_25266_1405# a_24327_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X192 VDD a_31354_508# a_31304_343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X193 a_30659_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X194 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X195 a_24434_6629# a_23315_6668# a_24352_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X196 a_27154_1405# a_28143_670# a_28103_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X197 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_43232_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X198 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X199 a_34643_6668# a_34191_6923# a_33792_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X200 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X201 a_21891_12573# a_21721_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X202 a_7765_6923# a_7489_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X203 VSS a_18138_507# a_18088_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X204 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X205 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 a_47687_18583# a_48692_18802# a_48632_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X207 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X208 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X209 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X210 VDD a_49512_13079# a_50035_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X211 VDD a_51400_13079# a_51923_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X212 VSS a_55405_6668# a_55928_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X213 VSS a_54004_507# a_53954_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X214 a_61090_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X215 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_44973_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X216 a_45243_6922# C[54] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X217 a_50948_12574# a_50672_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X218 a_26240_6629# a_26363_6923# a_27091_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X219 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X220 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X221 a_35803_6923# C[49] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X222 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X223 a_53351_18584# a_54356_18802# a_54296_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X224 a_57757_13117# a_57587_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X225 a_10798_6380# a_10628_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X226 VDD a_16815_671# a_16831_1080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X227 a_49762_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X228 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X229 a_25896_6924# a_25726_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X230 a_51177_6923# a_50901_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X231 a_1152_1106# a_1242_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X232 a_3561_518# a_3605_670# a_2616_1406# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 VSS a_9939_18040# a_9000_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X234 VDD a_60903_18584# a_63251_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X235 VSS a_17909_19374# a_17859_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X236 VSS a_9872_14117# a_10399_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X237 a_38415_5630# a_37967_6923# a_37568_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X238 a_36527_5630# a_35803_6923# a_35680_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X239 VSS a_17485_18583# a_16542_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X240 a_26240_5835# a_26363_6923# a_27087_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X241 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 a_40771_12573# a_40601_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X243 a_32755_6668# a_32027_6923# a_31904_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X244 a_20658_5835# a_19535_5630# a_20576_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X245 a_16771_519# a_16831_1080# a_15832_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X246 a_10569_13117# a_10399_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X247 a_24246_12574# C[107] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X248 a_39538_5835# a_38415_5630# a_39456_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X249 a_48340_507# a_47916_862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X250 VDD a_16021_18775# a_15971_18610# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X251 a_29042_861# a_30031_670# a_29987_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X252 VSS a_23573_19374# a_23523_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X253 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X254 VDD a_36527_5630# a_37054_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X255 a_1677_1557# a_1717_671# a_1242_317# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X256 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X257 a_53775_18776# a_53351_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X258 a_16233_13118# a_16063_13118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X259 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X260 VSS a_61069_6667# a_60189_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X261 a_31798_12574# C[111] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X262 a_17909_18776# a_17485_18039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X263 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X264 a_3017_13117# a_2847_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X265 VDD a_35466_19167# a_35482_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X266 VDD a_37354_19167# a_37370_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X267 a_43631_6923# a_43355_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X268 VSS a_49804_861# a_48861_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X269 VSS a_7152_19167# a_7168_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X270 a_48636_18261# a_48692_18802# a_47687_18583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X271 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X272 VSS a_8213_5630# a_8740_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X273 VSS a_42258_1405# a_41319_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X274 a_38253_18040# a_39242_19167# a_39202_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X275 a_6329_6668# a_5877_6923# a_5478_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X276 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 a_13652_13079# a_12924_12574# a_12801_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X278 a_59989_13913# a_58948_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X279 VDD a_20026_507# a_19976_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X280 a_44146_1405# a_45135_670# a_45095_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X281 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X282 VSS a_48340_1105# a_48290_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X283 VDD a_44570_507# a_44520_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X284 a_29237_18776# a_28813_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X285 a_24352_5835# a_24751_6923# a_25199_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X286 VSS C[77] a_33807_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X287 VSS a_42453_19374# a_42403_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X288 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X289 a_8681_12573# a_8511_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X290 a_45014_12575# C[118] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X291 VDD a_43247_670# a_43263_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X292 VDD a_36789_18776# a_36739_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X293 a_4212_13079# a_3484_12574# a_3361_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X294 a_12801_13118# a_12924_12574# a_13652_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X295 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_48661_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X296 a_17443_18859# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X297 VSS C[19] a_24138_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X298 a_36789_18776# a_36365_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X299 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_26322_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X300 a_45967_5629# a_45243_6922# a_45120_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X301 VSS a_45135_670# a_45151_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X302 a_45805_18584# a_46788_19166# a_46744_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X303 a_12883_13118# a_11764_13079# a_12801_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X304 a_3361_13118# a_3484_12574# a_4212_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X305 a_41426_5835# a_40303_5630# a_41344_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X306 a_57780_507# a_57356_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X307 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_7137_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X308 a_43232_6629# a_43355_6923# a_44083_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X309 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_47002_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X310 a_28975_5630# a_28527_6923# a_28128_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X311 a_8704_507# a_8280_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X312 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X313 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X314 a_8213_5630# a_7489_6923# a_7366_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X315 a_21914_1105# a_21490_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X316 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X317 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X318 VSS C[13] a_35466_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X319 a_4441_6668# a_3713_6923# a_3590_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X320 a_42888_6924# a_42718_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X321 VDD a_27087_5630# a_27614_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X322 a_27578_1105# a_27154_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X323 VDD C[2] a_56228_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X324 a_42216_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X325 VSS a_51692_861# a_50749_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X326 a_26215_1556# a_26255_670# a_25266_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X327 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X328 a_57127_18584# a_58116_19167# a_58072_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X329 VDD C[1] a_58116_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X330 VSS C[9] a_43018_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X331 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X332 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X333 VDD a_47620_14117# a_48147_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X334 a_4437_5630# a_3713_6923# a_3590_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X335 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_16882_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X336 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X337 a_31986_6629# a_30867_6667# a_31904_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X338 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X339 a_41344_6629# a_41743_6923# a_42195_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X340 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X341 a_25667_12573# a_25497_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X342 a_48784_12574# C[120] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X343 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X344 a_39309_13912# a_38186_14117# a_39227_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X345 a_53580_861# a_54585_1079# a_54525_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X346 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X347 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X348 VSS a_61065_5629# a_61592_6379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X349 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_60071_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X350 a_52641_1556# a_53580_1405# a_53538_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 a_3561_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X352 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X353 a_59181_6668# a_58729_6923# a_58330_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X354 a_23802_507# a_23378_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X355 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X356 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X357 a_41344_5835# a_41743_6923# a_42191_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X358 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X359 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X360 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X361 VSS a_13648_14117# a_14175_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X362 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X363 a_50901_6923# C[57] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X364 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_43314_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X365 a_44547_12573# a_44377_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X366 VSS a_57551_18776# a_57501_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X367 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_16653_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X368 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X369 VSS a_57289_5630# a_57816_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X370 a_25266_861# a_26271_1079# a_26211_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X371 a_24323_518# a_24383_1079# a_23378_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X372 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X373 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X374 a_61065_5629# a_60341_6922# a_60218_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X375 VDD a_46452_508# a_46402_343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X376 VSS a_6096_14117# a_6623_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X377 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_37650_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X378 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X379 a_50549_13912# a_50672_12574# a_51396_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X380 a_31331_13118# a_31161_13118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X381 a_54210_6924# a_54040_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X382 VDD a_44079_5630# a_44606_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X383 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 a_14889_518# a_15832_861# a_15790_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 VDD a_50564_19167# a_50580_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X386 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X387 a_57293_6668# a_56565_6923# a_56442_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X388 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_27981_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X389 a_56565_6923# C[60] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X390 VSS a_49999_19374# a_49949_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X391 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X392 a_3672_6629# a_1013_19128# a_3590_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X393 a_53351_18040# a_54340_19167# a_54300_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X394 a_20547_518# a_20607_1079# a_19602_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X395 a_56184_19299# a_56228_19167# a_55239_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X396 VDD a_21427_6668# a_21950_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X397 a_14889_518# a_14933_670# a_13944_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 VDD a_21685_19374# a_21635_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X399 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X400 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35533_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X401 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_33874_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X402 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X403 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X404 a_50434_6924# a_50264_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X405 a_57289_5630# a_56565_6923# a_56442_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X406 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X407 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X408 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X409 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X410 a_9876_13079# a_9148_12574# a_9025_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X411 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X412 VSS a_55892_1105# a_55842_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X413 a_12801_13912# a_11760_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X414 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_31675_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X415 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_14689_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X416 a_33792_5835# a_33915_6923# a_34639_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X417 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X418 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X419 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X420 a_49999_18776# a_49575_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X421 a_51887_18776# a_51463_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X422 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X423 a_37539_518# a_38482_861# a_38440_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X424 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X425 a_2616_1406# a_3605_670# a_3565_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X426 VDD a_33013_19374# a_32963_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X427 a_47687_18039# a_48692_18802# a_48636_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X428 a_9025_13118# a_9148_12574# a_9876_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X429 a_37568_5835# a_36527_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X430 VSS a_6816_507# a_6766_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X431 VDD a_34901_19374# a_34851_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X432 VSS C[90] a_9269_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X433 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X434 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X435 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X436 a_56213_13118# a_55176_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X437 a_56413_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X438 VDD a_40565_19374# a_40515_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X439 VSS C[5] a_50564_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X440 a_19331_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X441 a_53351_18040# a_54356_18802# a_54300_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X442 a_7219_13118# a_6100_13079# a_7137_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X443 VDD a_1488_19166# a_1504_18801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X444 VSS a_17422_13079# a_17945_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X445 a_31879_1557# a_31935_1080# a_30930_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X446 a_10363_19374# a_9939_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X447 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X448 a_33242_507# a_32818_862# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X449 a_37543_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X450 VSS a_15603_18584# a_14660_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X451 a_26883_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X452 a_15790_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X453 a_923_19373# a_1013_19128# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X454 a_46452_1106# a_46034_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X455 a_41315_518# a_41375_1079# a_40370_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X456 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X457 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X458 a_32547_18065# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X459 a_48743_13912# a_47620_14117# a_48661_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X460 VSS a_28750_13079# a_29273_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X461 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X462 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X463 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X464 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X465 VSS a_6163_18584# a_5220_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X466 VDD a_59668_507# a_59618_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X467 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_47084_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X468 VSS C[69] a_48905_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X469 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X470 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X471 a_34664_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X472 VDD a_58345_670# a_58361_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X473 a_18663_1556# a_18703_670# a_17714_862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X474 a_54407_13912# a_53284_14117# a_54325_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X475 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_5560_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X476 a_7366_6629# a_6329_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X477 VSS a_36302_13079# a_36825_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X478 a_59874_6924# a_59704_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X479 a_49737_5630# a_49289_6923# a_48890_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X480 a_6096_14117# a_5648_12574# a_5249_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X481 a_7984_14117# a_7536_12574# a_7137_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X482 a_20347_13118# a_20746_12574# a_21198_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X483 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X484 a_48632_19299# a_48692_18802# a_47687_18039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X485 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X486 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X487 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_52666_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X488 VSS a_21914_507# a_21864_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X489 a_45763_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X490 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X491 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X492 a_56524_6629# a_55405_6668# a_56442_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X493 VDD a_14368_1105# a_14318_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X494 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X495 a_9872_14117# a_9148_12574# a_9025_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X496 VDD a_47849_5630# a_48376_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X497 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X498 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X499 VSS a_15832_861# a_14889_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X500 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_10995_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X501 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_12883_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X502 a_16771_519# a_17714_862# a_17672_888# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X503 VSS a_2811_18776# a_2761_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X504 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X505 VDD a_23086_13079# a_23609_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X506 a_54953_6923# a_54677_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X507 a_38906_1105# a_38482_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X508 VSS a_14368_1105# a_14318_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X509 a_22634_12574# a_22358_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X510 a_57314_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X511 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_3443_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X512 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X513 a_29443_13117# a_29273_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X514 a_23779_12573# a_23609_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X515 a_39227_13118# a_39626_12574# a_40078_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X516 a_52748_6629# a_51629_6668# a_52666_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X517 a_55468_1405# a_56457_670# a_56417_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X518 a_25037_18584# a_26042_18802# a_25982_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X519 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X520 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_16571_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X521 a_20322_18261# a_21261_18040# a_21219_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X522 a_35107_13117# a_34937_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X523 a_36995_13117# a_36825_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X524 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_13030_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X525 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_11142_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X526 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X527 VDD a_48111_18776# a_48061_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X528 a_57127_18040# a_58116_19167# a_58076_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X529 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X530 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X531 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X532 VDD a_41966_13079# a_42489_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X533 a_54554_6629# a_54677_6923# a_55405_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X534 a_17714_862# a_18719_1079# a_18659_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X535 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X536 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X537 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X538 a_25461_18776# a_25037_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X539 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_29787_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X540 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_50631_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X541 a_42659_12573# a_42489_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X542 a_15041_6922# C[38] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X543 a_5453_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X544 a_31675_13118# a_31798_12574# a_32526_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X545 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X546 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X547 a_31125_18775# a_30701_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X548 VDD a_55663_18776# a_55613_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X549 a_39202_18261# a_40141_18040# a_40099_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X550 a_13429_6923# a_13153_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X551 a_19560_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X552 a_20347_13912# a_20746_12574# a_21194_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X553 a_56098_6380# a_55928_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X554 a_61069_6667# a_60341_6922# a_60218_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X555 VDD C[91] a_7381_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X556 a_31757_13118# a_30638_13080# a_31675_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X557 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_58412_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X558 VDD a_14704_19167# a_14720_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X559 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X560 a_7137_13912# a_6096_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X561 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_61959_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X562 a_48632_19299# a_49575_18584# a_49533_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X563 a_1473_13118# a_1242_317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X564 a_45120_5834# a_44079_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X565 VSS a_14139_19374# a_14089_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X566 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X567 a_44341_18776# a_43917_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X568 a_14139_19374# a_13715_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X569 a_7260_12574# C[98] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X570 a_52666_6629# a_53065_6923# a_53517_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X571 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X572 VDD C[23] a_16586_19166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X573 VSS a_30701_18584# a_29758_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_39227_13912# a_39626_12574# a_40074_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X575 a_44973_13119# a_43854_13079# a_44891_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X576 OUT a_63251_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X577 VSS a_31354_508# a_31304_343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X578 a_17485_18583# a_18474_19167# a_18430_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X579 a_10884_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X580 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X581 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X582 a_6587_19374# a_6163_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X583 a_44146_861# a_45135_670# a_45091_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X584 VSS a_19602_861# a_18659_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X585 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X586 a_54004_1105# a_53580_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X587 VSS a_12056_1405# a_11117_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X588 VDD a_16250_1106# a_16200_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X589 a_6816_1105# a_6392_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X590 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X591 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X592 a_52666_5835# a_53065_6923# a_53513_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X593 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X594 a_24522_12574# a_24246_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X595 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_39227_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X596 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X597 VSS a_18138_1105# a_18088_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X598 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X599 VSS C[24] a_14704_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X600 VSS a_49512_13079# a_50035_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X601 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X602 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X603 VSS a_51400_13079# a_51923_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X604 VDD a_38419_6668# a_38942_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X605 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_54636_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X606 VDD C[83] a_22479_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X607 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X608 a_26011_13118# a_26410_12574# a_26862_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X609 a_60861_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X610 VSS a_42195_6668# a_42718_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X611 a_50228_1105# a_49804_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X612 VDD a_35130_507# a_35080_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X613 a_36365_18584# a_37354_19167# a_37310_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X614 a_15765_5629# a_15041_6922# a_14918_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X615 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_60218_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X616 a_11224_5835# a_10101_5630# a_11142_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X617 VSS C[82] a_24367_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X618 a_39202_18261# a_39242_19167# a_38253_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X619 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X620 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X621 VSS a_60903_18584# a_63251_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X622 a_36552_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X623 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X624 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X625 a_43402_12574# a_43126_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X626 a_45095_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X627 VDD a_26862_13079# a_27385_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X628 a_12686_6924# a_12516_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X629 a_46977_1557# a_47033_1080# a_46034_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X630 a_48340_507# a_47916_862# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X631 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X632 a_28022_12574# C[109] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X633 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X634 VSS a_16021_18775# a_15971_18610# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X635 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X636 VSS a_21490_861# a_20547_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X637 a_36594_1405# a_37599_1079# a_37543_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X638 a_57064_13079# a_56612_12574# a_56213_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X639 VSS a_36527_5630# a_37054_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X640 a_26211_518# a_26255_670# a_25266_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X641 VDD a_34414_13079# a_34937_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X642 a_26639_6923# a_26363_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X643 a_17199_6923# a_16923_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X644 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X645 a_17909_18776# a_17485_18039# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X646 a_24098_18261# a_25037_18040# a_24995_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X647 a_25986_18261# a_26925_18040# a_26883_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X648 VSS a_11827_18040# a_10888_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X649 VSS a_45738_14118# a_46265_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X650 a_36365_18584# a_37370_18802# a_37310_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X651 a_50205_13117# a_50035_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X652 a_18138_1105# a_17714_1406# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X653 a_46748_18260# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X654 a_39350_12574# C[115] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X655 VDD a_56457_670# a_56473_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X656 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X657 a_16571_13912# a_16694_12574# a_17418_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X658 a_49762_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X659 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X660 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X661 a_48890_5835# a_47849_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X662 VSS a_20026_507# a_19976_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X663 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X664 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X665 a_11993_6668# a_11541_6923# a_11142_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X666 VSS a_44570_507# a_44520_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X667 a_29237_18776# a_28813_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X668 VDD a_9269_670# a_9285_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X669 a_16542_19298# a_16586_19166# a_15603_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X670 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X671 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_54407_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X672 VSS a_30863_5629# a_31390_6379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X673 a_6816_1105# a_6392_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X674 VSS a_36789_18776# a_36739_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X675 a_22235_13912# a_22358_12574# a_23082_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X676 a_8681_12573# a_8511_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X677 a_5453_1556# a_5493_670# a_4504_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X678 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X679 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X680 a_39427_518# a_40370_861# a_40328_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X681 a_59668_1105# a_59244_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X682 VSS a_35130_1105# a_35080_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X683 VDD a_24138_19167# a_24154_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X684 a_36789_18776# a_36365_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X685 a_44866_18261# a_45805_18040# a_45763_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X686 a_24123_13912# a_24522_12574# a_24970_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X687 a_31675_13912# a_30634_14118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X688 a_29869_13119# a_28750_13079# a_29787_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X689 a_48317_13117# a_48147_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X690 a_11142_5835# a_11541_6923# a_11989_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X691 a_26011_13912# a_26410_12574# a_26858_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X692 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X693 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X694 a_8704_507# a_8280_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X695 VDD a_29802_19167# a_29818_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X696 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_13112_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X697 a_52637_518# a_52697_1079# a_51692_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X698 a_31675_13912# a_32074_12574# a_32522_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X699 VDD a_53517_6668# a_54040_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X700 a_46034_861# a_47017_671# a_46973_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X701 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X702 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X703 VDD a_6329_6668# a_6852_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X704 a_50228_507# a_49804_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X705 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X706 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X707 a_44891_13913# a_43850_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X708 VSS a_27087_5630# a_27614_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X709 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X710 a_41115_13912# a_41238_12574# a_41962_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X711 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X712 a_43003_13912# a_43126_12574# a_43850_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X713 a_23573_18776# a_23149_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X714 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X715 a_60300_5834# a_59177_5630# a_60218_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X716 a_30930_861# a_31935_1080# a_31875_519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X717 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X718 VDD a_43018_19167# a_43034_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X719 VDD a_13877_5630# a_14404_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X720 a_14660_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X721 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X722 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X723 a_27091_6668# a_26363_6923# a_26240_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X724 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X725 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X726 VDD a_49741_6668# a_50264_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X727 a_26363_6923# C[44] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X728 a_61762_6923# a_61592_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X729 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X730 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X731 VSS C[68] a_50793_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X732 a_45095_1556# a_45151_1079# a_44146_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X733 VDD a_10592_507# a_10542_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X734 VDD a_12251_19374# a_12201_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X735 a_25037_18040# a_26042_18802# a_25986_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X736 a_26925_18040# a_27930_18802# a_27874_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X737 a_28298_12574# a_28022_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X738 VDD a_60233_670# a_60249_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X739 a_20551_1556# a_20591_670# a_19602_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X740 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X741 a_5220_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X742 a_7108_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X743 a_48865_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X744 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_54325_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X745 a_20232_6924# a_20062_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X746 a_27087_5630# a_26363_6923# a_26240_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X747 a_4504_861# a_5509_1079# a_5449_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X748 VSS C[16] a_29802_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X749 a_41962_14117# a_41514_12574# a_41115_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X750 VSS a_25690_1105# a_25640_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X751 a_42453_18776# a_42029_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X752 VSS a_11157_670# a_11173_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X753 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X754 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X755 a_7489_6923# C[34] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X756 a_23802_507# a_23378_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X757 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X758 a_36594_861# a_37583_670# a_37539_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X759 a_4699_19374# a_4275_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X760 a_51463_18584# a_52452_19167# a_52408_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X761 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X762 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X763 a_49512_13079# a_49060_12574# a_48661_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X764 a_39431_1556# a_40370_1405# a_40328_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X765 a_54300_18261# a_54340_19167# a_53351_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X766 a_26093_13912# a_24970_14117# a_26011_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_24352_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X768 a_27981_13912# a_26858_14117# a_27899_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X769 a_26211_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X770 a_28099_518# a_29042_861# a_29000_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X771 VSS a_21914_1105# a_21864_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X772 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X773 a_2324_13079# a_1872_12574# a_1473_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X774 VSS a_32818_1406# a_31879_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X775 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X776 VSS a_46452_508# a_46402_343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X777 VSS a_33807_670# a_33823_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X778 VDD a_55172_14117# a_55699_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X779 a_16250_1106# a_15832_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X780 a_37224_6924# a_37054_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X781 VSS a_44079_5630# a_44606_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X782 a_11113_518# a_11173_1079# a_10168_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X783 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X784 a_16923_6923# C[39] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X785 VDD a_59181_6668# a_59704_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X786 a_51463_18584# a_52468_18802# a_52408_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X787 a_55869_13117# a_55699_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X788 VSS a_60836_14118# a_61363_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X789 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X790 a_15769_6667# a_15041_6922# a_14918_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X791 VDD a_40794_1105# a_40744_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X792 a_19602_861# a_20607_1079# a_20547_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X793 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X794 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X795 a_44083_6668# a_43355_6923# a_43232_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X796 a_39198_19299# a_39258_18802# a_38253_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X797 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X798 a_17485_18039# a_18474_19167# a_18434_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X799 a_29672_6924# a_29502_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X800 a_43355_6923# C[53] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X801 a_19535_5630# a_19087_6923# a_18688_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X802 VSS a_17485_18039# a_16546_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X803 a_29787_13913# a_28746_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X804 a_60388_12575# a_60112_12575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X805 a_62000_12574# C[127] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X806 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X807 a_27899_13912# a_28022_12574# a_28746_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X808 a_22358_12574# C[106] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X809 a_41000_6380# a_40830_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X810 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_22464_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X811 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X812 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X813 a_33448_6924# a_33278_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X814 VSS a_21685_19374# a_21635_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X815 a_26322_6629# a_25203_6668# a_26240_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X816 a_49999_18776# a_49575_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X817 VDD a_17647_5630# a_18174_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X818 a_51887_18776# a_51463_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X819 a_59964_18261# a_60903_18040# a_60861_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X820 a_44079_5630# a_43355_6923# a_43232_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X821 VSS a_42682_1105# a_42632_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X822 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X823 a_33763_518# a_33807_670# a_32818_1406# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X824 a_46748_18260# a_46804_18801# a_45805_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X825 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X826 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X827 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X828 a_14345_12573# a_14175_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X829 a_24751_6923# a_24475_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X830 a_31354_1106# a_30930_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X831 VSS a_23378_1405# a_22439_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X832 VSS a_5264_19167# a_5280_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X833 VSS a_33013_19374# a_32963_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X834 VSS a_34901_19374# a_34851_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X835 VDD a_27349_18776# a_27299_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X836 a_36365_18040# a_37354_19167# a_37314_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X837 a_11764_13079# a_11036_12574# a_10913_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X838 a_39198_19299# a_39242_19167# a_38253_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X839 a_22546_6629# a_21427_6668# a_22464_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X840 a_25266_1405# a_26255_670# a_26215_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X841 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X842 a_41238_12574# C[116] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X843 a_27349_18776# a_26925_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X844 a_43203_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X845 VSS a_40565_19374# a_40515_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X846 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X847 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X848 a_6793_12573# a_6623_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X849 a_10913_13118# a_11036_12574# a_11764_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X850 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X851 a_29758_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X852 a_58076_18261# a_58132_18802# a_57127_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X853 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X854 a_2324_13079# a_1596_12574# a_1473_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X855 a_5877_6923# a_5601_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X856 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X857 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X858 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X859 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X860 VSS a_59668_507# a_59618_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X861 a_4928_1105# a_4504_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X862 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X863 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X864 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_5249_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X865 a_10995_13118# a_9876_13079# a_10913_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X866 a_24352_6629# a_24475_6923# a_25203_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X867 a_46748_18260# a_46788_19166# a_45805_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X868 a_33915_6923# C[48] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X869 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X870 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_58101_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X871 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X872 VDD C[6] a_48676_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X873 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X874 a_39227_13118# a_38190_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X875 a_59244_1405# a_60249_1079# a_60193_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X876 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X877 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X878 VSS C[14] a_33578_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X879 a_24008_6924# a_23838_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X880 VDD a_8475_19374# a_8425_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X881 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X882 a_5134_6924# a_4964_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X883 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X884 a_36527_5630# a_36079_6923# a_35680_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X885 VDD a_29466_1105# a_29416_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X886 VDD C[3] a_54340_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X887 VSS a_47849_5630# a_48376_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X888 a_47916_1406# a_48921_1079# a_48865_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X889 VSS C[10] a_41130_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X890 a_55239_18584# a_56228_19167# a_56184_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X891 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X892 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X893 a_58076_18261# a_58116_19167# a_57127_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X894 a_30139_6922# C[46] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X895 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_28210_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X896 a_20576_6629# a_20699_6923# a_21427_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X897 a_43314_6629# a_42195_6668# a_43232_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X898 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X899 a_59015_18040# a_60020_18802# a_59964_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 VDD a_34639_5630# a_35166_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X901 a_46664_6379# a_46494_6379# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X902 a_45120_5834# a_45519_6922# a_45967_5629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X903 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X904 VSS a_23086_13079# a_23609_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X905 a_62276_12574# a_62000_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X906 a_38906_507# a_38482_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X907 VDD RESET a_28116_9428# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X908 a_23779_12573# a_23609_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X909 a_46896_12574# C[119] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X910 a_22464_6629# a_22863_6923# a_23315_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X911 a_8213_5630# a_7765_6923# a_7366_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X912 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X913 a_11760_14117# a_11036_12574# a_10913_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X914 a_41743_6923# a_41467_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X915 VDD a_22479_670# a_22495_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X916 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X917 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X918 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X919 VDD a_58948_14117# a_59475_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X920 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X921 a_4441_6668# a_3989_6923# a_3590_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X922 a_20026_1105# a_19602_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X923 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X924 a_44570_1105# a_44146_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X925 a_42258_1405# a_43247_670# a_43207_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X926 VDD a_25690_507# a_25640_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X927 a_2320_14117# a_1596_12574# a_1473_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X928 a_51650_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X929 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X930 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X931 a_22464_5835# a_22863_6923# a_23311_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X932 VDD a_24367_670# a_24383_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X933 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X934 VSS a_48111_18776# a_48061_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X935 VSS a_41966_13079# a_42489_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X936 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X937 a_5601_6923# C[33] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X938 a_29987_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X939 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X940 VSS a_11760_14117# a_12287_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X941 a_60193_1556# a_61065_5629# a_61090_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X942 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X943 a_42659_12573# a_42489_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X944 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_24434_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X945 VSS a_26255_670# a_26271_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X946 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X947 a_58729_6923# a_58453_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X948 VSS a_55663_18776# a_55613_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X949 a_41344_6629# a_41467_6923# a_42195_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X950 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X951 a_20026_1105# a_19602_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X952 a_48865_1556# a_49804_1405# a_49762_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X953 a_16542_19298# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X954 a_7137_13118# a_7536_12574# a_7988_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X955 a_6325_5630# a_5601_6923# a_5478_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X956 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_30016_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X957 a_46973_519# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X958 VDD a_19797_18776# a_19747_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X959 VSS a_4208_14117# a_4735_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X960 a_9025_13118# a_9424_12574# a_9876_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X961 a_15000_5834# a_13877_5630# a_14918_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X962 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X963 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X964 a_9336_5835# a_8213_5630# a_9254_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X965 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X966 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X967 VDD a_25199_5630# a_25726_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X968 VDD C[75] a_37583_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X969 a_16250_508# a_15832_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X970 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X971 a_48632_19299# a_48676_19167# a_47687_18039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X972 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_26093_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X973 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X974 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X975 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X976 a_51463_18040# a_52452_19167# a_52412_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X977 VSS a_48905_670# a_48921_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X978 a_54296_19299# a_54340_19167# a_53351_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X979 a_61877_13912# a_62000_12574# a_60903_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X980 a_1448_18260# a_2387_18039# a_2345_18065# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X981 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_33645_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X982 a_30098_6628# a_28979_6668# a_30016_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X983 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X984 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X985 a_11117_1556# a_11173_1079# a_10168_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X986 VDD a_38677_18776# a_38627_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X987 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X988 a_7988_13079# a_7260_12574# a_7137_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X989 a_39456_6629# a_39855_6923# a_40307_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X990 a_42258_861# a_43263_1079# a_43203_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X991 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X992 a_7112_18261# a_8051_18040# a_8009_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X993 a_10913_13912# a_9872_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X994 VDD a_55892_1105# a_55842_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X995 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X996 a_48661_13118# a_47624_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X997 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X998 a_47084_6629# a_45971_6667# a_47002_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X999 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1000 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1001 a_18688_5835# a_17647_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1002 a_50753_1556# a_51692_1405# a_51650_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1003 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1004 a_57293_6668# a_56841_6923# a_56442_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1005 a_39456_5835# a_39855_6923# a_40303_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1006 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1007 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1008 a_54325_13118# a_53288_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1009 a_54525_518# a_54569_670# a_53580_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1010 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1011 a_29466_1105# a_29042_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1012 a_8910_6924# a_8740_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1013 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1014 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1015 VSS a_35130_507# a_35080_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1016 VSS a_30930_1405# a_29991_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1017 a_3336_18261# a_3376_19167# a_2387_18583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1018 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1019 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1020 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_41426_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1021 VSS a_13715_18584# a_12772_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1022 a_23107_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1023 a_24995_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1024 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1025 a_7137_13912# a_7536_12574# a_7984_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1026 a_46452_1106# a_46034_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1027 a_22435_518# a_22495_1079# a_21490_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1028 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1029 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1030 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1031 a_48632_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1032 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1033 a_46855_13912# a_45738_14118# a_46773_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1034 VSS a_26862_13079# a_27385_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1035 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1036 VSS a_4275_18584# a_3332_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1037 a_13648_14117# a_13200_12574# a_12801_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1038 a_52322_6924# a_52152_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1039 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1040 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1041 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1042 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1043 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1044 a_55405_6668# a_54677_6923# a_54554_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1045 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1046 a_52519_13912# a_51396_14117# a_52437_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1047 a_46223_19373# a_45805_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1048 VSS a_34414_13079# a_34937_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1049 a_54677_6923# C[59] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1050 a_46744_19298# a_46804_18801# a_45805_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1051 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1052 a_4208_14117# a_3760_12574# a_3361_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1053 a_10168_861# a_11157_670# a_11113_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1054 a_43875_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1055 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1056 VDD a_19539_6668# a_20062_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1057 a_14368_507# a_13944_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1058 a_13001_518# a_13045_670# a_12056_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1059 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1060 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1061 a_31560_6923# a_31390_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1062 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1063 a_6096_14117# a_5372_12574# a_5249_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1064 a_7984_14117# a_7260_12574# a_7137_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1065 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1066 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_48972_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1067 a_31904_5835# a_32027_6923# a_32751_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1068 a_58072_19299# a_58132_18802# a_57127_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1069 a_45120_6628# a_45519_6922# a_45971_6667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1070 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1071 VDD a_21198_13079# a_21721_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1072 a_37568_6629# a_36531_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1073 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1074 a_35680_5835# a_34639_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1075 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1555_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1076 a_20746_12574# a_20470_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1077 a_54525_518# a_55468_861# a_55426_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1078 a_27555_13117# a_27385_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1079 VSS C[87] a_14933_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1080 a_4233_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1081 a_23149_18584# a_24154_18802# a_24094_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1082 a_54525_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1083 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1084 a_30867_6667# a_30415_6922# a_30016_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1085 a_30701_18584# a_31706_18801# a_31646_19298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1086 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1087 a_33219_13117# a_33049_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1088 VDD a_32526_13079# a_33049_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1089 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1090 a_61762_6923# a_61592_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1091 VSS a_49575_18040# a_48636_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1092 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_7448_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1093 a_50228_507# a_49804_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1094 a_13902_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1095 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1096 VDD a_40078_13079# a_40601_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1097 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_54554_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1098 a_1677_1557# a_1733_1080# a_1242_317# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1099 a_23573_18776# a_23149_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1100 a_50749_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1101 a_13944_1405# a_14949_1079# a_14893_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1102 a_42029_18584# a_43034_18802# a_42974_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1103 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1104 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1105 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1106 VSS a_13877_5630# a_14404_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1107 a_43917_18584# a_44922_18802# a_44862_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1108 VDD a_53775_18776# a_53725_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1109 VDD a_28979_6668# a_29502_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1110 a_46435_12574# a_46265_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1111 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_3672_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1112 a_43207_1556# a_43247_670# a_42258_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1113 a_57986_6924# a_57816_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1114 a_47849_5630# a_47401_6923# a_47002_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1115 VSS a_10592_507# a_10542_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1116 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1117 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1118 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1119 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1120 VSS a_32755_6668# a_33278_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1121 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_52666_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1122 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_50778_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1123 VDD a_12816_19167# a_12832_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1124 a_13153_6923# C[37] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1125 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1126 a_14812_12575# C[102] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1127 VSS a_12251_19374# a_12201_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1128 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1129 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1130 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_44891_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1131 VSS a_13944_861# a_13001_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1132 a_42453_18776# a_42029_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1133 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18459_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1134 a_35655_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1135 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1136 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1137 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1138 a_5372_12574# C[97] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1139 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1140 VSS a_12480_1105# a_12430_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1141 a_15603_18584# a_16586_19166# a_16542_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1142 a_58072_19299# a_59015_18584# a_58973_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1143 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1144 a_16771_519# a_16815_671# a_15832_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1145 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1146 a_16970_12574# a_16694_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1147 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1148 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1149 a_4699_19374# a_4275_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1150 a_40794_507# a_40370_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1151 a_7341_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1152 VSS a_9939_18584# a_8996_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1153 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1154 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1155 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1156 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_11142_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1157 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_37339_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1158 a_48890_6629# a_49289_6923# a_49741_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 a_1242_317# a_1717_671# a_1673_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1160 a_14893_1556# a_15832_1405# a_15790_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1161 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1162 VDD C[17] a_27914_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1163 VSS C[25] a_12816_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1164 a_28813_18584# a_29802_19167# a_29758_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1165 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1166 a_9872_14117# a_9424_12574# a_9025_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1167 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1168 VDD a_19306_14117# a_19833_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1169 a_52666_6629# a_52789_6923# a_53517_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1170 VSS C[86] a_16815_671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1171 a_34477_18584# a_35466_19167# a_35422_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1172 VSS a_23315_6668# a_23838_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1173 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1174 a_35850_12574# a_35574_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1175 a_37314_18261# a_37354_19167# a_36365_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1176 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1177 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1178 a_18582_12574# C[104] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1179 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1180 a_41514_12574# a_41238_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 VDD a_24974_13079# a_25497_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1182 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1183 a_41000_6380# a_40830_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1184 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1185 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_56524_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1186 a_45120_6628# a_44083_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1187 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1188 a_55176_13079# a_54724_12574# a_54325_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1189 VSS a_17647_5630# a_18174_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1190 a_17714_1406# a_18719_1079# a_18663_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1191 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1192 a_28813_18584# a_29818_18802# a_29758_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1193 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1194 VDD a_38186_14117# a_38713_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1195 a_8704_1105# a_8280_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1196 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1197 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1198 a_22210_18261# a_23149_18040# a_23107_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1199 a_13112_6629# a_11993_6668# a_13030_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1200 a_56442_5835# a_56565_6923# a_57289_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1201 a_50860_5835# a_49737_5630# a_50778_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1202 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1203 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1204 a_16462_6379# a_16292_6379# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1205 a_50778_6629# a_51177_6923# a_51629_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1206 a_14345_12573# a_14175_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1207 a_37462_12574# C[114] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1208 VSS a_50793_670# a_50809_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1209 VSS a_27349_18776# a_27299_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1210 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1211 VDD a_43854_13079# a_44377_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1212 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1213 a_27349_18776# a_26925_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1214 a_43126_12574# C[117] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1215 a_11541_6923# a_11265_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1216 a_25266_861# a_26255_670# a_26211_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1217 VSS a_10168_1405# a_9229_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1218 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1219 a_20347_13912# a_20470_12574# a_21194_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1220 a_6793_12573# a_6623_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1221 a_29466_507# a_29042_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1222 VDD a_8704_1105# a_8654_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1223 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 a_12056_1405# a_13045_670# a_13005_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1225 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1226 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1227 a_41090_18261# a_42029_18040# a_41987_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1228 a_56188_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1229 a_58076_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1230 VDD a_22250_19167# a_22266_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1231 a_42978_18261# a_43917_18040# a_43875_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1232 a_22235_13912# a_22634_12574# a_23082_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1233 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1234 a_38211_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1235 a_61533_12574# a_61363_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1236 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1237 a_23149_18040# a_24138_19167# a_24098_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1238 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_60218_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1239 a_25982_19299# a_26026_19167# a_25037_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1240 a_35130_1105# a_34706_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1241 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1242 VSS a_40307_6668# a_40830_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1243 a_28527_6923# a_28251_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1244 a_30701_18040# a_31690_19166# a_31650_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1245 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1246 a_11142_6629# a_11265_6923# a_11993_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1247 VDD a_52116_507# a_52066_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1248 VSS a_58116_19167# a_58132_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1249 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_59989_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1250 a_59645_13117# a_59475_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1251 a_15790_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1252 a_5449_518# a_6392_861# a_6350_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1253 a_18663_1556# a_19602_1405# a_19560_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1254 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1255 a_39227_13912# a_39350_12574# a_40074_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1256 a_16771_519# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1257 a_34664_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1258 a_9148_12574# C[99] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1259 a_49512_13079# a_48784_12574# a_48661_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1260 a_35655_1556# a_35695_670# a_34706_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1261 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1262 a_21685_18776# a_21261_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1263 a_10798_6924# a_10628_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1264 VSS a_8475_19374# a_8425_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1265 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1266 a_58500_12574# a_58224_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1267 VDD a_4928_507# a_4878_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1268 VDD a_41130_19167# a_41146_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1269 a_17485_18039# a_18490_18802# a_18434_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1270 a_41115_13912# a_41514_12574# a_41962_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1271 a_43003_13912# a_43402_12574# a_43850_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1272 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1273 a_60617_6922# a_60341_6922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1274 a_34706_1405# a_35711_1079# a_35655_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1276 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1277 a_48661_13118# a_48784_12574# a_49512_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1278 VSS a_34639_5630# a_35166_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1279 VSS a_38482_861# a_37539_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1280 a_42029_18040# a_43018_19167# a_42978_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1281 a_26011_13118# a_24974_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1282 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1283 a_44862_19299# a_44906_19167# a_43917_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1284 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1285 a_27899_13118# a_26862_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1286 a_38906_507# a_38482_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1287 VDD a_10363_19374# a_10313_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1288 VSS C[21] a_20362_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1289 a_23149_18040# a_24154_18802# a_24098_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1290 a_32522_14117# a_32074_12574# a_31675_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1291 VDD a_23802_1105# a_23752_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1292 a_33013_18776# a_32589_18039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1293 VDD C[80] a_28143_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1294 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1295 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_52437_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1296 a_30701_18040# a_31706_18801# a_31650_18260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1297 a_9254_6629# a_9653_6923# a_10105_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1298 a_48890_6629# a_47853_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1299 a_40565_18776# a_40141_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1300 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1301 a_58305_1556# a_58345_670# a_57356_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1302 a_59668_1105# a_59244_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1303 VSS a_25690_507# a_25640_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1304 VSS a_34706_861# a_33763_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1305 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1306 a_18541_13912# a_17418_14117# a_18459_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1307 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1308 VSS C[27] a_9040_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1309 a_49575_18584# a_50564_19167# a_50520_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1310 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1311 a_45738_14118# a_45290_12575# a_44891_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1312 VDD a_8217_6668# a_8740_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1313 a_52412_18261# a_52452_19167# a_51463_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1314 VSS a_28116_9428# sky130_fd_sc_hd__buf_2_0/X VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1315 a_20551_1556# a_21490_1405# a_21448_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1316 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1317 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1318 a_27091_6668# a_26639_6923# a_26240_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1319 VSS a_33242_1105# a_33192_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1320 a_20547_518# a_21490_861# a_21448_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1321 VSS C[11] a_39242_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1322 a_42029_18040# a_43034_18802# a_42978_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1323 a_9254_5835# a_9653_6923# a_10101_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1324 a_43917_18040# a_44922_18802# a_44866_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 a_24205_13912# a_23082_14117# a_24123_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1326 a_24323_518# a_24367_670# a_23378_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1327 a_18430_19299# a_18490_18802# a_17485_18039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1328 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1329 a_15561_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1330 a_34706_861# a_35711_1079# a_35651_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1331 a_6350_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1332 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1333 VSS a_19797_18776# a_19747_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1334 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1335 a_37691_6923# C[50] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1336 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_11224_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1337 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1338 VDD a_53284_14117# a_53811_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1339 a_13877_5630# a_13429_6923# a_13030_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1340 a_15832_1405# a_16815_671# a_16775_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1341 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1342 VSS a_25199_5630# a_25726_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1343 a_55892_507# a_55468_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1344 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1345 a_16250_508# a_15832_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1346 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1347 a_6121_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1348 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1349 a_49575_18584# a_50580_18802# a_50520_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1350 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1351 a_52560_12574# C[122] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1352 a_22120_6924# a_21950_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1353 VDD a_11989_5630# a_12516_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1354 a_60218_6628# a_60341_6922# a_61069_6667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1355 a_43085_13912# a_41962_14117# a_43003_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1356 a_25203_6668# a_24475_6923# a_24352_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1357 a_15603_18040# a_16586_19166# a_16546_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1358 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1359 a_37310_19299# a_37370_18802# a_36365_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1360 a_10913_13118# a_11312_12574# a_11764_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1361 a_24475_6923# C[43] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1362 a_10592_1105# a_10168_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1363 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1364 a_26215_1556# a_26271_1079# a_25266_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1365 VSS a_38677_18776# a_38627_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1366 a_57356_861# a_58361_1079# a_58301_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1367 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1368 VDD C[94] a_1717_671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1369 a_17672_888# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1370 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1371 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 VDD a_26026_19167# a_26042_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1373 a_1473_13118# a_1872_12574# a_2324_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1374 a_50749_518# a_50809_1079# a_49804_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1375 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1376 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1377 a_25199_5630# a_24475_6923# a_24352_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1378 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1379 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1380 a_28813_18040# a_29802_19167# a_29762_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1381 a_17714_862# a_18703_670# a_18659_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1382 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1383 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1384 VSS a_3376_19167# a_3392_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1385 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1386 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1387 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_20429_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1388 a_12457_12573# a_12287_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1389 VDD a_25461_18776# a_25411_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1390 a_34477_18040# a_35466_19167# a_35426_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1391 VSS a_32589_18583# a_31646_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1392 a_44083_6668# a_43631_6923# a_43232_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1393 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1394 a_37310_19299# a_37354_19167# a_36365_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1395 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1396 a_3760_12574# a_3484_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1397 a_24323_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1398 VDD a_31125_18775# a_31075_18610# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1399 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1400 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1401 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1402 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1403 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_10913_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1404 a_4905_12573# a_4735_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1405 VDD C[74] a_39471_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1406 a_56188_18261# a_56244_18802# a_55239_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1407 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_12801_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1408 VSS a_38906_1105# a_38856_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1409 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1410 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1411 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1412 a_31560_6923# a_31390_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1413 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1414 a_18430_19299# a_19373_18584# a_19331_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1415 VDD a_14933_670# a_14949_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1416 VSS C[73] a_41359_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1417 a_59202_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1418 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1419 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1420 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1421 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_3361_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1422 VDD a_57293_6668# a_57816_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1423 VDD a_44341_18776# a_44291_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1424 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1425 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_60300_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1426 VSS a_31690_19166# a_31706_18801# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1427 VDD a_46788_19166# a_46804_18801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1428 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_56213_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1429 a_20547_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1430 a_14771_13119# a_13652_13079# a_14689_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1431 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1432 VDD a_6587_19374# a_6537_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1433 a_42195_6668# a_41467_6923# a_41344_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1434 a_49289_6923# a_49013_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1435 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1436 a_14368_507# a_13944_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1437 a_46223_19373# a_45805_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1438 a_27784_6924# a_27614_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1439 a_41467_6923# C[52] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1440 a_17647_5630# a_17199_6923# a_16800_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1441 a_32547_18859# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1442 a_53351_18584# a_54340_19167# a_54296_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1443 a_5331_13118# a_4212_13079# a_5249_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1444 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_22464_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1445 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1446 a_37310_19299# a_38253_18584# a_38211_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1447 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1448 a_60836_14118# a_60388_12575# a_59989_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1449 VDD a_61065_5629# a_61592_6379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1450 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_20576_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1451 a_56188_18261# a_56228_19167# a_55239_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1452 VDD a_37583_670# a_37599_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1453 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1454 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1455 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1456 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1457 VSS a_21198_13079# a_21721_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1458 VSS a_40794_1105# a_40744_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1459 VSS a_59244_861# a_58301_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1460 VDD a_3040_507# a_2990_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1461 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1462 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1463 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1464 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1465 a_22863_6923# a_22587_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1466 a_52641_1556# a_52697_1079# a_51692_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1467 VDD a_57060_14117# a_57587_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1468 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1469 VSS a_32526_13079# a_33049_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1470 a_20658_6629# a_19539_6668# a_20576_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1471 a_23378_1405# a_24367_670# a_24327_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1472 VSS a_2616_1406# a_1677_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1473 a_39538_6629# a_38419_6668# a_39456_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1474 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1475 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1476 a_13200_12574# a_12924_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1477 a_41315_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1478 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1479 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1480 a_56336_12574# C[124] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1481 VSS a_40078_13079# a_40601_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1482 a_3989_6923# a_3713_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1483 a_18688_6629# a_19087_6923# a_19539_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1484 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1485 a_45120_5834# a_45243_6922# a_45967_5629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1486 a_52408_19299# a_52468_18802# a_51463_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1487 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_48743_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1488 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1489 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_41344_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1490 VSS a_54004_1105# a_53954_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1491 a_31354_1106# a_30930_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1492 VSS a_53775_18776# a_53725_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1493 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1494 VSS a_15536_14118# a_16063_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1495 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1496 a_22464_6629# a_22587_6923# a_23315_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1497 a_32027_6923# C[47] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1498 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1499 a_21891_13117# a_21721_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1500 a_16546_18260# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1501 VSS a_2320_14117# a_2847_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1502 a_5249_13118# a_5648_12574# a_6100_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1503 a_46435_12574# a_46265_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1504 a_57085_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1505 a_58973_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1506 a_58453_6923# C[61] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1507 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_31986_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1508 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1509 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1510 a_15088_12575# a_14812_12575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1511 a_44776_6924# a_44606_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1512 a_34639_5630# a_34191_6923# a_33792_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1513 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1514 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1515 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_24205_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1516 a_18663_1556# a_18719_1079# a_17714_862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1517 VDD a_41359_670# a_41375_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1519 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_26322_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1520 VDD a_29237_18776# a_29187_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1521 a_54004_507# a_53580_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1522 VSS a_16586_19166# a_16602_18801# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1523 a_49575_18040# a_50564_19167# a_50524_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1524 VDD a_7988_13079# a_8511_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1525 a_45742_13080# a_45290_12575# a_44891_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1526 a_41426_6629# a_40307_6668# a_41344_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1528 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1529 a_14664_18261# a_15603_18040# a_15561_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1530 a_52408_19299# a_52452_19167# a_51463_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1531 a_18115_13117# a_17945_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1532 a_20003_13117# a_19833_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1533 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_31757_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1534 a_7536_12574# a_7260_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1535 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1536 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1537 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1538 a_51692_861# a_52681_670# a_52637_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1539 a_40771_13117# a_40601_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1540 a_35426_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1541 a_20576_6629# a_20975_6923# a_21427_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1542 a_40794_507# a_40370_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1543 a_5224_18261# a_6163_18040# a_6121_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1544 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1545 a_46773_13118# a_45742_13080# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1546 a_14689_13913# a_13648_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1547 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_43085_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1548 a_25690_1105# a_25266_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1549 a_12801_13912# a_12924_12574# a_13648_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1550 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1473_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1551 a_32751_5630# a_32027_6923# a_31904_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1552 a_52437_13118# a_51400_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1553 a_20576_5835# a_20975_6923# a_21423_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1554 a_60193_1556# a_60233_670# a_59244_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1555 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1556 a_38883_13117# a_38713_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1557 a_45091_518# a_46034_861# a_45992_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1558 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1559 a_5249_13912# a_4208_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1560 a_3713_6923# C[32] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1561 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1562 a_3361_13912# a_3484_12574# a_4208_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1563 a_49013_6923# C[56] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1564 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_22546_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1565 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1566 a_21219_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1567 a_58224_12574# C[125] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1568 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1569 VSS a_11827_18584# a_10884_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1570 a_52408_19299# a_53351_18584# a_53309_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1571 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1572 a_5249_13912# a_5648_12574# a_6096_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1573 a_39456_6629# a_39579_6923# a_40307_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1574 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_30016_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1575 VSS a_10105_6668# a_10628_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1576 a_37018_1105# a_36594_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1577 a_6325_5630# a_5877_6923# a_5478_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1578 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1579 VSS a_24974_13079# a_25497_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1580 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1581 a_11760_14117# a_11312_12574# a_10913_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1582 a_14918_6628# a_15041_6922# a_15769_6667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1583 a_7448_5835# a_6325_5630# a_7366_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1584 a_4504_861# a_5493_670# a_5449_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1585 a_12251_18776# a_11827_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1586 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1587 VDD C[85] a_18703_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1588 a_13005_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1589 a_34435_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1590 a_13648_14117# a_12924_12574# a_12801_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1591 VDD a_4437_5630# a_4964_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1592 VDD C[66] a_54569_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1593 a_29987_518# a_30047_1079# a_29042_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1594 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1595 a_56098_6924# a_55928_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1596 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1597 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1598 a_19310_13079# a_18858_12574# a_18459_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1599 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_43314_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1600 a_30415_6922# a_30139_6922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1601 a_40099_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1602 a_41987_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1603 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1604 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1605 VSS C[65] a_56457_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1606 a_4208_14117# a_3484_12574# a_3361_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1607 a_46973_519# a_47033_1080# a_46034_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1608 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 a_31650_18260# a_31690_19166# a_30701_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1610 a_43232_5835# a_43355_6923# a_44079_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1611 a_56413_518# a_56457_670# a_55468_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1612 a_56841_6923# a_56565_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1613 a_30016_5834# a_30415_6922# a_30863_5629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1614 VSS a_43854_13079# a_44377_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1615 a_47401_6923# a_47125_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1616 a_48546_6924# a_48376_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1617 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1618 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1619 a_57551_19374# a_57127_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1620 a_6163_18040# a_7168_18802# a_7112_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1621 a_56184_19299# a_56244_18802# a_55239_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1622 a_9424_12574# a_9148_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1623 a_59244_861# a_60249_1079# a_60189_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1624 a_18688_6629# a_17651_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1625 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1626 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_14771_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1627 a_16800_5835# a_15765_5629# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1628 a_29466_507# a_29042_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1629 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1630 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1631 a_38190_13079# a_37738_12574# a_37339_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1632 a_21261_18584# a_22266_18802# a_22206_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1633 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1634 a_25667_13117# a_25497_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1635 VSS a_30634_14118# a_31161_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1636 a_61533_12574# a_61363_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1637 a_52637_518# a_52681_670# a_51692_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1638 a_48865_1556# a_48905_670# a_47916_862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1639 a_27578_1105# a_27154_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1640 a_7022_6924# a_6852_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1641 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1642 a_30186_12575# a_29910_12575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1643 VSS a_52116_507# a_52066_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1644 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1645 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1646 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1647 a_34477_18584# a_35482_18802# a_35422_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1648 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1649 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1650 a_60840_13080# a_60388_12575# a_59989_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1651 a_39427_518# a_39487_1079# a_38482_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1652 a_29762_18261# a_30701_18040# a_30659_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1653 a_21685_18776# a_21261_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1654 VSS a_4928_507# a_4878_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1655 a_1673_519# a_1733_1080# a_1242_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1656 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1657 a_40141_18584# a_41146_18802# a_41086_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1658 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1659 a_44547_13117# a_44377_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1660 VDD a_51887_18776# a_51837_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1661 VSS a_59015_18040# a_58076_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1662 a_59177_5630# a_58729_6923# a_58330_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1663 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1664 a_53517_6668# a_52789_6923# a_52666_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1665 a_16546_18260# a_16602_18801# a_15603_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1666 VSS a_16815_671# a_16831_1080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1667 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1668 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1669 a_52789_6923# C[58] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1670 a_33013_18776# a_32589_18039# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1671 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1672 a_11036_12574# C[100] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1673 VDD a_36531_6668# a_37054_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1674 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1675 VSS a_10363_19374# a_10313_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1676 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1677 a_52093_13117# a_51923_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1678 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1679 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1680 a_40565_18776# a_40141_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1681 a_53981_13117# a_53811_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1682 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1683 a_7137_13912# a_7260_12574# a_7984_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1684 a_9229_1556# a_9269_670# a_8280_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1685 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1686 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1687 a_9025_13912# a_9148_12574# a_9872_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1688 a_3484_12574# C[96] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1689 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_47084_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1690 a_35680_6629# a_34643_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1691 VDD a_39471_670# a_39487_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1692 a_33792_5835# a_32751_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1693 VDD C[79] a_30031_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1694 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1695 VDD a_9040_19167# a_9056_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1696 a_35426_18261# a_35482_18802# a_34477_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1697 a_56184_19299# a_57127_18584# a_57085_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1698 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1699 a_16546_18260# a_16586_19166# a_15603_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1700 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_27899_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1701 VDD a_42682_507# a_42632_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1702 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1703 VDD C[22] a_18474_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1704 a_52641_1556# a_52681_670# a_51692_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1705 a_52637_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1706 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1707 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1708 a_5453_1556# a_5509_1079# a_4504_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1709 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1710 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35451_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1711 a_25037_18584# a_26026_19167# a_25982_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1712 VDD C[18] a_26026_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1713 VSS C[26] a_10928_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1714 a_26925_18584# a_27914_19167# a_27870_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1715 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_54554_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1716 VSS a_43247_670# a_43263_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1717 a_12014_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1718 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1719 a_27874_18261# a_27914_19167# a_26925_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1720 a_55892_507# a_55468_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1721 a_8475_18776# a_8051_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1722 a_29762_18261# a_29802_19167# a_28813_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1723 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1724 VDD C[15] a_31690_19166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1725 VDD a_17418_14117# a_17945_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1726 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1727 VSS C[31] a_1488_19166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1728 a_32589_18583# a_33578_19167# a_33534_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1729 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1730 a_32074_12574# a_31798_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1731 a_33962_12574# a_33686_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1732 a_35426_18261# a_35466_19167# a_34477_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1733 VSS a_11989_5630# a_12516_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1734 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1735 VDD C[12] a_37354_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1736 VDD a_27091_6668# a_27614_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1737 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1738 a_16694_12574# C[103] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1739 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_30098_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1740 a_2811_19374# a_2387_18583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1741 VSS C[28] a_7152_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1742 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1743 a_40328_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1744 a_24327_1556# a_24367_670# a_23378_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1745 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1746 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1747 a_47624_13079# a_47172_12574# a_46773_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1748 VDD a_28746_14117# a_29273_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1749 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_50778_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1750 VDD C[8] a_44906_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1751 a_19087_6923# a_18811_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1752 a_30930_861# a_31919_671# a_31875_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1753 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1754 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1755 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1756 a_45971_6667# a_45243_6922# a_45120_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1757 a_45290_12575# a_45014_12575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1758 a_11265_6923# C[36] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1759 a_26925_18584# a_27930_18802# a_27870_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1760 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1761 a_53288_13079# a_52836_12574# a_52437_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1762 VDD a_36298_14117# a_36825_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1763 VDD a_30863_5629# a_31390_6379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1764 a_29910_12575# C[110] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1765 a_5478_5835# a_4437_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1766 a_33767_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1767 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1768 a_20551_1556# a_20607_1079# a_19602_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1769 a_51692_861# a_52697_1079# a_52637_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1770 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1771 a_12457_12573# a_12287_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1772 a_35574_12574# C[113] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1773 VSS a_29042_861# a_28099_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1774 VSS a_10592_1105# a_10542_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1775 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1776 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1777 VSS a_25461_18776# a_25411_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1778 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1779 VSS a_31125_18775# a_31075_18610# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1780 VSS sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1781 VDD C[92] a_5493_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1782 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1783 a_4905_12573# a_4735_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1784 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1785 VSS a_53580_1405# a_52641_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1786 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1787 a_54300_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1788 a_47002_6629# a_47401_6923# a_47853_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1789 VDD a_20362_19167# a_20378_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1790 a_13005_1556# a_13944_1405# a_13902_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1791 a_36323_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1792 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1793 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1794 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_39309_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1795 VSS a_48676_19167# a_48692_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1796 a_21261_18040# a_22250_19167# a_22210_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1797 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1798 VDD a_37018_1105# a_36968_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1799 VSS a_44341_18776# a_44291_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1800 a_24094_19299# a_24138_19167# a_23149_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1801 a_31675_13912# a_31798_12574# a_32522_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1802 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1803 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1804 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1805 a_49060_12574# a_48784_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1806 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1807 a_57757_13117# a_57587_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1808 VDD a_44083_6668# a_44606_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1809 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1810 a_31646_19298# a_31690_19166# a_30701_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1811 a_13001_518# a_13944_861# a_13902_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1812 a_47624_13079# a_46896_12574# a_46773_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1813 VDD a_38906_1105# a_38856_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1814 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1815 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1816 a_21914_507# a_21490_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1817 a_51692_1405# a_52681_670# a_52641_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1818 VSS a_6587_19374# a_6537_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1819 a_18459_13118# a_17422_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1820 a_56612_12574# a_56336_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1821 a_28251_6923# C[45] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1822 a_39202_18261# a_39258_18802# a_38253_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1823 a_36079_6923# a_35803_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1824 a_18858_12574# a_18582_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1825 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_54636_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1826 a_19602_861# a_20591_670# a_20547_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1827 a_44891_13913# a_45014_12575# a_45738_14118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1828 a_14574_6924# a_14404_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1829 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1830 a_40141_18040# a_41130_19167# a_41090_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1831 a_24123_13118# a_23086_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1832 a_21261_18040# a_22266_18802# a_22210_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1833 a_42974_19299# a_43018_19167# a_42029_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1834 a_54554_5835# a_54677_6923# a_55401_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1835 VSS a_3040_507# a_2990_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1836 a_11224_6629# a_10105_6668# a_11142_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1837 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1838 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_7219_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1839 a_60341_6922# C[62] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1840 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1841 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1842 a_50778_6629# a_50901_6923# a_51629_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1843 a_58330_5835# a_57289_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1844 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1845 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_50549_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1846 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1847 VSS a_46034_861# a_45091_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1848 a_58101_13118# a_58224_12574# a_58952_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1849 a_35651_518# a_36594_861# a_36552_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1850 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1851 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1852 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1853 VDD a_1717_671# a_1733_1080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1854 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1855 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1856 a_34477_18040# a_35482_18802# a_35426_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1857 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1858 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1859 a_16653_13912# a_15536_14118# a_16571_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1860 a_37738_12574# a_37462_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1861 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1862 a_58183_13118# a_57064_13079# a_58101_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1863 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_61877_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1864 a_50778_5835# a_50901_6923# a_51625_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1865 a_10168_1405# a_11157_670# a_11117_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1866 VDD C[4] a_52452_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1867 a_50524_18261# a_50564_19167# a_49575_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1868 a_43003_13118# a_41966_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1869 a_40141_18040# a_41146_18802# a_41090_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1870 a_22317_13912# a_21194_14117# a_22235_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1871 a_45738_14118# a_45014_12575# a_44891_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1872 a_54554_5835# a_53513_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1873 a_16021_19373# a_15603_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1874 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1875 a_16542_19298# a_16602_18801# a_15603_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1876 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1877 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1878 a_59015_18584# a_60004_19167# a_59960_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1879 VDD C[0] a_60004_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1880 a_13673_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1881 VDD a_54569_670# a_54585_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1882 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1883 a_58952_13079# a_58500_12574# a_58101_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1884 a_18811_6923# C[40] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1885 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1886 a_52116_1105# a_51692_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1887 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1888 VDD a_49508_14117# a_50035_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1889 a_9254_6629# a_9377_6923# a_10105_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1890 a_35533_13912# a_34410_14117# a_35451_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1891 a_47620_14117# a_46896_12574# a_46773_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1892 VDD a_51396_14117# a_51923_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1893 VDD a_57780_507# a_57730_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1894 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1895 a_27870_19299# a_27930_18802# a_26925_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1896 a_29758_19299# a_29818_18802# a_28813_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1897 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1898 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1899 a_50672_12574# C[121] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1900 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1901 VSS a_29237_18776# a_29187_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1902 a_41197_13912# a_40074_14117# a_41115_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 a_54004_507# a_53580_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1904 VSS a_7988_13079# a_8511_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1905 VSS a_58345_670# a_58361_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1906 VSS a_36594_861# a_35651_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1907 a_32818_1406# a_33823_1079# a_33767_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1908 a_35422_19299# a_35482_18802# a_34477_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1909 VDD a_60903_18040# a_63251_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1910 VDD a_55401_5630# a_55928_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1911 VDD a_12480_1105# a_12430_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1912 a_58305_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1913 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_13112_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1914 VDD a_47853_6668# a_48376_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1915 VSS a_47620_14117# a_48147_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1916 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_50860_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1917 a_59015_18584# a_60020_18802# a_59960_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1918 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1919 VSS a_51629_6668# a_52152_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1920 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1921 VSS a_19373_18040# a_18434_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1922 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1923 a_51421_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1924 a_25037_18040# a_26026_19167# a_25986_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1925 a_18344_6924# a_18174_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1926 a_60300_6628# a_59181_6668# a_60218_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1927 a_55426_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1928 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1929 VDD a_17909_18776# a_17859_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1930 a_26925_18040# a_27914_19167# a_27874_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1931 VDD a_9876_13079# a_10399_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1932 a_27870_19299# a_27914_19167# a_26925_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1933 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1934 a_29758_19299# a_29802_19167# a_28813_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1935 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1936 a_10569_12573# a_10399_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1937 VSS a_45967_5629# a_46494_6379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1938 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1939 a_1444_19298# a_2387_18583# a_2345_18859# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1940 VDD a_23573_18776# a_23523_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1941 a_46748_18260# a_47687_18039# a_47645_18065# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1942 a_25203_6668# a_24751_6923# a_24352_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1943 a_37543_1556# a_38482_1405# a_38440_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1944 VSS a_32589_18039# a_31650_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1945 a_16233_12574# a_16063_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1946 a_22435_518# a_22479_670# a_21490_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1947 a_1872_12574# a_1596_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1948 VDD C[78] a_31919_671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1949 a_43207_1556# a_43263_1079# a_42258_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1950 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1951 a_8681_13117# a_8511_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1952 a_3017_12573# a_2847_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1953 VSS a_38253_18040# a_37314_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1954 a_54300_18261# a_54356_18802# a_53351_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1955 a_4462_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1956 a_35803_6923# C[49] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1957 VSS C[20] a_22250_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1958 a_12251_18776# a_11827_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1959 a_11989_5630# a_11541_6923# a_11142_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1960 a_33767_1556# a_34706_1405# a_34664_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1961 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1962 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1963 a_31875_519# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1964 a_4504_1405# a_5509_1079# a_5453_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1965 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1966 VSS a_4437_5630# a_4964_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1967 VSS a_8280_861# a_7337_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1968 VDD a_42453_18776# a_42403_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1969 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1970 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1971 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1972 a_39112_6924# a_38942_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1973 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1974 a_48636_18261# a_48676_19167# a_47687_18583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1975 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1976 a_23315_6668# a_22587_6923# a_22464_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1977 a_58101_13912# a_57060_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1978 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_31904_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1979 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1980 a_49575_18040# a_50580_18802# a_50524_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1981 a_3443_13118# a_2324_13079# a_3361_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1982 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1983 a_22587_6923# C[42] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1984 VSS C[91] a_7381_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1985 a_35422_19299# a_36365_18584# a_36323_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1986 a_52836_12574# a_52560_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1987 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1988 a_11113_518# a_12056_861# a_12014_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1989 VSS a_4504_861# a_3561_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1990 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1991 VSS a_49575_18584# a_48632_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1992 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1993 a_60836_14118# a_60112_12575# a_59989_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1994 a_43203_518# a_43247_670# a_42258_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1995 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1996 a_43631_6923# a_43355_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1997 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1998 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1999 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2000 a_34191_6923# a_33915_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2001 a_35336_6924# a_35166_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2002 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2003 VSS a_3040_1105# a_2990_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2004 a_57551_19374# a_57127_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2005 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2006 a_49508_14117# a_49060_12574# a_48661_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2007 a_42258_861# a_43247_670# a_43203_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2008 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2009 a_13030_6629# a_13429_6923# a_13881_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2010 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2011 a_50631_13912# a_49508_14117# a_50549_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2012 a_9897_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2013 a_11312_12574# a_11036_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2014 a_22435_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2015 a_45742_13080# a_45014_12575# a_44891_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2016 a_54448_12574# C[123] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2017 VDD C[84] a_20591_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2018 a_14368_1105# a_13944_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2019 VDD C[71] a_45135_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2020 a_12801_13118# a_13200_12574# a_13652_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2021 VDD a_33242_507# a_33192_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2022 a_50520_19299# a_50580_18802# a_49575_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2023 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2024 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_46855_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2025 a_44891_13119# a_45014_12575# a_45742_13080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2026 VSS C[83] a_22479_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2027 a_57314_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2028 a_49533_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2029 VSS a_51887_18776# a_51837_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2030 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2031 a_3361_13118# a_3760_12574# a_4212_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2032 a_57356_1405# a_58361_1079# a_58305_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2033 a_55197_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2034 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2035 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2036 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2037 VDD a_13652_13079# a_14175_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2038 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_58183_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2039 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2040 a_40307_6668# a_39579_6923# a_39456_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2041 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2042 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2043 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2044 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_22317_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2045 a_25896_6924# a_25726_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2046 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_20576_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2047 a_53538_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2048 a_28979_6668# a_28251_6923# a_28128_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2049 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_37568_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2050 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2051 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2052 VDD a_18703_670# a_18719_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2053 a_12776_18261# a_13715_18040# a_13673_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2054 VDD a_6100_13079# a_6623_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2055 a_50520_19299# a_50564_19167# a_49575_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2056 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_29869_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2057 a_5648_12574# a_5372_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2058 a_3040_1105# a_2616_1406# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2059 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2060 a_31331_12574# a_31161_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2061 a_54210_6380# a_54040_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2062 VSS a_57356_861# a_56413_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2063 a_53580_1405# a_54585_1079# a_54529_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2064 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2065 a_8051_18584# a_9056_18802# a_8996_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2066 a_31646_19298# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2067 VSS a_53351_18040# a_52412_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2068 a_33538_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2069 VSS a_56457_670# a_56473_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2070 VSS a_42682_507# a_42632_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2071 a_3336_18261# a_4275_18040# a_4233_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 a_20975_6923# a_20699_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2073 VDD a_7381_670# a_7397_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2074 VDD a_49999_18776# a_49949_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2075 a_59015_18040# a_60004_19167# a_59964_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2076 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2077 a_39855_6923# a_39579_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2078 a_3565_1556# a_3605_670# a_2616_862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2079 VSS a_27914_19167# a_27930_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2080 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_41197_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2081 a_29443_13117# a_29273_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2082 VDD a_27578_1105# a_27528_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2083 VSS a_8704_1105# a_8654_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2084 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2085 a_10913_13912# a_11036_12574# a_11760_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2086 a_19310_13079# a_18582_12574# a_18459_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2087 a_39427_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2088 VSS a_9269_670# a_9285_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2089 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2090 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2091 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2092 VDD a_10928_19167# a_10944_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2093 a_35107_13117# a_34937_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2094 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2095 a_50434_6380# a_50264_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2096 a_3361_13912# a_2320_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2097 a_12801_13912# a_13200_12574# a_13648_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2098 a_36995_13117# a_36825_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2099 a_8475_18776# a_8051_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2100 a_16800_6629# a_17199_6923# a_17651_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2101 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2102 a_18459_13118# a_18582_12574# a_19310_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2103 a_28099_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2104 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2105 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_41344_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2106 a_58305_1556# a_59244_1405# a_59202_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2107 VSS a_52116_1105# a_52066_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2108 a_1673_519# a_2616_862# a_2574_888# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2109 a_32755_6668# a_32303_6923# a_31904_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2110 a_50520_19299# a_51463_18584# a_51421_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2111 a_3361_13912# a_3760_12574# a_4208_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2112 a_18138_1105# a_17714_1406# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2113 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_22235_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2114 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2115 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2116 a_38190_13079# a_37462_12574# a_37339_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2117 VDD a_13881_6668# a_14404_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2118 a_2811_19374# a_2387_18583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2119 a_10363_18776# a_9939_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2120 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2121 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2122 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2123 a_47125_6923# C[55] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2124 a_56565_6923# C[60] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2125 VDD C[70] a_47017_671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2126 a_42888_6924# a_42718_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2127 a_32751_5630# a_32303_6923# a_31904_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2128 a_21490_1405# a_22479_670# a_22439_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2129 a_19373_18584# a_20362_19167# a_20318_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2130 a_923_18775# a_1013_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2131 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2132 a_15536_14118# a_15088_12575# a_14689_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2133 a_37339_13118# a_37462_12574# a_38190_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2134 a_22210_18261# a_22250_19167# a_21261_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2135 a_56184_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2136 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_24434_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2137 a_58072_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2138 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2139 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2140 a_13715_18040# a_14720_18802# a_14664_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2141 a_48111_19374# a_47687_18583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2142 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2143 a_24352_5835# a_24475_6923# a_25199_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2144 a_2616_862# a_3621_1079# a_3561_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2145 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2146 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2147 a_37421_13118# a_36302_13079# a_37339_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2148 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_41115_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2149 a_60840_13080# a_60112_12575# a_59989_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2150 VSS a_60233_670# a_60249_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2151 a_61959_13912# a_60836_14118# a_61877_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2152 a_15000_6628# a_13881_6668# a_14918_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2153 a_37650_5835# a_36527_5630# a_37568_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2154 a_9336_6629# a_8217_6668# a_9254_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2155 a_37568_6629# a_37967_6923# a_38419_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2156 a_28128_5835# a_27087_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2157 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2158 a_59874_6380# a_59704_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2159 a_34706_861# a_35695_670# a_35651_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2160 a_55663_19374# a_55239_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2161 a_54296_19299# a_54356_18802# a_53351_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2162 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2163 VDD a_23082_14117# a_23609_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2164 a_59989_13119# a_60112_12575# a_60840_13080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2165 a_45967_5629# a_45519_6922# a_45120_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2166 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2167 a_41090_18261# a_41130_19167# a_40141_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2168 a_23779_13117# a_23609_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2169 a_36302_13079# a_35850_12574# a_35451_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2170 a_8238_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2171 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2172 a_19373_18584# a_20378_18802# a_20318_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2173 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2174 a_18434_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2175 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2176 a_20576_5835# a_20699_6923# a_21423_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2177 a_26211_518# a_27154_861# a_27112_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2178 a_1152_1106# a_1242_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2179 VSS a_40370_1405# a_39431_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2180 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2181 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2182 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2183 a_33792_6629# a_34191_6923# a_34643_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2184 a_24352_5835# a_23311_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2185 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2186 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2187 a_32589_18583# a_33594_18802# a_33534_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2188 a_57356_861# a_58345_670# a_58301_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2189 VDD a_41962_14117# a_42489_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2190 a_4437_5630# a_3989_6923# a_3590_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2191 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_45120_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2192 a_21914_507# a_21490_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2193 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2194 a_42659_13117# a_42489_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2195 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2196 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2197 a_37314_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2198 VSS a_57127_18040# a_56188_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2199 VDD a_1152_1106# a_1102_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2200 a_11117_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2201 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2202 a_9000_18261# a_9939_18040# a_9897_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2203 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_41426_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2204 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2205 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2206 a_41000_6924# a_40830_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2207 VDD a_48340_507# a_48290_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2208 VDD a_923_19373# a_873_19154# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2209 a_14893_1556# a_14933_670# a_13944_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2210 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2211 VDD a_17651_6668# a_18174_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2212 a_23336_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2213 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_20658_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2214 a_41344_5835# a_41467_6923# a_42191_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2215 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2216 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2217 a_54953_6923# a_54677_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2218 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2219 a_25986_18261# a_26042_18802# a_25037_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2220 a_50205_13117# a_50035_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2221 VSS a_21427_6668# a_21950_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2222 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2223 a_5249_13912# a_5372_12574# a_6096_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2224 VSS a_56228_19167# a_56244_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2225 a_1596_12574# C[95] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2226 a_39626_12574# a_39350_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2227 a_16800_6629# a_15769_6667# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2228 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2229 VDD a_7152_19167# a_7168_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2230 a_33538_18261# a_33594_18802# a_32589_18583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2231 a_54296_19299# a_55239_18584# a_55197_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2232 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2233 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2234 a_9025_13912# a_9424_12574# a_9872_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2235 VDD a_14139_18776# a_14089_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2236 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_26011_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2237 a_29987_518# a_30930_861# a_30888_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2238 a_8051_18040# a_9040_19167# a_9000_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2239 VSS a_15765_5629# a_16292_6379# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2240 a_61065_5629# a_60617_6922# a_60218_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2241 a_50749_518# a_50793_670# a_49804_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2242 a_14139_18776# a_13715_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2243 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2244 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2245 a_12480_507# a_12056_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2246 VDD a_46223_19373# a_46173_19154# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2247 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2248 a_16021_19373# a_15603_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2249 a_44866_18261# a_44922_18802# a_43917_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2250 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_33563_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2251 VDD a_5493_670# a_5509_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2252 a_23149_18584# a_24138_19167# a_24094_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2253 VDD C[19] a_24138_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2254 a_63421_12573# a_63251_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2255 a_25986_18261# a_26026_19167# a_25037_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2256 a_30634_14118# a_30186_12575# a_29787_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2257 a_52437_13118# a_52560_12574# a_53288_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2258 VSS a_57780_507# a_57730_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2259 a_6587_18776# a_6163_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2260 a_60189_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2261 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2262 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2263 a_37339_13912# a_36298_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2264 a_30701_18584# a_31690_19166# a_31646_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2265 a_13429_6923# a_13153_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2266 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2267 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2268 VDD C[13] a_35466_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2269 VDD a_59439_19374# a_59389_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2270 a_57289_5630# a_56841_6923# a_56442_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2271 a_52637_518# a_53580_861# a_53538_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2272 VSS C[29] a_5264_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2273 a_8051_18040# a_9056_18802# a_9000_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2274 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2275 a_53517_6668# a_53065_6923# a_52666_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2276 a_51629_6668# a_50901_6923# a_50778_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2277 VSS a_55401_5630# a_55928_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2278 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2279 a_17485_18583# a_18490_18802# a_18430_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2280 a_59439_19374# a_59015_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2281 a_45202_5834# a_44079_5630# a_45120_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2282 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2283 VDD a_26858_14117# a_27385_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2284 a_35655_1556# a_35711_1079# a_34706_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2285 a_42029_18584# a_43018_19167# a_42974_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2286 VDD C[9] a_43018_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2287 a_43917_18584# a_44906_19167# a_44862_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2288 VDD a_42191_5630# a_42718_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2289 a_44866_18261# a_44906_19167# a_43917_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2290 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2291 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2292 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2293 a_51400_13079# a_50948_12574# a_50549_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2294 VDD a_34643_6668# a_35166_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2295 a_46664_6923# a_46494_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2296 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2297 a_26134_12574# C[108] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2298 VDD a_34410_14117# a_34937_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2299 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2300 VSS a_9876_13079# a_10399_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2301 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2302 VSS a_17909_18776# a_17859_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2303 a_37539_518# a_37599_1079# a_36594_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2304 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18541_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2305 a_10569_12573# a_10399_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2306 a_33686_12574# C[112] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2307 a_33792_6629# a_32755_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2308 VDD a_20591_670# a_20607_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2309 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2310 VSS a_23573_18776# a_23523_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2311 a_9107_13912# a_7984_14117# a_9025_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2312 a_31904_5835# a_30863_5629# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2313 a_55401_5630# a_54677_6923# a_54554_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2314 a_42682_1105# a_42258_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2315 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2316 a_58305_1556# a_58361_1079# a_57356_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2317 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2318 a_16233_12574# a_16063_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2319 VSS a_22479_670# a_22495_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2320 VDD C[88] a_13045_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2321 a_58330_6629# a_58729_6923# a_59181_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2322 a_28771_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2323 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2324 a_3017_12573# a_2847_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2325 a_46773_13118# a_47172_12574# a_47624_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2326 a_18659_518# a_19602_861# a_19560_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2327 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2328 VDD a_45742_13080# a_46265_12574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2329 a_45971_6667# a_45519_6922# a_45120_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2330 a_52412_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2331 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2332 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2333 a_9225_518# a_9285_1079# a_8280_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2334 a_18434_18261# a_18490_18802# a_17485_18583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2335 VSS a_24367_670# a_24383_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2336 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2337 a_19373_18040# a_20362_19167# a_20322_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2338 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_37421_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2339 a_37018_507# a_36594_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2340 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2341 a_15540_13080# a_15088_12575# a_14689_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2342 VSS a_61065_5629# a_60193_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2343 VSS a_42453_18776# a_42403_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2344 a_22206_19299# a_22250_19167# a_21261_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2345 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2346 VSS a_55172_14117# a_55699_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2347 a_27112_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2348 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2349 a_55869_13117# a_55699_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2350 a_47172_12574# a_46896_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2351 a_48317_12573# a_48147_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2352 VDD a_25203_6668# a_25726_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2353 VDD C[76] a_35695_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2354 VSS a_49804_1405# a_48865_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2355 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2356 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2357 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2358 a_27154_1405# a_28159_1079# a_28103_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2359 a_32589_18039# a_33578_19167# a_33538_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2360 a_16571_13118# a_15540_13080# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2361 a_35422_19299# a_35466_19167# a_34477_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2362 a_54724_12574# a_54448_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2363 a_17199_6923# a_16923_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2364 a_10105_6668# a_9377_6923# a_9254_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2365 VSS C[75] a_37583_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2366 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2367 a_37314_18261# a_37370_18802# a_36365_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2368 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2369 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_48661_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2370 a_22235_13118# a_21198_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2371 a_5478_6629# a_4441_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2372 a_23336_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2373 a_41086_19299# a_41130_19167# a_40141_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2374 a_44891_13913# a_45290_12575# a_45738_14118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2375 a_3590_5835# a_1013_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2376 a_57064_13079# a_56336_12574# a_56213_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2377 a_58952_13079# a_58224_12574# a_58101_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2378 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2379 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2380 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_5331_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2381 a_40370_861# a_41375_1079# a_41315_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2382 a_48972_5835# a_47849_5630# a_48890_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2383 VSS a_27154_861# a_26211_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2384 a_23378_1405# a_24383_1079# a_24327_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2385 a_56213_13118# a_56336_12574# a_57064_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2386 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2387 a_35451_13118# a_34414_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2388 a_32589_18039# a_33594_18802# a_33538_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2389 VDD a_4699_19374# a_4649_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2390 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2391 a_56295_13118# a_55176_13079# a_56213_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2392 VSS a_51692_1405# a_50753_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2393 a_41115_13118# a_40078_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2394 VDD C[5] a_50564_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2395 a_9225_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2396 a_20429_13912# a_19306_14117# a_20347_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2397 a_50860_6629# a_49741_6668# a_50778_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2398 VSS a_33242_507# a_33192_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2399 a_53580_1405# a_54569_670# a_54529_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2400 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2401 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2402 a_20232_6380# a_20062_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2403 a_61069_6667# a_60617_6922# a_60218_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2404 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2405 VDD a_18138_1105# a_18088_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2406 a_11785_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2407 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2408 a_28103_1556# a_29042_1405# a_29000_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2409 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2410 a_59964_18261# a_60004_19167# a_59015_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2411 VSS a_38419_6668# a_38942_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2412 VDD a_54004_1105# a_53954_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2413 a_44104_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2414 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2415 a_35422_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2416 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2417 a_2345_18065# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2418 a_33645_13912# a_32522_14117# a_33563_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2419 VSS a_13652_13079# a_14175_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2420 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2421 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2422 a_25982_19299# a_26042_18802# a_25037_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2423 a_49804_1405# a_50793_670# a_50753_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2424 a_44146_1405# a_45151_1079# a_45095_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2425 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2426 a_59244_861# a_60233_670# a_60189_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2427 a_26363_6923# C[44] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2428 a_3565_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2429 a_48890_5835# a_49289_6923# a_49737_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2430 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2431 VSS a_6100_13079# a_6623_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2432 a_12686_6924# a_12516_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2433 a_34901_19374# a_34477_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2434 a_33534_19299# a_33594_18802# a_32589_18039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2435 a_57060_14117# a_56336_12574# a_56213_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2436 a_31331_12574# a_31161_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2437 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2438 a_54210_6380# a_54040_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2439 a_52666_5835# a_52789_6923# a_53513_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2440 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2441 VDD a_60840_13080# a_61363_12574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2442 a_58330_6629# a_57293_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2443 a_56442_5835# a_55401_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2444 VSS a_49999_18776# a_49949_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2445 a_60112_12575# C[126] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2446 VSS a_44146_861# a_43203_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2447 VDD a_50228_507# a_50178_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2448 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2449 a_44862_19299# a_44922_18802# a_43917_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2450 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2451 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_52519_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2452 a_30638_13080# a_30186_12575# a_29787_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2453 a_29672_6380# a_29502_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2454 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2455 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2456 VSS a_58948_14117# a_59475_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2457 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2458 a_50434_6380# a_50264_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2459 a_15765_5629# a_15317_6922# a_14918_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2460 a_14345_13117# a_14175_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2461 a_11827_18584# a_12832_18802# a_12772_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2462 VDD a_21685_18776# a_21635_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2463 a_54554_6629# a_53517_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2464 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2465 a_52666_5835# a_51625_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2466 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2467 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2468 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2469 VSS a_36365_18040# a_35426_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2470 a_6793_13117# a_6623_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2471 a_50778_5835# a_51177_6923# a_51625_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2472 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2473 a_52412_18261# a_52468_18802# a_51463_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2474 a_14889_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2475 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2476 a_45095_1556# a_46034_1405# a_45992_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2477 VDD a_33013_18776# a_32963_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2478 a_43917_18040# a_44906_19167# a_44866_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2479 a_16923_6923# C[39] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2480 VDD a_34901_18776# a_34851_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2481 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_46773_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2482 a_57780_1105# a_57356_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2483 VDD C[89] a_11157_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2484 a_10363_18776# a_9939_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2485 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_14689_13913# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2486 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_52748_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2487 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_9107_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2488 a_59989_13913# a_60388_12575# a_60836_14118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2489 VSS a_53517_6668# a_54040_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2490 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_14918_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2491 a_9229_1556# a_9285_1079# a_8280_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2492 a_30888_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2493 VDD a_40565_18776# a_40515_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2494 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2495 VSS a_6329_6668# a_6852_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2496 a_41319_1556# a_41359_670# a_40370_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2497 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2498 a_1473_13118# a_1596_12574# a_2324_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2499 a_43355_6923# C[53] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2500 a_923_18775# a_1013_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2501 a_48661_13912# a_48784_12574# a_49508_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2502 a_27870_19299# a_28813_18584# a_28771_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2503 a_56213_13912# a_55172_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2504 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2505 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2506 VSS a_33578_19167# a_33594_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2507 a_50549_13118# a_49512_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2508 a_56417_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2509 a_47874_1682# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2510 a_1555_13118# a_1242_317# a_1473_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2511 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_11224_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2512 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2513 a_50948_12574# a_50672_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2514 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2515 a_60189_518# a_60249_1079# a_59244_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2516 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2517 a_33534_19299# a_34477_18584# a_34435_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2518 VSS a_49741_6668# a_50264_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2519 a_32818_862# a_33823_1079# a_33763_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2520 a_48111_19374# a_47687_18583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2521 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2522 a_59874_6380# a_59704_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2523 a_11142_5835# a_11265_6923# a_11989_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2524 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2525 a_24751_6923# a_24475_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2526 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2527 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2528 a_19797_19374# a_19373_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2529 a_55663_19374# a_55239_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2530 a_19539_6668# a_18811_6923# a_18688_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2531 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2532 a_38440_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2533 a_1152_508# a_1242_317# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2534 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2535 VSS a_59015_18584# a_58072_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2536 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2537 a_49508_14117# a_48784_12574# a_48661_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2538 a_35655_1556# a_36594_1405# a_36552_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2539 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2540 a_8009_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2541 VSS a_47916_862# a_46973_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2542 a_24327_1556# a_24383_1079# a_23378_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2543 a_39427_518# a_39471_670# a_38482_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2544 a_20547_518# a_20591_670# a_19602_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2545 a_55468_861# a_56473_1079# a_56413_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2546 VDD C[24] a_14704_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2547 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_9025_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2548 a_60193_1556# a_60249_1079# a_59244_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2549 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2550 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2551 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2552 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2553 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2554 a_23086_13079# a_22634_12574# a_22235_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2555 a_33915_6923# C[48] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2556 VSS a_46452_1106# a_46402_887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2557 a_57780_1105# a_57356_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2558 a_8280_861# a_9269_670# a_9225_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2559 VSS a_15832_1405# a_14893_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2560 a_38677_19374# a_38253_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2561 a_24974_13079# a_24522_12574# a_24123_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2562 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2563 a_60071_13913# a_58948_14117# a_59989_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2564 a_6163_18584# a_7152_19167# a_7108_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2565 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2566 VSS a_6392_861# a_5449_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2567 a_2616_1406# a_3621_1079# a_3565_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2568 a_9000_18261# a_9040_19167# a_8051_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2569 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2570 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2571 a_18659_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2572 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2573 a_53309_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2574 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2575 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2576 a_37224_6924# a_37054_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2577 a_27087_5630# a_26639_6923# a_26240_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2578 a_59960_19299# a_60020_18802# a_59015_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2579 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_56295_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2580 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_31904_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2581 VSS a_59181_6668# a_59704_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2582 VSS a_48340_507# a_48290_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2583 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2584 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2585 VDD a_11764_13079# a_12287_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2586 a_23315_6668# a_22863_6923# a_22464_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2587 a_30139_6922# C[46] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2588 a_21427_6668# a_20699_6923# a_20576_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2589 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2590 a_12924_12574# C[101] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2591 a_20699_6923# C[41] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2592 a_39579_6923# C[51] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2593 VSS a_923_19373# a_873_19154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2594 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2595 a_43854_13079# a_43402_12574# a_43003_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2596 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_18688_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2597 a_25986_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2598 VDD a_4212_13079# a_4735_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2599 a_16462_6923# a_16292_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2600 VDD a_47017_671# a_47033_1080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2601 a_31875_519# a_31935_1080# a_30930_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2602 a_10888_18261# a_11827_18040# a_11785_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2603 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2604 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_60300_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2605 a_41315_518# a_41359_670# a_40370_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2606 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2607 a_41743_6923# a_41467_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2608 a_32303_6923# a_32027_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2609 a_33448_6924# a_33278_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2610 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2611 VSS a_18474_19167# a_18490_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2612 a_6163_18584# a_7168_18802# a_7108_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2613 a_31650_18260# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2614 a_7341_1556# a_8280_1405# a_8238_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2615 VSS a_51463_18040# a_50524_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2616 VSS a_14139_18776# a_14089_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2617 a_23378_861# a_24367_670# a_24323_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2618 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2619 VDD a_6816_1105# a_6766_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2620 a_14139_18776# a_13715_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2621 a_59960_19299# a_60004_19167# a_59015_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2622 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2623 a_27555_13117# a_27385_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2624 a_12480_507# a_12056_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2625 a_27578_507# a_27154_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2626 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2627 a_17422_13079# a_16694_12574# a_16571_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2628 a_5601_6923# C[33] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2629 VDD C[63] a_60233_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2630 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2631 a_63421_12573# a_63251_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2632 a_28128_6629# a_28527_6923# a_28979_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2633 a_26410_12574# a_26134_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2634 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2635 VSS a_46223_19373# a_46173_19154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2636 a_44866_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2637 a_1473_13912# a_1242_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2638 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_44973_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2639 a_33219_13117# a_33049_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2640 a_48784_12574# C[120] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2641 a_15769_6667# a_15317_6922# a_14918_5834# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2642 a_3565_1556# a_4504_1405# a_4462_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2643 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2644 a_6587_18776# a_6163_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2645 a_10913_13912# a_11312_12574# a_11760_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2646 a_1673_519# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2647 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2648 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2649 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2650 a_46664_6923# a_46494_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2651 a_33242_1105# a_32818_1406# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2652 VSS a_39242_19167# a_39258_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2653 a_48865_1556# a_48921_1079# a_47916_862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2654 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2655 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2656 a_55426_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2657 a_1473_13912# a_1872_12574# a_2320_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2658 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_39456_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2659 a_13902_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2660 a_61877_13118# a_60840_13080# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2661 VSS a_44906_19167# a_44922_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2662 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_20347_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2663 a_33767_1556# a_33807_670# a_32818_862# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2664 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2665 a_46034_1405# a_47017_671# a_46977_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2666 VSS a_59439_19374# a_59389_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2667 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2668 a_36302_13079# a_35574_12574# a_35451_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2669 a_44079_5630# a_43631_6923# a_43232_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2670 a_55468_1405# a_56473_1079# a_56417_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2671 a_8910_6380# a_8740_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2672 VSS a_19602_1405# a_18663_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2673 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2674 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2675 VSS a_42191_5630# a_42718_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2676 a_59439_19374# a_59015_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2677 a_30659_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2678 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2679 a_24008_6924# a_23838_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2680 a_35451_13118# a_35574_12574# a_36302_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2681 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_37568_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2682 a_20322_18261# a_20362_19167# a_19373_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2683 VSS C[7] a_46788_19166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2684 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_39227_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2685 a_5134_6924# a_4964_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2686 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_35680_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2687 VDD a_21914_1105# a_21864_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2688 a_54296_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2689 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2690 a_15536_14118# a_14812_12575# a_14689_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2691 VDD C[81] a_26255_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2692 a_11827_18040# a_12832_18802# a_12776_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2693 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2694 a_31875_519# a_32818_862# a_32776_888# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2695 a_52322_6380# a_52152_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2696 VSS a_55468_861# a_54525_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2697 a_51692_1405# a_52697_1079# a_52641_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2698 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2699 VDD C[16] a_29802_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2700 VSS C[80] a_28143_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2701 a_56417_1556# a_56457_670# a_55468_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2702 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2703 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_31986_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2704 a_18770_5835# a_17647_5630# a_18688_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2705 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2706 a_28750_13079# a_28298_12574# a_27899_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2707 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2708 a_53775_19374# a_53351_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2709 a_37967_6923# a_37691_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2710 a_42191_5630# a_41467_6923# a_41344_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2711 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2712 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2713 VDD a_21194_14117# a_21721_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2714 VSS a_45742_13080# a_46265_12574# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2715 VSS a_6816_1105# a_6766_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2716 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2717 a_20470_12574# C[105] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2718 VSS a_21490_1405# a_20551_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2719 a_1242_861# a_1717_671# a_1677_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2720 a_37018_507# a_36594_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2721 a_12883_13912# a_11760_14117# a_12801_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2722 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2723 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2724 VDD a_32522_14117# a_33049_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2725 a_56417_1556# a_57356_1405# a_57314_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2726 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2727 VSS a_19306_14117# a_19833_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2728 a_48317_12573# a_48147_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2729 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2730 VDD a_40074_14117# a_40601_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2731 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2732 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2733 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2734 VDD a_11993_6668# a_12516_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2735 a_54677_6923# C[59] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2736 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_7366_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2737 VSS a_55239_18040# a_54300_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2738 a_19602_1405# a_20591_670# a_20551_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2739 a_46435_13118# a_46265_13118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2740 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_22546_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2741 a_18688_5835# a_19087_6923# a_19535_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2742 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2743 a_16546_18260# a_17485_18039# a_17443_18065# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2744 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2745 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2746 VSS a_38186_14117# a_38713_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2747 a_9653_6923# a_9377_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2748 a_22464_5835# a_22587_6923# a_23311_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2749 VSS C[94] a_1717_671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2750 a_24098_18261# a_24154_18802# a_23149_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2751 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_60071_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2752 a_28128_6629# a_27091_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2753 a_35762_5835# a_34639_5630# a_35680_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2754 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2755 a_7448_6629# a_6329_6668# a_7366_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2756 a_35680_6629# a_36079_6923# a_36531_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2757 a_26240_5835# a_25199_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2758 a_37568_6629# a_37691_6923# a_38419_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2759 a_57986_6380# a_57816_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2760 VSS a_52452_19167# a_52468_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2761 VDD a_32751_5630# a_33278_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2762 VSS a_54340_19167# a_54356_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2763 VDD a_31354_1106# a_31304_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2764 VDD a_5264_19167# a_5280_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2765 a_31650_18260# a_31706_18801# a_30701_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2766 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2767 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2768 a_53065_6923# a_52789_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2769 VSS a_4699_19374# a_4649_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2770 VDD a_12251_18776# a_12201_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2771 VSS a_60004_19167# a_60020_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2772 a_6163_18040# a_7152_19167# a_7112_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2773 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_24123_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2774 a_20232_6380# a_20062_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2775 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2776 a_8996_19299# a_9040_19167# a_8051_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2777 a_24352_6629# a_23315_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2778 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2779 a_18434_18261# a_18474_19167# a_17485_18583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2780 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2781 a_51400_13079# a_50672_12574# a_50549_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2782 VDD a_14368_507# a_14318_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2783 a_22464_5835# a_21423_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2784 a_40370_1405# a_41359_670# a_41319_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2785 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2786 a_42978_18261# a_43034_18802# a_42029_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2787 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2788 a_21261_18584# a_22250_19167# a_22206_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2789 a_19373_18040# a_20378_18802# a_20322_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2790 VDD a_13045_670# a_13061_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2791 a_22634_12574# a_22358_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2792 VSS C[74] a_39471_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2793 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2794 a_24098_18261# a_24138_19167# a_23149_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2795 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_54325_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2796 a_50549_13118# a_50672_12574# a_51400_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2797 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_45120_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2798 a_8280_861# a_9285_1079# a_9225_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2799 a_4699_18776# a_4275_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2800 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2801 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2802 VSS a_19373_18584# a_18430_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2803 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2804 a_30634_14118# a_29910_12575# a_29787_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2805 VSS a_14933_670# a_14949_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2806 a_39309_13118# a_38190_13079# a_39227_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2807 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_43003_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2808 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2809 VDD C[14] a_33578_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2810 VDD a_57551_19374# a_57501_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2811 a_9025_13118# a_7988_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2812 VSS C[30] a_3376_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2813 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2814 a_19306_14117# a_18858_12574# a_18459_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2815 a_13153_6923# C[37] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2816 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2817 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2818 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2819 VDD a_24970_14117# a_25497_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2820 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2821 VDD a_61069_6667# a_61592_6923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2822 a_48340_1105# a_47916_1406# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2823 a_40141_18584# a_41130_19167# a_41086_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2824 VDD C[10] a_41130_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2825 VSS a_60840_13080# a_61363_12574# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2826 a_45519_6922# a_45243_6922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2827 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2828 a_34901_19374# a_34477_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2829 a_7366_6629# a_7765_6923# a_8217_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2830 VDD a_23311_5630# a_23838_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2831 VDD a_35695_670# a_35711_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2832 a_26215_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2833 a_17672_1682# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2834 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2835 a_42978_18261# a_43018_19167# a_42029_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2836 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2837 a_15540_13080# a_14812_12575# a_14689_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2838 a_24246_12574# C[107] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2839 a_39456_5835# a_39579_6923# a_40303_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2840 VSS a_50228_507# a_50178_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2841 a_29000_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2842 VSS a_38253_18584# a_37310_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2843 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2844 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2845 VSS a_19539_6668# a_20062_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2846 VSS a_37583_670# a_37599_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2847 a_43232_5835# a_42191_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2848 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2849 a_29672_6380# a_29502_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2850 a_18659_518# a_18719_1079# a_17714_1406# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2851 a_20318_19299# a_20378_18802# a_19373_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2852 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2853 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_16653_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2854 a_14689_13119# a_14812_12575# a_15540_13080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2855 a_38186_14117# a_37738_12574# a_37339_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2856 a_31798_12574# C[111] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2857 a_7366_5835# a_7765_6923# a_8213_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2858 a_19331_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2859 a_7219_13912# a_6096_14117# a_7137_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2860 VDD a_20026_1105# a_19976_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2861 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2862 VSS a_21685_18776# a_21635_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2863 a_60903_18584# a_62276_12574# a_61877_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2864 a_3590_6629# a_3989_6923# a_4441_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2865 VDD a_44570_1105# a_44520_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2866 VDD a_43850_14117# a_44377_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2867 a_23378_861# a_24383_1079# a_24323_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2868 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2869 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_9336_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2870 a_26883_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2871 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_27981_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2872 a_46973_519# a_47916_862# a_47874_888# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2873 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2874 VSS a_17714_862# a_16771_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2875 a_4928_1105# a_4504_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2876 VSS a_33013_18776# a_32963_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2877 a_50524_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2878 a_45014_12575# C[118] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2879 a_55405_6668# a_54953_6923# a_54554_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2880 VSS a_34901_18776# a_34851_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2881 a_61533_13118# a_61363_13118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2882 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2883 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35533_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2884 a_8704_1105# a_8280_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2885 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2886 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2887 a_46744_19298# a_47687_18583# a_47645_18859# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2888 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2889 VSS a_16250_1106# a_16200_887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2890 a_20318_19299# a_20362_19167# a_19373_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2891 a_56213_13118# a_56612_12574# a_57064_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2892 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2893 VSS a_40565_18776# a_40515_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2894 VSS a_53284_14117# a_53811_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2895 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2896 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2897 a_55401_5630# a_54953_6923# a_54554_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2898 a_27874_18261# a_27930_18802# a_26925_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2899 a_29762_18261# a_29818_18802# a_28813_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2900 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2901 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2902 a_45763_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2903 a_51629_6668# a_51177_6923# a_50778_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2904 VDD a_16250_508# a_16200_343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2905 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2906 a_45120_6628# a_45243_6922# a_45971_6667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2907 VSS a_28979_6668# a_29502_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2908 a_33534_19299# a_33578_19167# a_32589_18039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2909 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_10995_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2910 a_47916_862# a_48921_1079# a_48861_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2911 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_12883_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2912 VDD a_40303_5630# a_40830_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2913 a_43207_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2914 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2915 a_20347_13118# a_19310_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2916 VSS a_41359_670# a_41375_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2917 a_59645_12573# a_59475_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2918 a_55176_13079# a_54448_12574# a_54325_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2919 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2920 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_3443_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2921 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_30098_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2922 a_35651_518# a_35711_1079# a_34706_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2923 a_11113_518# a_11157_670# a_10168_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2924 VDD a_8475_18776# a_8425_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2925 a_11541_6923# a_11265_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2926 a_31904_6629# a_30867_6667# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2927 a_19797_19374# a_19373_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2928 a_30016_5834# a_28975_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2929 a_1152_508# a_1242_317# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2930 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2931 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2932 a_28022_12574# C[109] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2933 a_54325_13118# a_54448_12574# a_55176_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2934 a_60903_18584# a_62000_12574# a_61877_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2935 a_53513_5630# a_52789_6923# a_52666_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2936 a_20318_19299# a_21261_18584# a_21219_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2937 a_39227_13912# a_38186_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2938 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_58101_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2939 a_48743_13118# a_47624_13079# a_48661_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2940 a_23802_1105# a_23378_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2941 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2942 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2943 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2944 a_33563_13118# a_32526_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2945 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2946 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2947 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2948 a_56442_6629# a_56841_6923# a_57293_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2949 VDD a_2811_19374# a_2761_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2950 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2951 a_47002_5835# a_45967_5629# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2952 a_43203_518# a_44146_861# a_44104_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2953 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2954 a_54407_13118# a_53288_13079# a_54325_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2955 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2956 a_7337_518# a_7397_1079# a_6392_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2957 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2958 a_39350_12574# C[115] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2959 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2960 a_2574_888# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2961 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2962 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2963 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2964 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2965 a_18138_507# a_17714_862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2966 a_38677_19374# a_38253_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2967 a_16462_6923# a_16292_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2968 a_44570_1105# a_44146_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2969 VDD a_46452_1106# a_46402_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2970 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2971 a_39198_19299# a_40141_18584# a_40099_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2972 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2973 a_25224_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2974 VSS a_53351_18584# a_52408_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2975 a_2616_862# a_3605_670# a_3561_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2976 a_33534_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2977 a_31757_13912# a_30634_14118# a_31675_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2978 VSS a_11764_13079# a_12287_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2979 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2980 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2981 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2982 a_60617_6922# a_60341_6922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2983 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_45202_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2984 a_24094_19299# a_24154_18802# a_23149_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2985 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2986 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2987 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2988 VDD a_4441_6668# a_4964_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2989 VDD C[67] a_52681_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2990 a_6816_507# a_6392_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2991 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2992 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2993 a_25461_19374# a_25037_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2994 a_25266_1405# a_26271_1079# a_26215_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2995 a_53284_14117# a_52836_12574# a_52437_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2996 a_29787_13119# a_29910_12575# a_30638_13080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2997 VSS C[85] a_18703_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2998 a_31125_19373# a_30701_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2999 VSS a_4212_13079# a_4735_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3000 VDD a_28143_670# a_28159_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3001 a_31646_19298# a_31706_18801# a_30701_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3002 VSS C[66] a_54569_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3003 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3004 a_55172_14117# a_54448_12574# a_54325_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3005 a_3590_6629# a_1013_19128# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3006 a_21448_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3007 VDD a_45967_5629# a_46494_6379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3008 a_29991_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3009 a_44973_13913# a_43850_14117# a_44891_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3010 a_48661_13118# a_49060_12574# a_49512_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3011 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3012 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3013 a_18430_19299# a_18474_19167# a_17485_18039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3014 a_60903_18040# a_62000_12574# a_61877_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3015 a_22120_6380# a_21950_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3016 a_48890_6629# a_49013_6923# a_49741_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3017 VSS a_25266_861# a_24323_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3018 a_21490_1405# a_22495_1079# a_22439_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3019 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3020 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3021 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3022 a_42974_19299# a_43034_18802# a_42029_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3023 a_27578_507# a_27154_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3024 a_46977_1557# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3025 a_44341_19374# a_43917_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3026 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3027 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_50631_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3028 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3029 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3030 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3031 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3032 VSS a_57060_14117# a_57587_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3033 a_27112_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3034 a_12457_13117# a_12287_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3035 a_9939_18584# a_10944_18802# a_10884_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3036 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3037 a_48890_5835# a_49013_6923# a_49737_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3038 VSS a_28813_18040# a_27874_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3039 a_30016_6628# a_30415_6922# a_30867_6667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3040 a_60861_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3041 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_61959_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3042 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3043 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3044 a_1013_19128# a_1504_18801# a_1444_19298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3045 a_48636_18261# a_49575_18040# a_49533_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3046 a_4905_13117# a_4735_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3047 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3048 a_50524_18261# a_50580_18802# a_49575_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3049 VSS a_34477_18040# a_33538_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3050 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3051 a_26215_1556# a_27154_1405# a_27112_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3052 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3053 VSS a_20026_1105# a_19976_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3054 a_42216_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3055 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3056 VDD a_59668_1105# a_59618_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3057 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3058 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3059 a_21891_13117# a_21721_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3060 a_8910_6380# a_8740_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3061 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3062 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3063 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3064 a_48661_13912# a_47620_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3065 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3066 a_48340_1105# a_47916_1406# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3067 a_42258_1405# a_43263_1079# a_43207_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3068 a_24475_6923# C[43] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3069 a_24094_19299# a_25037_18584# a_24995_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3070 a_25982_19299# a_26925_18584# a_26883_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3071 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3072 a_47002_5835# a_47401_6923# a_47849_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3073 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3074 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3075 a_54325_13912# a_53284_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3076 a_10798_6924# a_10628_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3077 a_18430_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3078 a_48661_13912# a_49060_12574# a_49508_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3079 a_52322_6380# a_52152_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3080 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3081 VDD a_16021_19373# a_15971_19154# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3082 a_56442_6629# a_55405_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3083 a_58101_13912# a_58224_12574# a_58948_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3084 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3085 a_40771_13117# a_40601_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3086 VSS a_42258_861# a_41315_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3087 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3088 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3089 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3090 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3091 a_17909_19374# a_17485_18583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3092 a_59989_13119# a_58952_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3093 a_39431_1556# a_39487_1079# a_38482_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3094 a_46223_18775# a_45805_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3095 a_27784_6380# a_27614_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3096 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3097 a_53775_19374# a_53351_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3098 a_29869_13913# a_28746_14117# a_29787_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3099 a_60388_12575# a_60112_12575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3100 a_62000_12574# C[127] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3101 VDD a_40794_507# a_40744_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3102 a_44862_19299# a_45805_18584# a_45763_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3103 VSS a_39471_670# a_39487_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3104 a_50753_1556# a_50793_670# a_49804_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3105 VSS a_57127_18584# a_56184_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3106 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3107 VSS C[79] a_30031_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3108 a_37310_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3109 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_50860_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3110 a_52666_6629# a_51629_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3111 a_3565_1556# a_3621_1079# a_2616_862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3112 VSS a_29466_1105# a_29416_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3113 a_29237_19374# a_28813_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3114 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3115 VSS a_8217_6668# a_8740_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3116 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3117 VDD C[25] a_12816_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3118 VDD a_36789_19374# a_36739_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3119 a_57060_14117# a_56612_12574# a_56213_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3120 a_58948_14117# a_58500_12574# a_58101_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3121 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_7137_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3122 a_13715_18584# a_14704_19167# a_14660_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3123 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3124 a_43207_1556# a_44146_1405# a_44104_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3125 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3126 a_36789_19374# a_36365_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3127 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3128 a_21198_13079# a_20746_12574# a_20347_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3129 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3130 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_14918_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3131 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3132 a_61762_6379# a_61592_6379# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3133 a_4275_18584# a_5264_19167# a_5220_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3134 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3135 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3136 a_7112_18261# a_7152_19167# a_6163_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3137 a_31354_508# a_30930_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3138 a_58301_518# a_59244_861# a_59202_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3139 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3140 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3141 a_41467_6923# C[52] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3142 a_34414_13079# a_33962_12574# a_33563_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3143 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_54407_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3144 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3145 a_54529_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3146 sky130_fd_sc_hd__buf_2_0/X a_28116_9428# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3147 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3148 VDD a_30867_6667# a_31390_6923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3149 a_13715_18584# a_14720_18802# a_14660_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3150 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3151 VDD a_15540_13080# a_16063_12574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3152 a_40078_13079# a_39626_12574# a_39227_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3153 a_41966_13079# a_41514_12574# a_41115_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3154 a_15317_6922# a_15041_6922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3155 a_38482_861# a_39471_670# a_39427_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3156 a_22210_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3157 VDD a_2324_13079# a_2847_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3158 a_24098_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3159 VDD a_7984_14117# a_8511_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3160 VSS a_32751_5630# a_33278_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3161 a_57986_6380# a_57816_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3162 a_9254_5835# a_9377_6923# a_10101_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3163 a_4928_507# a_4504_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3164 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3165 a_22863_6923# a_22587_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3166 a_49804_861# a_50809_1079# a_50749_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3167 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3168 a_4275_18584# a_5280_18802# a_5220_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3169 a_13030_5835# a_11989_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3170 a_7260_12574# C[98] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3171 a_44776_6380# a_44606_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3172 a_50753_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3173 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3174 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3175 VSS a_12251_18776# a_12201_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3176 a_59989_13913# a_60112_12575# a_60836_14118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3177 VDD C[93] a_3605_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3178 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3179 a_19560_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3180 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3181 a_25667_13117# a_25497_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3182 VDD a_29466_507# a_29416_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3183 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3184 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3185 a_18115_12573# a_17945_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3186 a_20003_12573# a_19833_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3187 VSS a_14368_507# a_14318_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3188 VSS C[92] a_5493_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3189 a_37539_518# a_37583_670# a_36594_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3190 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3191 VSS a_61069_6667# a_61592_6923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3192 a_42978_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3193 a_24522_12574# a_24246_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3194 a_46896_12574# C[119] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3195 a_4699_18776# a_4275_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3196 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3197 VDD a_35130_1105# a_35080_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3198 a_55892_1105# a_55468_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3199 VSS a_13944_1405# a_13005_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3200 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3201 VSS a_35466_19167# a_35482_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3202 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3203 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18459_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3204 a_32027_6923# C[47] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3205 VSS a_37354_19167# a_37370_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3206 a_9939_18040# a_10928_19167# a_10888_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3207 a_10884_19299# a_10928_19167# a_9939_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3208 a_14689_13913# a_15088_12575# a_15536_14118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3209 a_12772_19299# a_12816_19167# a_11827_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3210 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3211 a_28750_13079# a_28022_12574# a_27899_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3212 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3213 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3214 VDD a_58116_19167# a_58132_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3215 a_1013_18584# a_1488_19166# a_1448_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3216 a_44547_13117# a_44377_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3217 a_20026_507# a_19602_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3218 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3219 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3220 VSS a_57551_19374# a_57501_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3221 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3222 a_38883_12573# a_38713_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3223 a_25199_5630# a_24751_6923# a_24352_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3224 a_44570_507# a_44146_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3225 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3226 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3227 a_34414_13079# a_33686_12574# a_33563_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3228 a_27899_13118# a_28022_12574# a_28750_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3229 VSS a_57293_6668# a_57816_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3230 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3231 a_21427_6668# a_20975_6923# a_20576_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3232 VSS a_23311_5630# a_23838_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3233 a_38419_6668# a_37691_6923# a_37568_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3234 a_46977_1557# a_47916_1406# a_47874_1682# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3235 a_43402_12574# a_43126_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3236 a_59960_19299# a_60903_18584# a_60861_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3237 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_18688_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3238 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_37339_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3239 a_26093_13118# a_24974_13079# a_26011_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3240 a_33563_13118# a_33686_12574# a_34414_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3241 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_16800_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3242 VDD C[21] a_20362_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3243 a_52408_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3244 a_27981_13118# a_26862_13079# a_27899_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3245 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_31675_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3246 VDD a_10101_5630# a_10628_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3247 a_12801_13118# a_11764_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3248 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3249 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3250 a_9939_18040# a_10944_18802# a_10888_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3251 a_14893_1556# a_14949_1079# a_13944_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3252 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3253 a_2320_14117# a_1872_12574# a_1473_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3254 a_21423_5630# a_20975_6923# a_20576_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3255 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3256 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3257 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3258 VDD a_30031_670# a_30047_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3259 a_5453_1556# a_6392_1405# a_6350_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3260 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3261 a_1013_18584# a_1504_18801# a_1448_18260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3262 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3263 a_49999_19374# a_49575_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3264 a_26862_13079# a_26410_12574# a_26011_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3265 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3266 a_9225_518# a_9269_670# a_8280_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3267 a_51887_19374# a_51463_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3268 VSS C[2] a_56228_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3269 VSS C[1] a_58116_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3270 a_23311_5630# a_22587_6923# a_22464_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3271 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3272 VSS a_1717_671# a_1733_1080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3273 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3274 a_8051_18584# a_9040_19167# a_8996_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3275 VDD C[27] a_9040_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3276 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3277 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3278 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3279 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3280 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3281 VDD C[11] a_39242_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3282 a_3713_6923# C[32] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3283 a_26240_6629# a_26639_6923# a_27091_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3284 a_37539_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3285 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3286 a_48546_6380# a_48376_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3287 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3288 a_10995_13912# a_9872_14117# a_10913_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3289 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3290 a_42195_6668# a_41743_6923# a_41344_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3291 VDD a_52681_670# a_52697_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3292 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3293 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3294 a_50228_1105# a_49804_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3295 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3296 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_39456_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3297 VSS a_17418_14117# a_17945_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3298 VDD a_55892_507# a_55842_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3299 VDD a_30638_13080# a_31161_12574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3300 VSS a_16250_508# a_16200_343# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3301 VSS a_54569_670# a_54585_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3302 a_27874_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3303 a_34410_14117# a_33686_12574# a_33563_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3304 a_13030_5835# a_13429_6923# a_13877_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3305 a_30888_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3306 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3307 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3308 a_9377_6923# C[35] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3309 a_42191_5630# a_41743_6923# a_41344_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3310 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3311 a_7022_6380# a_6852_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3312 a_30930_1405# a_31919_671# a_31879_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3313 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3314 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3315 a_30415_6922# a_30139_6922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3316 VSS a_40303_5630# a_40830_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3317 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_15000_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3318 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3319 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3320 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3321 VSS a_28746_14117# a_29273_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3322 VDD a_55405_6668# a_55928_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3323 a_59645_12573# a_59475_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3324 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_35680_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3325 VDD a_10592_1105# a_10542_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3326 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_33792_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3327 a_7108_19299# a_7168_18802# a_6163_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3328 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3329 a_47401_6923# a_47125_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3330 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3331 VSS a_36298_14117# a_36825_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3332 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3333 VSS a_8475_18776# a_8425_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3334 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3335 VDD a_15765_5629# a_16292_6379# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3336 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3337 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3338 a_28298_12574# a_28022_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3339 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3340 a_46452_508# a_46034_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3341 a_22210_18261# a_22266_18802# a_21261_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3342 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3343 a_16882_5835# a_15765_5629# a_16800_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3344 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3345 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3346 a_18688_6629# a_18811_6923# a_19539_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3347 VSS a_50564_19167# a_50580_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3348 a_13715_18040# a_14704_19167# a_14664_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3349 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_16571_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3350 a_40303_5630# a_39579_6923# a_39456_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3351 a_16775_1557# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3352 a_39431_1556# a_39471_670# a_38482_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3353 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3354 VDD a_3376_19167# a_3392_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3355 a_29787_13913# a_30186_12575# a_30634_14118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3356 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3357 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3358 VSS a_2811_19374# a_2761_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3359 VDD a_10363_18776# a_10313_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3360 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3361 a_43232_6629# a_43631_6923# a_44083_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3362 a_28975_5630# a_28251_6923# a_28128_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3363 VSS a_2387_18583# a_1444_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3364 a_4275_18040# a_5264_19167# a_5224_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3365 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3366 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3367 a_52093_12573# a_51923_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3368 a_41319_1556# a_41375_1079# a_40370_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3369 a_7108_19299# a_7152_19167# a_6163_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3370 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3371 a_53981_12573# a_53811_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3372 a_18688_5835# a_18811_6923# a_19535_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3373 VSS a_38482_1405# a_37543_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3374 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3375 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_9254_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3376 a_18138_507# a_17714_862# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3377 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3378 a_26011_13912# a_24970_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3379 a_27899_13912# a_26858_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3380 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_29787_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3381 a_37650_6629# a_36531_6668# a_37568_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3382 a_54529_1556# a_55468_1405# a_55426_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3383 a_41090_18261# a_41146_18802# a_40141_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3384 VSS C[78] a_31919_671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3385 a_5449_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3386 a_20746_12574# a_20470_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3387 VDD a_48111_19374# a_48061_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3388 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_52437_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3389 a_6816_507# a_6392_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3390 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3391 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3392 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3393 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_7366_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3394 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3395 VDD a_31690_19166# a_31706_18801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3396 a_52789_6923# C[58] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3397 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_5478_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3398 VSS a_34706_1405# a_33767_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3399 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3400 VDD a_55663_19374# a_55613_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3401 a_7137_13118# a_6100_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3402 a_6350_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3403 VSS a_1488_19166# a_1504_18801# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3404 a_25461_19374# a_25037_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3405 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3406 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3407 a_61877_13118# a_62000_12574# a_60903_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3408 a_36594_1405# a_37583_670# a_37543_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3409 a_12056_1405# a_13061_1079# a_13005_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3410 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3411 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3412 a_16800_5835# a_17199_6923# a_17647_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3413 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3414 a_31125_19373# a_30701_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3415 a_19306_14117# a_18582_12574# a_18459_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3416 a_60189_518# a_61069_6667# a_61090_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3417 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3418 a_2345_18859# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3419 a_56098_6924# a_55928_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3420 a_9225_518# a_10168_861# a_10126_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3421 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3422 a_7108_19299# a_8051_18584# a_8009_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3423 a_47645_18065# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3424 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3425 a_7765_6923# a_7489_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3426 a_22120_6380# a_21950_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3427 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3428 VSS a_36365_18584# a_35422_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3429 a_22358_12574# C[106] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3430 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_18770_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3431 a_38482_861# a_39487_1079# a_39427_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3432 a_26240_6629# a_25203_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3433 a_45243_6922# C[54] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3434 a_33874_5835# a_32751_5630# a_33792_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3435 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3436 a_35680_6629# a_35803_6923# a_36531_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3437 VSS a_12056_861# a_11113_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3438 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3439 a_40370_861# a_41359_670# a_41315_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3440 a_44341_19374# a_43917_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3441 a_36298_14117# a_35850_12574# a_35451_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3442 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3443 a_60189_518# a_60233_670# a_59244_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3444 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3445 a_51177_6923# a_50901_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3446 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3447 a_38186_14117# a_37462_12574# a_37339_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3448 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3449 a_23107_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3450 a_35680_5835# a_35803_6923# a_36527_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3451 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3452 a_24995_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3453 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_26093_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3454 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_20658_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3455 a_22464_6629# a_21427_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3456 a_41238_12574# C[116] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3457 a_7366_6629# a_7489_6923# a_8217_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3458 a_20576_5835# a_19535_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3459 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3460 a_39456_5835# a_38415_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3461 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3462 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3463 VSS C[84] a_20591_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3464 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_33645_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3465 a_37568_5835# a_37967_6923# a_38415_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3466 VSS C[71] a_45135_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3467 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3468 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3469 VSS a_49508_14117# a_50035_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3470 VSS a_51396_14117# a_51923_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3471 a_54325_13118# a_54724_12574# a_55176_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3472 a_45091_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3473 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3474 a_31560_6379# a_31390_6379# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3475 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_39538_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3476 a_30016_5834# a_30139_6922# a_30863_5629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3477 VSS a_21261_18040# a_20322_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3478 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3479 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3480 a_43875_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3481 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3482 a_61877_13118# a_62276_12574# a_60903_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3483 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_58330_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3484 a_35130_1105# a_34706_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3485 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3486 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3487 a_11265_6923# C[36] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3488 a_33792_5835# a_34191_6923# a_34639_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3489 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3490 VSS a_60903_18040# a_63251_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3491 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3492 a_5478_6629# a_5877_6923# a_6329_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3493 a_5560_5835# a_4437_5630# a_5478_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3494 a_24327_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3495 VDD a_16586_19166# a_16602_18801# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3496 VDD C[72] a_43247_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3497 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3498 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3499 a_57757_12573# a_57587_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3500 a_54210_6924# a_54040_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3501 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_35762_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3502 a_38906_1105# a_38482_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3503 VSS a_16021_19373# a_15971_19154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3504 a_18582_12574# C[104] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3505 a_53288_13079# a_52560_12574# a_52437_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3506 a_43232_6629# a_42195_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3507 VSS a_18703_670# a_18719_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3508 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3509 a_46773_13118# a_46896_12574# a_47624_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3510 VSS a_36531_6668# a_37054_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3511 a_41344_5835# a_40303_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3512 a_15832_1405# a_16831_1080# a_16775_1557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3513 a_46223_18775# a_45805_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3514 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1555_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3515 a_62276_12574# a_62000_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3516 a_27784_6380# a_27614_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3517 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3518 VSS a_40794_507# a_40744_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3519 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3520 VDD a_6587_18776# a_6537_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3521 VSS a_40141_18040# a_39202_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3522 a_17909_19374# a_17485_18583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3523 a_45202_6628# a_44083_6668# a_45120_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3524 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3525 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_56213_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3526 a_46855_13118# a_45742_13080# a_46773_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3527 a_14574_6380# a_14404_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3528 a_20551_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3529 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3530 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3531 a_31675_13118# a_30638_13080# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3532 VDD a_25690_1105# a_25640_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3533 VSS a_14704_19167# a_14720_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3534 VSS a_7381_670# a_7397_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3535 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3536 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3537 a_49741_6668# a_49013_6923# a_48890_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3538 VDD a_31919_671# a_31935_1080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3539 a_33767_1556# a_33823_1079# a_32818_862# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3540 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3541 a_50434_6924# a_50264_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3542 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3543 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3544 a_52519_13118# a_51400_13079# a_52437_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3545 a_13944_861# a_14949_1079# a_14889_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3546 a_29237_19374# a_28813_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3547 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3548 a_37462_12574# C[114] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3549 a_8681_13117# a_8511_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3550 VSS a_30867_6667# a_31390_6923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3551 VSS a_36789_19374# a_36739_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3552 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3553 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3554 VSS C[23] a_16586_19166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3555 a_25982_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3556 a_44891_13119# a_43854_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3557 a_49737_5630# a_49013_6923# a_48890_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3558 a_25690_1105# a_25266_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3559 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3560 a_36789_19374# a_36365_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3561 a_43126_12574# C[117] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3562 a_31354_508# a_30930_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3563 VSS a_59244_1405# a_58305_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3564 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3565 a_53513_5630# a_53065_6923# a_52666_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3566 VSS a_51463_18584# a_50520_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3567 a_61877_13912# a_62276_12574# a_60903_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3568 a_16250_1106# a_15832_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3569 a_56417_1556# a_56473_1079# a_55468_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3570 VDD a_8704_507# a_8654_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3571 a_23573_19374# a_23149_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3572 a_22206_19299# a_22266_18802# a_21261_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3573 VSS a_27091_6668# a_27614_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3574 a_4233_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3575 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3576 a_51396_14117# a_50948_12574# a_50549_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3577 VSS a_15540_13080# a_16063_12574# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3578 a_48861_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3579 a_16775_1557# a_17714_1406# a_17672_1682# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3580 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3581 VSS C[70] a_47017_671# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3582 a_41319_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3583 a_32776_1682# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3584 VSS a_2324_13079# a_2847_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3585 a_32776_888# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3586 a_4928_507# a_4504_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3587 a_16775_1557# a_16815_671# a_15832_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3588 a_44862_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3589 a_53284_14117# a_52560_12574# a_52437_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3590 a_60341_6922# C[62] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3591 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3592 a_58412_5835# a_57289_5630# a_58330_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3593 a_50901_6923# C[57] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3594 a_35130_507# a_34706_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3595 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3596 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3597 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3598 a_30016_6628# a_28979_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3599 a_44776_6380# a_44606_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3600 a_33763_518# a_33823_1079# a_32818_1406# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3601 a_58500_12574# a_58224_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3602 a_59874_6924# a_59704_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3603 a_32818_862# a_33807_670# a_33763_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3604 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3605 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3606 a_51625_5630# a_50901_6923# a_50778_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3607 VSS a_29466_507# a_29416_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3608 a_42453_19374# a_42029_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3609 a_41086_19299# a_41146_18802# a_40141_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3610 a_18115_12573# a_17945_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3611 VDD a_9872_14117# a_10399_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3612 a_20003_12573# a_19833_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3613 a_58101_13118# a_58500_12574# a_58952_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3614 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3615 VDD a_47624_13079# a_48147_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3616 a_47002_6629# a_45971_6667# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3617 a_54636_5835# a_53513_5630# a_54554_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3618 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3619 a_10569_13117# a_10399_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3620 a_24323_518# a_25266_861# a_25224_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3621 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3622 a_9876_13079# a_9424_12574# a_9025_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3623 VDD a_51625_5630# a_52152_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3624 VSS a_25037_18040# a_24098_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3625 VSS a_26925_18040# a_25986_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3626 VSS a_32818_862# a_31875_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3627 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3628 a_48972_6629# a_47853_6668# a_48890_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3629 VDD a_23802_507# a_23752_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3630 a_16233_13118# a_16063_13118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3631 a_18344_6380# a_18174_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3632 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3633 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3634 a_3017_13117# a_2847_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3635 a_42682_1105# a_42258_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3636 a_55468_861# a_56457_670# a_56413_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3637 VSS a_31354_1106# a_31304_887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3638 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3639 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3640 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3641 a_38883_12573# a_38713_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3642 a_20026_507# a_19602_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3643 a_59668_507# a_59244_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3644 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3645 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3646 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3647 a_44570_507# a_44146_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3648 a_59244_1405# a_60233_670# a_60193_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3649 a_15832_861# a_16831_1080# a_16771_519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3650 a_58076_18261# a_59015_18040# a_58973_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3651 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3652 a_46773_13912# a_45738_14118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3653 a_58330_5835# a_58729_6923# a_59177_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3654 VSS a_24138_19167# a_24154_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3655 a_29787_13119# a_28750_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3656 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3657 a_47916_1406# a_48905_670# a_48865_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3658 a_59964_18261# a_60020_18802# a_59015_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3659 VSS a_45805_18040# a_44866_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3660 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_1473_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3661 VSS a_44083_6668# a_44606_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3662 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3663 a_22206_19299# a_23149_18584# a_23107_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3664 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3665 VSS a_10101_5630# a_10628_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3666 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3667 a_14368_1105# a_13944_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3668 a_52437_13912# a_51396_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3669 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3670 a_30016_6628# a_30139_6922# a_30867_6667# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3671 a_13005_1556# a_13045_670# a_12056_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3672 a_5449_518# a_5509_1079# a_4504_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3673 VSS a_29802_19167# a_29818_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3674 a_46773_13912# a_47172_12574# a_47620_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3675 a_21448_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3676 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3677 a_45992_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3678 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3679 a_56213_13912# a_56336_12574# a_57060_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3680 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3681 a_52560_12574# C[122] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3682 a_47002_6629# a_47125_6923# a_47853_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3683 a_19602_1405# a_20607_1079# a_20551_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3684 a_39112_6380# a_38942_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3685 VSS a_23378_861# a_22435_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3686 a_38482_1405# a_39487_1079# a_39431_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3687 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3688 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3689 a_20347_13118# a_20470_12574# a_21198_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3690 a_58101_13912# a_58500_12574# a_58948_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3691 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3692 VSS a_43018_19167# a_43034_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3693 a_49999_19374# a_49575_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3694 a_51887_19374# a_51463_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3695 a_41086_19299# a_42029_18584# a_41987_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3696 a_42974_19299# a_43917_18584# a_43875_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3697 a_10101_5630# a_9377_6923# a_9254_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3698 a_48546_6380# a_48376_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3699 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3700 VDD a_27349_19374# a_27299_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3701 VSS a_55239_18584# a_54296_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3702 VDD C[64] a_58345_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3703 a_10592_507# a_10168_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3704 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3705 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3706 a_27349_19374# a_26925_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3707 a_35336_6380# a_35166_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3708 VDD a_3605_670# a_3621_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3709 a_55172_14117# a_54724_12574# a_54325_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3710 VDD C[26] a_10928_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3711 a_57551_18776# a_57127_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3712 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_5249_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3713 VSS a_30638_13080# a_31161_12574# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3714 VSS a_55892_507# a_55842_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3715 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3716 a_11827_18584# a_12816_19167# a_12772_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3717 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3718 a_39227_13118# a_39350_12574# a_40078_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3719 a_24327_1556# a_25266_1405# a_25224_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3720 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3721 a_14664_18261# a_14704_19167# a_13715_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3722 VSS a_5493_670# a_5509_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3723 a_58948_14117# a_58224_12574# a_58101_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3724 a_40328_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3725 VDD C[31] a_1488_19166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3726 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3727 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3728 a_7022_6380# a_6852_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3729 a_50749_518# a_51692_861# a_51650_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3730 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3731 a_2387_18583# a_3376_19167# a_3332_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3732 a_12056_861# a_13061_1079# a_13001_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3733 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3734 a_3760_12574# a_3484_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3735 VDD C[28] a_7152_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3736 a_5224_18261# a_5264_19167# a_4275_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3737 a_40370_1405# a_41375_1079# a_41319_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3738 a_22587_6923# C[42] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3739 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3740 a_32526_13079# a_32074_12574# a_31675_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3741 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3742 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3743 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3744 VDD a_42195_6668# a_42718_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3745 VDD a_13648_14117# a_14175_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3746 a_46452_508# a_46034_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3747 a_58301_518# a_58361_1079# a_57356_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3748 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3749 a_34191_6923# a_33915_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3750 a_38211_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3751 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_52748_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3752 a_20322_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3753 VDD a_6096_14117# a_6623_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3754 a_14812_12575# C[102] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3755 VSS a_47853_6668# a_48376_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3756 a_31331_13118# a_31161_13118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3757 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3758 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3759 a_15041_6922# C[38] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3760 a_16542_19298# a_17485_18583# a_17443_18859# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3761 a_5372_12574# C[97] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3762 VSS a_10363_18776# a_10313_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3763 a_25896_6380# a_25726_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3764 a_40794_1105# a_40370_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3765 VSS a_23082_14117# a_23609_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3766 VSS a_20591_670# a_20607_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3767 a_52093_12573# a_51923_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3768 a_53981_12573# a_53811_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3769 a_16970_12574# a_16694_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3770 a_47874_888# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3771 a_29987_518# a_30031_670# a_29042_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3772 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3773 a_23779_13117# a_23609_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3774 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3775 a_15561_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3776 a_33563_13118# a_33962_12574# a_34414_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3777 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3778 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3779 VSS C[88] a_13045_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3780 a_18659_518# a_18703_670# a_17714_1406# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3781 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3782 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3783 a_39202_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3784 a_41090_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3785 VSS a_60903_18040# a_59964_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3786 a_47916_862# a_48905_670# a_48861_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3787 a_46973_519# a_47017_671# a_46034_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3788 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3789 a_41319_1556# a_42258_1405# a_42216_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3790 a_6121_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3791 VDD a_48676_19167# a_48692_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3792 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3793 VSS a_48111_19374# a_48061_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3794 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3795 a_29443_12573# a_29273_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3796 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3797 a_26862_13079# a_26134_12574# a_26011_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3798 VSS a_41962_14117# a_42489_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3799 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3800 a_1473_13912# a_1596_12574# a_2320_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3801 a_44891_13119# a_45290_12575# a_45742_13080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3802 VDD C[77] a_33807_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3803 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3804 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3805 a_35850_12574# a_35574_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3806 VDD a_19797_19374# a_19747_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3807 a_42659_13117# a_42489_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3808 a_35107_12573# a_34937_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3809 a_56336_12574# C[124] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3810 a_1444_19298# a_1488_19166# a_1013_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3811 a_36995_12573# a_36825_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3812 VSS a_55663_19374# a_55613_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3813 a_24123_13118# a_24246_12574# a_24974_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3814 a_26011_13118# a_26134_12574# a_26862_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3815 a_32526_13079# a_31798_12574# a_31675_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3816 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_27899_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3817 a_18541_13118# a_17422_13079# a_18459_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3818 VSS C[76] a_35695_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3819 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3820 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3821 a_41514_12574# a_41238_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3822 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_28128_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3823 VDD a_45135_670# a_45151_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3824 a_52641_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3825 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3826 a_9000_18261# a_9056_18802# a_8051_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3827 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3828 a_24205_13118# a_23086_13079# a_24123_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3829 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3830 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_35451_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3831 a_50520_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3832 a_10913_13118# a_9876_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3833 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3834 a_17422_13079# a_16970_12574# a_16571_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3835 a_2811_18776# a_2387_18039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3836 VSS C[6] a_48676_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3837 a_20975_6923# a_20699_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3838 a_13030_6629# a_11993_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3839 a_39855_6923# a_39579_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3840 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3841 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3842 VDD a_38677_19374# a_38627_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3843 a_11142_5835# a_10101_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3844 a_1673_519# a_1717_671# a_1242_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3845 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3846 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3847 a_15088_12575# a_14812_12575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3848 a_42888_6380# a_42718_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3849 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3850 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3851 VSS C[3] a_54340_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3852 a_44104_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3853 a_29466_1105# a_29042_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3854 a_28103_1556# a_28143_670# a_27154_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3855 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3856 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3857 a_4275_18040# a_5280_18802# a_5224_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3858 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3859 a_7536_12574# a_7260_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3860 a_43085_13118# a_41966_13079# a_43003_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3861 VSS a_30930_861# a_29987_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3862 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3863 a_20232_6924# a_20062_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3864 a_35651_518# a_35695_670# a_34706_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3865 a_26639_6923# a_26363_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3866 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3867 VDD a_52116_1105# a_52066_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3868 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3869 a_14771_13913# a_13648_14117# a_14689_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3870 a_18459_13118# a_18858_12574# a_19310_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3871 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3872 a_19535_5630# a_18811_6923# a_18688_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3873 a_13944_1405# a_14933_670# a_14893_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3874 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3875 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3876 a_47125_6923# C[55] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3877 VSS a_29042_1405# a_28103_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3878 a_32522_14117# a_31798_12574# a_31675_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3879 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3880 a_5331_13912# a_4208_14117# a_5249_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3881 a_23311_5630# a_22863_6923# a_22464_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3882 a_25690_507# a_25266_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3883 VDD a_4928_1105# a_4878_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3884 a_14660_19299# a_14720_18802# a_13715_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3885 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3886 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_20429_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3887 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3888 a_9148_12574# C[99] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3889 a_38419_6668# a_37967_6923# a_37568_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3890 VSS a_26858_14117# a_27385_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3891 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_16800_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3892 a_57757_12573# a_57587_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3893 a_13030_6629# a_13153_6923# a_13881_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3894 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3895 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3896 a_5220_19299# a_5280_18802# a_4275_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3897 VSS a_34410_14117# a_34937_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3898 a_37339_13118# a_37738_12574# a_38190_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3899 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3900 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3901 VSS a_6587_18776# a_6537_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3902 a_28210_5835# a_27087_5630# a_28128_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3903 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3904 a_27154_861# a_28159_1079# a_28099_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3905 a_18434_18261# a_19373_18040# a_19331_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3906 a_20322_18261# a_20378_18802# a_19373_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3907 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3908 a_14689_13913# a_14812_12575# a_15536_14118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3909 a_14574_6380# a_14404_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3910 a_29672_6924# a_29502_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3911 a_13030_5835# a_13153_6923# a_13877_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3912 a_11827_18040# a_12816_19167# a_12776_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3913 a_7337_518# a_7381_670# a_6392_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3914 a_14660_19299# a_14704_19167# a_13715_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3915 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3916 a_21423_5630# a_20699_6923# a_20576_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3917 a_60218_5834# a_59177_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3918 a_31650_18260# a_32589_18039# a_32547_18065# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3919 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3920 a_18459_13912# a_17418_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3921 a_59989_13119# a_60388_12575# a_60840_13080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3922 a_24352_6629# a_24751_6923# a_25203_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3923 a_36531_6668# a_35803_6923# a_35680_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3924 a_24434_5835# a_23311_5630# a_24352_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3925 a_2387_18039# a_3376_19167# a_3336_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3926 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_48743_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3927 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3928 VSS a_2387_18039# a_1448_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3929 a_50205_12573# a_50035_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3930 VDD a_21423_5630# a_21950_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3931 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3932 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3933 a_5220_19299# a_5264_19167# a_4275_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3934 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3935 a_24123_13912# a_23082_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3936 a_40307_6668# a_39855_6923# a_39456_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3937 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3938 a_37314_18261# a_38253_18040# a_38211_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3939 a_18459_13912# a_18858_12574# a_19306_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3940 a_18770_6629# a_17651_6668# a_18688_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3941 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3942 VSS a_8051_18040# a_7112_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3943 OUT a_63251_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3944 VDD C[90] a_9269_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3945 a_28979_6668# a_28527_6923# a_28128_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3946 a_55892_1105# a_55468_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3947 a_12480_1105# a_12056_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3948 VDD C[20] a_22250_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3949 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3950 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_50549_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3951 VSS a_46034_1405# a_45095_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3952 a_8217_6668# a_7489_6923# a_7366_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3953 VSS a_8704_507# a_8654_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3954 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3955 VSS C[89] a_11157_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3956 a_7341_1556# a_7397_1079# a_6392_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3957 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3958 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3959 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3960 a_7489_6923# C[34] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3961 a_40303_5630# a_39855_6923# a_39456_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3962 a_29042_1405# a_30031_670# a_29991_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3963 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3964 VDD a_53775_19374# a_53725_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3965 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3966 a_16021_18775# a_15603_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3967 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3968 a_35451_13912# a_35574_12574# a_36298_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3969 a_28128_5835# a_28527_6923# a_28975_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3970 a_3561_518# a_4504_861# a_4462_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3971 a_23573_19374# a_23149_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3972 a_14660_19299# a_15603_18584# a_15561_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3973 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3974 a_30186_12575# a_29910_12575# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3975 a_17714_1406# a_18703_670# a_18663_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3976 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3977 a_33538_18261# a_33578_19167# a_32589_18583# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3978 a_43003_13912# a_41962_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3979 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_61877_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3980 VSS a_13881_6668# a_14404_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3981 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_33792_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3982 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3983 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3984 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_44891_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3985 a_35130_507# a_34706_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X3986 a_35651_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3987 VSS a_28813_18584# a_27870_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3988 a_17418_14117# a_16694_12574# a_16571_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3989 a_37339_13912# a_37738_12574# a_38186_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3990 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3991 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3992 a_30863_5629# a_30139_6922# a_30016_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3993 a_5220_19299# a_6163_18584# a_6121_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3994 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3995 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3996 VSS a_34477_18584# a_33534_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3997 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_48890_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3998 VDD C[69] a_48905_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3999 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4000 a_28746_14117# a_28298_12574# a_27899_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4001 a_51650_1681# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4002 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4003 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4004 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4005 a_16800_6629# a_16923_6923# a_17651_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4006 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4007 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4008 VSS a_47624_13079# a_48147_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4009 a_7337_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4010 a_42453_19374# a_42029_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4011 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4012 a_34410_14117# a_33962_12574# a_33563_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4013 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4014 a_36552_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4015 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4016 VSS a_51625_5630# a_52152_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4017 a_57085_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4018 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4019 a_58973_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4020 a_36298_14117# a_35574_12574# a_35451_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4021 a_18344_6380# a_18174_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4022 a_22439_1556# a_22495_1079# a_21490_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4023 VSS a_23802_507# a_23752_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4024 a_21219_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4025 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4026 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_9254_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4027 a_16800_5835# a_16923_6923# a_17647_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4028 VSS a_36594_1405# a_35655_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4029 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4030 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_24205_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4031 VDD a_45738_14118# a_46265_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4032 a_38253_18040# a_39258_18802# a_39202_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4033 a_35762_6629# a_34643_6668# a_35680_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4034 a_6392_861# a_7381_670# a_7337_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4035 a_38482_1405# a_39471_670# a_39431_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4036 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4037 a_59668_507# a_59244_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4038 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4039 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4040 a_11764_13079# a_11312_12574# a_10913_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4041 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4042 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4043 a_8996_19299# a_9056_18802# a_8051_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4044 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_31757_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4045 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4046 a_59202_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4047 a_34435_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4048 a_52437_13118# a_52836_12574# a_53288_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4049 a_10126_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4050 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_5478_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4051 a_49804_861# a_50793_670# a_50749_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4052 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4053 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_3590_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4054 VSS a_50228_1105# a_50178_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4055 a_59964_18261# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4056 a_40099_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4057 a_45805_18584# a_46804_18801# a_46744_19298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4058 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4059 a_48317_13117# a_48147_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4060 a_41987_18860# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4061 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4062 a_29787_13913# a_29910_12575# a_30634_14118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4063 a_34706_1405# a_35695_670# a_35655_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4064 a_10168_1405# a_11173_1079# a_11117_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4065 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4066 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4067 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_43085_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4068 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4069 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4070 VDD a_55176_13079# a_55699_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4071 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4072 a_5877_6923# a_5601_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4073 a_41000_6924# a_40830_6924# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4074 a_39112_6380# a_38942_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4075 VDD a_3040_1105# a_2990_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4076 a_28099_518# a_28159_1079# a_27154_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4077 a_57127_18584# a_58132_18802# a_58072_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4078 a_12776_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4079 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4080 a_16694_12574# C[103] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4081 a_55869_12573# a_55699_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4082 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_16882_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4083 a_37568_5835# a_37691_6923# a_38415_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4084 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_14771_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4085 a_31986_5835# a_30863_5629# a_31904_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4086 VSS a_47017_671# a_47033_1080# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4087 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4088 VSS a_17651_6668# a_18174_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4089 a_33792_6629# a_33915_6923# a_34643_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4090 VSS a_10168_861# a_9225_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4091 a_52412_18261# a_53351_18040# a_53309_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4092 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4093 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4094 a_21490_861# a_22479_670# a_22435_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4095 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4096 a_1444_19298# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4097 a_31879_1557# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4098 a_3336_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4099 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4100 VSS a_8280_1405# a_7341_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4101 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4102 VDD a_27914_19167# a_27930_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4103 a_10592_507# a_10168_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4104 VSS a_12816_19167# a_12832_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4105 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4106 a_14345_13117# a_14175_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4107 a_35336_6380# a_35166_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4108 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4109 VSS a_27349_19374# a_27299_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4110 a_29910_12575# C[110] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4111 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4112 a_20576_6629# a_19539_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4113 a_57551_18776# a_57127_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4114 a_13200_12574# a_12924_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4115 a_39456_6629# a_38419_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4116 VSS C[63] a_60233_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4117 a_27349_19374# a_26925_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4118 a_35574_12574# C[113] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4119 a_29991_1556# a_30031_670# a_29042_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4120 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4121 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4122 a_6793_13117# a_6623_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4123 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4124 a_29758_19299# a_30701_18584# a_30659_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4125 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4126 VSS a_59668_1105# a_59618_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4127 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_59989_13119# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4128 a_35680_5835# a_36079_6923# a_36527_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4129 VSS a_4504_1405# a_3565_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4130 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4131 a_22206_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4132 a_52437_13912# a_52836_12574# a_53284_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4133 a_12014_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4134 a_11117_1556# a_12056_1405# a_12014_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4135 a_24094_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4136 a_31904_6629# a_32303_6923# a_32755_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4137 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4138 a_6392_1405# a_7381_670# a_7341_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4139 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4140 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_37650_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4141 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4142 a_8910_6924# a_8740_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4143 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_9336_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4144 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4145 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_58330_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4146 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_56442_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4147 a_33242_1105# a_32818_1406# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4148 a_21685_19374# a_21261_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4149 a_49741_6668# a_49289_6923# a_48890_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4150 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4151 VSS C[17] a_27914_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4152 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4153 a_31904_5835# a_32303_6923# a_32751_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4154 a_54004_1105# a_53580_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4155 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4156 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4157 a_3672_5835# a_1013_18584# a_3590_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4158 a_22439_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4159 a_7137_13118# a_7260_12574# a_7988_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4160 a_5478_6629# a_5601_6923# a_6329_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4161 VDD a_38415_5630# a_38942_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4162 VDD C[82] a_24367_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4163 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4164 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4165 a_42974_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4166 a_51396_14117# a_50672_12574# a_50549_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4167 a_49060_12574# a_48784_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4168 a_52322_6924# a_52152_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4169 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_33874_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4170 a_45091_518# a_45151_1079# a_44146_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4171 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4172 a_41344_6629# a_40307_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4173 VDD a_37018_507# a_36968_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4174 a_33013_19374# a_32589_18583# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4175 VSS a_34643_6668# a_35166_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4176 a_58729_6923# a_58453_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4177 VSS C[81] a_26255_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4178 a_54529_1556# a_54569_670# a_53580_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4179 VDD a_60836_14118# a_61363_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4180 a_25896_6380# a_25726_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4181 a_60903_18040# a_62276_12574# a_61877_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4182 a_30867_6667# a_30139_6922# a_30016_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4183 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4184 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4185 a_56612_12574# a_56336_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4186 a_5478_5835# a_5601_6923# a_6325_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4187 a_40565_19374# a_40141_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4188 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4189 a_14918_5834# a_13877_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4190 VDD a_38906_507# a_38856_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4191 a_12686_6380# a_12516_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4192 a_9254_5835# a_8213_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4193 a_29042_861# a_30047_1079# a_29987_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4194 a_47853_6668# a_47125_6923# a_47002_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4195 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4196 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4197 a_6100_13079# a_5648_12574# a_5249_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4198 VSS a_23149_18040# a_22210_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4199 a_7988_13079# a_7536_12574# a_7137_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4200 a_50753_1556# a_50809_1079# a_49804_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4201 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4202 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4203 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4204 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4205 a_29443_12573# a_29273_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4206 a_47849_5630# a_47125_6923# a_47002_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4207 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4208 VDD a_58952_13079# a_59475_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4209 a_23802_1105# a_23378_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4210 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4211 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4212 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4213 VSS a_57356_1405# a_56417_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4214 a_35107_12573# a_34937_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4215 a_36995_12573# a_36825_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4216 a_58224_12574# C[125] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4217 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4218 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4219 a_2387_18583# a_3392_18802# a_3332_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4220 a_3590_5835# a_3989_6923# a_4437_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4221 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4222 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4223 VSS a_19797_19374# a_19747_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4224 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4225 a_7341_1556# a_7381_670# a_6392_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4226 a_56188_18261# a_57127_18040# a_57085_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4227 VSS a_42029_18040# a_41090_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4228 VSS a_22250_19167# a_22266_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4229 VSS a_43917_18040# a_42978_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4230 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_5560_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4231 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4232 a_9000_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4233 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4234 VSS a_25203_6668# a_25726_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4235 a_39431_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4236 a_56524_5835# a_55401_5630# a_56442_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4237 a_2811_18776# a_2387_18039# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4238 a_45805_18040# a_46788_19166# a_46748_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4239 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4240 a_58330_6629# a_58453_6923# a_59181_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4241 a_28103_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4242 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4243 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4244 VDD a_53513_5630# a_54040_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4245 a_30930_1405# a_31935_1080# a_31879_1557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4246 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4247 VDD a_6325_5630# a_6852_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4248 a_42888_6380# a_42718_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4249 a_52116_507# a_51692_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4250 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4251 a_54325_13912# a_54448_12574# a_55172_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4252 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4253 a_10888_18261# a_10944_18802# a_9939_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4254 a_12776_18261# a_12832_18802# a_11827_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4255 a_50672_12574# C[121] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4256 VDD a_32755_6668# a_33278_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4257 a_57986_6924# a_57816_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4258 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_45202_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4259 VSS a_38677_19374# a_38627_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4260 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4261 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4262 VDD a_56228_19167# a_56244_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4263 a_56213_13912# a_56612_12574# a_57060_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4264 a_51625_5630# a_51177_6923# a_50778_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4265 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4266 VSS a_41130_19167# a_41146_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4267 a_27870_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4268 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_22235_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4269 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4270 a_48861_518# a_48921_1079# a_47916_1406# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4271 a_9424_12574# a_9148_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4272 a_58330_5835# a_58453_6923# a_59177_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4273 VDD C[68] a_50793_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4274 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4275 a_52748_5835# a_51625_5630# a_52666_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4276 a_3336_18261# a_3392_18802# a_2387_18583# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4277 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_10913_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4278 a_30638_13080# a_29910_12575# a_29787_13913# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4279 VDD a_49737_5630# a_50264_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4280 VDD a_25461_19374# a_25411_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4281 a_48111_18776# a_47687_18039# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4282 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4283 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_39309_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4284 a_47620_14117# a_47172_12574# a_46773_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4285 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_12801_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4286 a_61762_6379# a_61592_6379# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4287 a_60218_5834# a_60617_6922# a_61065_5629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4288 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4289 VDD a_12480_507# a_12430_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4290 VDD a_31125_19373# a_31075_19154# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4291 a_45805_18040# a_46804_18801# a_46748_18260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4292 VDD a_11157_670# a_11173_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4293 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4294 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4295 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4296 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_3361_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4297 a_10105_6668# a_9653_6923# a_9254_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4298 a_40794_1105# a_40370_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4299 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4300 a_9939_18584# a_10928_19167# a_10884_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4301 a_55663_18776# a_55239_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4302 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4303 a_6392_861# a_7397_1079# a_7337_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4304 a_10888_18261# a_10928_19167# a_9939_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4305 a_12776_18261# a_12816_19167# a_11827_18584# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4306 a_17443_18065# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4307 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_41115_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4308 VSS a_13045_670# a_13061_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4309 a_25690_507# a_25266_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4310 a_1013_19128# a_1488_19166# a_1444_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4311 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4312 a_2574_1682# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4313 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4314 a_57127_18040# a_58132_18802# a_58076_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4315 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4316 a_1872_12574# a_1596_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4317 a_56442_5835# a_56841_6923# a_57289_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4318 VDD a_44341_19374# a_44291_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4319 a_10101_5630# a_9653_6923# a_9254_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4320 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4321 VDD C[29] a_5264_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4322 a_61090_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4323 a_31879_1557# a_32818_1406# a_32776_1682# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4324 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4325 VDD a_11760_14117# a_12287_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4326 VDD a_23315_6668# a_23838_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4327 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_58412_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4328 VDD a_33807_670# a_33823_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4329 a_10126_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4330 a_3561_518# a_3621_1079# a_2616_1406# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4331 a_36323_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4332 a_11036_12574# C[100] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4333 VSS a_35695_670# a_35711_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4334 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4335 VDD a_4208_14117# a_4735_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4336 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4337 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4338 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4339 a_37224_6380# a_37054_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4340 VDD a_59177_5630# a_59704_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4341 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4342 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4343 a_58183_13912# a_57060_14117# a_58101_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4344 VSS a_2616_862# a_1673_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4345 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4346 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4347 a_3484_12574# C[96] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4348 a_24123_13118# a_24522_12574# a_24974_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4349 VDD a_42682_1105# a_42632_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4350 a_21490_861# a_22495_1079# a_22435_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4351 VSS a_21194_14117# a_21721_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4352 VDD a_923_18775# a_873_18610# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4353 a_50205_12573# a_50035_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4354 VSS a_21423_5630# a_21950_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4355 VSS a_1152_1106# a_1102_887# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4356 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4357 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4358 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4359 a_11142_6629# a_11541_6923# a_11993_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4360 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4361 a_13673_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4362 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4363 a_31675_13118# a_32074_12574# a_32526_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4364 VSS a_26026_19167# a_26042_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4365 a_33448_6380# a_33278_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4366 VSS a_32522_14117# a_33049_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4367 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4368 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4369 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4370 a_22439_1556# a_23378_1405# a_23336_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4371 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4372 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4373 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_7219_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4374 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4375 a_27555_12573# a_27385_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4376 a_23086_13079# a_22358_12574# a_22235_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4377 a_16571_13118# a_16694_12574# a_17422_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4378 VSS a_40074_14117# a_40601_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4379 a_16021_18775# a_15603_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4380 VSS a_47687_18583# a_46744_19298# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4381 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4382 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4383 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4384 a_24974_13079# a_24246_12574# a_24123_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4385 a_32074_12574# a_31798_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4386 a_33962_12574# a_33686_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4387 a_54448_12574# C[123] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4388 VDD a_46223_18775# a_46173_18610# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4389 a_33219_12573# a_33049_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4390 a_20699_6923# C[41] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4391 a_8238_1681# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4392 VSS a_53775_19374# a_53725_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4393 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4394 a_22235_13118# a_22358_12574# a_23086_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4395 a_39579_6923# C[51] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4396 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4397 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4398 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_26011_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4399 a_16653_13118# a_15540_13080# a_16571_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4400 a_46435_13118# a_46265_13118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4401 VDD a_40307_6668# a_40830_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4402 a_7112_18261# a_7168_18802# a_6163_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4403 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4404 a_8280_1405# a_9285_1079# a_9229_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4405 a_56413_518# a_56473_1079# a_55468_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4406 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4407 VDD a_29237_19374# a_29187_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4408 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_33563_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4409 a_22317_13118# a_21198_13079# a_22235_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4410 a_32303_6923# a_32027_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4411 a_45290_12575# a_45014_12575# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4412 a_13944_861# a_14933_670# a_14889_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4413 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4414 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4415 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4416 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4417 VDD a_59439_18776# a_59389_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4418 a_43854_13079# a_43126_12574# a_43003_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4419 a_60193_1556# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4420 VSS a_46788_19166# a_46804_18801# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4421 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4422 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4423 a_13881_6668# a_13153_6923# a_13030_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4424 a_59439_18776# a_59015_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4425 a_14689_13119# a_13652_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4426 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4427 a_41115_13118# a_41238_12574# a_41966_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4428 a_24008_6380# a_23838_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4429 a_35533_13118# a_34414_13079# a_35451_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4430 a_43003_13118# a_43126_12574# a_43854_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4431 a_47645_18859# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4432 a_5134_6380# a_4964_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4433 VSS a_21261_18584# a_20318_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4434 a_5249_13118# a_4212_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4435 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4436 a_41315_518# a_42258_861# a_42216_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4437 a_2387_18039# a_3392_18802# a_3336_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4438 a_5648_12574# a_5372_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4439 a_41197_13118# a_40078_13079# a_41115_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4440 NBR128half_0/sky130_fd_sc_hd__inv_16_4/A sky130_fd_sc_hd__inv_8_0/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4441 a_13877_5630# a_13153_6923# a_13030_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4442 a_21194_14117# a_20746_12574# a_20347_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4443 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4444 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4445 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4446 a_60218_6628# a_60617_6922# a_61069_6667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4447 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4448 a_3040_507# a_2616_862# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4449 a_23082_14117# a_22358_12574# a_22235_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4450 a_50778_5835# a_49737_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4451 a_24970_14117# a_24246_12574# a_24123_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4452 a_16571_13118# a_16970_12574# a_17422_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4453 VSS a_40141_18584# a_39198_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4454 a_51421_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4455 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4456 a_13001_518# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4457 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4458 a_21914_1105# a_21490_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4459 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4460 a_3443_13912# a_2320_14117# a_3361_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4461 VSS RESET a_28116_9428# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4462 VDD a_27578_507# a_27528_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4463 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4464 a_12251_19374# a_11827_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4465 a_10884_19299# a_10944_18802# a_9939_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4466 a_12772_19299# a_12832_18802# a_11827_18040# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4467 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_28128_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4468 a_40074_14117# a_39626_12574# a_39227_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4469 VSS a_55176_13079# a_55699_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4470 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4471 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_26240_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4472 VDD a_26255_670# a_26271_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4473 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4474 VSS a_24970_14117# a_25497_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4475 a_19539_6668# a_19087_6923# a_18688_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4476 VSS C[67] a_52681_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4477 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4478 a_22439_1556# a_22479_670# a_21490_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4479 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4480 VDD a_19310_13079# a_19833_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4481 a_55869_12573# a_55699_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4482 VDD a_45971_6667# a_46494_6923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4483 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4484 a_18858_12574# a_18582_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4485 a_3332_19299# a_3392_18802# a_2387_18039# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4486 a_43850_14117# a_43126_12574# a_43003_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4487 VSS a_28143_670# a_28159_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4488 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4489 a_35451_13118# a_35850_12574# a_36302_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4490 a_22120_6924# a_21950_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4491 a_14889_518# a_14949_1079# a_13944_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4492 a_11142_6629# a_10105_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4493 a_28527_6923# a_28251_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4494 a_37967_6923# a_37691_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4495 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4496 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4497 a_9897_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4498 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4499 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4500 VSS a_43850_14117# a_44377_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4501 VDD a_48905_670# a_48921_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4502 a_25224_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4503 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4504 a_14918_5834# a_15317_6922# a_15765_5629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4505 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4506 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4507 VDD a_38190_13079# a_38713_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4508 a_16571_13912# a_15536_14118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4509 a_37738_12574# a_37462_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4510 a_17651_6668# a_16923_6923# a_16800_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4511 a_15832_861# a_16815_671# a_16771_519# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4512 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4513 VSS a_15603_18040# a_14664_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4514 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_46855_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4515 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4516 a_35426_18261# a_36365_18040# a_36323_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4517 a_22235_13912# a_21194_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4518 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4519 a_16571_13912# a_16970_12574# a_17418_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4520 a_61533_13118# a_61363_13118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4521 VSS a_6163_18040# a_5224_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4522 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4523 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4524 a_17647_5630# a_16923_6923# a_16800_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4525 VDD a_57780_1105# a_57730_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4526 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4527 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_58183_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4528 VDD a_4699_18776# a_4649_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4529 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4530 VSS a_27154_1405# a_26215_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4531 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4532 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4533 a_35451_13912# a_34410_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4534 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4535 a_29991_1556# a_30930_1405# a_30888_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4536 VDD a_51887_19374# a_51837_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4537 a_33563_13912# a_33686_12574# a_34410_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4538 VSS a_38415_5630# a_38942_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4539 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_43232_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4540 a_21685_19374# a_21261_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4541 a_36531_6668# a_36079_6923# a_35680_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4542 a_12772_19299# a_13715_18584# a_13673_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4543 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4544 VDD a_33578_19167# a_33594_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4545 a_41115_13912# a_40074_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4546 a_50631_13118# a_49512_13079# a_50549_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4547 a_9653_6923# a_9377_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4548 VSS a_37018_507# a_36968_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4549 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4550 VSS a_25037_18584# a_24094_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4551 VSS a_26925_18584# a_25982_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4552 a_35451_13912# a_35850_12574# a_36298_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4553 a_9229_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4554 a_3332_19299# a_4275_18584# a_4233_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4555 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4556 a_26322_5835# a_25199_5630# a_26240_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4557 a_28128_6629# a_28251_6923# a_28979_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4558 a_33013_19374# a_32589_18583# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4559 a_26858_14117# a_26410_12574# a_26011_13118# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4560 a_37691_6923# C[50] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4561 a_12686_6380# a_12516_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4562 a_37543_1556# a_37599_1079# a_36594_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4563 VSS a_38906_507# a_38856_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4564 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4565 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4566 a_49533_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4567 a_27784_6924# a_27614_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4568 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_15000_6628# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4569 a_31879_1557# a_31919_671# a_30930_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4570 a_28746_14117# a_28022_12574# a_27899_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4571 a_53065_6923# a_52789_6923# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4572 a_60218_6628# a_59181_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4573 a_5449_518# a_5493_670# a_4504_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4574 a_40565_19374# a_40141_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4575 a_38415_5630# a_37691_6923# a_37568_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4576 VDD a_1152_508# a_1102_343# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4577 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4578 a_34901_18776# a_34477_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4579 a_33763_518# a_34706_861# a_34664_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4580 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4581 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4582 a_28128_5835# a_28251_6923# a_28975_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4583 a_12056_861# a_13045_670# a_13001_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4584 VSS a_45805_18584# a_44862_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4585 a_55197_18066# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4586 a_34643_6668# a_33915_6923# a_33792_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4587 a_22546_5835# a_21423_5630# a_22464_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4588 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4589 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4590 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4591 VDD a_19535_5630# a_20062_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4592 a_31560_6379# a_31390_6379# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4593 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_22317_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4594 VSS a_58952_13079# a_59475_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4595 a_30863_5629# a_30415_6922# a_30016_6628# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4596 a_36365_18040# a_37370_18802# a_37314_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4597 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4598 a_39626_12574# a_39350_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4599 a_16882_6629# a_15769_6667# a_16800_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4600 a_34639_5630# a_33915_6923# a_33792_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4601 VDD C[87] a_14933_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4602 a_10592_1105# a_10168_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4603 a_8475_19374# a_8051_18584# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4604 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_29869_13119# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4605 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4606 a_8217_6668# a_7765_6923# a_7366_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4607 a_6329_6668# a_5601_6923# a_5478_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4608 VSS a_44146_1405# a_43207_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4609 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4610 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4611 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4612 a_50549_13118# a_50948_12574# a_51400_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4613 a_56413_518# a_57356_861# a_57314_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4614 a_45519_6922# a_45243_6922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4615 a_26240_5835# a_26639_6923# a_27087_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4616 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_41197_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4617 VSS a_11993_6668# a_12516_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4618 a_46034_861# a_47033_1080# a_46973_519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4619 a_33763_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4620 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4621 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4622 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4623 a_37421_13912# a_36298_14117# a_37339_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4624 VSS a_53513_5630# a_54040_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4625 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_28210_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4626 VDD a_53288_13079# a_53811_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4627 VSS a_6325_5630# a_6852_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4628 a_52116_507# a_51692_861# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4629 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4630 a_52836_12574# a_52560_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4631 sky130_fd_sc_hd__buf_2_0/X a_28116_9428# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4632 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_48890_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4633 a_43314_5835# a_42191_5630# a_43232_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4634 a_16775_1557# a_16831_1080# a_15832_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4635 a_14893_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4636 a_10888_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4637 VSS a_30701_18040# a_29762_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4638 a_18459_13912# a_18582_12574# a_19306_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4639 a_59645_13117# a_59475_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4640 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_47002_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4641 a_55239_18584# a_56244_18802# a_56184_19299# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4642 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4643 VDD a_18474_19167# a_18490_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4644 VSS NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_46773_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4645 a_44776_6924# a_44606_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4646 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4647 a_50524_18261# a_51463_18040# a_51421_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4648 VDD a_28975_5630# a_29502_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4649 a_1448_18260# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4650 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4651 a_49804_1405# a_50809_1079# a_50753_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4652 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4653 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4654 VSS a_49737_5630# a_50264_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4655 a_45095_1556# a_45135_670# a_44146_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4656 VSS a_53580_861# a_52637_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4657 a_48111_18776# a_47687_18039# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4658 a_14689_13119# a_15088_12575# a_15540_13080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4659 VSS a_12480_507# a_12430_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4660 a_53538_887# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4661 a_58301_518# a_58345_670# a_57356_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4662 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4663 a_12457_13117# a_12287_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4664 a_26134_12574# C[108] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4665 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4666 a_49289_6923# a_49013_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4667 VSS C[93] a_3605_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4668 VSS a_25461_19374# a_25411_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4669 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4670 a_50549_13912# a_49508_14117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4671 a_55663_18776# a_55239_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4672 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y a_18770_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4673 VSS a_4928_1105# a_4878_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4674 a_37339_13912# a_37462_12574# a_38186_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4675 a_11312_12574# a_11036_12574# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4676 a_14918_6628# a_15317_6922# a_15769_6667# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4677 VDD a_33242_1105# a_33192_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4678 VSS a_31125_19373# a_31075_19154# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4679 a_19797_18776# a_19373_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4680 a_33686_12574# C[112] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4681 a_33874_6629# a_32755_6668# a_33792_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4682 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4683 a_4905_13117# a_4735_13117# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4684 VDD a_39242_19167# a_39258_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4685 a_20318_19299# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4686 a_50549_13912# a_50948_12574# a_51396_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4687 VSS a_9040_19167# a_9056_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4688 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4689 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4690 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4691 a_8996_19299# a_9939_18584# a_9897_18860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4692 a_61959_13118# a_60840_13080# a_61877_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4693 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_3590_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4694 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4695 VSS C[22] a_18474_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4696 VDD a_44906_19167# a_44922_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4697 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4698 a_42682_507# a_42258_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4699 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4700 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4701 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4702 VSS a_44341_19374# a_44291_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4703 a_43232_5835# a_43631_6923# a_44079_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4704 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4705 a_32818_1406# a_33807_670# a_33767_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4706 a_6100_13079# a_5372_12574# a_5249_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4707 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4708 VSS C[18] a_26026_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4709 VSS a_47916_1406# a_46977_1557# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4710 a_38677_18776# a_38253_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4711 NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4712 VDD a_10105_6668# a_10628_6924# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4713 VDD C[86] a_16815_671# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4714 VDD C[7] a_46788_19166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4715 VSS C[15] a_31690_19166# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4716 a_39198_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4717 a_5249_13118# a_5372_12574# a_6100_13079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4718 a_47687_18583# a_48676_19167# a_48632_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4719 a_41086_19299# NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4720 VSS a_60903_18584# a_59960_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4721 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_9025_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4722 a_47172_12574# a_46896_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4723 a_3989_6923# a_3713_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4724 a_37224_6380# a_37054_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4725 a_13005_1556# a_13061_1079# a_12056_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4726 a_26211_518# a_26271_1079# a_25266_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4727 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4728 VSS a_59177_5630# a_59704_6380# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4729 a_30098_5834# a_28975_5630# a_30016_5834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4730 a_44146_861# a_45151_1079# a_45091_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4731 VSS C[12] a_37354_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4732 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4733 a_31904_6629# a_32027_6923# a_32755_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4734 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_39538_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4735 a_51463_18040# a_52468_18802# a_52412_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4736 VSS a_923_18775# a_873_18610# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4737 a_54724_12574# a_54448_12574# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4738 sky130_fd_sc_hd__inv_8_0/Y sky130_fd_sc_hd__buf_2_0/X VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4739 VSS a_30031_670# a_30047_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4740 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4741 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4742 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4743 NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4744 a_13652_13079# a_13200_12574# a_12801_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4745 a_59181_6668# a_58453_6923# a_58330_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4746 a_47084_5835# a_45967_5629# a_47002_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4747 VSS a_6392_1405# a_5453_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4748 VSS C[8] a_44906_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4749 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4750 a_5560_6629# a_4441_6668# a_5478_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4751 a_58453_6923# C[61] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4752 a_18663_1556# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4753 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4754 a_33448_6380# a_33278_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4755 a_8280_1405# a_9269_670# a_9229_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4756 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4757 a_4212_13079# a_3760_12574# a_3361_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4758 a_48546_6924# a_48376_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4759 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y a_35762_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4760 a_59177_5630# a_58453_6923# a_58330_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4761 VDD a_50793_670# a_50809_1079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4762 a_27555_12573# a_27385_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4763 VSS a_57780_1105# a_57730_886# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4764 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4765 a_46977_1557# a_47017_671# a_46034_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4766 a_9229_1556# a_10168_1405# a_10126_1681# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4767 VDD a_57064_13079# a_57587_12573# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4768 VSS a_52681_670# a_52697_1079# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4769 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4770 a_4504_1405# a_5493_670# a_5453_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4771 a_33219_12573# a_33049_12573# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4772 a_48861_518# a_49804_861# a_49762_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4773 VSS a_46223_18775# a_46173_18610# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4774 a_14664_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4775 a_27154_861# a_28143_670# a_28099_518# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4776 a_7022_6924# a_6852_6924# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4777 a_46664_6379# a_46494_6379# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4778 VSS NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_56442_6629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4779 a_58301_518# NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4780 a_54300_18261# a_55239_18040# a_55197_18066# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4781 a_47853_6668# a_47401_6923# a_47002_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4782 VSS a_20362_19167# a_20378_18802# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4783 a_5224_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4784 a_7366_5835# a_7489_6923# a_8213_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4785 a_7112_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4786 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4787 a_29787_13119# a_30186_12575# a_30638_13080# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4788 a_3590_6629# a_3713_6923# a_4441_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4789 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4790 VSS a_59439_18776# a_59389_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4791 a_46773_13912# a_46896_12574# a_47620_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4792 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4793 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_18541_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4794 VDD a_15769_6667# a_16292_6923# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4795 a_43203_518# a_43263_1079# a_42258_1405# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4796 a_1677_1557# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4797 VSS a_29237_19374# a_29187_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4798 a_21891_12573# a_21721_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4799 VDD a_18138_507# a_18088_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4800 a_59439_18776# a_59015_18040# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4801 VSS a_7984_14117# a_8511_13117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4802 a_49013_6923# C[56] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4803 NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4804 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4805 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4806 a_46744_19298# a_46788_19166# a_45805_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4807 a_24008_6380# a_23838_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4808 VDD a_54004_507# a_53954_342# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4809 a_52437_13912# a_52560_12574# a_53284_14117# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4810 a_5134_6380# a_4964_6380# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4811 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_48972_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4812 a_7337_518# a_8280_861# a_8238_887# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4813 VSS NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4814 a_14918_6628# a_13881_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4815 a_3590_5835# a_3713_6923# a_4437_5630# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4816 VDD a_52452_19167# a_52468_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4817 VDD a_54340_19167# a_54356_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4818 a_61877_13912# a_60836_14118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4819 a_37543_1556# a_37583_670# a_36594_861# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4820 VDD a_17909_19374# a_17859_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4821 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4822 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4823 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_20347_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4824 a_54325_13912# a_54724_12574# a_55172_14117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4825 a_10798_6380# a_10628_6380# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4826 a_9254_6629# a_8217_6668# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4827 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4828 a_7366_5835# a_6325_5630# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4829 a_1448_18260# a_1504_18801# a_1013_19128# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4830 a_55239_18040# a_56228_19167# a_56188_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4831 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4832 VDD a_60004_19167# a_60020_18802# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4833 a_58072_19299# a_58116_19167# a_57127_18040# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4834 a_58412_6629# a_57293_6668# a_58330_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4835 a_5478_5835# a_5877_6923# a_6325_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4836 VDD a_23573_19374# a_23523_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4837 NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4838 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y a_37421_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4839 a_40771_12573# a_40601_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4840 a_60112_12575# C[126] VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4841 a_3040_507# a_2616_862# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4842 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4843 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4844 VSS a_45971_6667# a_46494_6923# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4845 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_7448_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4846 a_31875_519# a_31919_671# a_30930_1405# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4847 NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4848 a_53775_18776# a_53351_18040# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4849 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4850 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4851 a_56841_6923# a_56565_6923# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4852 VSS a_55468_1405# a_54529_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4853 VDD a_28116_9428# sky130_fd_sc_hd__buf_2_0/X VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4854 a_3040_1105# a_2616_1406# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4855 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4856 VSS a_27578_507# a_27528_342# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4857 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4858 NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4859 a_54636_6629# a_53517_6668# a_54554_6629# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4860 a_57356_1405# a_58345_670# a_58305_1556# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4861 a_58101_13118# a_57064_13079# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4862 a_1448_18260# a_1488_19166# a_1013_19128# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4863 NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4864 VDD a_8213_5630# a_8740_6380# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4865 a_4462_887# NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4866 VDD a_42453_19374# a_42403_19155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4867 VSS C[4] a_52452_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4868 a_55239_18040# a_56244_18802# a_56188_18261# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4869 a_9107_13118# a_7988_13079# a_9025_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4870 VDD C[30] a_3376_19167# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4871 a_12251_19374# a_11827_18584# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4872 VSS a_19310_13079# a_19833_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4873 VDD NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_3672_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4874 a_60218_5834# a_60341_6922# a_61065_5629# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4875 VDD a_48340_1105# a_48290_886# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4876 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4877 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y a_13030_5835# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4878 VSS a_4441_6668# a_4964_6924# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4879 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4880 VSS C[0] a_60004_19167# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4881 a_28771_18066# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4882 a_56442_6629# a_56565_6923# a_57293_6668# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4883 a_36594_861# a_37599_1079# a_37539_518# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4884 a_29042_1405# a_30047_1079# a_29991_1556# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4885 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4886 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4887 VDD a_15536_14118# a_16063_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4888 VSS a_8051_18584# a_7108_19299# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4889 a_57780_507# a_57356_861# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4890 VDD a_2320_14117# a_2847_13117# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4891 a_46034_1405# a_47033_1080# a_46977_1557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4892 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4893 a_56295_13912# a_55172_14117# a_56213_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4894 VSS a_38190_13079# a_38713_12573# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4895 a_1596_12574# C[95] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4896 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4897 a_22235_13118# a_22634_12574# a_23086_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4898 a_29762_18261# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4899 a_12480_1105# a_12056_1405# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4900 a_15603_18584# a_16602_18801# a_16542_19298# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4901 a_18115_13117# a_17945_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4902 a_28103_1556# a_28159_1079# a_27154_861# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4903 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4904 NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4905 a_11785_18860# NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4906 NBR128half_0/nbrhalf_3/sky130_fd_sc_hd__inv_16_3/Y NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4907 a_20003_13117# a_19833_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4908 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4909 a_54554_6629# a_54953_6923# a_55405_6668# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4910 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4911 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4912 VSS a_4699_18776# a_4649_18611# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4913 a_31646_19298# a_32589_18583# a_32547_18859# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4914 VDD NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y a_5331_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4915 a_25667_12573# a_25497_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4916 a_21198_13079# a_20470_12574# a_20347_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4917 a_41115_13118# a_41514_12574# a_41966_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4918 a_43003_13118# a_43402_12574# a_43854_13079# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4919 NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4920 a_47687_18039# a_48676_19167# a_48636_18261# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4921 VSS a_47687_18039# a_46748_18260# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4922 a_54554_5835# a_54953_6923# a_55401_5630# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4923 a_14664_18261# a_14720_18802# a_13715_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4924 NBR128half_0/sky130_fd_sc_hd__inv_16_4/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4925 VSS a_51887_19374# a_51837_19155# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4926 a_38883_13117# a_38713_13117# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4927 VDD sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__inv_8_0/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4928 VDD sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4929 VDD NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_1/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4930 VSS NBR128half_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y a_24123_13912# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4931 a_15317_6922# a_15041_6922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4932 a_1242_861# a_1733_1080# a_1677_1557# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4933 VDD NBR128half_bottom_0/nbrhalf_2/sky130_fd_sc_hd__inv_16_3/Y a_56524_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4934 VDD C[73] a_41359_670# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4935 a_3332_19299# a_3376_19167# a_2387_18039# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4936 VSS NBR128half_0/sky130_fd_sc_hd__inv_16_4/A NBR128half_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4937 VSS sky130_fd_sc_hd__inv_8_0/Y NBR128half_0/sky130_fd_sc_hd__inv_16_4/A VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4938 a_5224_18261# a_5280_18802# a_4275_18584# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4939 a_20429_13118# a_19310_13079# a_20347_13118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4940 a_52116_1105# a_51692_1405# VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X4941 VDD NBR128half_0/nbrhalf_1/sky130_fd_sc_hd__inv_16_3/Y a_52519_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4942 a_44547_12573# a_44377_12573# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4943 VSS C[72] a_43247_670# VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4944 VSS NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_3/A NBR128half_bottom_0/nbrhalf_128_0/sky130_fd_sc_hd__inv_16_1/Y VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4945 a_40078_13079# a_39350_12574# a_39227_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4946 a_13112_5835# a_11989_5630# a_13030_5835# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4947 VDD NBR128half_bottom_0/sky130_fd_sc_hd__inv_16_1/Y NBR128half_bottom_0/nbrhalf_0/sky130_fd_sc_hd__inv_16_3/Y VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4948 VDD a_57551_18776# a_57501_18611# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X4949 a_41966_13079# a_41238_12574# a_41115_13912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

