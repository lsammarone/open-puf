magic
tech sky130A
magscale 1 2
timestamp 1654402208
<< metal3 >>
rect 24564 17620 51004 17720
rect 24556 11447 51008 11730
rect 24556 11383 31005 11447
rect 31069 11383 31085 11447
rect 31149 11383 51008 11447
rect 24556 11172 51008 11383
rect 24556 11170 51002 11172
rect 24554 5376 51000 5380
rect 24554 4820 51012 5376
rect 50894 4818 51012 4820
rect 24546 -1480 51004 -920
rect 41002 -7514 41126 -7512
rect 27598 -7532 47866 -7514
rect 27598 -7534 41032 -7532
rect 27598 -7598 27628 -7534
rect 27692 -7598 34332 -7534
rect 34396 -7596 41032 -7534
rect 41096 -7534 47866 -7532
rect 41096 -7596 47772 -7534
rect 34396 -7598 47772 -7596
rect 47836 -7598 47866 -7534
rect 27598 -7618 47866 -7598
<< via3 >>
rect 31005 11383 31069 11447
rect 31085 11383 31149 11447
rect 27628 -7598 27692 -7534
rect 34332 -7598 34396 -7534
rect 41032 -7596 41096 -7532
rect 47772 -7598 47836 -7534
<< metal4 >>
rect 26628 -7516 26782 17949
rect 31002 11485 31156 17871
rect 31001 11447 31156 11485
rect 31001 11383 31005 11447
rect 31069 11383 31085 11447
rect 31149 11383 31156 11447
rect 31001 11345 31156 11383
rect 27608 -7513 27712 -7380
rect 26628 -7735 26778 -7516
rect 27607 -7534 27713 -7513
rect 27607 -7598 27628 -7534
rect 27692 -7598 27713 -7534
rect 27607 -7619 27713 -7598
rect 31002 -7741 31156 11345
rect 34312 -7513 34416 -7378
rect 41012 -7511 41116 -7362
rect 34311 -7534 34417 -7513
rect 34311 -7598 34332 -7534
rect 34396 -7598 34417 -7534
rect 34311 -7619 34417 -7598
rect 41011 -7532 41117 -7511
rect 47752 -7513 47856 -7360
rect 41011 -7596 41032 -7532
rect 41096 -7596 41117 -7532
rect 41011 -7617 41117 -7596
rect 47751 -7534 47857 -7513
rect 47751 -7598 47772 -7534
rect 47836 -7598 47857 -7534
rect 47751 -7619 47857 -7598
use sky130_fd_pr__cap_mim_m3_1_5F9S4M  sky130_fd_pr__cap_mim_m3_1_5F9S4M_0
timestamp 1654402208
transform 1 0 27710 0 1 5116
box -3150 -12600 3149 12600
use sky130_fd_pr__cap_mim_m3_1_5F9S4M  sky130_fd_pr__cap_mim_m3_1_5F9S4M_1
timestamp 1654402208
transform 1 0 34414 0 1 5118
box -3150 -12600 3149 12600
use sky130_fd_pr__cap_mim_m3_1_5F9S4M  sky130_fd_pr__cap_mim_m3_1_5F9S4M_2
timestamp 1654402208
transform 1 0 41114 0 1 5134
box -3150 -12600 3149 12600
use sky130_fd_pr__cap_mim_m3_1_5F9S4M  sky130_fd_pr__cap_mim_m3_1_5F9S4M_3
timestamp 1654402208
transform 1 0 47854 0 1 5136
box -3150 -12600 3149 12600
<< labels >>
flabel metal4 s 31016 -7548 31140 -7286 1 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal4 s 26634 -7542 26758 -7280 1 FreeSans 2000 0 0 0 VDD
port 2 nsew
<< end >>
