VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO decap
  CLASS BLOCK ;
  FOREIGN decap ;
  ORIGIN -122.730 38.705 ;
  SIZE 132.330 BY 128.450 ;
  PIN VSS
    PORT
      LAYER met4 ;
        RECT 155.010 -38.705 155.780 56.915 ;
    END
  END VSS
  PIN VDD
    PORT
      LAYER met4 ;
        RECT 133.170 -37.710 133.790 -36.400 ;
    END
  END VDD
  OBS
      LAYER met3 ;
        RECT 122.730 -38.090 255.060 88.600 ;
      LAYER met4 ;
        RECT 123.495 57.315 254.995 89.745 ;
        RECT 123.495 -36.000 154.610 57.315 ;
        RECT 123.495 -38.110 132.770 -36.000 ;
        RECT 134.190 -38.110 154.610 -36.000 ;
        RECT 123.495 -38.675 154.610 -38.110 ;
        RECT 156.180 -38.675 254.995 57.315 ;
  END
END decap
END LIBRARY

