magic
tech sky130B
timestamp 1648127584
<< properties >>
string GDS_END 27743366
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27742082
<< end >>
