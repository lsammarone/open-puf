magic
tech sky130A
timestamp 1648127584
<< properties >>
string GDS_END 31254382
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31252138
<< end >>
