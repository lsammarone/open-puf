/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__res_high_po_5p73.model.spice