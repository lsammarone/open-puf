magic
tech sky130A
magscale 1 2
timestamp 1654658503
<< nwell >>
rect 31643 4383 32021 5502
rect 31376 4354 32021 4383
rect 31376 4062 31912 4354
rect 15656 3686 16038 4007
rect 45798 3846 46180 4167
<< nsubdiff >>
rect 45923 4019 46057 4038
rect 45923 3985 45995 4019
rect 46029 3985 46057 4019
rect 45923 3968 46057 3985
rect 15781 3859 15915 3878
rect 15781 3825 15853 3859
rect 15887 3825 15915 3859
rect 15781 3808 15915 3825
<< nsubdiffcont >>
rect 45995 3985 46029 4019
rect 15853 3825 15887 3859
<< locali >>
rect 30618 4060 30974 4066
rect 30618 4026 30665 4060
rect 30699 4026 30753 4060
rect 30787 4026 30974 4060
rect 30618 4016 30974 4026
rect 45720 4019 46263 4039
rect 45720 3985 45995 4019
rect 46029 3985 46263 4019
rect 45720 3967 46263 3985
rect 15578 3859 16121 3879
rect 15578 3825 15853 3859
rect 15887 3825 16121 3859
rect 15578 3807 16121 3825
<< viali >>
rect 30665 4026 30699 4060
rect 30753 4026 30787 4060
rect 31330 4058 31364 4092
rect 31601 4022 31635 4056
rect 31689 4022 31723 4056
rect 31777 4022 31811 4056
rect 31865 4022 31899 4056
rect 31953 4022 31987 4056
rect 32041 4022 32075 4056
rect 32129 4022 32163 4056
rect 32217 4022 32251 4056
rect 31330 3978 31364 4012
rect 31955 3920 31989 3954
rect 32121 3916 32155 3950
rect 32289 3922 32323 3956
rect 32456 3920 32490 3954
rect 32626 3921 32660 3955
rect 32790 3922 32824 3956
rect 44421 3899 44455 3944
rect 44589 3906 44623 3951
rect 44757 3896 44791 3941
rect 44925 3908 44959 3953
rect 45091 3906 45125 3951
rect 45257 3908 45291 3953
rect 45425 3908 45459 3953
rect 45599 3906 45633 3951
rect 46355 3900 46389 3945
rect 46517 3904 46551 3949
rect 46687 3908 46721 3953
rect 46851 3904 46885 3949
rect 47021 3904 47055 3949
rect 47189 3900 47223 3945
rect 47357 3904 47391 3949
rect 47531 3900 47565 3945
rect 44621 3808 44655 3842
rect 44721 3808 44755 3842
rect 44821 3808 44855 3842
rect 44921 3808 44955 3842
rect 45021 3808 45055 3842
rect 45121 3808 45155 3842
rect 45221 3808 45255 3842
rect 45321 3808 45355 3842
rect 46281 3808 46315 3842
rect 46381 3808 46415 3842
rect 46481 3808 46515 3842
rect 46581 3808 46615 3842
rect 46681 3808 46715 3842
rect 46781 3808 46815 3842
rect 46881 3808 46915 3842
rect 46981 3808 47015 3842
rect 14279 3739 14313 3784
rect 14447 3746 14481 3791
rect 14615 3736 14649 3781
rect 14783 3748 14817 3793
rect 14949 3746 14983 3791
rect 15115 3748 15149 3793
rect 15283 3748 15317 3793
rect 15457 3746 15491 3791
rect 16213 3740 16247 3785
rect 16375 3744 16409 3789
rect 16545 3748 16579 3793
rect 16709 3744 16743 3789
rect 16879 3744 16913 3789
rect 17047 3740 17081 3785
rect 17215 3744 17249 3789
rect 17389 3740 17423 3785
rect 14479 3648 14513 3682
rect 14579 3648 14613 3682
rect 14679 3648 14713 3682
rect 14779 3648 14813 3682
rect 14879 3648 14913 3682
rect 14979 3648 15013 3682
rect 15079 3648 15113 3682
rect 15179 3648 15213 3682
rect 16139 3648 16173 3682
rect 16239 3648 16273 3682
rect 16339 3648 16373 3682
rect 16439 3648 16473 3682
rect 16539 3648 16573 3682
rect 16639 3648 16673 3682
rect 16739 3648 16773 3682
rect 16839 3648 16873 3682
<< metal1 >>
rect 15330 4977 15585 5333
rect 31266 5000 31600 5324
rect 15330 4925 15350 4977
rect 15402 4925 15428 4977
rect 15480 4925 15521 4977
rect 15573 4925 15585 4977
rect 15330 4895 15585 4925
rect 31266 4948 31309 5000
rect 31361 4948 31422 5000
rect 31474 4948 31523 5000
rect 31575 4948 31600 5000
rect 31266 4904 31600 4948
rect 45470 4977 45697 5345
rect 45470 4925 45501 4977
rect 45553 4925 45584 4977
rect 45636 4925 45697 4977
rect 45470 4891 45697 4925
rect 7986 4760 8522 4844
rect 23020 4769 23628 4827
rect 38124 4777 38748 4835
rect 53130 4783 53863 4841
rect 31394 4380 31502 4393
rect 31394 4328 31424 4380
rect 31476 4328 31502 4380
rect 31394 4297 31502 4328
rect 32934 4297 32969 4393
rect 0 4161 18000 4227
rect 17934 4075 18000 4161
rect 45639 4153 46306 4162
rect 31315 4092 31394 4120
rect 45649 4104 46306 4153
rect 17934 4060 30881 4075
rect 17934 4026 30665 4060
rect 30699 4026 30753 4060
rect 30787 4026 30881 4060
rect 17934 4009 30881 4026
rect 31315 4058 31330 4092
rect 31364 4064 31394 4092
rect 31364 4058 32313 4064
rect 31315 4056 32313 4058
rect 31315 4022 31601 4056
rect 31635 4022 31689 4056
rect 31723 4022 31777 4056
rect 31811 4022 31865 4056
rect 31899 4022 31953 4056
rect 31987 4022 32041 4056
rect 32075 4022 32129 4056
rect 32163 4022 32217 4056
rect 32251 4022 32313 4056
rect 31315 4016 32313 4022
rect 31315 4012 31397 4016
rect 15549 3948 16198 3998
rect 31315 3978 31330 4012
rect 31364 3978 31397 4012
rect 31315 3960 31397 3978
rect 31886 3971 32831 3984
rect 15497 3940 16198 3948
rect 31886 3954 32102 3971
rect 31886 3920 31955 3954
rect 31989 3920 32102 3954
rect 32154 3950 32262 3971
rect 32314 3956 32395 3971
rect 31886 3919 32102 3920
rect 32155 3919 32262 3950
rect 32323 3922 32395 3956
rect 32314 3919 32395 3922
rect 32447 3954 32508 3971
rect 32447 3920 32456 3954
rect 32490 3920 32508 3954
rect 32447 3919 32508 3920
rect 32560 3956 32831 3971
rect 32560 3955 32790 3956
rect 32560 3921 32626 3955
rect 32660 3922 32790 3955
rect 32824 3922 32831 3956
rect 32660 3921 32831 3922
rect 32560 3919 32831 3921
rect 31886 3916 32121 3919
rect 32155 3916 32831 3919
rect 31886 3901 32831 3916
rect 38288 3953 53723 3963
rect 38288 3951 44925 3953
rect 38288 3944 44589 3951
rect 38288 3943 38470 3944
rect 38288 3891 38367 3943
rect 38419 3892 38470 3943
rect 38522 3899 44421 3944
rect 44455 3906 44589 3944
rect 44623 3941 44925 3951
rect 44623 3906 44757 3941
rect 44455 3899 44757 3906
rect 38522 3896 44757 3899
rect 44791 3908 44925 3941
rect 44959 3951 45257 3953
rect 44959 3908 45091 3951
rect 44791 3906 45091 3908
rect 45125 3908 45257 3951
rect 45291 3908 45425 3953
rect 45459 3951 46687 3953
rect 45459 3908 45599 3951
rect 45125 3906 45599 3908
rect 45633 3949 46687 3951
rect 45633 3945 46517 3949
rect 45633 3906 46355 3945
rect 44791 3900 46355 3906
rect 46389 3904 46517 3945
rect 46551 3908 46687 3949
rect 46721 3949 53723 3953
rect 46721 3908 46851 3949
rect 46551 3904 46851 3908
rect 46885 3904 47021 3949
rect 47055 3945 47357 3949
rect 47055 3904 47189 3945
rect 46389 3900 47189 3904
rect 47223 3904 47357 3945
rect 47391 3945 53723 3949
rect 47391 3904 47531 3945
rect 47223 3900 47531 3904
rect 47565 3944 53723 3945
rect 47565 3939 53571 3944
rect 47565 3900 53480 3939
rect 44791 3896 53480 3900
rect 38522 3892 53480 3896
rect 38419 3891 53480 3892
rect 38288 3887 53480 3891
rect 53532 3892 53571 3939
rect 53623 3892 53723 3944
rect 53532 3887 53723 3892
rect 38288 3882 53723 3887
rect 31394 3830 31497 3849
rect 31394 3827 31484 3830
rect 8131 3793 23497 3803
rect 8131 3791 14783 3793
rect 8131 3788 14447 3791
rect 8131 3736 8172 3788
rect 8224 3736 8268 3788
rect 8320 3784 14447 3788
rect 8320 3739 14279 3784
rect 14313 3746 14447 3784
rect 14481 3781 14783 3791
rect 14481 3746 14615 3781
rect 14313 3739 14615 3746
rect 8320 3736 14615 3739
rect 14649 3748 14783 3781
rect 14817 3791 15115 3793
rect 14817 3748 14949 3791
rect 14649 3746 14949 3748
rect 14983 3748 15115 3791
rect 15149 3748 15283 3793
rect 15317 3791 16545 3793
rect 15317 3748 15457 3791
rect 14983 3746 15457 3748
rect 15491 3789 16545 3791
rect 15491 3785 16375 3789
rect 15491 3746 16213 3785
rect 14649 3740 16213 3746
rect 16247 3744 16375 3785
rect 16409 3748 16545 3789
rect 16579 3789 23497 3793
rect 16579 3748 16709 3789
rect 16409 3744 16709 3748
rect 16743 3744 16879 3789
rect 16913 3785 17215 3789
rect 16913 3744 17047 3785
rect 16247 3740 17047 3744
rect 17081 3744 17215 3785
rect 17249 3786 23497 3789
rect 17249 3785 23382 3786
rect 17249 3744 17389 3785
rect 17081 3740 17389 3744
rect 17423 3779 23382 3785
rect 17423 3740 23283 3779
rect 14649 3736 23283 3740
rect 8131 3727 23283 3736
rect 23335 3734 23382 3779
rect 23434 3734 23497 3786
rect 31425 3778 31484 3827
rect 31425 3775 31497 3778
rect 31394 3753 31497 3775
rect 32934 3753 32969 3849
rect 44589 3842 47192 3848
rect 44589 3808 44621 3842
rect 44655 3808 44721 3842
rect 44755 3808 44821 3842
rect 44855 3808 44921 3842
rect 44955 3808 45021 3842
rect 45055 3808 45121 3842
rect 45155 3808 45221 3842
rect 45255 3808 45321 3842
rect 45355 3808 46281 3842
rect 46315 3808 46381 3842
rect 46415 3808 46481 3842
rect 46515 3808 46581 3842
rect 46615 3808 46681 3842
rect 46715 3808 46781 3842
rect 46815 3808 46881 3842
rect 46915 3808 46981 3842
rect 47015 3808 47192 3842
rect 44589 3803 47192 3808
rect 44589 3800 46035 3803
rect 45885 3799 46035 3800
rect 23335 3727 23497 3734
rect 8131 3722 23497 3727
rect 45885 3747 45930 3799
rect 45982 3751 46035 3799
rect 46087 3800 47192 3803
rect 46087 3751 46113 3800
rect 45982 3747 46113 3751
rect 45885 3708 46113 3747
rect 14447 3682 17050 3688
rect 14447 3648 14479 3682
rect 14513 3648 14579 3682
rect 14613 3648 14679 3682
rect 14713 3648 14779 3682
rect 14813 3648 14879 3682
rect 14913 3648 14979 3682
rect 15013 3648 15079 3682
rect 15113 3648 15179 3682
rect 15213 3648 16139 3682
rect 16173 3648 16239 3682
rect 16273 3648 16339 3682
rect 16373 3648 16439 3682
rect 16473 3648 16539 3682
rect 16573 3648 16639 3682
rect 16673 3648 16739 3682
rect 16773 3648 16839 3682
rect 16873 3648 17050 3682
rect 14447 3643 17050 3648
rect 14447 3640 15893 3643
rect 15743 3639 15893 3640
rect 15743 3587 15788 3639
rect 15840 3591 15893 3639
rect 15945 3640 17050 3643
rect 15945 3591 15971 3640
rect 15840 3587 15971 3591
rect 15743 3548 15971 3587
rect 45639 3556 46391 3614
rect 14109 3378 14160 3474
rect 15497 3402 16178 3460
rect 20628 3405 46139 3449
rect 20628 3403 46027 3405
rect 14109 3377 14159 3378
rect 20628 3351 32091 3403
rect 32143 3351 32235 3403
rect 32287 3351 32379 3403
rect 32431 3402 46027 3403
rect 32431 3351 45938 3402
rect 20628 3350 45938 3351
rect 45990 3353 46027 3402
rect 46079 3353 46139 3405
rect 45990 3350 46139 3353
rect 20628 3326 46139 3350
rect 20628 3319 45938 3326
rect 20628 3267 32090 3319
rect 32142 3267 32234 3319
rect 32286 3267 32378 3319
rect 32430 3274 45938 3319
rect 45990 3274 46031 3326
rect 46083 3274 46139 3326
rect 32430 3267 46139 3274
rect 15755 3243 46139 3267
rect 15755 3222 20834 3243
rect 15755 3170 15792 3222
rect 15844 3217 20834 3222
rect 15844 3170 15886 3217
rect 15755 3165 15886 3170
rect 15938 3165 20834 3217
rect 15755 3144 20834 3165
rect 15755 3142 15886 3144
rect 7922 3068 8585 3126
rect 15755 3090 15792 3142
rect 15844 3092 15886 3142
rect 15938 3092 20834 3144
rect 15844 3090 20834 3092
rect 15755 3061 20834 3090
rect 23020 3080 23648 3138
rect 38032 3080 38795 3138
rect 53222 3071 53873 3129
rect 61289 1010 61511 1088
<< via1 >>
rect 8171 4991 8223 5043
rect 8252 4990 8304 5042
rect 23287 4988 23339 5040
rect 23382 4988 23434 5040
rect 15350 4925 15402 4977
rect 15428 4925 15480 4977
rect 15521 4925 15573 4977
rect 31309 4948 31361 5000
rect 31422 4948 31474 5000
rect 31523 4948 31575 5000
rect 38364 4990 38416 5042
rect 38466 4990 38518 5042
rect 45501 4925 45553 4977
rect 45584 4925 45636 4977
rect 53482 4963 53534 5015
rect 53577 4963 53629 5015
rect 7179 4769 7231 4821
rect 7286 4771 7338 4823
rect 7388 4771 7440 4823
rect 7488 4772 7540 4824
rect 22209 4775 22261 4827
rect 22312 4775 22364 4827
rect 22395 4775 22447 4827
rect 22496 4775 22548 4827
rect 22583 4775 22635 4827
rect 37341 4771 37393 4823
rect 37429 4771 37481 4823
rect 37514 4776 37566 4828
rect 54257 4768 54309 4820
rect 54351 4768 54403 4820
rect 54428 4768 54480 4820
rect 54508 4767 54560 4819
rect 54582 4768 54634 4820
rect 31321 4325 31373 4377
rect 31424 4328 31476 4380
rect 31525 4328 31577 4380
rect 45507 4100 45559 4152
rect 45597 4101 45649 4153
rect 15374 3948 15426 4000
rect 15497 3948 15549 4000
rect 32102 3950 32154 3971
rect 32262 3956 32314 3971
rect 32102 3919 32121 3950
rect 32121 3919 32154 3950
rect 32262 3922 32289 3956
rect 32289 3922 32314 3956
rect 32262 3919 32314 3922
rect 32395 3919 32447 3971
rect 32508 3919 32560 3971
rect 38367 3891 38419 3943
rect 38470 3892 38522 3944
rect 53480 3887 53532 3939
rect 53571 3892 53623 3944
rect 8172 3736 8224 3788
rect 8268 3736 8320 3788
rect 23283 3727 23335 3779
rect 23382 3734 23434 3786
rect 31277 3773 31329 3825
rect 31373 3775 31425 3827
rect 31484 3778 31536 3830
rect 31576 3775 31628 3827
rect 45930 3747 45982 3799
rect 46035 3751 46087 3803
rect 15788 3587 15840 3639
rect 15893 3591 15945 3643
rect 46942 3560 46994 3612
rect 47034 3561 47086 3613
rect 47124 3560 47176 3612
rect 47212 3559 47264 3611
rect 14587 3399 14639 3451
rect 14671 3399 14723 3451
rect 14764 3400 14816 3452
rect 32091 3351 32143 3403
rect 32235 3351 32287 3403
rect 32379 3351 32431 3403
rect 45938 3350 45990 3402
rect 46027 3353 46079 3405
rect 32090 3267 32142 3319
rect 32234 3267 32286 3319
rect 32378 3267 32430 3319
rect 45938 3274 45990 3326
rect 46031 3274 46083 3326
rect 15792 3170 15844 3222
rect 15886 3165 15938 3217
rect 7173 3071 7225 3123
rect 7271 3071 7323 3123
rect 7366 3071 7418 3123
rect 7471 3071 7523 3123
rect 15792 3090 15844 3142
rect 15886 3092 15938 3144
rect 22223 3076 22275 3128
rect 22323 3076 22375 3128
rect 22422 3076 22474 3128
rect 22525 3076 22577 3128
rect 37331 3070 37383 3122
rect 37419 3070 37471 3122
rect 37517 3066 37569 3118
rect 54253 3067 54305 3119
rect 54341 3067 54393 3119
rect 54424 3067 54476 3119
rect 54511 3067 54563 3119
rect 8172 2853 8224 2905
rect 8252 2851 8304 2903
rect 23288 2868 23340 2920
rect 23371 2868 23423 2920
rect 38366 2858 38418 2910
rect 38457 2858 38509 2910
rect 53483 2843 53535 2895
rect 53566 2843 53618 2895
<< metal2 >>
rect 2297 6878 2341 8034
rect 4185 6878 4229 8034
rect 6073 6878 6117 8034
rect 7961 6878 8005 8034
rect 9849 6878 9893 8034
rect 11737 6878 11781 8034
rect 13625 6878 13669 8034
rect 15513 6878 15557 8034
rect 17401 6878 17445 8034
rect 19289 6878 19333 8034
rect 21177 6878 21221 8034
rect 23065 6878 23109 8034
rect 24953 6878 24997 8034
rect 26841 6878 26885 8034
rect 28729 6878 28773 8034
rect 30617 6878 30661 8034
rect 32505 6878 32549 8034
rect 34393 6878 34437 8034
rect 36281 6878 36325 8034
rect 38169 6878 38213 8034
rect 40057 6878 40101 8034
rect 41945 6878 41989 8034
rect 43833 6878 43877 8034
rect 45721 6878 45765 8034
rect 47609 6878 47653 8034
rect 49497 6878 49541 8034
rect 51385 6878 51429 8034
rect 53273 6878 53317 8034
rect 55161 6878 55205 8034
rect 57049 6878 57093 8034
rect 58937 6878 58981 8034
rect 60825 6878 60869 8034
rect 61398 6196 61512 6243
rect 271 6160 513 6196
rect 60845 6160 61512 6196
rect 271 6106 387 6160
rect 278 1740 368 6106
rect 8147 5043 8336 5073
rect 8147 4991 8171 5043
rect 8223 5042 8336 5043
rect 8223 4991 8252 5042
rect 8147 4990 8252 4991
rect 8304 4990 8336 5042
rect 7115 4824 7599 4949
rect 7115 4823 7488 4824
rect 7115 4821 7286 4823
rect 7115 4769 7179 4821
rect 7231 4771 7286 4821
rect 7338 4771 7388 4823
rect 7440 4772 7488 4823
rect 7540 4772 7599 4824
rect 7440 4771 7599 4772
rect 7231 4769 7599 4771
rect 7115 3602 7599 4769
rect 7115 3546 7182 3602
rect 7238 3546 7296 3602
rect 7352 3546 7410 3602
rect 7466 3546 7599 3602
rect 7115 3487 7599 3546
rect 7115 3431 7182 3487
rect 7238 3431 7296 3487
rect 7352 3431 7410 3487
rect 7466 3431 7599 3487
rect 7115 3372 7599 3431
rect 7115 3316 7182 3372
rect 7238 3316 7296 3372
rect 7352 3316 7410 3372
rect 7466 3316 7599 3372
rect 7115 3123 7599 3316
rect 7115 3071 7173 3123
rect 7225 3071 7271 3123
rect 7323 3071 7366 3123
rect 7418 3071 7471 3123
rect 7523 3071 7599 3123
rect 7115 2959 7599 3071
rect 8147 3788 8336 4990
rect 15330 4977 15590 5048
rect 15330 4925 15350 4977
rect 15402 4925 15428 4977
rect 15480 4925 15521 4977
rect 15573 4925 15590 4977
rect 23258 5040 23447 5063
rect 23258 4988 23287 5040
rect 23339 4988 23382 5040
rect 23434 4988 23447 5040
rect 15330 4000 15590 4925
rect 15330 3948 15374 4000
rect 15426 3948 15497 4000
rect 15549 3948 15590 4000
rect 15330 3904 15590 3948
rect 22171 4827 22638 4927
rect 22171 4775 22209 4827
rect 22261 4775 22312 4827
rect 22364 4775 22395 4827
rect 22447 4775 22496 4827
rect 22548 4775 22583 4827
rect 22635 4775 22638 4827
rect 8147 3736 8172 3788
rect 8224 3736 8268 3788
rect 8320 3736 8336 3788
rect 8147 2905 8336 3736
rect 15755 3643 15961 3688
rect 15755 3639 15893 3643
rect 15755 3587 15788 3639
rect 15840 3591 15893 3639
rect 15945 3591 15961 3643
rect 15840 3587 15961 3591
rect 8147 2853 8172 2905
rect 8224 2903 8336 2905
rect 8224 2853 8252 2903
rect 8147 2851 8252 2853
rect 8304 2851 8336 2903
rect 14536 3452 14889 3498
rect 14536 3451 14764 3452
rect 14536 3399 14587 3451
rect 14639 3399 14671 3451
rect 14723 3400 14764 3451
rect 14816 3400 14889 3452
rect 14723 3399 14889 3400
rect 14536 3041 14889 3399
rect 15755 3222 15961 3587
rect 15755 3170 15792 3222
rect 15844 3217 15961 3222
rect 15844 3170 15886 3217
rect 15755 3165 15886 3170
rect 15938 3165 15961 3217
rect 15755 3144 15961 3165
rect 15755 3142 15886 3144
rect 15755 3090 15792 3142
rect 15844 3092 15886 3142
rect 15938 3092 15961 3144
rect 15844 3090 15961 3092
rect 15755 3061 15961 3090
rect 22171 3512 22638 4775
rect 22171 3456 22221 3512
rect 22277 3456 22325 3512
rect 22381 3456 22429 3512
rect 22485 3456 22533 3512
rect 22589 3456 22638 3512
rect 22171 3396 22638 3456
rect 22171 3340 22221 3396
rect 22277 3340 22325 3396
rect 22381 3340 22429 3396
rect 22485 3340 22533 3396
rect 22589 3340 22638 3396
rect 22171 3280 22638 3340
rect 22171 3224 22221 3280
rect 22277 3224 22325 3280
rect 22381 3224 22429 3280
rect 22485 3224 22533 3280
rect 22589 3224 22638 3280
rect 22171 3128 22638 3224
rect 22171 3076 22223 3128
rect 22275 3076 22323 3128
rect 22375 3076 22422 3128
rect 22474 3076 22525 3128
rect 22577 3076 22638 3128
rect 14536 2985 14576 3041
rect 14632 2985 14684 3041
rect 14740 2985 14792 3041
rect 14848 2985 14889 3041
rect 14536 2947 14889 2985
rect 22171 2976 22638 3076
rect 23258 3786 23447 4988
rect 31263 5000 31598 5043
rect 31263 4948 31309 5000
rect 31361 4948 31422 5000
rect 31474 4948 31523 5000
rect 31575 4948 31598 5000
rect 31263 4380 31598 4948
rect 38349 5042 38536 5061
rect 38349 4990 38364 5042
rect 38416 4990 38466 5042
rect 38518 4990 38536 5042
rect 31263 4377 31424 4380
rect 31263 4325 31321 4377
rect 31373 4328 31424 4377
rect 31476 4328 31525 4380
rect 31577 4328 31598 4380
rect 31373 4325 31598 4328
rect 31263 4293 31598 4325
rect 37287 4828 37587 4925
rect 37287 4823 37514 4828
rect 37287 4771 37341 4823
rect 37393 4771 37429 4823
rect 37481 4776 37514 4823
rect 37566 4776 37587 4828
rect 37481 4771 37587 4776
rect 32034 3971 32573 3994
rect 32034 3919 32102 3971
rect 32154 3919 32262 3971
rect 32314 3919 32395 3971
rect 32447 3919 32508 3971
rect 32560 3919 32573 3971
rect 23258 3779 23382 3786
rect 23258 3727 23283 3779
rect 23335 3734 23382 3779
rect 23434 3734 23447 3786
rect 23335 3727 23447 3734
rect 14536 2891 14576 2947
rect 14632 2891 14684 2947
rect 14740 2891 14792 2947
rect 14848 2891 14889 2947
rect 14536 2865 14889 2891
rect 23258 2920 23447 3727
rect 31225 3830 31650 3848
rect 31225 3827 31484 3830
rect 31225 3825 31373 3827
rect 31225 3773 31277 3825
rect 31329 3775 31373 3825
rect 31425 3778 31484 3827
rect 31536 3827 31650 3830
rect 31536 3778 31576 3827
rect 31425 3775 31576 3778
rect 31628 3775 31650 3827
rect 31329 3773 31650 3775
rect 31225 3161 31650 3773
rect 32034 3403 32573 3919
rect 32034 3351 32091 3403
rect 32143 3351 32235 3403
rect 32287 3351 32379 3403
rect 32431 3351 32573 3403
rect 32034 3319 32573 3351
rect 32034 3267 32090 3319
rect 32142 3267 32234 3319
rect 32286 3267 32378 3319
rect 32430 3267 32573 3319
rect 32034 3193 32573 3267
rect 37287 3861 37587 4771
rect 37287 3805 37308 3861
rect 37364 3805 37402 3861
rect 37458 3805 37496 3861
rect 37552 3805 37587 3861
rect 37287 3773 37587 3805
rect 37287 3717 37308 3773
rect 37364 3717 37402 3773
rect 37458 3717 37496 3773
rect 37552 3717 37587 3773
rect 37287 3685 37587 3717
rect 37287 3629 37308 3685
rect 37364 3629 37402 3685
rect 37458 3629 37496 3685
rect 37552 3629 37587 3685
rect 31225 3105 31271 3161
rect 31327 3105 31396 3161
rect 31452 3105 31521 3161
rect 31577 3105 31650 3161
rect 31225 3065 31650 3105
rect 31225 3009 31271 3065
rect 31327 3009 31396 3065
rect 31452 3009 31521 3065
rect 31577 3009 31650 3065
rect 31225 2977 31650 3009
rect 37287 3122 37587 3629
rect 37287 3070 37331 3122
rect 37383 3070 37419 3122
rect 37471 3118 37587 3122
rect 37471 3070 37517 3118
rect 37287 3066 37517 3070
rect 37569 3066 37587 3118
rect 37287 2973 37587 3066
rect 38349 3944 38536 4990
rect 45478 4977 45697 5030
rect 45478 4925 45501 4977
rect 45553 4925 45584 4977
rect 45636 4925 45697 4977
rect 45478 4153 45697 4925
rect 45478 4152 45597 4153
rect 45478 4100 45507 4152
rect 45559 4101 45597 4152
rect 45649 4101 45697 4153
rect 45559 4100 45697 4101
rect 45478 4065 45697 4100
rect 53453 5015 53642 5038
rect 53453 4963 53482 5015
rect 53534 4963 53577 5015
rect 53629 4963 53642 5015
rect 38349 3943 38470 3944
rect 38349 3891 38367 3943
rect 38419 3892 38470 3943
rect 38522 3892 38536 3944
rect 38419 3891 38536 3892
rect 23258 2868 23288 2920
rect 23340 2868 23371 2920
rect 23423 2868 23447 2920
rect 23258 2855 23447 2868
rect 38349 2910 38536 3891
rect 53453 3944 53642 4963
rect 53453 3939 53571 3944
rect 53453 3887 53480 3939
rect 53532 3892 53571 3939
rect 53623 3892 53642 3944
rect 53532 3887 53642 3892
rect 45897 3803 46103 3848
rect 45897 3799 46035 3803
rect 45897 3747 45930 3799
rect 45982 3751 46035 3799
rect 46087 3751 46103 3803
rect 45982 3747 46103 3751
rect 45897 3405 46103 3747
rect 45897 3402 46027 3405
rect 45897 3350 45938 3402
rect 45990 3353 46027 3402
rect 46079 3353 46103 3405
rect 45990 3350 46103 3353
rect 45897 3326 46103 3350
rect 45897 3274 45938 3326
rect 45990 3274 46031 3326
rect 46083 3274 46103 3326
rect 45897 3231 46103 3274
rect 46905 3613 47319 3635
rect 46905 3612 47034 3613
rect 46905 3560 46942 3612
rect 46994 3561 47034 3612
rect 47086 3612 47319 3613
rect 47086 3561 47124 3612
rect 46994 3560 47124 3561
rect 47176 3611 47319 3612
rect 47176 3560 47212 3611
rect 46905 3559 47212 3560
rect 47264 3559 47319 3611
rect 38349 2858 38366 2910
rect 38418 2858 38457 2910
rect 38509 2858 38536 2910
rect 8147 2833 8336 2851
rect 38349 2850 38536 2858
rect 46905 3014 47319 3559
rect 46905 2958 46942 3014
rect 46998 2958 47035 3014
rect 47091 2958 47128 3014
rect 47184 2958 47221 3014
rect 47277 2958 47319 3014
rect 46905 2932 47319 2958
rect 46905 2876 46942 2932
rect 46998 2876 47035 2932
rect 47091 2876 47128 2932
rect 47184 2876 47221 2932
rect 47277 2876 47319 2932
rect 46905 2839 47319 2876
rect 53453 2895 53642 3887
rect 54218 4820 54639 4925
rect 54218 4768 54257 4820
rect 54309 4768 54351 4820
rect 54403 4768 54428 4820
rect 54480 4819 54582 4820
rect 54480 4768 54508 4819
rect 54218 4767 54508 4768
rect 54560 4768 54582 4819
rect 54634 4768 54639 4820
rect 54560 4767 54639 4768
rect 54218 3406 54639 4767
rect 54218 3350 54255 3406
rect 54311 3350 54359 3406
rect 54415 3350 54463 3406
rect 54519 3350 54567 3406
rect 54623 3350 54639 3406
rect 54218 3316 54639 3350
rect 54218 3260 54255 3316
rect 54311 3260 54359 3316
rect 54415 3260 54463 3316
rect 54519 3260 54567 3316
rect 54623 3260 54639 3316
rect 54218 3119 54639 3260
rect 54218 3067 54253 3119
rect 54305 3067 54341 3119
rect 54393 3067 54424 3119
rect 54476 3067 54511 3119
rect 54563 3067 54639 3119
rect 54218 2975 54639 3067
rect 53453 2843 53483 2895
rect 53535 2843 53566 2895
rect 53618 2843 53642 2895
rect 53453 2830 53642 2843
rect 61398 1818 61512 6160
rect 61355 1740 61549 1818
rect 273 1704 958 1740
rect 61283 1704 61549 1740
rect 278 1621 368 1704
rect 927 124 971 1022
rect 2815 124 2859 1022
rect 4703 124 4747 1022
rect 6591 124 6635 1022
rect 8479 124 8523 1022
rect 10367 124 10411 1022
rect 12255 124 12299 1022
rect 14143 124 14187 1022
rect 16031 124 16075 1022
rect 17919 124 17963 1022
rect 19807 124 19851 1022
rect 21695 124 21739 1022
rect 23583 124 23627 1022
rect 25471 124 25515 1022
rect 27359 24 27403 1022
rect 29247 124 29291 1022
rect 31135 124 31179 1022
rect 33023 124 33067 1022
rect 34911 124 34955 1022
rect 36799 124 36843 1022
rect 38687 124 38731 1022
rect 40575 0 40619 1022
rect 42463 124 42507 1022
rect 44351 124 44395 1022
rect 46239 124 46283 1022
rect 48127 124 48171 1022
rect 50015 124 50059 1022
rect 51903 124 51947 1022
rect 53791 124 53835 1022
rect 55679 124 55723 1022
rect 57567 902 57611 1022
rect 57567 124 57613 902
rect 59455 124 59499 1022
rect 57569 4 57613 124
<< via2 >>
rect 7182 3546 7238 3602
rect 7296 3546 7352 3602
rect 7410 3546 7466 3602
rect 7182 3431 7238 3487
rect 7296 3431 7352 3487
rect 7410 3431 7466 3487
rect 7182 3316 7238 3372
rect 7296 3316 7352 3372
rect 7410 3316 7466 3372
rect 22221 3456 22277 3512
rect 22325 3456 22381 3512
rect 22429 3456 22485 3512
rect 22533 3456 22589 3512
rect 22221 3340 22277 3396
rect 22325 3340 22381 3396
rect 22429 3340 22485 3396
rect 22533 3340 22589 3396
rect 22221 3224 22277 3280
rect 22325 3224 22381 3280
rect 22429 3224 22485 3280
rect 22533 3224 22589 3280
rect 14576 2985 14632 3041
rect 14684 2985 14740 3041
rect 14792 2985 14848 3041
rect 14576 2891 14632 2947
rect 14684 2891 14740 2947
rect 14792 2891 14848 2947
rect 37308 3805 37364 3861
rect 37402 3805 37458 3861
rect 37496 3805 37552 3861
rect 37308 3717 37364 3773
rect 37402 3717 37458 3773
rect 37496 3717 37552 3773
rect 37308 3629 37364 3685
rect 37402 3629 37458 3685
rect 37496 3629 37552 3685
rect 31271 3105 31327 3161
rect 31396 3105 31452 3161
rect 31521 3105 31577 3161
rect 31271 3009 31327 3065
rect 31396 3009 31452 3065
rect 31521 3009 31577 3065
rect 46942 2958 46998 3014
rect 47035 2958 47091 3014
rect 47128 2958 47184 3014
rect 47221 2958 47277 3014
rect 46942 2876 46998 2932
rect 47035 2876 47091 2932
rect 47128 2876 47184 2932
rect 47221 2876 47277 2932
rect 54255 3350 54311 3406
rect 54359 3350 54415 3406
rect 54463 3350 54519 3406
rect 54567 3350 54623 3406
rect 54255 3260 54311 3316
rect 54359 3260 54415 3316
rect 54463 3260 54519 3316
rect 54567 3260 54623 3316
<< metal3 >>
rect 37285 3861 37589 3875
rect 37285 3805 37308 3861
rect 37364 3805 37402 3861
rect 37458 3805 37496 3861
rect 37552 3805 37589 3861
rect 37285 3773 37589 3805
rect 37285 3717 37308 3773
rect 37364 3762 37402 3773
rect 37458 3763 37496 3773
rect 37552 3763 37589 3773
rect 37458 3717 37475 3763
rect 37285 3685 37321 3717
rect 37408 3685 37475 3717
rect 7181 3628 7523 3661
rect 37285 3629 37308 3685
rect 37458 3651 37475 3685
rect 37562 3651 37589 3763
rect 37364 3629 37402 3650
rect 37458 3629 37496 3651
rect 37552 3629 37589 3651
rect 7113 3602 7602 3628
rect 37285 3609 37589 3629
rect 7113 3546 7182 3602
rect 7238 3546 7296 3602
rect 7352 3546 7410 3602
rect 7466 3546 7602 3602
rect 7113 3487 7602 3546
rect 7113 3459 7182 3487
rect 7238 3459 7296 3487
rect 7352 3465 7410 3487
rect 7466 3465 7602 3487
rect 7113 3368 7179 3459
rect 7265 3431 7296 3459
rect 7466 3431 7475 3465
rect 7265 3374 7330 3431
rect 7416 3374 7475 3431
rect 7561 3374 7602 3465
rect 7265 3372 7602 3374
rect 7265 3368 7296 3372
rect 7113 3316 7182 3368
rect 7238 3316 7296 3368
rect 7352 3316 7410 3372
rect 7466 3316 7602 3372
rect 7113 3261 7602 3316
rect 22171 3512 22638 3566
rect 22171 3469 22221 3512
rect 22277 3469 22325 3512
rect 22171 3385 22219 3469
rect 22312 3456 22325 3469
rect 22381 3469 22429 3512
rect 22381 3456 22386 3469
rect 22485 3456 22533 3512
rect 22589 3456 22638 3512
rect 22312 3396 22386 3456
rect 22479 3396 22638 3456
rect 22312 3385 22325 3396
rect 22171 3340 22221 3385
rect 22277 3340 22325 3385
rect 22381 3385 22386 3396
rect 22381 3340 22429 3385
rect 22485 3340 22533 3396
rect 22589 3340 22638 3396
rect 22171 3308 22638 3340
rect 22171 3224 22219 3308
rect 22312 3280 22386 3308
rect 22479 3280 22638 3308
rect 22312 3224 22325 3280
rect 22381 3224 22386 3280
rect 22485 3224 22533 3280
rect 22589 3224 22638 3280
rect 54218 3413 54640 3434
rect 54218 3406 54262 3413
rect 54346 3406 54383 3413
rect 54467 3406 54521 3413
rect 54605 3406 54640 3413
rect 54218 3350 54255 3406
rect 54346 3350 54359 3406
rect 54519 3350 54521 3406
rect 54623 3350 54640 3406
rect 54218 3316 54262 3350
rect 54346 3316 54383 3350
rect 54467 3316 54521 3350
rect 54605 3316 54640 3350
rect 54218 3260 54255 3316
rect 54346 3260 54359 3316
rect 54519 3260 54521 3316
rect 54623 3260 54640 3316
rect 54218 3255 54262 3260
rect 54346 3255 54383 3260
rect 54467 3255 54521 3260
rect 54605 3255 54640 3260
rect 54218 3226 54640 3255
rect 22171 3180 22638 3224
rect 31223 3161 31648 3199
rect 31223 3122 31271 3161
rect 31327 3122 31396 3161
rect 31452 3122 31521 3161
rect 31577 3122 31648 3161
rect 14536 3041 14889 3064
rect 14536 2993 14576 3041
rect 14632 2993 14684 3041
rect 14740 2993 14792 3041
rect 14536 2924 14560 2993
rect 14637 2924 14663 2993
rect 14740 2924 14766 2993
rect 14848 2985 14889 3041
rect 14843 2947 14889 2985
rect 31223 3010 31269 3122
rect 31356 3010 31388 3122
rect 31475 3010 31507 3122
rect 31594 3010 31648 3122
rect 31223 3009 31271 3010
rect 31327 3009 31396 3010
rect 31452 3009 31521 3010
rect 31577 3009 31648 3010
rect 31223 2972 31648 3009
rect 46905 3038 47320 3081
rect 46905 3037 47083 3038
rect 46905 3014 46943 3037
rect 47027 3014 47083 3037
rect 47167 3014 47211 3038
rect 14536 2891 14576 2924
rect 14632 2891 14684 2924
rect 14740 2891 14792 2924
rect 14848 2891 14889 2947
rect 14536 2865 14889 2891
rect 46905 2958 46942 3014
rect 47027 2958 47035 3014
rect 47184 2958 47211 3014
rect 46905 2932 46943 2958
rect 47027 2932 47083 2958
rect 47167 2932 47211 2958
rect 46905 2876 46942 2932
rect 47027 2879 47035 2932
rect 47184 2880 47211 2932
rect 47295 2880 47320 3038
rect 46998 2876 47035 2879
rect 47091 2876 47128 2880
rect 47184 2876 47221 2880
rect 47277 2876 47320 2880
rect 46905 2840 47320 2876
<< via3 >>
rect 3425 7441 3531 7619
rect 3634 7440 3740 7618
rect 3800 7440 3906 7618
rect 3980 7442 4086 7620
rect 20054 7458 20160 7636
rect 20270 7458 20376 7636
rect 20486 7458 20592 7636
rect 28546 7457 28652 7635
rect 28762 7457 28868 7635
rect 28978 7457 29084 7635
rect 42074 7463 42180 7641
rect 42290 7463 42396 7641
rect 42506 7463 42612 7641
rect 58559 7456 58665 7634
rect 58775 7456 58881 7634
rect 58991 7456 59097 7634
rect 2191 5323 2297 5501
rect 2363 5324 2469 5502
rect 2537 5323 2643 5501
rect 18519 5344 18625 5522
rect 18735 5344 18841 5522
rect 18951 5344 19057 5522
rect 27027 5336 27133 5514
rect 27243 5336 27349 5514
rect 27459 5336 27565 5514
rect 40499 5331 40605 5509
rect 40715 5331 40821 5509
rect 40931 5331 41037 5509
rect 57050 5323 57156 5501
rect 57266 5323 57372 5501
rect 57482 5323 57588 5501
rect 37321 3717 37364 3762
rect 37364 3717 37402 3762
rect 37402 3717 37408 3762
rect 37475 3717 37496 3763
rect 37496 3717 37552 3763
rect 37552 3717 37562 3763
rect 37321 3685 37408 3717
rect 37475 3685 37562 3717
rect 37321 3650 37364 3685
rect 37364 3650 37402 3685
rect 37402 3650 37408 3685
rect 37475 3651 37496 3685
rect 37496 3651 37552 3685
rect 37552 3651 37562 3685
rect 7179 3431 7182 3459
rect 7182 3431 7238 3459
rect 7238 3431 7265 3459
rect 7330 3431 7352 3465
rect 7352 3431 7410 3465
rect 7410 3431 7416 3465
rect 7179 3372 7265 3431
rect 7330 3374 7416 3431
rect 7475 3374 7561 3465
rect 7179 3368 7182 3372
rect 7182 3368 7238 3372
rect 7238 3368 7265 3372
rect 22219 3456 22221 3469
rect 22221 3456 22277 3469
rect 22277 3456 22312 3469
rect 22386 3456 22429 3469
rect 22429 3456 22479 3469
rect 22219 3396 22312 3456
rect 22386 3396 22479 3456
rect 22219 3385 22221 3396
rect 22221 3385 22277 3396
rect 22277 3385 22312 3396
rect 22386 3385 22429 3396
rect 22429 3385 22479 3396
rect 22219 3280 22312 3308
rect 22386 3280 22479 3308
rect 22219 3224 22221 3280
rect 22221 3224 22277 3280
rect 22277 3224 22312 3280
rect 22386 3224 22429 3280
rect 22429 3224 22479 3280
rect 54262 3406 54346 3413
rect 54383 3406 54467 3413
rect 54521 3406 54605 3413
rect 54262 3350 54311 3406
rect 54311 3350 54346 3406
rect 54383 3350 54415 3406
rect 54415 3350 54463 3406
rect 54463 3350 54467 3406
rect 54521 3350 54567 3406
rect 54567 3350 54605 3406
rect 54262 3316 54346 3350
rect 54383 3316 54467 3350
rect 54521 3316 54605 3350
rect 54262 3260 54311 3316
rect 54311 3260 54346 3316
rect 54383 3260 54415 3316
rect 54415 3260 54463 3316
rect 54463 3260 54467 3316
rect 54521 3260 54567 3316
rect 54567 3260 54605 3316
rect 54262 3255 54346 3260
rect 54383 3255 54467 3260
rect 54521 3255 54605 3260
rect 14560 2985 14576 2993
rect 14576 2985 14632 2993
rect 14632 2985 14637 2993
rect 14560 2947 14637 2985
rect 14560 2924 14576 2947
rect 14576 2924 14632 2947
rect 14632 2924 14637 2947
rect 14663 2985 14684 2993
rect 14684 2985 14740 2993
rect 14663 2947 14740 2985
rect 14663 2924 14684 2947
rect 14684 2924 14740 2947
rect 14766 2985 14792 2993
rect 14792 2985 14843 2993
rect 14766 2947 14843 2985
rect 31269 3105 31271 3122
rect 31271 3105 31327 3122
rect 31327 3105 31356 3122
rect 31269 3065 31356 3105
rect 31269 3010 31271 3065
rect 31271 3010 31327 3065
rect 31327 3010 31356 3065
rect 31388 3105 31396 3122
rect 31396 3105 31452 3122
rect 31452 3105 31475 3122
rect 31388 3065 31475 3105
rect 31388 3010 31396 3065
rect 31396 3010 31452 3065
rect 31452 3010 31475 3065
rect 31507 3105 31521 3122
rect 31521 3105 31577 3122
rect 31577 3105 31594 3122
rect 31507 3065 31594 3105
rect 31507 3010 31521 3065
rect 31521 3010 31577 3065
rect 31577 3010 31594 3065
rect 46943 3014 47027 3037
rect 47083 3014 47167 3038
rect 47211 3014 47295 3038
rect 14766 2924 14792 2947
rect 14792 2924 14843 2947
rect 46943 2958 46998 3014
rect 46998 2958 47027 3014
rect 47083 2958 47091 3014
rect 47091 2958 47128 3014
rect 47128 2958 47167 3014
rect 47211 2958 47221 3014
rect 47221 2958 47277 3014
rect 47277 2958 47295 3014
rect 46943 2932 47027 2958
rect 47083 2932 47167 2958
rect 47211 2932 47295 2958
rect 46943 2879 46998 2932
rect 46998 2879 47027 2932
rect 47083 2880 47091 2932
rect 47091 2880 47128 2932
rect 47128 2880 47167 2932
rect 47211 2880 47221 2932
rect 47221 2880 47277 2932
rect 47277 2880 47295 2932
rect 2193 2375 2299 2553
rect 2398 2377 2504 2555
rect 2597 2377 2703 2555
rect 18510 2393 18616 2571
rect 18726 2393 18832 2571
rect 18942 2393 19048 2571
rect 27032 2388 27138 2566
rect 27248 2388 27354 2566
rect 27464 2388 27570 2566
rect 40535 2390 40641 2568
rect 40751 2390 40857 2568
rect 40967 2390 41073 2568
rect 57030 2401 57136 2579
rect 57246 2401 57352 2579
rect 57462 2401 57568 2579
rect 3439 264 3545 442
rect 3660 264 3766 442
rect 3869 264 3975 442
rect 4043 264 4149 442
rect 7167 296 7253 387
rect 7315 296 7401 387
rect 7463 296 7549 387
rect 14686 370 14763 439
rect 14709 251 14786 320
rect 20072 263 20178 441
rect 20288 263 20394 441
rect 20504 263 20610 441
rect 22224 291 22320 399
rect 22357 291 22453 399
rect 22490 291 22586 399
rect 28501 268 28607 446
rect 28717 268 28823 446
rect 28933 268 29039 446
rect 31290 278 31377 390
rect 31413 278 31500 390
rect 31545 278 31632 390
rect 37319 275 37406 387
rect 37488 275 37575 387
rect 42019 258 42125 436
rect 42235 258 42341 436
rect 42451 258 42557 436
rect 46945 262 47029 420
rect 47058 262 47142 420
rect 47173 262 47257 420
rect 54268 272 54352 430
rect 54387 272 54471 430
rect 54516 272 54600 430
rect 58531 253 58637 431
rect 58747 253 58853 431
rect 58963 253 59069 431
<< metal4 >>
rect 2047 5502 2853 7801
rect 2047 5501 2363 5502
rect 2047 5323 2191 5501
rect 2297 5324 2363 5501
rect 2469 5501 2853 5502
rect 2469 5324 2537 5501
rect 2297 5323 2537 5324
rect 2643 5323 2853 5501
rect 2047 2555 2853 5323
rect 2047 2553 2398 2555
rect 2047 2375 2193 2553
rect 2299 2377 2398 2553
rect 2504 2377 2597 2555
rect 2703 2377 2853 2555
rect 2299 2375 2853 2377
rect 2047 95 2853 2375
rect 3390 7620 4196 7802
rect 3390 7619 3980 7620
rect 3390 7441 3425 7619
rect 3531 7618 3980 7619
rect 3531 7441 3634 7618
rect 3390 7440 3634 7441
rect 3740 7440 3800 7618
rect 3906 7442 3980 7618
rect 4086 7442 4196 7620
rect 3906 7440 4196 7442
rect 3390 442 4196 7440
rect 18390 5522 19196 7802
rect 18390 5344 18519 5522
rect 18625 5344 18735 5522
rect 18841 5344 18951 5522
rect 19057 5344 19196 5522
rect 3390 264 3439 442
rect 3545 264 3660 442
rect 3766 264 3869 442
rect 3975 264 4043 442
rect 4149 264 4196 442
rect 3390 96 4196 264
rect 7121 3465 7590 3580
rect 7121 3459 7330 3465
rect 7121 3368 7179 3459
rect 7265 3374 7330 3459
rect 7416 3374 7475 3465
rect 7561 3374 7590 3465
rect 7265 3368 7590 3374
rect 7121 387 7590 3368
rect 14536 2993 14890 3065
rect 14536 2924 14560 2993
rect 14637 2924 14663 2993
rect 14740 2924 14766 2993
rect 14843 2924 14890 2993
rect 14536 2864 14890 2924
rect 7121 296 7167 387
rect 7253 296 7315 387
rect 7401 296 7463 387
rect 7549 296 7590 387
rect 7121 197 7590 296
rect 14612 439 14813 2864
rect 14612 370 14686 439
rect 14763 370 14813 439
rect 14612 320 14813 370
rect 14612 251 14709 320
rect 14786 251 14813 320
rect 14612 172 14813 251
rect 18390 2571 19196 5344
rect 18390 2393 18510 2571
rect 18616 2393 18726 2571
rect 18832 2393 18942 2571
rect 19048 2393 19196 2571
rect 18390 96 19196 2393
rect 19890 7636 20696 7802
rect 19890 7458 20054 7636
rect 20160 7458 20270 7636
rect 20376 7458 20486 7636
rect 20592 7458 20696 7636
rect 19890 441 20696 7458
rect 26890 5514 27696 7802
rect 26890 5336 27027 5514
rect 27133 5336 27243 5514
rect 27349 5336 27459 5514
rect 27565 5336 27696 5514
rect 19890 263 20072 441
rect 20178 263 20288 441
rect 20394 263 20504 441
rect 20610 263 20696 441
rect 19890 96 20696 263
rect 22171 3469 22638 3594
rect 22171 3385 22219 3469
rect 22312 3385 22386 3469
rect 22479 3385 22638 3469
rect 22171 3308 22638 3385
rect 22171 3224 22219 3308
rect 22312 3224 22386 3308
rect 22479 3224 22638 3308
rect 22171 399 22638 3224
rect 22171 291 22224 399
rect 22320 291 22357 399
rect 22453 291 22490 399
rect 22586 291 22638 399
rect 22171 222 22638 291
rect 26890 2566 27696 5336
rect 26890 2388 27032 2566
rect 27138 2388 27248 2566
rect 27354 2388 27464 2566
rect 27570 2388 27696 2566
rect 26890 96 27696 2388
rect 28390 7635 29196 7802
rect 28390 7457 28546 7635
rect 28652 7457 28762 7635
rect 28868 7457 28978 7635
rect 29084 7457 29196 7635
rect 28390 446 29196 7457
rect 40390 5509 41196 7802
rect 40390 5331 40499 5509
rect 40605 5331 40715 5509
rect 40821 5331 40931 5509
rect 41037 5331 41196 5509
rect 37285 3763 37590 3920
rect 37285 3762 37475 3763
rect 37285 3650 37321 3762
rect 37408 3651 37475 3762
rect 37562 3651 37590 3763
rect 37408 3650 37590 3651
rect 28390 268 28501 446
rect 28607 268 28717 446
rect 28823 268 28933 446
rect 29039 268 29196 446
rect 28390 96 29196 268
rect 31223 3122 31648 3201
rect 31223 3010 31269 3122
rect 31356 3010 31388 3122
rect 31475 3010 31507 3122
rect 31594 3010 31648 3122
rect 31223 390 31648 3010
rect 31223 278 31290 390
rect 31377 278 31413 390
rect 31500 278 31545 390
rect 31632 278 31648 390
rect 31223 236 31648 278
rect 37285 387 37590 3650
rect 37285 275 37319 387
rect 37406 275 37488 387
rect 37575 275 37590 387
rect 37285 227 37590 275
rect 40390 2568 41196 5331
rect 40390 2390 40535 2568
rect 40641 2390 40751 2568
rect 40857 2390 40967 2568
rect 41073 2390 41196 2568
rect 40390 96 41196 2390
rect 41890 7641 42696 7802
rect 41890 7463 42074 7641
rect 42180 7463 42290 7641
rect 42396 7463 42506 7641
rect 42612 7463 42696 7641
rect 41890 436 42696 7463
rect 56890 5501 57696 7802
rect 56890 5323 57050 5501
rect 57156 5323 57266 5501
rect 57372 5323 57482 5501
rect 57588 5323 57696 5501
rect 54218 3413 54643 3436
rect 54218 3255 54262 3413
rect 54346 3255 54383 3413
rect 54467 3255 54521 3413
rect 54605 3255 54643 3413
rect 41890 258 42019 436
rect 42125 258 42235 436
rect 42341 258 42451 436
rect 42557 258 42696 436
rect 41890 96 42696 258
rect 46905 3038 47319 3127
rect 46905 3037 47083 3038
rect 46905 2879 46943 3037
rect 47027 2880 47083 3037
rect 47167 2880 47211 3038
rect 47295 2880 47319 3038
rect 47027 2879 47319 2880
rect 46905 420 47319 2879
rect 46905 262 46945 420
rect 47029 262 47058 420
rect 47142 262 47173 420
rect 47257 262 47319 420
rect 46905 174 47319 262
rect 54218 430 54643 3255
rect 54218 272 54268 430
rect 54352 272 54387 430
rect 54471 272 54516 430
rect 54600 272 54643 430
rect 54218 186 54643 272
rect 56890 2579 57696 5323
rect 56890 2401 57030 2579
rect 57136 2401 57246 2579
rect 57352 2401 57462 2579
rect 57568 2401 57696 2579
rect 56890 96 57696 2401
rect 58390 7634 59196 7802
rect 58390 7456 58559 7634
rect 58665 7456 58775 7634
rect 58881 7456 58991 7634
rect 59097 7456 59196 7634
rect 58390 431 59196 7456
rect 58390 253 58531 431
rect 58637 253 58747 431
rect 58853 253 58963 431
rect 59069 253 59196 431
rect 58390 96 59196 253
use brbufhalf  brbufhalf_0
timestamp 1654657656
transform 1 0 4459 0 1 -2298
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_1
timestamp 1654657656
transform 1 0 34661 0 1 -2298
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_2
timestamp 1654657656
transform -1 0 57337 0 -1 10198
box -3552 2527 26658 5446
use brbufhalf  brbufhalf_3
timestamp 1654657656
transform -1 0 27135 0 -1 10198
box -3552 2527 26658 5446
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1653697408
transform 1 0 30934 0 1 3801
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654402208
transform 1 0 16076 0 1 3425
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654402208
transform 1 0 14146 0 1 3425
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_2
timestamp 1654402208
transform 1 0 31482 0 1 3801
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_3
timestamp 1654402208
transform 1 0 46218 0 1 3585
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_4
timestamp 1654402208
transform 1 0 44288 0 1 3585
box -38 -48 1510 592
<< labels >>
flabel metal1 61289 1010 61511 1088 1 FreeSans 1600 0 0 0 OUT
port 3 n
flabel metal1 0 4161 254 4227 1 FreeSans 1600 0 0 0 RESET
port 68 n
flabel metal4 2047 95 2853 7801 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 3390 96 4196 7802 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 18390 96 19196 7802 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 19890 96 20696 7802 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 26890 96 27696 7802 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 28390 96 29196 7802 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 40390 96 41196 7802 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 41890 96 42696 7802 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal4 56890 96 57696 7802 1 FreeSans 1600 0 0 0 VDD
port 69 n
flabel metal4 58390 96 59196 7802 1 FreeSans 1600 0 0 0 VSS
port 70 n
flabel metal2 60825 6878 60869 8034 1 FreeSans 1600 0 0 0 C[0]
port 134 n
flabel metal2 58937 6878 58981 8034 1 FreeSans 1600 0 0 0 C[1]
port 133 n
flabel metal2 57049 6878 57093 8034 1 FreeSans 1600 0 0 0 C[2]
port 132 n
flabel metal2 55161 6878 55205 8034 1 FreeSans 1600 0 0 0 C[3]
port 131 n
flabel metal2 53273 6878 53317 8034 1 FreeSans 1600 0 0 0 C[4]
port 130 n
flabel metal2 51385 6878 51429 8034 1 FreeSans 1600 0 0 0 C[5]
port 129 n
flabel metal2 49497 6878 49541 8034 1 FreeSans 1600 0 0 0 C[6]
port 128 n
flabel metal2 47609 6878 47653 8034 1 FreeSans 1600 0 0 0 C[7]
port 127 n
flabel metal2 45721 6878 45765 8034 1 FreeSans 1600 0 0 0 C[8]
port 126 n
flabel metal2 43833 6878 43877 8034 1 FreeSans 1600 0 0 0 C[9]
port 125 n
flabel metal2 41945 6878 41989 8034 1 FreeSans 1600 0 0 0 C[10]
port 124 n
flabel metal2 40057 6878 40101 8034 1 FreeSans 1600 0 0 0 C[11]
port 123 n
flabel metal2 38169 6878 38213 8034 1 FreeSans 1600 0 0 0 C[12]
port 122 n
flabel metal2 36281 6878 36325 8034 1 FreeSans 1600 0 0 0 C[13]
port 121 n
flabel metal2 34393 6878 34437 8034 1 FreeSans 1600 0 0 0 C[14]
port 120 n
flabel metal2 32505 6878 32549 8034 1 FreeSans 1600 0 0 0 C[15]
port 119 n
flabel metal2 30617 6878 30661 8034 1 FreeSans 1600 0 0 0 C[16]
port 118 n
flabel metal2 26841 6878 26885 8034 1 FreeSans 1600 0 0 0 C[18]
port 116 n
flabel metal2 24953 6878 24997 8034 1 FreeSans 1600 0 0 0 C[19]
port 115 n
flabel metal2 23065 6878 23109 8034 1 FreeSans 1600 0 0 0 C[20]
port 114 n
flabel metal2 21177 6878 21221 8034 1 FreeSans 1600 0 0 0 C[21]
port 113 n
flabel metal2 19289 6878 19333 8034 1 FreeSans 1600 0 0 0 C[22]
port 112 n
flabel metal2 17401 6878 17445 8034 1 FreeSans 1600 0 0 0 C[23]
port 111 n
flabel metal2 15513 6878 15557 8034 1 FreeSans 1600 0 0 0 C[24]
port 110 n
flabel metal2 13625 6878 13669 8034 1 FreeSans 1600 0 0 0 C[25]
port 109 n
flabel metal2 11737 6878 11781 8034 1 FreeSans 1600 0 0 0 C[26]
port 108 n
flabel metal2 9849 6878 9893 8034 1 FreeSans 1600 0 0 0 C[27]
port 107 n
flabel metal2 7961 6878 8005 8034 1 FreeSans 1600 0 0 0 C[28]
port 106 n
flabel metal2 6073 6878 6117 8034 1 FreeSans 1600 0 0 0 C[29]
port 105 n
flabel metal2 4185 6878 4229 8034 1 FreeSans 1600 0 0 0 C[30]
port 104 n
flabel metal2 2297 6878 2341 8034 1 FreeSans 1600 0 0 0 C[31]
port 103 n
flabel metal2 927 124 971 1022 1 FreeSans 1600 0 0 0 C[32]
port 102 n
flabel metal2 2815 124 2859 1022 1 FreeSans 1600 0 0 0 C[33]
port 101 n
flabel metal2 4703 124 4747 1022 1 FreeSans 1600 0 0 0 C[34]
port 100 n
flabel metal2 6591 124 6635 1022 1 FreeSans 1600 0 0 0 C[35]
port 99 n
flabel metal2 8479 124 8523 1022 1 FreeSans 1600 0 0 0 C[36]
port 98 n
flabel metal2 10367 124 10411 1022 1 FreeSans 1600 0 0 0 C[37]
port 97 n
flabel metal2 12255 124 12299 1022 1 FreeSans 1600 0 0 0 C[38]
port 96 n
flabel metal2 14143 124 14187 1022 1 FreeSans 1600 0 0 0 C[39]
port 95 n
flabel metal2 16031 124 16075 1022 1 FreeSans 1600 0 0 0 C[40]
port 94 n
flabel metal2 17919 124 17963 1022 1 FreeSans 1600 0 0 0 C[41]
port 93 n
flabel metal2 19807 124 19851 1022 1 FreeSans 1600 0 0 0 C[42]
port 92 n
flabel metal2 21695 124 21739 1022 1 FreeSans 1600 0 0 0 C[43]
port 91 n
flabel metal2 23583 124 23627 1022 1 FreeSans 1600 0 0 0 C[44]
port 90 n
flabel metal2 29247 124 29291 1022 1 FreeSans 1600 0 0 0 C[47]
port 87 n
flabel metal2 31135 124 31179 1022 1 FreeSans 1600 0 0 0 C[48]
port 86 n
flabel metal2 33023 124 33067 1022 1 FreeSans 1600 0 0 0 C[49]
port 85 n
flabel metal2 34911 124 34955 1022 1 FreeSans 1600 0 0 0 C[50]
port 84 n
flabel metal2 36799 124 36843 1022 1 FreeSans 1600 0 0 0 C[51]
port 83 n
flabel metal2 38687 124 38731 1022 1 FreeSans 1600 0 0 0 C[52]
port 82 n
flabel metal2 42463 124 42507 1022 1 FreeSans 1600 0 0 0 C[54]
port 80 n
flabel metal2 44351 124 44395 1022 1 FreeSans 1600 0 0 0 C[55]
port 79 n
flabel metal2 46239 124 46283 1022 1 FreeSans 1600 0 0 0 C[56]
port 78 n
flabel metal2 48127 124 48171 1022 1 FreeSans 1600 0 0 0 C[57]
port 77 n
flabel metal2 50015 124 50059 1022 1 FreeSans 1600 0 0 0 C[58]
port 76 n
flabel metal2 51903 124 51947 1022 1 FreeSans 1600 0 0 0 C[59]
port 75 n
flabel metal2 53791 124 53835 1022 1 FreeSans 1600 0 0 0 C[60]
port 74 n
flabel metal2 55679 124 55723 1022 1 FreeSans 1600 0 0 0 C[61]
port 73 n
flabel metal2 59455 124 59499 1022 1 FreeSans 1600 0 0 0 C[63]
port 71 n
flabel metal2 25471 124 25515 1022 1 FreeSans 1600 0 0 0 C[45]
port 89 n
flabel metal2 28729 6878 28773 8034 1 FreeSans 1600 0 0 0 C[17]
port 117 n
flabel metal2 27359 24 27403 922 1 FreeSans 1600 0 0 0 C[46]
port 135 n
flabel metal2 40575 0 40619 898 1 FreeSans 1600 0 0 0 C[53]
port 136 n
flabel metal2 57569 4 57613 902 1 FreeSans 1600 0 0 0 C[62]
port 137 n
<< end >>
