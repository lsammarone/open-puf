magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect 25 4633 324 4865
rect 376 4576 1284 4770
rect 5946 4576 6819 4670
rect 12433 241 12603 4576
<< pdiff >>
rect 6858 6772 12565 6784
rect 3004 5002 3020 5318
rect 4208 5002 4226 5318
rect 3004 4976 3008 5002
rect 2970 4738 3008 4976
rect 4228 4738 4260 4976
<< poly >>
rect 13335 4597 13469 4613
rect 13335 4563 13351 4597
rect 13385 4563 13419 4597
rect 13453 4563 13469 4597
rect 13335 4547 13469 4563
rect 13335 4479 13455 4547
<< polycont >>
rect 13351 4563 13385 4597
rect 13419 4563 13453 4597
<< locali >>
rect 1508 6962 1546 6996
rect 13332 4597 13901 4644
rect 13332 4563 13351 4597
rect 13385 4563 13419 4597
rect 13453 4563 13901 4597
rect 271 4054 305 4100
rect 271 3974 305 4020
rect 271 3893 305 3940
rect 271 3812 305 3859
rect 13847 3585 13901 4563
rect 12366 1420 12400 1458
rect 12366 1348 12400 1386
rect 12700 1044 12734 1087
rect 12700 967 12734 1010
rect 12700 889 12734 933
rect 12700 811 12734 855
rect 12700 733 12734 777
<< viali >>
rect 1474 6962 1508 6996
rect 1546 6962 1580 6996
rect 271 4100 305 4134
rect 271 4020 305 4054
rect 271 3940 305 3974
rect 271 3859 305 3893
rect 271 3778 305 3812
rect 12366 1458 12400 1492
rect 12366 1386 12400 1420
rect 12366 1314 12400 1348
rect 12700 1087 12734 1121
rect 12700 1010 12734 1044
rect 12700 933 12734 967
rect 12700 855 12734 889
rect 12700 777 12734 811
rect 12700 699 12734 733
<< metal1 >>
rect 1462 6953 1468 7005
rect 1520 6953 1534 7005
rect 1586 6953 1592 7005
rect 5095 6957 5128 6995
rect 5854 6502 5967 6850
rect 7271 6574 7277 6626
rect 7329 6574 7341 6626
rect 7393 6574 9428 6626
rect 9480 6574 9492 6626
rect 9544 6574 9550 6626
rect 14736 6434 14788 6440
rect 14854 6410 14989 6527
rect 14736 6370 14788 6382
rect 14736 6298 14788 6318
tri 14736 6297 14737 6298 ne
rect 14737 6297 14788 6298
tri 14788 6297 14803 6312 sw
tri 14737 6247 14787 6297 ne
rect 14787 6247 14803 6297
tri 14787 6231 14803 6247 ne
tri 14803 6231 14869 6297 sw
tri 14803 6211 14823 6231 ne
rect 14823 6141 14869 6231
rect 14824 6126 14868 6141
rect 288 5857 328 6059
rect 13102 5787 13142 5989
rect 13170 5809 13337 5965
tri 6699 5642 6713 5656 ne
rect 6713 5642 6735 5656
rect -370 5625 -318 5642
tri 6713 5631 6724 5642 ne
rect 6724 5631 6735 5642
tri 6724 5620 6735 5631 ne
tri 6831 5622 6865 5656 nw
rect 11679 5626 11685 5678
rect 11737 5626 11749 5678
rect 11801 5626 12949 5678
rect 13001 5626 13013 5678
rect 13065 5626 13071 5678
rect 13425 5630 13492 5674
rect -370 5561 -318 5573
rect 6870 5546 6876 5598
rect 6928 5546 6940 5598
rect 6992 5546 12200 5598
rect 12252 5546 12264 5598
rect 12316 5546 12322 5598
rect -370 5503 -318 5509
rect -18 5498 34 5504
rect -194 5492 -142 5498
rect -194 5406 -142 5440
tri 7432 5466 7449 5483 se
rect 7449 5480 8435 5483
tri 8435 5480 8438 5483 sw
rect 7449 5466 8438 5480
tri 8438 5466 8452 5480 sw
rect -18 5426 34 5446
tri 7395 5429 7432 5466 se
rect 7432 5445 8452 5466
rect 7432 5429 7449 5445
tri 7449 5429 7465 5445 nw
tri 8419 5429 8435 5445 ne
rect 8435 5429 8452 5445
tri 7378 5412 7395 5429 se
rect 7395 5412 7432 5429
tri 7432 5412 7449 5429 nw
tri 8435 5412 8452 5429 ne
tri 8452 5428 8490 5466 sw
rect 9422 5428 9428 5480
rect 9480 5428 9492 5480
rect 9544 5428 11573 5480
rect 11625 5428 11637 5480
rect 11689 5428 11695 5480
rect 12073 5443 12079 5495
rect 12131 5443 12143 5495
rect 12195 5443 12990 5495
tri 12910 5428 12925 5443 ne
rect 12925 5428 12990 5443
rect 8452 5412 8490 5428
tri 8490 5412 8506 5428 sw
tri 12925 5412 12941 5428 ne
rect 12941 5412 12990 5428
tri 7341 5375 7378 5412 se
rect 7378 5375 7395 5412
tri 7395 5375 7432 5412 nw
tri 8452 5375 8489 5412 ne
rect 8489 5409 8506 5412
tri 8506 5409 8509 5412 sw
tri 12941 5409 12944 5412 ne
rect 8489 5398 8509 5409
tri 8509 5398 8520 5409 sw
rect 8489 5375 8520 5398
rect -18 5368 34 5374
tri 7334 5368 7341 5375 se
rect 7341 5368 7378 5375
tri 7324 5358 7334 5368 se
rect 7334 5358 7378 5368
tri 7378 5358 7395 5375 nw
tri 8489 5358 8506 5375 ne
rect 8506 5368 8520 5375
tri 8520 5368 8550 5398 sw
rect 8506 5358 8550 5368
tri 8550 5358 8560 5368 sw
rect -194 5348 -142 5354
tri 7314 5348 7324 5358 se
rect 7324 5348 7341 5358
tri 7298 5332 7314 5348 se
rect 7314 5332 7341 5348
rect 715 5280 721 5332
rect 773 5280 785 5332
rect 837 5326 847 5332
tri 847 5326 853 5332 sw
tri 7292 5326 7298 5332 se
rect 7298 5326 7341 5332
rect 837 5280 6876 5326
rect 715 5274 6876 5280
rect 6928 5274 6940 5326
rect 6992 5274 6998 5326
tri 7287 5321 7292 5326 se
rect 7292 5321 7341 5326
tri 7341 5321 7378 5358 nw
tri 8506 5321 8543 5358 ne
rect 8543 5348 8560 5358
tri 8560 5348 8570 5358 sw
rect 8543 5346 8570 5348
tri 8570 5346 8572 5348 sw
rect 12194 5346 12200 5398
rect 12252 5346 12264 5398
rect 12316 5346 12863 5398
rect 8543 5332 8572 5346
tri 8572 5332 8586 5346 sw
tri 12777 5332 12791 5346 ne
rect 12791 5332 12863 5346
rect 8543 5326 8586 5332
tri 8586 5326 8592 5332 sw
tri 12791 5326 12797 5332 ne
rect 12797 5326 12863 5332
rect 8543 5321 8592 5326
tri 7270 5304 7287 5321 se
rect 7287 5304 7324 5321
tri 7324 5304 7341 5321 nw
tri 8543 5304 8560 5321 ne
rect 8560 5318 8592 5321
tri 8592 5318 8600 5326 sw
tri 12797 5318 12805 5326 ne
rect 12805 5318 12863 5326
rect 8560 5312 8600 5318
tri 8600 5312 8606 5318 sw
tri 9429 5312 9435 5318 se
rect 9435 5312 9441 5318
rect 8560 5304 8606 5312
tri 8606 5304 8614 5312 sw
tri 9421 5304 9429 5312 se
rect 9429 5304 9441 5312
tri 7240 5274 7270 5304 se
rect 7270 5274 7287 5304
tri 7233 5267 7240 5274 se
rect 7240 5267 7287 5274
tri 7287 5267 7324 5304 nw
tri 8560 5267 8597 5304 ne
rect 8597 5267 9441 5304
tri 7211 5245 7233 5267 se
rect 7233 5245 7265 5267
tri 7265 5245 7287 5267 nw
tri 8597 5266 8598 5267 ne
rect 8598 5266 9441 5267
rect 9493 5266 9505 5318
rect 9557 5266 9563 5318
tri 12805 5312 12811 5318 ne
rect 12811 5305 12863 5318
rect 12944 5351 12990 5412
tri 12990 5351 13024 5385 sw
tri 12863 5305 12869 5311 sw
rect 12944 5305 13136 5351
tri 13705 5305 13711 5311 se
rect 12811 5277 12869 5305
tri 12869 5277 12897 5305 sw
tri 13677 5277 13705 5305 se
rect 13705 5277 13711 5305
rect 14478 5304 14522 5348
rect 15042 5345 15116 5380
rect 5228 5239 7244 5245
rect 5280 5224 7244 5239
tri 7244 5224 7265 5245 nw
rect 5280 5207 7227 5224
tri 7227 5207 7244 5224 nw
rect 7411 5218 7463 5224
rect 12811 5219 13711 5277
rect 5228 5175 5280 5187
tri 5280 5134 5353 5207 nw
rect 7411 5154 7463 5166
rect 5228 5117 5280 5123
tri 7463 5148 7497 5182 sw
rect 7463 5102 8333 5148
rect 7411 5096 8333 5102
rect -12 4743 328 4945
rect 524 4938 564 5068
rect 12900 4938 12940 5068
rect 13335 4987 13341 4991
rect 13251 4939 13341 4987
rect 13393 4939 13413 4991
rect 13465 4939 13484 4991
rect 13536 4939 13555 4991
rect 13607 4939 13626 4991
rect 13678 4939 13684 4991
rect 13251 4916 13684 4939
rect 288 4708 328 4743
rect 823 4858 829 4910
rect 881 4858 894 4910
rect 946 4858 959 4910
rect 1011 4858 1024 4910
rect 1076 4858 1089 4910
rect 1141 4858 1153 4910
rect 1205 4858 1217 4910
rect 1269 4858 1281 4910
rect 1333 4858 1345 4910
rect 1397 4858 1409 4910
rect 1461 4858 1473 4910
rect 1525 4858 1531 4910
rect 823 4835 1531 4858
rect 823 4783 829 4835
rect 881 4783 894 4835
rect 946 4783 959 4835
rect 1011 4783 1024 4835
rect 1076 4783 1089 4835
rect 1141 4783 1153 4835
rect 1205 4783 1217 4835
rect 1269 4783 1281 4835
rect 1333 4783 1345 4835
rect 1397 4783 1409 4835
rect 1461 4783 1473 4835
rect 1525 4783 1531 4835
rect 823 4760 1531 4783
rect 823 4708 829 4760
rect 881 4708 894 4760
rect 946 4708 959 4760
rect 1011 4708 1024 4760
rect 1076 4708 1089 4760
rect 1141 4708 1153 4760
rect 1205 4708 1217 4760
rect 1269 4708 1281 4760
rect 1333 4708 1345 4760
rect 1397 4708 1409 4760
rect 1461 4708 1473 4760
rect 1525 4708 1531 4760
rect 12991 4708 13031 4910
rect 13251 4864 13341 4916
rect 13393 4864 13413 4916
rect 13465 4864 13484 4916
rect 13536 4864 13555 4916
rect 13607 4864 13626 4916
rect 13678 4864 13684 4916
rect 13251 4841 13684 4864
rect 13251 4812 13341 4841
rect 13335 4789 13341 4812
rect 13393 4789 13413 4841
rect 13465 4789 13484 4841
rect 13536 4789 13555 4841
rect 13607 4789 13626 4841
rect 13678 4789 13684 4841
rect 9930 4626 9936 4678
rect 9988 4626 10000 4678
rect 10052 4626 10190 4678
rect 10242 4626 10254 4678
rect 10306 4626 10312 4678
rect 11615 4544 11621 4596
rect 11673 4544 11685 4596
rect 11737 4585 12071 4596
tri 12071 4585 12082 4596 sw
rect 12153 4585 12159 4637
rect 12211 4585 12224 4637
rect 12276 4585 14690 4637
rect 14742 4585 14754 4637
rect 14806 4585 14812 4637
rect 11737 4557 12082 4585
tri 12082 4557 12110 4585 sw
rect 11737 4544 14591 4557
tri 12049 4505 12088 4544 ne
rect 12088 4505 14591 4544
rect 14643 4505 14655 4557
rect 14707 4505 14713 4557
tri 323 4338 327 4342 se
rect 327 4338 4286 4342
tri 4286 4338 4290 4342 sw
tri 253 4268 323 4338 se
rect 323 4290 4290 4338
rect 323 4268 327 4290
tri 327 4268 349 4290 nw
tri 4264 4268 4286 4290 ne
rect 4286 4268 4290 4290
tri 249 4264 253 4268 se
rect 253 4264 323 4268
tri 323 4264 327 4268 nw
tri 4286 4264 4290 4268 ne
tri 4290 4264 4364 4338 sw
tri 231 4246 249 4264 se
rect 249 4246 305 4264
tri 305 4246 323 4264 nw
tri 4290 4246 4308 4264 ne
rect 4308 4246 5178 4264
rect 92 4200 259 4246
tri 259 4200 305 4246 nw
tri 4308 4212 4342 4246 ne
rect 4342 4212 5178 4246
rect 5230 4212 5242 4264
rect 5294 4212 5301 4264
rect 14840 4258 15007 4414
rect 238 4140 311 4146
rect 290 4134 311 4140
rect 305 4100 311 4134
rect 290 4088 311 4100
rect 238 4061 311 4088
rect 290 4054 311 4061
rect 305 4020 311 4054
rect 290 4009 311 4020
rect 238 3982 311 4009
rect 290 3979 311 3982
tri 311 3979 324 3992 sw
rect 470 3979 512 4181
rect 1698 4129 1704 4181
rect 1756 4129 1773 4181
rect 1825 4129 1842 4181
rect 1894 4129 1911 4181
rect 1963 4129 1980 4181
rect 2032 4129 2038 4181
rect 1698 4106 2038 4129
rect 1698 4054 1704 4106
rect 1756 4054 1773 4106
rect 1825 4054 1842 4106
rect 1894 4054 1911 4106
rect 1963 4054 1980 4106
rect 2032 4054 2038 4106
rect 1698 4031 2038 4054
rect 1698 3979 1704 4031
rect 1756 3979 1773 4031
rect 1825 3979 1842 4031
rect 1894 3979 1911 4031
rect 1963 3979 1980 4031
rect 2032 3979 2038 4031
rect 3150 4129 3156 4181
rect 3208 4129 3220 4181
rect 3272 4129 3284 4181
rect 3336 4129 3348 4181
rect 3400 4129 3412 4181
rect 3464 4129 3476 4181
rect 3528 4129 3540 4181
rect 3592 4129 3598 4181
rect 3150 4106 3598 4129
rect 3150 4054 3156 4106
rect 3208 4054 3220 4106
rect 3272 4054 3284 4106
rect 3336 4054 3348 4106
rect 3400 4054 3412 4106
rect 3464 4054 3476 4106
rect 3528 4054 3540 4106
rect 3592 4054 3598 4106
rect 3150 4031 3598 4054
rect 3150 3979 3156 4031
rect 3208 3979 3220 4031
rect 3272 3979 3284 4031
rect 3336 3979 3348 4031
rect 3400 3979 3412 4031
rect 3464 3979 3476 4031
rect 3528 3979 3540 4031
rect 3592 3979 3598 4031
rect 9029 3979 9071 4181
rect 290 3974 324 3979
rect 305 3951 324 3974
tri 324 3951 352 3979 sw
rect 305 3940 352 3951
rect 290 3934 352 3940
tri 352 3934 369 3951 sw
rect 290 3930 1248 3934
rect 238 3923 1248 3930
rect 238 3903 829 3923
rect 290 3893 829 3903
rect 305 3871 829 3893
rect 881 3871 902 3923
rect 954 3871 974 3923
rect 1026 3871 1046 3923
rect 1098 3871 1118 3923
rect 1170 3871 1190 3923
rect 1242 3871 1248 3923
rect 8031 3899 8037 3951
rect 8089 3899 8101 3951
rect 8153 3945 10053 3951
rect 8153 3923 10001 3945
rect 8153 3899 8522 3923
tri 8522 3899 8546 3923 nw
tri 9528 3899 9552 3923 ne
rect 9552 3899 10001 3923
tri 9552 3879 9572 3899 ne
rect 9572 3893 10001 3899
rect 9572 3881 10053 3893
rect 9572 3879 10001 3881
rect 305 3861 1248 3871
tri 9945 3861 9963 3879 ne
rect 9963 3861 10001 3879
rect 305 3859 343 3861
rect 290 3851 343 3859
rect 238 3824 343 3851
rect 290 3823 343 3824
tri 343 3823 381 3861 nw
tri 9963 3823 10001 3861 ne
rect 10001 3823 10053 3829
rect 290 3812 311 3823
rect 305 3778 311 3812
tri 311 3791 343 3823 nw
rect 290 3772 311 3778
rect 238 3766 311 3772
tri 12928 3710 12931 3713 se
rect 12931 3710 12965 3713
tri 12873 3655 12928 3710 se
rect 12928 3655 12965 3710
rect 13337 3704 13683 3710
rect 941 3654 1531 3655
rect 941 3602 947 3654
rect 999 3602 1013 3654
rect 1065 3602 1079 3654
rect 1131 3602 1145 3654
rect 1197 3602 1211 3654
rect 1263 3602 1277 3654
rect 1329 3602 1343 3654
rect 1395 3602 1408 3654
rect 1460 3602 1473 3654
rect 1525 3602 1531 3654
rect 941 3580 1531 3602
rect 941 3528 947 3580
rect 999 3528 1013 3580
rect 1065 3528 1079 3580
rect 1131 3528 1145 3580
rect 1197 3528 1211 3580
rect 1263 3528 1277 3580
rect 1329 3528 1343 3580
rect 1395 3528 1408 3580
rect 1460 3528 1473 3580
rect 1525 3528 1531 3580
rect 941 3506 1531 3528
rect 941 3454 947 3506
rect 999 3454 1013 3506
rect 1065 3454 1079 3506
rect 1131 3454 1145 3506
rect 1197 3454 1211 3506
rect 1263 3454 1277 3506
rect 1329 3454 1343 3506
rect 1395 3454 1408 3506
rect 1460 3454 1473 3506
rect 1525 3454 1531 3506
rect 12634 3566 13026 3655
rect 13337 3652 13338 3704
rect 13390 3652 13411 3704
rect 13463 3652 13484 3704
rect 13536 3652 13557 3704
rect 13609 3652 13630 3704
rect 13682 3652 13683 3704
rect 13337 3638 13683 3652
rect 13337 3586 13338 3638
rect 13390 3586 13411 3638
rect 13463 3586 13484 3638
rect 13536 3586 13557 3638
rect 13609 3586 13630 3638
rect 13682 3586 13683 3638
rect 13337 3572 13683 3586
rect 12634 3560 13216 3566
rect 12634 3508 12887 3560
rect 12939 3508 12956 3560
rect 13008 3508 13025 3560
rect 13077 3508 13094 3560
rect 13146 3508 13163 3560
rect 13215 3508 13216 3560
rect 12634 3490 13216 3508
rect 12634 3456 12887 3490
rect 941 3453 1531 3454
tri 12544 3453 12547 3456 ne
rect 12547 3453 12887 3456
tri 12547 3311 12689 3453 ne
rect 12689 3355 12749 3453
rect 12689 3311 12743 3355
tri 12743 3349 12749 3355 ne
rect 12886 3438 12887 3453
rect 12939 3438 12956 3490
rect 13008 3438 13025 3490
rect 13077 3438 13094 3490
rect 13146 3438 13163 3490
rect 13215 3438 13216 3490
rect 12886 3420 13216 3438
rect 12886 3368 12887 3420
rect 12939 3368 12956 3420
rect 13008 3368 13025 3420
rect 13077 3368 13094 3420
rect 13146 3368 13163 3420
rect 13215 3368 13216 3420
rect 12886 3349 13216 3368
rect 12886 3297 12887 3349
rect 12939 3297 12956 3349
rect 13008 3297 13025 3349
rect 13077 3297 13094 3349
rect 13146 3297 13163 3349
rect 13215 3297 13216 3349
rect 2367 3240 2373 3292
rect 2425 3240 2437 3292
rect 2489 3240 7005 3292
rect 7057 3240 7069 3292
rect 7121 3240 7127 3292
rect 12886 3278 13216 3297
rect 12886 3226 12887 3278
rect 12939 3226 12956 3278
rect 13008 3226 13025 3278
rect 13077 3226 13094 3278
rect 13146 3226 13163 3278
rect 13215 3226 13216 3278
rect 12886 3220 13216 3226
rect 13337 3520 13338 3572
rect 13390 3520 13411 3572
rect 13463 3520 13484 3572
rect 13536 3520 13557 3572
rect 13609 3520 13630 3572
rect 13682 3520 13683 3572
rect 13337 3506 13683 3520
rect 13337 3454 13338 3506
rect 13390 3454 13411 3506
rect 13463 3454 13484 3506
rect 13536 3454 13557 3506
rect 13609 3454 13630 3506
rect 13682 3454 13683 3506
rect 13337 3440 13683 3454
rect 13337 3388 13338 3440
rect 13390 3388 13411 3440
rect 13463 3388 13484 3440
rect 13536 3388 13557 3440
rect 13609 3388 13630 3440
rect 13682 3388 13683 3440
rect 13337 3374 13683 3388
rect 13337 3322 13338 3374
rect 13390 3322 13411 3374
rect 13463 3322 13484 3374
rect 13536 3322 13557 3374
rect 13609 3322 13630 3374
rect 13682 3322 13683 3374
rect 13337 3308 13683 3322
rect 13337 3256 13338 3308
rect 13390 3256 13411 3308
rect 13463 3256 13484 3308
rect 13536 3256 13557 3308
rect 13609 3256 13630 3308
rect 13682 3256 13683 3308
rect 13337 3242 13683 3256
rect 14697 3248 15008 3480
rect 13337 3190 13338 3242
rect 13390 3190 13411 3242
rect 13463 3190 13484 3242
rect 13536 3190 13557 3242
rect 13609 3190 13630 3242
rect 13682 3190 13683 3242
rect 13337 3176 13683 3190
rect 238 3126 290 3132
rect 13337 3124 13338 3176
rect 13390 3124 13411 3176
rect 13463 3124 13484 3176
rect 13536 3124 13557 3176
rect 13609 3124 13630 3176
rect 13682 3124 13683 3176
rect 13337 3118 13683 3124
rect 238 3054 290 3074
rect 238 2982 290 3002
rect 238 2909 290 2930
rect 1264 2928 1306 3058
rect 1698 3005 1704 3057
rect 1756 3005 1773 3057
rect 1825 3005 1842 3057
rect 1894 3005 1911 3057
rect 1963 3005 1980 3057
rect 2032 3005 2038 3057
rect 1698 2981 2038 3005
rect 1698 2929 1704 2981
rect 1756 2929 1773 2981
rect 1825 2929 1842 2981
rect 1894 2929 1911 2981
rect 1963 2929 1980 2981
rect 2032 2929 2038 2981
rect 3150 3005 3156 3057
rect 3208 3005 3220 3057
rect 3272 3005 3284 3057
rect 3336 3005 3348 3057
rect 3400 3005 3412 3057
rect 3464 3005 3476 3057
rect 3528 3005 3540 3057
rect 3592 3005 3598 3057
rect 3150 2981 3598 3005
rect 3150 2929 3156 2981
rect 3208 2929 3220 2981
rect 3272 2929 3284 2981
rect 3336 2929 3348 2981
rect 3400 2929 3412 2981
rect 3464 2929 3476 2981
rect 3528 2929 3540 2981
rect 3592 2929 3598 2981
rect 12123 2928 12182 3058
rect 238 2836 290 2857
rect 10167 2848 10173 2900
rect 10225 2848 10237 2900
rect 10289 2894 12125 2900
rect 10289 2854 12073 2894
rect 10289 2848 10295 2854
tri 10295 2848 10301 2854 nw
tri 12039 2848 12045 2854 ne
rect 12045 2848 12073 2854
tri 12045 2820 12073 2848 ne
rect 12073 2830 12125 2842
rect 238 2763 290 2784
rect 12073 2772 12125 2778
rect 238 2690 290 2711
rect 238 2617 290 2638
rect 238 2559 290 2565
rect 11863 2475 11928 2502
rect 1264 2312 1306 2442
rect 1698 2390 1704 2442
rect 1756 2390 1773 2442
rect 1825 2390 1842 2442
rect 1894 2390 1911 2442
rect 1963 2390 1980 2442
rect 2032 2390 2038 2442
rect 1698 2364 2038 2390
rect 1698 2312 1704 2364
rect 1756 2312 1773 2364
rect 1825 2312 1842 2364
rect 1894 2312 1911 2364
rect 1963 2312 1980 2364
rect 2032 2312 2038 2364
rect 3150 2390 3156 2442
rect 3208 2390 3220 2442
rect 3272 2390 3284 2442
rect 3336 2390 3348 2442
rect 3400 2390 3412 2442
rect 3464 2390 3476 2442
rect 3528 2390 3540 2442
rect 3592 2390 3598 2442
rect 3150 2364 3598 2390
rect 3150 2312 3156 2364
rect 3208 2312 3220 2364
rect 3272 2312 3284 2364
rect 3336 2312 3348 2364
rect 3400 2312 3412 2364
rect 3464 2312 3476 2364
rect 3528 2312 3540 2364
rect 3592 2312 3598 2364
rect 12258 2312 12300 2442
rect 14840 2226 15007 2382
rect 951 1828 993 2030
rect 1698 2029 2038 2030
rect 1698 1977 1704 2029
rect 1756 1977 1773 2029
rect 1825 1977 1842 2029
rect 1894 1977 1911 2029
rect 1963 1977 1980 2029
rect 2032 1977 2038 2029
rect 1698 1955 2038 1977
rect 1698 1903 1704 1955
rect 1756 1903 1773 1955
rect 1825 1903 1842 1955
rect 1894 1903 1911 1955
rect 1963 1903 1980 1955
rect 2032 1903 2038 1955
rect 1698 1881 2038 1903
rect 1698 1829 1704 1881
rect 1756 1829 1773 1881
rect 1825 1829 1842 1881
rect 1894 1829 1911 1881
rect 1963 1829 1980 1881
rect 2032 1829 2038 1881
rect 1698 1828 2038 1829
rect 3150 2029 3598 2030
rect 3150 1977 3156 2029
rect 3208 1977 3220 2029
rect 3272 1977 3284 2029
rect 3336 1977 3348 2029
rect 3400 1977 3412 2029
rect 3464 1977 3476 2029
rect 3528 1977 3540 2029
rect 3592 1977 3598 2029
rect 3150 1955 3598 1977
rect 3150 1903 3156 1955
rect 3208 1903 3220 1955
rect 3272 1903 3284 1955
rect 3336 1903 3348 1955
rect 3400 1903 3412 1955
rect 3464 1903 3476 1955
rect 3528 1903 3540 1955
rect 3592 1903 3598 1955
rect 3150 1881 3598 1903
rect 3150 1829 3156 1881
rect 3208 1829 3220 1881
rect 3272 1829 3284 1881
rect 3336 1829 3348 1881
rect 3400 1829 3412 1881
rect 3464 1829 3476 1881
rect 3528 1829 3540 1881
rect 3592 1829 3598 1881
rect 3150 1828 3598 1829
rect 12158 1828 12200 2030
rect 8535 1772 12799 1800
rect 8535 1758 8685 1772
tri 8685 1758 8699 1772 nw
tri 12779 1758 12793 1772 ne
rect 12793 1758 12799 1772
tri 12799 1758 12841 1800 sw
rect 8535 1726 8665 1758
tri 8665 1738 8685 1758 nw
tri 12793 1752 12799 1758 ne
rect 12799 1752 12841 1758
tri 12799 1738 12813 1752 ne
rect 706 1654 758 1660
tri 672 1578 706 1612 se
tri 758 1606 764 1612 sw
rect 7828 1606 7997 1658
rect 8049 1606 8061 1658
rect 8113 1606 8119 1658
rect 758 1602 764 1606
rect 706 1590 764 1602
rect 758 1578 764 1590
tri 764 1578 792 1606 sw
rect 706 1532 758 1538
rect 288 1302 330 1504
rect 986 1503 1531 1504
rect 986 1451 992 1503
rect 1044 1451 1061 1503
rect 1113 1451 1130 1503
rect 1182 1451 1199 1503
rect 1251 1451 1268 1503
rect 1320 1451 1337 1503
rect 1389 1451 1405 1503
rect 1457 1451 1473 1503
rect 1525 1451 1531 1503
rect 986 1429 1531 1451
rect 986 1377 992 1429
rect 1044 1377 1061 1429
rect 1113 1377 1130 1429
rect 1182 1377 1199 1429
rect 1251 1377 1268 1429
rect 1320 1377 1337 1429
rect 1389 1377 1405 1429
rect 1457 1377 1473 1429
rect 1525 1377 1531 1429
rect 986 1355 1531 1377
rect 986 1303 992 1355
rect 1044 1303 1061 1355
rect 1113 1303 1130 1355
rect 1182 1303 1199 1355
rect 1251 1303 1268 1355
rect 1320 1303 1337 1355
rect 1389 1303 1405 1355
rect 1457 1303 1473 1355
rect 1525 1303 1531 1355
rect 986 1302 1531 1303
rect 12360 1492 12406 1504
rect 12360 1458 12366 1492
rect 12400 1458 12406 1492
rect 12360 1420 12406 1458
rect 12360 1386 12366 1420
rect 12400 1386 12406 1420
rect 12360 1348 12406 1386
rect 12360 1314 12366 1348
rect 12400 1314 12406 1348
rect 12626 1489 12676 1504
tri 12676 1489 12691 1504 sw
rect 12813 1496 12841 1752
tri 12813 1489 12820 1496 ne
rect 12820 1489 12841 1496
tri 12841 1489 12875 1523 sw
tri 14792 1489 14826 1523 se
rect 12626 1468 12691 1489
tri 12691 1468 12712 1489 sw
tri 12820 1468 12841 1489 ne
rect 12841 1468 14872 1489
rect 12626 1461 12712 1468
tri 12712 1461 12719 1468 sw
tri 12841 1461 12848 1468 ne
rect 12848 1461 14872 1468
rect 12626 1423 12719 1461
tri 12719 1423 12757 1461 sw
rect 12626 1322 12817 1423
rect 12360 1302 12406 1314
tri 12579 1302 12599 1322 ne
rect 12599 1302 12817 1322
tri 12599 1274 12627 1302 ne
rect 12627 1274 12817 1302
rect 6054 1228 6094 1274
rect 6190 1228 6231 1274
tri 12627 1237 12664 1274 ne
rect 12664 1237 12817 1274
tri 12287 1228 12296 1237 sw
tri 12664 1228 12673 1237 ne
rect 12673 1228 12817 1237
rect 12287 1203 12296 1228
tri 12296 1203 12321 1228 sw
tri 12673 1203 12698 1228 ne
rect 12698 1203 12817 1228
rect 7956 1148 7996 1194
rect 12287 1179 12499 1203
tri 12499 1179 12523 1203 sw
tri 12698 1179 12722 1203 ne
rect 12722 1179 12817 1203
rect 12287 1151 12523 1179
rect 12287 1148 12304 1151
tri 12304 1148 12307 1151 nw
tri 12477 1148 12480 1151 ne
rect 12480 1148 12523 1151
tri 12287 1131 12304 1148 nw
tri 12480 1131 12497 1148 ne
rect 12497 1131 12523 1148
tri 12497 1121 12507 1131 ne
rect 12507 1121 12523 1131
tri 12523 1121 12581 1179 sw
tri 12722 1133 12768 1179 ne
rect 12768 1133 12817 1179
rect 12694 1121 12740 1133
tri 12507 1118 12510 1121 ne
rect 12510 1118 12581 1121
rect 8148 1030 8194 1076
rect 9390 1030 9436 1076
rect 10362 1072 10402 1118
tri 12510 1105 12523 1118 ne
rect 12523 1105 12581 1118
tri 12581 1105 12597 1121 sw
tri 12523 1096 12532 1105 ne
rect 12532 1096 12597 1105
rect 12153 1090 12205 1096
tri 12532 1087 12541 1096 ne
rect 12541 1087 12597 1096
tri 12541 1084 12544 1087 ne
rect 12544 1084 12597 1087
tri 12544 1083 12545 1084 ne
rect 12153 1026 12205 1038
tri 12147 968 12153 974 se
rect 12153 968 12205 974
tri 12146 967 12147 968 se
rect 12147 967 12205 968
tri 12119 940 12146 967 se
rect 12146 940 12205 967
rect 10737 888 10743 940
rect 10795 888 10807 940
rect 10859 898 12205 940
rect 10859 889 10866 898
tri 10866 889 10875 898 nw
rect 10859 888 10865 889
tri 10865 888 10866 889 nw
rect 288 644 325 790
rect 986 738 992 790
rect 1044 738 1061 790
rect 1113 738 1130 790
rect 1182 738 1199 790
rect 1251 738 1268 790
rect 1320 738 1337 790
rect 1389 738 1405 790
rect 1457 738 1473 790
rect 1525 738 1531 790
rect 986 696 1531 738
tri 12322 699 12350 727 se
rect 12350 699 12406 727
rect 986 644 992 696
rect 1044 644 1061 696
rect 1113 644 1130 696
rect 1182 644 1199 696
rect 1251 644 1268 696
rect 1320 644 1337 696
rect 1389 644 1405 696
rect 1457 644 1473 696
rect 1525 644 1531 696
tri 12271 648 12322 699 se
rect 12322 648 12406 699
rect 12271 642 12406 648
rect 12271 610 12323 642
tri 12323 610 12355 642 nw
rect 12271 415 12321 610
tri 12321 608 12323 610 nw
rect 12359 592 12427 598
rect 12359 540 12363 592
rect 12415 540 12427 592
rect 12545 571 12597 1084
rect 12694 1087 12700 1121
rect 12734 1087 12740 1121
tri 12768 1096 12805 1133 ne
rect 12805 1096 12817 1133
rect 12694 1074 12740 1087
tri 12805 1084 12817 1096 ne
rect 12886 1415 13216 1421
rect 12886 1363 12887 1415
rect 12939 1363 12956 1415
rect 13008 1363 13025 1415
rect 13077 1363 13094 1415
rect 13146 1363 13163 1415
rect 13215 1363 13216 1415
rect 12886 1345 13216 1363
rect 12886 1293 12887 1345
rect 12939 1293 12956 1345
rect 13008 1293 13025 1345
rect 13077 1293 13094 1345
rect 13146 1293 13163 1345
rect 13215 1293 13216 1345
rect 12886 1275 13216 1293
rect 12886 1223 12887 1275
rect 12939 1223 12956 1275
rect 13008 1223 13025 1275
rect 13077 1223 13094 1275
rect 13146 1223 13163 1275
rect 13215 1223 13216 1275
rect 12886 1204 13216 1223
rect 12886 1152 12887 1204
rect 12939 1152 12956 1204
rect 13008 1152 13025 1204
rect 13077 1152 13094 1204
rect 13146 1152 13163 1204
rect 13215 1152 13216 1204
rect 12886 1133 13216 1152
rect 14697 1137 15008 1369
rect 12886 1081 12887 1133
rect 12939 1081 12956 1133
rect 13008 1081 13025 1133
rect 13077 1081 13094 1133
rect 13146 1081 13163 1133
rect 13215 1081 13216 1133
rect 12886 1075 13216 1081
rect 12657 1044 12859 1074
rect 12657 1010 12700 1044
rect 12734 1010 12859 1044
rect 12657 1003 12859 1010
tri 12859 1003 12930 1074 nw
rect 12657 967 12832 1003
tri 12832 976 12859 1003 nw
rect 14823 997 14875 1003
rect 12657 933 12700 967
rect 12734 933 12832 967
rect 12657 889 12832 933
rect 12657 855 12700 889
rect 12734 855 12832 889
rect 14823 931 14875 945
rect 14823 873 14875 879
rect 12657 811 12832 855
tri 12636 790 12657 811 se
rect 12657 790 12700 811
rect 12636 777 12700 790
rect 12734 777 12832 811
rect 12636 733 12832 777
rect 12636 699 12700 733
rect 12734 699 12832 733
rect 12636 644 12832 699
tri 12752 610 12786 644 ne
tri 12545 540 12576 571 ne
rect 12576 540 12597 571
tri 12597 540 12650 593 sw
rect 12359 528 12427 540
rect 12359 476 12363 528
rect 12415 476 12427 528
tri 12576 519 12597 540 ne
rect 12597 519 12675 540
tri 12597 488 12628 519 ne
rect 12628 516 12675 519
tri 12675 516 12699 540 sw
tri 14711 516 14735 540 se
rect 14735 516 14753 540
rect 12628 488 14753 516
rect 14805 488 14817 540
rect 14869 488 14875 540
rect 12359 472 12427 476
tri 12427 472 12439 484 sw
rect 12359 470 12439 472
tri 12359 423 12406 470 ne
rect 12406 423 12439 470
tri 12439 423 12488 472 sw
tri 12321 415 12329 423 sw
tri 12406 415 12414 423 ne
rect 12414 415 12488 423
tri 12488 415 12496 423 sw
tri 12245 389 12271 415 se
rect 12271 389 12329 415
tri 12329 389 12355 415 sw
tri 12414 390 12439 415 ne
rect 12439 389 12496 415
tri 12496 389 12522 415 sw
rect 12439 355 12522 389
tri 12522 355 12556 389 sw
tri 12412 307 12439 334 se
rect 12439 307 12556 355
tri 12406 301 12412 307 se
rect 12412 301 12434 307
rect 12428 255 12434 301
rect 12486 255 12498 307
rect 12550 255 12556 307
rect 14840 260 15007 416
<< via1 >>
rect 1468 6996 1520 7005
rect 1468 6962 1474 6996
rect 1474 6962 1508 6996
rect 1508 6962 1520 6996
rect 1468 6953 1520 6962
rect 1534 6996 1586 7005
rect 1534 6962 1546 6996
rect 1546 6962 1580 6996
rect 1580 6962 1586 6996
rect 1534 6953 1586 6962
rect 7277 6574 7329 6626
rect 7341 6574 7393 6626
rect 9428 6574 9480 6626
rect 9492 6574 9544 6626
rect 14736 6382 14788 6434
rect 14736 6318 14788 6370
rect -370 5573 -318 5625
rect 11685 5626 11737 5678
rect 11749 5626 11801 5678
rect 12949 5626 13001 5678
rect 13013 5626 13065 5678
rect -370 5509 -318 5561
rect 6876 5546 6928 5598
rect 6940 5546 6992 5598
rect 12200 5546 12252 5598
rect 12264 5546 12316 5598
rect -194 5440 -142 5492
rect -194 5354 -142 5406
rect -18 5446 34 5498
rect -18 5374 34 5426
rect 9428 5428 9480 5480
rect 9492 5428 9544 5480
rect 11573 5428 11625 5480
rect 11637 5428 11689 5480
rect 12079 5443 12131 5495
rect 12143 5443 12195 5495
rect 721 5280 773 5332
rect 785 5280 837 5332
rect 6876 5274 6928 5326
rect 6940 5274 6992 5326
rect 12200 5346 12252 5398
rect 12264 5346 12316 5398
rect 9441 5266 9493 5318
rect 9505 5266 9557 5318
rect 5228 5187 5280 5239
rect 5228 5123 5280 5175
rect 7411 5166 7463 5218
rect 7411 5102 7463 5154
rect 13341 4939 13393 4991
rect 13413 4939 13465 4991
rect 13484 4939 13536 4991
rect 13555 4939 13607 4991
rect 13626 4939 13678 4991
rect 829 4858 881 4910
rect 894 4858 946 4910
rect 959 4858 1011 4910
rect 1024 4858 1076 4910
rect 1089 4858 1141 4910
rect 1153 4858 1205 4910
rect 1217 4858 1269 4910
rect 1281 4858 1333 4910
rect 1345 4858 1397 4910
rect 1409 4858 1461 4910
rect 1473 4858 1525 4910
rect 829 4783 881 4835
rect 894 4783 946 4835
rect 959 4783 1011 4835
rect 1024 4783 1076 4835
rect 1089 4783 1141 4835
rect 1153 4783 1205 4835
rect 1217 4783 1269 4835
rect 1281 4783 1333 4835
rect 1345 4783 1397 4835
rect 1409 4783 1461 4835
rect 1473 4783 1525 4835
rect 829 4708 881 4760
rect 894 4708 946 4760
rect 959 4708 1011 4760
rect 1024 4708 1076 4760
rect 1089 4708 1141 4760
rect 1153 4708 1205 4760
rect 1217 4708 1269 4760
rect 1281 4708 1333 4760
rect 1345 4708 1397 4760
rect 1409 4708 1461 4760
rect 1473 4708 1525 4760
rect 13341 4864 13393 4916
rect 13413 4864 13465 4916
rect 13484 4864 13536 4916
rect 13555 4864 13607 4916
rect 13626 4864 13678 4916
rect 13341 4789 13393 4841
rect 13413 4789 13465 4841
rect 13484 4789 13536 4841
rect 13555 4789 13607 4841
rect 13626 4789 13678 4841
rect 9936 4626 9988 4678
rect 10000 4626 10052 4678
rect 10190 4626 10242 4678
rect 10254 4626 10306 4678
rect 11621 4544 11673 4596
rect 11685 4544 11737 4596
rect 12159 4585 12211 4637
rect 12224 4585 12276 4637
rect 14690 4585 14742 4637
rect 14754 4585 14806 4637
rect 14591 4505 14643 4557
rect 14655 4505 14707 4557
rect 5178 4212 5230 4264
rect 5242 4212 5294 4264
rect 238 4134 290 4140
rect 238 4100 271 4134
rect 271 4100 290 4134
rect 238 4088 290 4100
rect 238 4054 290 4061
rect 238 4020 271 4054
rect 271 4020 290 4054
rect 238 4009 290 4020
rect 238 3974 290 3982
rect 1704 4129 1756 4181
rect 1773 4129 1825 4181
rect 1842 4129 1894 4181
rect 1911 4129 1963 4181
rect 1980 4129 2032 4181
rect 1704 4054 1756 4106
rect 1773 4054 1825 4106
rect 1842 4054 1894 4106
rect 1911 4054 1963 4106
rect 1980 4054 2032 4106
rect 1704 3979 1756 4031
rect 1773 3979 1825 4031
rect 1842 3979 1894 4031
rect 1911 3979 1963 4031
rect 1980 3979 2032 4031
rect 3156 4129 3208 4181
rect 3220 4129 3272 4181
rect 3284 4129 3336 4181
rect 3348 4129 3400 4181
rect 3412 4129 3464 4181
rect 3476 4129 3528 4181
rect 3540 4129 3592 4181
rect 3156 4054 3208 4106
rect 3220 4054 3272 4106
rect 3284 4054 3336 4106
rect 3348 4054 3400 4106
rect 3412 4054 3464 4106
rect 3476 4054 3528 4106
rect 3540 4054 3592 4106
rect 3156 3979 3208 4031
rect 3220 3979 3272 4031
rect 3284 3979 3336 4031
rect 3348 3979 3400 4031
rect 3412 3979 3464 4031
rect 3476 3979 3528 4031
rect 3540 3979 3592 4031
rect 238 3940 271 3974
rect 271 3940 290 3974
rect 238 3930 290 3940
rect 238 3893 290 3903
rect 238 3859 271 3893
rect 271 3859 290 3893
rect 829 3871 881 3923
rect 902 3871 954 3923
rect 974 3871 1026 3923
rect 1046 3871 1098 3923
rect 1118 3871 1170 3923
rect 1190 3871 1242 3923
rect 8037 3899 8089 3951
rect 8101 3899 8153 3951
rect 10001 3893 10053 3945
rect 238 3851 290 3859
rect 238 3812 290 3824
rect 10001 3829 10053 3881
rect 238 3778 271 3812
rect 271 3778 290 3812
rect 238 3772 290 3778
rect 947 3602 999 3654
rect 1013 3602 1065 3654
rect 1079 3602 1131 3654
rect 1145 3602 1197 3654
rect 1211 3602 1263 3654
rect 1277 3602 1329 3654
rect 1343 3602 1395 3654
rect 1408 3602 1460 3654
rect 1473 3602 1525 3654
rect 947 3528 999 3580
rect 1013 3528 1065 3580
rect 1079 3528 1131 3580
rect 1145 3528 1197 3580
rect 1211 3528 1263 3580
rect 1277 3528 1329 3580
rect 1343 3528 1395 3580
rect 1408 3528 1460 3580
rect 1473 3528 1525 3580
rect 947 3454 999 3506
rect 1013 3454 1065 3506
rect 1079 3454 1131 3506
rect 1145 3454 1197 3506
rect 1211 3454 1263 3506
rect 1277 3454 1329 3506
rect 1343 3454 1395 3506
rect 1408 3454 1460 3506
rect 1473 3454 1525 3506
rect 13338 3652 13390 3704
rect 13411 3652 13463 3704
rect 13484 3652 13536 3704
rect 13557 3652 13609 3704
rect 13630 3652 13682 3704
rect 13338 3586 13390 3638
rect 13411 3586 13463 3638
rect 13484 3586 13536 3638
rect 13557 3586 13609 3638
rect 13630 3586 13682 3638
rect 12887 3508 12939 3560
rect 12956 3508 13008 3560
rect 13025 3508 13077 3560
rect 13094 3508 13146 3560
rect 13163 3508 13215 3560
rect 12887 3438 12939 3490
rect 12956 3438 13008 3490
rect 13025 3438 13077 3490
rect 13094 3438 13146 3490
rect 13163 3438 13215 3490
rect 12887 3368 12939 3420
rect 12956 3368 13008 3420
rect 13025 3368 13077 3420
rect 13094 3368 13146 3420
rect 13163 3368 13215 3420
rect 12887 3297 12939 3349
rect 12956 3297 13008 3349
rect 13025 3297 13077 3349
rect 13094 3297 13146 3349
rect 13163 3297 13215 3349
rect 2373 3240 2425 3292
rect 2437 3240 2489 3292
rect 7005 3240 7057 3292
rect 7069 3240 7121 3292
rect 12887 3226 12939 3278
rect 12956 3226 13008 3278
rect 13025 3226 13077 3278
rect 13094 3226 13146 3278
rect 13163 3226 13215 3278
rect 13338 3520 13390 3572
rect 13411 3520 13463 3572
rect 13484 3520 13536 3572
rect 13557 3520 13609 3572
rect 13630 3520 13682 3572
rect 13338 3454 13390 3506
rect 13411 3454 13463 3506
rect 13484 3454 13536 3506
rect 13557 3454 13609 3506
rect 13630 3454 13682 3506
rect 13338 3388 13390 3440
rect 13411 3388 13463 3440
rect 13484 3388 13536 3440
rect 13557 3388 13609 3440
rect 13630 3388 13682 3440
rect 13338 3322 13390 3374
rect 13411 3322 13463 3374
rect 13484 3322 13536 3374
rect 13557 3322 13609 3374
rect 13630 3322 13682 3374
rect 13338 3256 13390 3308
rect 13411 3256 13463 3308
rect 13484 3256 13536 3308
rect 13557 3256 13609 3308
rect 13630 3256 13682 3308
rect 13338 3190 13390 3242
rect 13411 3190 13463 3242
rect 13484 3190 13536 3242
rect 13557 3190 13609 3242
rect 13630 3190 13682 3242
rect 238 3074 290 3126
rect 13338 3124 13390 3176
rect 13411 3124 13463 3176
rect 13484 3124 13536 3176
rect 13557 3124 13609 3176
rect 13630 3124 13682 3176
rect 238 3002 290 3054
rect 238 2930 290 2982
rect 1704 3005 1756 3057
rect 1773 3005 1825 3057
rect 1842 3005 1894 3057
rect 1911 3005 1963 3057
rect 1980 3005 2032 3057
rect 1704 2929 1756 2981
rect 1773 2929 1825 2981
rect 1842 2929 1894 2981
rect 1911 2929 1963 2981
rect 1980 2929 2032 2981
rect 3156 3005 3208 3057
rect 3220 3005 3272 3057
rect 3284 3005 3336 3057
rect 3348 3005 3400 3057
rect 3412 3005 3464 3057
rect 3476 3005 3528 3057
rect 3540 3005 3592 3057
rect 3156 2929 3208 2981
rect 3220 2929 3272 2981
rect 3284 2929 3336 2981
rect 3348 2929 3400 2981
rect 3412 2929 3464 2981
rect 3476 2929 3528 2981
rect 3540 2929 3592 2981
rect 238 2857 290 2909
rect 10173 2848 10225 2900
rect 10237 2848 10289 2900
rect 238 2784 290 2836
rect 12073 2842 12125 2894
rect 12073 2778 12125 2830
rect 238 2711 290 2763
rect 238 2638 290 2690
rect 238 2565 290 2617
rect 1704 2390 1756 2442
rect 1773 2390 1825 2442
rect 1842 2390 1894 2442
rect 1911 2390 1963 2442
rect 1980 2390 2032 2442
rect 1704 2312 1756 2364
rect 1773 2312 1825 2364
rect 1842 2312 1894 2364
rect 1911 2312 1963 2364
rect 1980 2312 2032 2364
rect 3156 2390 3208 2442
rect 3220 2390 3272 2442
rect 3284 2390 3336 2442
rect 3348 2390 3400 2442
rect 3412 2390 3464 2442
rect 3476 2390 3528 2442
rect 3540 2390 3592 2442
rect 3156 2312 3208 2364
rect 3220 2312 3272 2364
rect 3284 2312 3336 2364
rect 3348 2312 3400 2364
rect 3412 2312 3464 2364
rect 3476 2312 3528 2364
rect 3540 2312 3592 2364
rect 1704 1977 1756 2029
rect 1773 1977 1825 2029
rect 1842 1977 1894 2029
rect 1911 1977 1963 2029
rect 1980 1977 2032 2029
rect 1704 1903 1756 1955
rect 1773 1903 1825 1955
rect 1842 1903 1894 1955
rect 1911 1903 1963 1955
rect 1980 1903 2032 1955
rect 1704 1829 1756 1881
rect 1773 1829 1825 1881
rect 1842 1829 1894 1881
rect 1911 1829 1963 1881
rect 1980 1829 2032 1881
rect 3156 1977 3208 2029
rect 3220 1977 3272 2029
rect 3284 1977 3336 2029
rect 3348 1977 3400 2029
rect 3412 1977 3464 2029
rect 3476 1977 3528 2029
rect 3540 1977 3592 2029
rect 3156 1903 3208 1955
rect 3220 1903 3272 1955
rect 3284 1903 3336 1955
rect 3348 1903 3400 1955
rect 3412 1903 3464 1955
rect 3476 1903 3528 1955
rect 3540 1903 3592 1955
rect 3156 1829 3208 1881
rect 3220 1829 3272 1881
rect 3284 1829 3336 1881
rect 3348 1829 3400 1881
rect 3412 1829 3464 1881
rect 3476 1829 3528 1881
rect 3540 1829 3592 1881
rect 706 1602 758 1654
rect 7997 1606 8049 1658
rect 8061 1606 8113 1658
rect 706 1538 758 1590
rect 992 1451 1044 1503
rect 1061 1451 1113 1503
rect 1130 1451 1182 1503
rect 1199 1451 1251 1503
rect 1268 1451 1320 1503
rect 1337 1451 1389 1503
rect 1405 1451 1457 1503
rect 1473 1451 1525 1503
rect 992 1377 1044 1429
rect 1061 1377 1113 1429
rect 1130 1377 1182 1429
rect 1199 1377 1251 1429
rect 1268 1377 1320 1429
rect 1337 1377 1389 1429
rect 1405 1377 1457 1429
rect 1473 1377 1525 1429
rect 992 1303 1044 1355
rect 1061 1303 1113 1355
rect 1130 1303 1182 1355
rect 1199 1303 1251 1355
rect 1268 1303 1320 1355
rect 1337 1303 1389 1355
rect 1405 1303 1457 1355
rect 1473 1303 1525 1355
rect 12153 1038 12205 1090
rect 12153 974 12205 1026
rect 10743 888 10795 940
rect 10807 888 10859 940
rect 992 738 1044 790
rect 1061 738 1113 790
rect 1130 738 1182 790
rect 1199 738 1251 790
rect 1268 738 1320 790
rect 1337 738 1389 790
rect 1405 738 1457 790
rect 1473 738 1525 790
rect 992 644 1044 696
rect 1061 644 1113 696
rect 1130 644 1182 696
rect 1199 644 1251 696
rect 1268 644 1320 696
rect 1337 644 1389 696
rect 1405 644 1457 696
rect 1473 644 1525 696
rect 12363 540 12415 592
rect 12887 1363 12939 1415
rect 12956 1363 13008 1415
rect 13025 1363 13077 1415
rect 13094 1363 13146 1415
rect 13163 1363 13215 1415
rect 12887 1293 12939 1345
rect 12956 1293 13008 1345
rect 13025 1293 13077 1345
rect 13094 1293 13146 1345
rect 13163 1293 13215 1345
rect 12887 1223 12939 1275
rect 12956 1223 13008 1275
rect 13025 1223 13077 1275
rect 13094 1223 13146 1275
rect 13163 1223 13215 1275
rect 12887 1152 12939 1204
rect 12956 1152 13008 1204
rect 13025 1152 13077 1204
rect 13094 1152 13146 1204
rect 13163 1152 13215 1204
rect 12887 1081 12939 1133
rect 12956 1081 13008 1133
rect 13025 1081 13077 1133
rect 13094 1081 13146 1133
rect 13163 1081 13215 1133
rect 14823 945 14875 997
rect 14823 879 14875 931
rect 12363 476 12415 528
rect 14753 488 14805 540
rect 14817 488 14869 540
rect 12434 255 12486 307
rect 12498 255 12550 307
<< metal2 >>
tri 1301 6953 1353 7005 se
rect 1353 6953 1468 7005
rect 1520 6953 1534 7005
rect 1586 6953 1592 7005
tri 1273 6925 1301 6953 se
rect 1301 6925 1347 6953
tri 1347 6925 1375 6953 nw
tri 1221 6873 1273 6925 se
rect 1221 5703 1273 6873
tri 1273 6851 1347 6925 nw
rect 3354 6878 3400 6924
rect 3827 6885 3879 6924
rect 7271 6574 7277 6626
rect 7329 6574 7341 6626
rect 7393 6574 7399 6626
tri 7271 6498 7347 6574 ne
tri 1221 5701 1223 5703 ne
rect 1223 5701 1273 5703
tri 1273 5701 1297 5725 sw
tri 1223 5678 1246 5701 ne
rect 1246 5678 1297 5701
tri 1297 5678 1320 5701 sw
tri 1246 5651 1273 5678 ne
rect 1273 5651 1320 5678
tri 1273 5631 1293 5651 ne
rect 1293 5631 1320 5651
rect -370 5625 -318 5631
tri 1293 5627 1297 5631 ne
rect 1297 5627 1320 5631
tri 1320 5627 1371 5678 sw
tri 1297 5626 1298 5627 ne
rect 1298 5626 1371 5627
tri 1371 5626 1372 5627 sw
tri 1298 5598 1326 5626 ne
rect 1326 5598 1372 5626
tri 1372 5598 1400 5626 sw
rect -370 5561 -318 5573
tri 1326 5553 1371 5598 ne
rect 1371 5553 1400 5598
tri 1400 5553 1445 5598 sw
tri 1371 5546 1378 5553 ne
rect 1378 5546 1445 5553
tri 1445 5546 1452 5553 sw
rect 6870 5546 6876 5598
rect 6928 5546 6940 5598
rect 6992 5546 6998 5598
tri -374 696 -370 700 se
rect -370 696 -318 5509
tri 1378 5504 1420 5546 ne
rect 1420 5512 1452 5546
tri 1452 5512 1486 5546 sw
tri 6874 5512 6908 5546 ne
rect 1420 5504 1486 5512
rect -18 5498 34 5504
rect -194 5492 -142 5498
rect -194 5406 -142 5440
rect -194 4885 -142 5354
tri 1420 5495 1429 5504 ne
rect 1429 5495 1486 5504
tri 1486 5495 1503 5512 sw
tri 1429 5480 1444 5495 ne
rect 1444 5480 1503 5495
tri 1503 5480 1518 5495 sw
tri 1444 5479 1445 5480 ne
rect 1445 5479 1518 5480
tri 1518 5479 1519 5480 sw
rect -18 5426 34 5446
tri 1445 5428 1496 5479 ne
rect 1496 5428 1519 5479
tri 1519 5428 1570 5479 sw
tri 1496 5405 1519 5428 ne
rect 1519 5405 1570 5428
tri 1570 5405 1593 5428 sw
tri 1519 5398 1526 5405 ne
rect 1526 5398 1593 5405
tri 1593 5398 1600 5405 sw
tri -142 4885 -136 4891 sw
rect -194 4869 -136 4885
tri -194 4858 -183 4869 ne
rect -183 4858 -136 4869
tri -136 4858 -109 4885 sw
tri -183 4841 -166 4858 ne
rect -166 4841 -109 4858
tri -109 4841 -92 4858 sw
tri -166 4835 -160 4841 ne
rect -160 4835 -92 4841
tri -92 4835 -86 4841 sw
tri -160 4827 -152 4835 ne
rect -152 4827 -86 4835
tri -86 4827 -78 4835 sw
tri -152 4817 -142 4827 ne
rect -142 4817 -78 4827
tri -142 4805 -130 4817 ne
tri -144 4544 -130 4558 se
rect -130 4544 -78 4817
rect -18 4708 34 5374
tri 1526 5346 1578 5398 ne
rect 1578 5360 1600 5398
tri 1600 5360 1638 5398 sw
rect 1578 5346 1638 5360
tri 1638 5346 1652 5360 sw
tri 6894 5346 6908 5360 se
rect 6908 5346 6960 5546
tri 6960 5512 6994 5546 nw
tri 6960 5346 6974 5360 sw
tri 1578 5332 1592 5346 ne
rect 1592 5332 1652 5346
tri 1652 5332 1666 5346 sw
tri 6880 5332 6894 5346 se
rect 6894 5332 6974 5346
rect 715 5280 721 5332
rect 773 5280 785 5332
rect 837 5280 843 5332
tri 1592 5331 1593 5332 ne
rect 1593 5331 1666 5332
tri 1666 5331 1667 5332 sw
tri 6879 5331 6880 5332 se
rect 6880 5331 6974 5332
tri 1593 5326 1598 5331 ne
rect 1598 5326 1667 5331
tri 1667 5326 1672 5331 sw
tri 6874 5326 6879 5331 se
rect 6879 5326 6974 5331
tri 6974 5326 6994 5346 sw
tri 7339 5326 7347 5334 se
rect 7347 5326 7399 6574
rect 9422 6574 9428 6626
rect 9480 6574 9492 6626
rect 9544 6574 9550 6626
tri 13110 6574 13136 6600 se
rect 13136 6574 14739 6600
tri 14739 6574 14765 6600 sw
tri 9422 6536 9460 6574 ne
tri 9437 5495 9460 5518 se
rect 9460 5512 9512 6574
tri 9512 6536 9550 6574 nw
tri 13087 6551 13110 6574 se
rect 13110 6551 14765 6574
tri 14765 6551 14788 6574 sw
tri 13072 6536 13087 6551 se
rect 13087 6548 14788 6551
rect 13087 6536 13136 6548
tri 13062 6526 13072 6536 se
rect 13072 6526 13136 6536
tri 13136 6526 13158 6548 nw
tri 14701 6526 14723 6548 ne
rect 14723 6526 14788 6548
tri 12988 6452 13062 6526 se
tri 13062 6452 13136 6526 nw
tri 14723 6513 14736 6526 ne
tri 12981 6445 12988 6452 se
rect 12988 6445 13055 6452
tri 13055 6445 13062 6452 nw
rect 12981 6434 13044 6445
tri 13044 6434 13055 6445 nw
rect 14736 6434 14788 6526
tri 12943 5678 12981 5716 se
rect 12981 5678 13033 6434
tri 13033 6423 13044 6434 nw
rect 14736 6370 14788 6382
rect 14736 6312 14788 6318
tri 13033 5678 13071 5716 sw
rect 11679 5626 11685 5678
rect 11737 5626 11749 5678
rect 11801 5626 11807 5678
rect 12943 5626 12949 5678
rect 13001 5626 13013 5678
rect 13065 5626 13071 5678
tri 11676 5598 11679 5601 se
rect 11679 5598 11774 5626
tri 11774 5598 11802 5626 nw
tri 11624 5546 11676 5598 se
rect 11676 5546 11722 5598
tri 11722 5546 11774 5598 nw
rect 12194 5546 12200 5598
rect 12252 5546 12264 5598
rect 12316 5546 12322 5598
tri 11597 5519 11624 5546 se
rect 11624 5519 11695 5546
tri 11695 5519 11722 5546 nw
tri 12198 5519 12225 5546 ne
rect 12225 5519 12284 5546
tri 11596 5518 11597 5519 se
rect 11597 5518 11695 5519
tri 9512 5512 9518 5518 sw
tri 11590 5512 11596 5518 se
rect 11596 5512 11695 5518
tri 12225 5512 12232 5519 ne
rect 9460 5495 9518 5512
tri 9518 5495 9535 5512 sw
tri 11573 5495 11590 5512 se
rect 11590 5495 11695 5512
tri 9422 5480 9437 5495 se
rect 9437 5480 9535 5495
tri 9535 5480 9550 5495 sw
rect 9422 5428 9428 5480
rect 9480 5428 9492 5480
rect 9544 5428 9550 5480
tri 11567 5489 11573 5495 se
rect 11573 5489 11695 5495
rect 11567 5480 11695 5489
rect 11567 5428 11573 5480
rect 11625 5428 11637 5480
rect 11689 5428 11695 5480
rect 12073 5443 12079 5495
rect 12131 5443 12143 5495
rect 12195 5443 12201 5495
tri 1598 5280 1644 5326 ne
rect 1644 5280 1672 5326
tri 1672 5280 1718 5326 sw
rect 715 5274 795 5280
tri 795 5274 801 5280 nw
tri 1644 5274 1650 5280 ne
rect 1650 5274 1718 5280
tri 1718 5274 1724 5280 sw
rect 6870 5274 6876 5326
rect 6928 5274 6940 5326
rect 6992 5274 6998 5326
tri 7331 5318 7339 5326 se
rect 7339 5318 7399 5326
tri 7287 5274 7331 5318 se
rect 7331 5312 7399 5318
rect 7331 5274 7353 5312
rect 715 5266 787 5274
tri 787 5266 795 5274 nw
tri 1650 5266 1658 5274 ne
rect 1658 5266 1724 5274
tri 1724 5266 1732 5274 sw
tri 7279 5266 7287 5274 se
rect 7287 5266 7353 5274
tri 7353 5266 7399 5312 nw
rect 9435 5266 9441 5318
rect 9493 5266 9505 5318
rect 9557 5266 9563 5318
tri 688 4858 715 4885 se
rect 715 4862 767 5266
tri 767 5246 787 5266 nw
tri 1658 5257 1667 5266 ne
rect 1667 5257 1732 5266
tri 1732 5257 1741 5266 sw
tri 7273 5260 7279 5266 se
rect 7279 5260 7347 5266
tri 7347 5260 7353 5266 nw
tri 9435 5260 9441 5266 ne
rect 9441 5260 9557 5266
tri 9557 5260 9563 5266 nw
tri 7270 5257 7273 5260 se
rect 7273 5257 7315 5260
tri 1667 5246 1678 5257 ne
rect 1678 5246 1741 5257
tri 1741 5246 1752 5257 sw
tri 7259 5246 7270 5257 se
rect 7270 5246 7315 5257
tri 1678 5239 1685 5246 ne
rect 1685 5239 1752 5246
tri 1752 5239 1759 5246 sw
tri 7258 5245 7259 5246 se
rect 7259 5245 7315 5246
rect 5228 5239 5280 5245
tri 1685 5187 1737 5239 ne
rect 1737 5187 1759 5239
tri 1759 5187 1811 5239 sw
tri 1737 5183 1741 5187 ne
rect 1741 5183 1811 5187
tri 1811 5183 1815 5187 sw
tri 1741 5175 1749 5183 ne
rect 1749 5175 1815 5183
tri 1815 5175 1823 5183 sw
rect 5228 5175 5280 5187
tri 1749 5123 1801 5175 ne
rect 1801 5123 1823 5175
tri 1823 5123 1875 5175 sw
tri 1801 5109 1815 5123 ne
rect 1815 5109 1875 5123
tri 1875 5109 1889 5123 sw
tri 1815 5102 1822 5109 ne
rect 1822 5102 1889 5109
tri 1889 5102 1896 5109 sw
tri 1822 5035 1889 5102 ne
rect 1889 5035 1896 5102
tri 1896 5035 1963 5102 sw
tri 1889 5013 1911 5035 ne
rect 715 4858 763 4862
tri 763 4858 767 4862 nw
rect 823 4858 829 4910
rect 881 4858 894 4910
rect 946 4858 959 4910
rect 1011 4858 1024 4910
rect 1076 4858 1089 4910
rect 1141 4858 1153 4910
rect 1205 4858 1217 4910
rect 1269 4858 1281 4910
rect 1333 4858 1345 4910
rect 1397 4858 1409 4910
rect 1461 4858 1473 4910
rect 1525 4858 1531 4910
tri 677 4847 688 4858 se
rect 688 4847 752 4858
tri 752 4847 763 4858 nw
rect 677 4841 746 4847
tri 746 4841 752 4847 nw
rect 677 4835 740 4841
tri 740 4835 746 4841 nw
rect 823 4835 1531 4858
tri 34 4708 45 4719 sw
rect -18 4697 45 4708
tri -18 4678 1 4697 ne
rect 1 4678 45 4697
tri 45 4678 75 4708 sw
tri 1 4649 30 4678 ne
rect 30 4649 75 4678
tri 75 4649 104 4678 sw
tri 30 4645 34 4649 ne
rect 34 4645 104 4649
tri 34 4627 52 4645 ne
tri -183 4505 -144 4544 se
rect -144 4518 -78 4544
rect -144 4505 -91 4518
tri -91 4505 -78 4518 nw
tri -193 4495 -183 4505 se
rect -183 4495 -101 4505
tri -101 4495 -91 4505 nw
tri -267 4365 -193 4439 se
rect -193 4417 -141 4495
tri -141 4455 -101 4495 nw
tri -193 4365 -141 4417 nw
rect -374 687 -318 696
rect -374 607 -318 631
rect -374 541 -318 551
tri -277 4355 -267 4365 se
rect -267 4355 -203 4365
tri -203 4355 -193 4365 nw
tri -351 379 -277 453 se
rect -277 431 -225 4355
tri -225 4333 -203 4355 nw
tri 20 3454 52 3486 se
rect 52 3464 104 4645
rect 52 3454 94 3464
tri 94 3454 104 3464 nw
rect 238 4140 290 4146
rect 238 4061 290 4088
rect 238 3982 290 4009
rect 238 3903 290 3930
rect 238 3824 290 3851
tri 4 3438 20 3454 se
rect 20 3438 78 3454
tri 78 3438 94 3454 nw
tri -14 3420 4 3438 se
rect 4 3420 60 3438
tri 60 3420 78 3438 nw
tri -22 3412 -14 3420 se
rect -14 3412 52 3420
tri 52 3412 60 3420 nw
tri -66 3368 -22 3412 se
rect -22 3368 8 3412
tri 8 3368 52 3412 nw
tri -85 3349 -66 3368 se
rect -66 3349 -11 3368
tri -11 3349 8 3368 nw
tri -96 3338 -85 3349 se
rect -85 3338 -22 3349
tri -22 3338 -11 3349 nw
tri -105 3329 -96 3338 se
rect -96 3329 -31 3338
tri -31 3329 -22 3338 nw
tri -277 379 -225 431 nw
tri -126 2101 -105 2122 se
rect -105 2101 -53 3329
tri -53 3307 -31 3329 nw
rect 238 3126 290 3772
rect 238 3054 290 3074
rect 238 2982 290 3002
rect 238 2909 290 2930
rect 677 2947 729 4835
tri 729 4824 740 4835 nw
rect 823 4783 829 4835
rect 881 4783 894 4835
rect 946 4783 959 4835
rect 1011 4783 1024 4835
rect 1076 4783 1089 4835
rect 1141 4783 1153 4835
rect 1205 4783 1217 4835
rect 1269 4783 1281 4835
rect 1333 4783 1345 4835
rect 1397 4783 1409 4835
rect 1461 4783 1473 4835
rect 1525 4783 1531 4835
rect 1911 4806 1963 5035
tri 1963 4806 1975 4818 sw
rect 1911 4796 1975 4806
tri 1911 4789 1918 4796 ne
rect 1918 4789 1975 4796
tri 1975 4789 1992 4806 sw
rect 823 4760 1531 4783
rect 823 4708 829 4760
rect 881 4708 894 4760
rect 946 4708 959 4760
rect 1011 4708 1024 4760
rect 1076 4708 1089 4760
rect 1141 4708 1153 4760
rect 1205 4708 1217 4760
rect 1269 4708 1281 4760
rect 1333 4708 1345 4760
rect 1397 4708 1409 4760
rect 1461 4708 1473 4760
rect 1525 4708 1531 4760
tri 1918 4732 1975 4789 ne
rect 1975 4732 1992 4789
tri 1992 4732 2049 4789 sw
rect 823 3923 1531 4708
tri 1975 4678 2029 4732 ne
rect 2029 4678 2049 4732
tri 2049 4678 2103 4732 sw
tri 2029 4658 2049 4678 ne
rect 2049 4658 2103 4678
tri 2103 4658 2123 4678 sw
tri 2049 4626 2081 4658 ne
rect 2081 4626 2123 4658
tri 2123 4626 2155 4658 sw
tri 2081 4596 2111 4626 ne
rect 2111 4596 2155 4626
tri 2155 4596 2185 4626 sw
tri 2111 4584 2123 4596 ne
rect 2123 4584 2185 4596
tri 2185 4584 2197 4596 sw
tri 2123 4544 2163 4584 ne
rect 2163 4544 2197 4584
tri 2197 4544 2237 4584 sw
tri 2163 4510 2197 4544 ne
rect 2197 4510 2237 4544
tri 2237 4510 2271 4544 sw
tri 2197 4505 2202 4510 ne
rect 2202 4505 2271 4510
tri 2271 4505 2276 4510 sw
tri 2202 4436 2271 4505 ne
rect 2271 4436 2276 4505
tri 2276 4436 2345 4505 sw
tri 2271 4362 2345 4436 ne
tri 2345 4362 2419 4436 sw
tri 2345 4340 2367 4362 ne
rect 823 3871 829 3923
rect 881 3871 902 3923
rect 954 3871 974 3923
rect 1026 3871 1046 3923
rect 1098 3871 1118 3923
rect 1170 3871 1190 3923
rect 1242 3871 1531 3923
rect 823 3654 1531 3871
rect 823 3602 947 3654
rect 999 3602 1013 3654
rect 1065 3602 1079 3654
rect 1131 3602 1145 3654
rect 1197 3602 1211 3654
rect 1263 3602 1277 3654
rect 1329 3602 1343 3654
rect 1395 3602 1408 3654
rect 1460 3602 1473 3654
rect 1525 3602 1531 3654
rect 823 3580 1531 3602
rect 823 3528 947 3580
rect 999 3528 1013 3580
rect 1065 3528 1079 3580
rect 1131 3528 1145 3580
rect 1197 3528 1211 3580
rect 1263 3528 1277 3580
rect 1329 3528 1343 3580
rect 1395 3528 1408 3580
rect 1460 3528 1473 3580
rect 1525 3528 1531 3580
rect 823 3506 1531 3528
rect 823 3454 947 3506
rect 999 3454 1013 3506
rect 1065 3454 1079 3506
rect 1131 3454 1145 3506
rect 1197 3454 1211 3506
rect 1263 3454 1277 3506
rect 1329 3454 1343 3506
rect 1395 3454 1408 3506
rect 1460 3454 1473 3506
rect 1525 3454 1531 3506
rect 823 3445 1531 3454
tri 823 3438 830 3445 ne
rect 830 3438 1531 3445
tri 830 3420 848 3438 ne
rect 848 3420 1531 3438
tri 848 3368 900 3420 ne
rect 900 3368 1531 3420
tri 900 3349 919 3368 ne
rect 919 3349 1531 3368
tri 919 3297 971 3349 ne
rect 971 3297 1531 3349
tri 971 3292 976 3297 ne
rect 976 3292 1531 3297
tri 976 3282 986 3292 ne
tri 729 2947 751 2969 sw
tri 677 2929 695 2947 ne
rect 695 2940 751 2947
tri 751 2940 758 2947 sw
rect 695 2929 758 2940
tri 695 2918 706 2929 ne
rect 238 2836 290 2857
rect 238 2763 290 2784
rect 238 2690 290 2711
rect 238 2617 290 2638
rect 238 2559 290 2565
rect -126 2100 -53 2101
tri -129 405 -126 408 se
rect -126 405 -74 2100
tri -74 2079 -53 2100 nw
rect 706 1654 758 2929
rect 706 1590 758 1602
rect 706 1532 758 1538
rect 986 2718 1531 3292
rect 1698 4129 1704 4181
rect 1756 4129 1773 4181
rect 1825 4129 1842 4181
rect 1894 4129 1911 4181
rect 1963 4129 1980 4181
rect 2032 4129 2038 4181
rect 1698 4106 2038 4129
rect 1698 4054 1704 4106
rect 1756 4054 1773 4106
rect 1825 4054 1842 4106
rect 1894 4054 1911 4106
rect 1963 4054 1980 4106
rect 2032 4054 2038 4106
rect 1698 4031 2038 4054
rect 1698 3979 1704 4031
rect 1756 3979 1773 4031
rect 1825 3979 1842 4031
rect 1894 3979 1911 4031
rect 1963 3979 1980 4031
rect 2032 3979 2038 4031
rect 1698 3057 2038 3979
rect 2367 3297 2419 4362
tri 5193 4284 5228 4319 se
rect 5228 4284 5280 5123
tri 7241 5228 7258 5245 se
rect 7258 5228 7315 5245
tri 7315 5228 7347 5260 nw
tri 9441 5244 9457 5260 ne
rect 9457 5244 9541 5260
tri 9541 5244 9557 5260 nw
tri 9457 5242 9459 5244 ne
rect 9459 5242 9541 5244
tri 9459 5228 9473 5242 ne
rect 9473 5228 9541 5242
tri 10508 5228 10522 5242 se
rect 10522 5228 11301 5242
tri 11301 5228 11315 5242 sw
rect 7241 5224 7311 5228
tri 7311 5224 7315 5228 nw
tri 9473 5224 9477 5228 ne
rect 9477 5224 9541 5228
tri 10504 5224 10508 5228 se
rect 10508 5224 11315 5228
tri 11315 5224 11319 5228 sw
rect 7241 5218 7305 5224
tri 7305 5218 7311 5224 nw
rect 7411 5218 7463 5224
tri 7212 4544 7241 4573 se
rect 7241 4551 7293 5218
tri 7293 5206 7305 5218 nw
rect 7241 4544 7286 4551
tri 7286 4544 7293 4551 nw
tri 9477 5208 9493 5224 ne
rect 7411 5154 7463 5166
tri 7178 4510 7212 4544 se
rect 7212 4510 7247 4544
tri 7173 4505 7178 4510 se
rect 7178 4505 7247 4510
tri 7247 4505 7286 4544 nw
tri 7389 4508 7411 4530 se
rect 7411 4508 7463 5102
rect 7960 5168 8051 5176
tri 8051 5168 8059 5176 nw
rect 7960 5133 8016 5168
tri 8016 5133 8051 5168 nw
tri 7957 4544 7960 4547 se
rect 7960 4544 8012 5133
tri 8012 5129 8016 5133 nw
tri 7386 4505 7389 4508 se
rect 7389 4505 7460 4508
tri 7460 4505 7463 4508 nw
tri 7918 4505 7957 4544 se
rect 7957 4525 8012 4544
rect 7957 4505 7992 4525
tri 7992 4505 8012 4525 nw
tri 7167 4499 7173 4505 se
rect 7173 4499 7241 4505
tri 7241 4499 7247 4505 nw
tri 7380 4499 7386 4505 se
rect 7386 4499 7454 4505
tri 7454 4499 7460 4505 nw
tri 7912 4499 7918 4505 se
rect 7918 4499 7986 4505
tri 7986 4499 7992 4505 nw
tri 7104 4436 7167 4499 se
tri 7093 4425 7104 4436 se
rect 7104 4425 7167 4436
tri 7167 4425 7241 4499 nw
tri 7360 4479 7380 4499 se
rect 7380 4479 7412 4499
tri 7082 4414 7093 4425 se
rect 7093 4414 7156 4425
tri 7156 4414 7167 4425 nw
tri 7019 4351 7082 4414 se
rect 7082 4351 7093 4414
tri 7093 4351 7156 4414 nw
tri 7010 4342 7019 4351 se
rect 7019 4342 7084 4351
tri 7084 4342 7093 4351 nw
tri 5173 4264 5193 4284 se
rect 5193 4264 5280 4284
tri 5280 4264 5300 4284 sw
rect 5172 4212 5178 4264
rect 5230 4212 5242 4264
rect 5294 4212 5300 4264
rect 3150 4129 3156 4181
rect 3208 4129 3220 4181
rect 3272 4129 3284 4181
rect 3336 4129 3348 4181
rect 3400 4129 3412 4181
rect 3464 4129 3476 4181
rect 3528 4129 3540 4181
rect 3592 4129 3598 4181
rect 3150 4106 3598 4129
rect 3150 4054 3156 4106
rect 3208 4054 3220 4106
rect 3272 4054 3284 4106
rect 3336 4054 3348 4106
rect 3400 4054 3412 4106
rect 3464 4054 3476 4106
rect 3528 4054 3540 4106
rect 3592 4054 3598 4106
rect 3150 4031 3598 4054
rect 3150 3987 3156 4031
rect 3208 3987 3220 4031
rect 3272 3987 3284 4031
rect 3336 3987 3348 4031
rect 3400 3987 3412 4031
rect 3464 3987 3476 4031
rect 3528 3987 3540 4031
rect 3592 3987 3598 4031
rect 3150 3931 3154 3987
rect 3210 3979 3220 3987
rect 3336 3979 3346 3987
rect 3402 3979 3412 3987
rect 3528 3979 3538 3987
rect 3210 3931 3250 3979
rect 3306 3931 3346 3979
rect 3402 3931 3442 3979
rect 3498 3931 3538 3979
rect 3594 3931 3598 3987
rect 3150 3906 3598 3931
rect 3150 3850 3154 3906
rect 3210 3850 3250 3906
rect 3306 3850 3346 3906
rect 3402 3850 3442 3906
rect 3498 3850 3538 3906
rect 3594 3850 3598 3906
rect 3150 3825 3598 3850
rect 3150 3769 3154 3825
rect 3210 3769 3250 3825
rect 3306 3769 3346 3825
rect 3402 3769 3442 3825
rect 3498 3769 3538 3825
rect 3594 3769 3598 3825
rect 3150 3744 3598 3769
rect 3150 3688 3154 3744
rect 3210 3688 3250 3744
rect 3306 3688 3346 3744
rect 3402 3688 3442 3744
rect 3498 3688 3538 3744
rect 3594 3688 3598 3744
rect 3150 3663 3598 3688
rect 3150 3607 3154 3663
rect 3210 3607 3250 3663
rect 3306 3607 3346 3663
rect 3402 3607 3442 3663
rect 3498 3607 3538 3663
rect 3594 3607 3598 3663
rect 3150 3582 3598 3607
rect 3150 3526 3154 3582
rect 3210 3526 3250 3582
rect 3306 3526 3346 3582
rect 3402 3526 3442 3582
rect 3498 3526 3538 3582
rect 3594 3526 3598 3582
rect 3150 3501 3598 3526
rect 3150 3445 3154 3501
rect 3210 3445 3250 3501
rect 3306 3445 3346 3501
rect 3402 3445 3442 3501
rect 3498 3445 3538 3501
rect 3594 3445 3598 3501
rect 3150 3420 3598 3445
rect 3150 3364 3154 3420
rect 3210 3364 3250 3420
rect 3306 3364 3346 3420
rect 3402 3364 3442 3420
rect 3498 3364 3538 3420
rect 3594 3364 3598 3420
rect 3150 3339 3598 3364
tri 2419 3297 2448 3326 sw
rect 2367 3292 2448 3297
tri 2448 3292 2453 3297 sw
rect 2367 3240 2373 3292
rect 2425 3240 2437 3292
rect 2489 3240 2495 3292
rect 3150 3283 3154 3339
rect 3210 3283 3250 3339
rect 3306 3283 3346 3339
rect 3402 3283 3442 3339
rect 3498 3283 3538 3339
rect 3594 3283 3598 3339
rect 7010 3349 7062 4342
tri 7062 4320 7084 4342 nw
tri 7062 3349 7070 3357 sw
rect 7010 3303 7070 3349
tri 7070 3303 7116 3349 sw
tri 7004 3297 7010 3303 se
rect 7010 3297 7116 3303
tri 7116 3297 7122 3303 sw
rect 3150 3258 3598 3283
rect 1698 3005 1704 3057
rect 1756 3005 1773 3057
rect 1825 3005 1842 3057
rect 1894 3005 1911 3057
rect 1963 3005 1980 3057
rect 2032 3005 2038 3057
rect 1698 2981 2038 3005
rect 1698 2929 1704 2981
rect 1756 2929 1773 2981
rect 1825 2929 1842 2981
rect 1894 2929 1911 2981
rect 1963 2929 1980 2981
rect 2032 2929 2038 2981
rect 986 2034 1279 2718
tri 1279 2555 1442 2718 nw
rect 1698 2442 2038 2929
rect 1698 2390 1704 2442
rect 1756 2390 1773 2442
rect 1825 2390 1842 2442
rect 1894 2390 1911 2442
rect 1963 2390 1980 2442
rect 2032 2390 2038 2442
rect 1698 2364 2038 2390
rect 1698 2312 1704 2364
rect 1756 2312 1773 2364
rect 1825 2312 1842 2364
rect 1894 2312 1911 2364
rect 1963 2312 1980 2364
rect 2032 2312 2038 2364
tri 1279 2034 1422 2177 sw
rect 986 1503 1531 2034
rect 1698 2029 2038 2312
rect 1698 1977 1704 2029
rect 1756 1977 1773 2029
rect 1825 1977 1842 2029
rect 1894 1977 1911 2029
rect 1963 1977 1980 2029
rect 2032 1977 2038 2029
rect 1698 1955 2038 1977
rect 1698 1903 1704 1955
rect 1756 1903 1773 1955
rect 1825 1903 1842 1955
rect 1894 1903 1911 1955
rect 1963 1903 1980 1955
rect 2032 1903 2038 1955
rect 1698 1881 2038 1903
rect 1698 1829 1704 1881
rect 1756 1829 1773 1881
rect 1825 1829 1842 1881
rect 1894 1829 1911 1881
rect 1963 1829 1980 1881
rect 2032 1829 2038 1881
rect 1698 1828 2038 1829
rect 3150 3202 3154 3258
rect 3210 3202 3250 3258
rect 3306 3202 3346 3258
rect 3402 3202 3442 3258
rect 3498 3202 3538 3258
rect 3594 3202 3598 3258
tri 6999 3292 7004 3297 se
rect 7004 3292 7122 3297
tri 7122 3292 7127 3297 sw
rect 6999 3240 7005 3292
rect 7057 3240 7069 3292
rect 7121 3240 7127 3292
rect 3150 3177 3598 3202
rect 3150 3121 3154 3177
rect 3210 3121 3250 3177
rect 3306 3121 3346 3177
rect 3402 3121 3442 3177
rect 3498 3121 3538 3177
rect 3594 3121 3598 3177
rect 3150 3096 3598 3121
rect 3150 3040 3154 3096
rect 3210 3057 3250 3096
rect 3306 3057 3346 3096
rect 3402 3057 3442 3096
rect 3498 3057 3538 3096
rect 3210 3040 3220 3057
rect 3336 3040 3346 3057
rect 3402 3040 3412 3057
rect 3528 3040 3538 3057
rect 3594 3040 3598 3096
rect 3150 3015 3156 3040
rect 3208 3015 3220 3040
rect 3272 3015 3284 3040
rect 3336 3015 3348 3040
rect 3400 3015 3412 3040
rect 3464 3015 3476 3040
rect 3528 3015 3540 3040
rect 3592 3015 3598 3040
rect 3150 2959 3154 3015
rect 3210 3005 3220 3015
rect 3336 3005 3346 3015
rect 3402 3005 3412 3015
rect 3528 3005 3538 3015
rect 3210 2981 3250 3005
rect 3306 2981 3346 3005
rect 3402 2981 3442 3005
rect 3498 2981 3538 3005
rect 3210 2959 3220 2981
rect 3336 2959 3346 2981
rect 3402 2959 3412 2981
rect 3528 2959 3538 2981
rect 3594 2959 3598 3015
rect 3150 2934 3156 2959
rect 3208 2934 3220 2959
rect 3272 2934 3284 2959
rect 3336 2934 3348 2959
rect 3400 2934 3412 2959
rect 3464 2934 3476 2959
rect 3528 2934 3540 2959
rect 3592 2934 3598 2959
tri 7359 2947 7360 2948 se
rect 7360 2947 7412 4479
tri 7412 4457 7454 4499 nw
tri 7886 4473 7912 4499 se
rect 7912 4473 7960 4499
tri 7960 4473 7986 4499 nw
tri 7871 4458 7886 4473 se
rect 7886 4458 7945 4473
tri 7945 4458 7960 4473 nw
tri 7870 4457 7871 4458 se
rect 7871 4457 7902 4458
tri 7828 4415 7870 4457 se
rect 7870 4415 7902 4457
tri 7902 4415 7945 4458 nw
tri 7794 4261 7828 4295 se
rect 7828 4261 7880 4415
tri 7880 4393 7902 4415 nw
rect 9493 4393 9541 5224
tri 10487 5207 10504 5224 se
rect 10504 5207 11319 5224
tri 11319 5207 11336 5224 sw
tri 10448 5168 10487 5207 se
rect 10487 5190 11336 5207
rect 10487 5168 10522 5190
tri 10522 5168 10544 5190 nw
tri 11279 5168 11301 5190 ne
rect 11301 5168 11336 5190
tri 10413 5133 10448 5168 se
rect 10448 5133 10487 5168
tri 10487 5133 10522 5168 nw
tri 11301 5133 11336 5168 ne
tri 11336 5133 11410 5207 sw
tri 10374 5094 10413 5133 se
rect 10413 5094 10448 5133
tri 10448 5094 10487 5133 nw
tri 11336 5094 11375 5133 ne
rect 11375 5094 11410 5133
tri 10339 5059 10374 5094 se
rect 10374 5059 10413 5094
tri 10413 5059 10448 5094 nw
tri 11375 5059 11410 5094 ne
tri 11410 5059 11484 5133 sw
tri 10300 5020 10339 5059 se
rect 10339 5020 10374 5059
tri 10374 5020 10413 5059 nw
tri 11410 5020 11449 5059 ne
rect 11449 5020 11484 5059
tri 10271 4991 10300 5020 se
rect 10300 4991 10345 5020
tri 10345 4991 10374 5020 nw
tri 11449 4991 11478 5020 ne
rect 11478 4991 11484 5020
tri 11484 4991 11552 5059 sw
tri 10265 4985 10271 4991 se
rect 10271 4985 10339 4991
tri 10339 4985 10345 4991 nw
tri 11478 4985 11484 4991 ne
rect 11484 4985 11552 4991
tri 11552 4985 11558 4991 sw
tri 10237 4957 10265 4985 se
rect 10265 4957 10311 4985
tri 10311 4957 10339 4985 nw
tri 11484 4957 11512 4985 ne
rect 11512 4957 11558 4985
rect 10237 4939 10293 4957
tri 10293 4939 10311 4957 nw
tri 11512 4939 11530 4957 ne
rect 11530 4939 11558 4957
tri 11558 4939 11604 4985 sw
tri 10184 4678 10237 4731 se
rect 10237 4678 10289 4939
tri 10289 4935 10293 4939 nw
tri 11530 4935 11534 4939 ne
rect 11534 4935 11604 4939
tri 11534 4916 11553 4935 ne
rect 11553 4916 11604 4935
tri 11604 4916 11627 4939 sw
tri 11553 4911 11558 4916 ne
rect 11558 4911 11627 4916
tri 11627 4911 11632 4916 sw
tri 11558 4889 11580 4911 ne
tri 10289 4678 10312 4701 sw
rect 9930 4626 9936 4678
rect 9988 4626 10000 4678
rect 10052 4626 10058 4678
rect 10184 4626 10190 4678
rect 10242 4626 10254 4678
rect 10306 4626 10312 4678
rect 11580 4637 11632 4911
tri 11632 4637 11636 4641 sw
rect 11580 4626 11636 4637
tri 11636 4626 11647 4637 sw
rect 9930 4529 10058 4626
rect 11580 4596 11647 4626
tri 11647 4596 11677 4626 sw
rect 11580 4544 11621 4596
rect 11673 4544 11685 4596
rect 11737 4544 11743 4596
tri 9930 4505 9954 4529 ne
rect 9954 4505 10058 4529
tri 9954 4499 9960 4505 ne
rect 9960 4499 10058 4505
tri 9960 4458 10001 4499 ne
rect 10001 4426 10058 4499
tri 9541 4393 9543 4395 sw
rect 9493 4391 9543 4393
tri 9543 4391 9545 4393 sw
rect 9493 4375 9545 4391
tri 9493 4323 9545 4375 ne
tri 9545 4323 9613 4391 sw
tri 9545 4261 9607 4323 ne
rect 9607 4261 9613 4323
tri 9613 4261 9675 4323 sw
tri 9607 4255 9613 4261 ne
rect 9613 4255 9675 4261
tri 9675 4255 9681 4261 sw
tri 9613 4187 9681 4255 ne
tri 9681 4187 9749 4255 sw
tri 9681 4119 9749 4187 ne
tri 9749 4119 9817 4187 sw
tri 9749 4051 9817 4119 ne
tri 9817 4051 9885 4119 sw
tri 9817 4031 9837 4051 ne
rect 8031 3899 8037 3951
rect 8089 3899 8101 3951
rect 8153 3899 8159 3951
tri 8031 3897 8033 3899 ne
rect 8033 3897 8157 3899
tri 8157 3897 8159 3899 nw
rect 3150 2878 3154 2934
rect 3210 2929 3220 2934
rect 3336 2929 3346 2934
rect 3402 2929 3412 2934
rect 3528 2929 3538 2934
rect 3210 2878 3250 2929
rect 3306 2878 3346 2929
rect 3402 2878 3442 2929
rect 3498 2878 3538 2929
rect 3594 2878 3598 2934
tri 7326 2914 7359 2947 se
rect 7359 2914 7412 2947
rect 3150 2853 3598 2878
rect 3150 2797 3154 2853
rect 3210 2797 3250 2853
rect 3306 2797 3346 2853
rect 3402 2797 3442 2853
rect 3498 2797 3538 2853
rect 3594 2797 3598 2853
rect 3150 2772 3598 2797
rect 3150 2716 3154 2772
rect 3210 2716 3250 2772
rect 3306 2716 3346 2772
rect 3402 2716 3442 2772
rect 3498 2716 3538 2772
rect 3594 2716 3598 2772
rect 3150 2691 3598 2716
rect 3150 2635 3154 2691
rect 3210 2635 3250 2691
rect 3306 2635 3346 2691
rect 3402 2635 3442 2691
rect 3498 2635 3538 2691
rect 3594 2635 3598 2691
rect 7163 2862 7412 2914
rect 8033 3893 8153 3897
tri 8153 3893 8157 3897 nw
rect 8033 3881 8141 3893
tri 8141 3881 8153 3893 nw
rect 8033 3829 8089 3881
tri 8089 3829 8141 3881 nw
rect 7163 2848 7235 2862
tri 7235 2848 7249 2862 nw
rect 7163 2842 7229 2848
tri 7229 2842 7235 2848 nw
rect 7163 2830 7217 2842
tri 7217 2830 7229 2842 nw
tri 7129 2656 7163 2690 se
rect 7163 2656 7215 2830
tri 7215 2828 7217 2830 nw
rect 3150 2610 3598 2635
rect 3150 2554 3154 2610
rect 3210 2554 3250 2610
rect 3306 2554 3346 2610
rect 3402 2554 3442 2610
rect 3498 2554 3538 2610
rect 3594 2554 3598 2610
rect 3150 2529 3598 2554
rect 3150 2473 3154 2529
rect 3210 2473 3250 2529
rect 3306 2473 3346 2529
rect 3402 2473 3442 2529
rect 3498 2473 3538 2529
rect 3594 2473 3598 2529
rect 3150 2447 3598 2473
rect 3150 2391 3154 2447
rect 3210 2442 3250 2447
rect 3306 2442 3346 2447
rect 3402 2442 3442 2447
rect 3498 2442 3538 2447
rect 3210 2391 3220 2442
rect 3336 2391 3346 2442
rect 3402 2391 3412 2442
rect 3528 2391 3538 2442
rect 3594 2391 3598 2447
rect 3150 2390 3156 2391
rect 3208 2390 3220 2391
rect 3272 2390 3284 2391
rect 3336 2390 3348 2391
rect 3400 2390 3412 2391
rect 3464 2390 3476 2391
rect 3528 2390 3540 2391
rect 3592 2390 3598 2391
rect 3150 2365 3598 2390
rect 3150 2309 3154 2365
rect 3210 2364 3250 2365
rect 3306 2364 3346 2365
rect 3402 2364 3442 2365
rect 3498 2364 3538 2365
rect 3210 2312 3220 2364
rect 3336 2312 3346 2364
rect 3402 2312 3412 2364
rect 3528 2312 3538 2364
rect 3210 2309 3250 2312
rect 3306 2309 3346 2312
rect 3402 2309 3442 2312
rect 3498 2309 3538 2312
rect 3594 2309 3598 2365
rect 3150 2283 3598 2309
rect 3150 2227 3154 2283
rect 3210 2227 3250 2283
rect 3306 2227 3346 2283
rect 3402 2227 3442 2283
rect 3498 2227 3538 2283
rect 3594 2227 3598 2283
rect 3150 2201 3598 2227
rect 3150 2145 3154 2201
rect 3210 2145 3250 2201
rect 3306 2145 3346 2201
rect 3402 2145 3442 2201
rect 3498 2145 3538 2201
rect 3594 2145 3598 2201
rect 3150 2119 3598 2145
rect 3150 2063 3154 2119
rect 3210 2063 3250 2119
rect 3306 2063 3346 2119
rect 3402 2063 3442 2119
rect 3498 2063 3538 2119
rect 3594 2063 3598 2119
rect 3150 2037 3598 2063
rect 3150 1981 3154 2037
rect 3210 2029 3250 2037
rect 3306 2029 3346 2037
rect 3402 2029 3442 2037
rect 3498 2029 3538 2037
rect 3210 1981 3220 2029
rect 3336 1981 3346 2029
rect 3402 1981 3412 2029
rect 3528 1981 3538 2029
rect 3594 1981 3598 2037
rect 3150 1977 3156 1981
rect 3208 1977 3220 1981
rect 3272 1977 3284 1981
rect 3336 1977 3348 1981
rect 3400 1977 3412 1981
rect 3464 1977 3476 1981
rect 3528 1977 3540 1981
rect 3592 1977 3598 1981
rect 3150 1955 3598 1977
rect 3150 1899 3154 1955
rect 3210 1903 3220 1955
rect 3336 1903 3346 1955
rect 3402 1903 3412 1955
rect 3528 1903 3538 1955
rect 3210 1899 3250 1903
rect 3306 1899 3346 1903
rect 3402 1899 3442 1903
rect 3498 1899 3538 1903
rect 3594 1899 3598 1955
rect 3150 1881 3598 1899
rect 3150 1873 3156 1881
rect 3208 1873 3220 1881
rect 3272 1873 3284 1881
rect 3336 1873 3348 1881
rect 3400 1873 3412 1881
rect 3464 1873 3476 1881
rect 3528 1873 3540 1881
rect 3592 1873 3598 1881
rect 3150 1817 3154 1873
rect 3210 1829 3220 1873
rect 3336 1829 3346 1873
rect 3402 1829 3412 1873
rect 3528 1829 3538 1873
rect 3210 1817 3250 1829
rect 3306 1817 3346 1829
rect 3402 1817 3442 1829
rect 3498 1817 3538 1829
rect 3594 1817 3598 1873
rect 3150 1791 3598 1817
rect 3150 1735 3154 1791
rect 3210 1735 3250 1791
rect 3306 1735 3346 1791
rect 3402 1735 3442 1791
rect 3498 1735 3538 1791
rect 3594 1735 3598 1791
rect 3150 1709 3598 1735
rect 3150 1653 3154 1709
rect 3210 1653 3250 1709
rect 3306 1653 3346 1709
rect 3402 1653 3442 1709
rect 3498 1653 3538 1709
rect 3594 1653 3598 1709
rect 3150 1644 3598 1653
tri 7991 1658 8033 1700 se
rect 8033 1658 8084 3829
tri 8084 3824 8089 3829 nw
rect 9837 3769 9885 4051
rect 10001 3945 10053 4426
tri 10053 4421 10058 4426 nw
rect 10001 3881 10053 3893
rect 10001 3823 10053 3829
tri 9837 3758 9848 3769 ne
rect 9848 3758 9885 3769
tri 9885 3758 9909 3782 sw
tri 9848 3721 9885 3758 ne
rect 9885 3721 9909 3758
tri 9885 3704 9902 3721 ne
rect 9902 3704 9909 3721
tri 9909 3704 9963 3758 sw
tri 9902 3697 9909 3704 ne
rect 9909 3697 9963 3704
tri 9963 3697 9970 3704 sw
tri 9909 3652 9954 3697 ne
rect 9954 3652 9970 3697
tri 9970 3652 10015 3697 sw
tri 9954 3638 9968 3652 ne
rect 9968 3638 10015 3652
tri 10015 3638 10029 3652 sw
tri 9968 3636 9970 3638 ne
rect 9970 3636 10029 3638
tri 10029 3636 10031 3638 sw
tri 9970 3623 9983 3636 ne
rect 9983 3048 10031 3636
tri 9983 3020 10011 3048 ne
rect 10011 3020 10031 3048
tri 10031 3020 10079 3068 sw
tri 10011 3000 10031 3020 ne
rect 10031 3000 10140 3020
tri 10031 2993 10038 3000 ne
rect 10038 2993 10140 3000
tri 10140 2993 10167 3020 sw
tri 10038 2972 10059 2993 ne
rect 10059 2972 10167 2993
tri 10120 2925 10167 2972 ne
tri 10167 2925 10235 2993 sw
rect 10167 2900 10235 2925
tri 10235 2900 10260 2925 sw
rect 10167 2848 10173 2900
rect 10225 2848 10237 2900
rect 10289 2848 10295 2900
rect 12073 2894 12125 5443
tri 12125 5409 12159 5443 nw
tri 12209 5409 12232 5432 se
rect 12232 5409 12284 5519
tri 12284 5512 12318 5546 nw
tri 12284 5409 12307 5432 sw
tri 12198 5398 12209 5409 se
rect 12209 5398 12307 5409
tri 12307 5398 12318 5409 sw
rect 12194 5346 12200 5398
rect 12252 5346 12264 5398
rect 12316 5346 12322 5398
rect 13335 4939 13341 4991
rect 13393 4939 13413 4991
rect 13465 4939 13484 4991
rect 13536 4939 13555 4991
rect 13607 4939 13626 4991
rect 13678 4939 13684 4991
rect 13335 4916 13684 4939
rect 13335 4864 13341 4916
rect 13393 4864 13413 4916
rect 13465 4864 13484 4916
rect 13536 4864 13555 4916
rect 13607 4864 13626 4916
rect 13678 4864 13684 4916
rect 13335 4841 13684 4864
rect 13335 4789 13341 4841
rect 13393 4789 13413 4841
rect 13465 4789 13484 4841
rect 13536 4789 13555 4841
rect 13607 4789 13626 4841
rect 13678 4789 13684 4841
rect 12073 2830 12125 2842
rect 12073 2772 12125 2778
rect 12153 4585 12159 4637
rect 12211 4585 12224 4637
rect 12276 4585 12282 4637
rect 12153 4557 12214 4585
tri 12214 4557 12242 4585 nw
rect 10919 2470 10967 2522
rect 11401 2065 11449 2117
tri 8084 1658 8119 1693 sw
rect 7991 1606 7997 1658
rect 8049 1606 8061 1658
rect 8113 1606 8119 1658
rect 986 1451 992 1503
rect 1044 1451 1061 1503
rect 1113 1451 1130 1503
rect 1182 1451 1199 1503
rect 1251 1451 1268 1503
rect 1320 1451 1337 1503
rect 1389 1451 1405 1503
rect 1457 1451 1473 1503
rect 1525 1451 1531 1503
rect 986 1429 1531 1451
rect 986 1377 992 1429
rect 1044 1377 1061 1429
rect 1113 1377 1130 1429
rect 1182 1377 1199 1429
rect 1251 1377 1268 1429
rect 1320 1377 1337 1429
rect 1389 1377 1405 1429
rect 1457 1377 1473 1429
rect 1525 1377 1531 1429
rect 986 1355 1531 1377
rect 986 1303 992 1355
rect 1044 1303 1061 1355
rect 1113 1303 1130 1355
rect 1182 1303 1199 1355
rect 1251 1303 1268 1355
rect 1320 1303 1337 1355
rect 1389 1303 1405 1355
rect 1457 1303 1473 1355
rect 1525 1303 1531 1355
rect 986 790 1531 1303
rect 12153 1090 12205 4557
tri 12205 4548 12214 4557 nw
rect 13335 3704 13684 4789
rect 14684 4585 14690 4637
rect 14742 4585 14754 4637
rect 14806 4585 14812 4637
tri 14726 4557 14754 4585 ne
rect 14754 4557 14812 4585
rect 14585 4505 14591 4557
rect 14643 4505 14655 4557
rect 14707 4505 14713 4557
tri 14754 4551 14760 4557 ne
tri 14604 4474 14635 4505 ne
rect 14635 4100 14687 4505
tri 14687 4479 14713 4505 nw
tri 14726 3866 14760 3900 se
rect 14760 3866 14812 4557
rect 13335 3652 13338 3704
rect 13390 3652 13411 3704
rect 13463 3652 13484 3704
rect 13536 3652 13557 3704
rect 13609 3652 13630 3704
rect 13682 3652 13684 3704
rect 13335 3638 13684 3652
rect 13335 3586 13338 3638
rect 13390 3586 13411 3638
rect 13463 3586 13484 3638
rect 13536 3586 13557 3638
rect 13609 3586 13630 3638
rect 13682 3586 13684 3638
rect 13335 3572 13684 3586
rect 12886 3560 13216 3566
rect 12886 3508 12887 3560
rect 12939 3508 12956 3560
rect 13008 3508 13025 3560
rect 13077 3508 13094 3560
rect 13146 3508 13163 3560
rect 13215 3508 13216 3560
rect 12886 3490 13216 3508
rect 12886 3438 12887 3490
rect 12939 3438 12956 3490
rect 13008 3438 13025 3490
rect 13077 3438 13094 3490
rect 13146 3438 13163 3490
rect 13215 3438 13216 3490
rect 12886 3420 13216 3438
rect 12886 3368 12887 3420
rect 12939 3368 12956 3420
rect 13008 3368 13025 3420
rect 13077 3368 13094 3420
rect 13146 3368 13163 3420
rect 13215 3368 13216 3420
rect 12886 3349 13216 3368
rect 12886 3297 12887 3349
rect 12939 3297 12956 3349
rect 13008 3297 13025 3349
rect 13077 3297 13094 3349
rect 13146 3297 13163 3349
rect 13215 3297 13216 3349
rect 12886 3278 13216 3297
rect 12886 3226 12887 3278
rect 12939 3226 12956 3278
rect 13008 3226 13025 3278
rect 13077 3226 13094 3278
rect 13146 3226 13163 3278
rect 13215 3226 13216 3278
rect 12886 1415 13216 3226
rect 13335 3520 13338 3572
rect 13390 3520 13411 3572
rect 13463 3520 13484 3572
rect 13536 3520 13557 3572
rect 13609 3520 13630 3572
rect 13682 3520 13684 3572
rect 13335 3506 13684 3520
rect 13335 3454 13338 3506
rect 13390 3454 13411 3506
rect 13463 3454 13484 3506
rect 13536 3454 13557 3506
rect 13609 3454 13630 3506
rect 13682 3454 13684 3506
rect 13335 3440 13684 3454
rect 13335 3388 13338 3440
rect 13390 3388 13411 3440
rect 13463 3388 13484 3440
rect 13536 3388 13557 3440
rect 13609 3388 13630 3440
rect 13682 3388 13684 3440
rect 13335 3374 13684 3388
rect 13335 3322 13338 3374
rect 13390 3322 13411 3374
rect 13463 3322 13484 3374
rect 13536 3322 13557 3374
rect 13609 3322 13630 3374
rect 13682 3322 13684 3374
rect 13335 3308 13684 3322
rect 13335 3256 13338 3308
rect 13390 3256 13411 3308
rect 13463 3256 13484 3308
rect 13536 3256 13557 3308
rect 13609 3256 13630 3308
rect 13682 3256 13684 3308
rect 13335 3242 13684 3256
rect 13335 3190 13338 3242
rect 13390 3190 13411 3242
rect 13463 3190 13484 3242
rect 13536 3190 13557 3242
rect 13609 3190 13630 3242
rect 13682 3190 13684 3242
rect 13335 3176 13684 3190
rect 13335 3124 13338 3176
rect 13390 3124 13411 3176
rect 13463 3124 13484 3176
rect 13536 3124 13557 3176
rect 13609 3124 13630 3176
rect 13682 3124 13684 3176
rect 13335 3118 13684 3124
rect 14554 3814 14812 3866
rect 14554 3038 14606 3814
tri 14606 3780 14640 3814 nw
rect 12886 1363 12887 1415
rect 12939 1363 12956 1415
rect 13008 1363 13025 1415
rect 13077 1363 13094 1415
rect 13146 1363 13163 1415
rect 13215 1363 13216 1415
rect 12886 1345 13216 1363
rect 12886 1293 12887 1345
rect 12939 1293 12956 1345
rect 13008 1293 13025 1345
rect 13077 1293 13094 1345
rect 13146 1293 13163 1345
rect 13215 1293 13216 1345
rect 12886 1275 13216 1293
rect 12886 1223 12887 1275
rect 12939 1223 12956 1275
rect 13008 1223 13025 1275
rect 13077 1223 13094 1275
rect 13146 1223 13163 1275
rect 13215 1223 13216 1275
rect 12886 1204 13216 1223
rect 12886 1152 12887 1204
rect 12939 1152 12956 1204
rect 13008 1152 13025 1204
rect 13077 1152 13094 1204
rect 13146 1152 13163 1204
rect 13215 1152 13216 1204
rect 12886 1133 13216 1152
rect 12886 1081 12887 1133
rect 12939 1081 12956 1133
rect 13008 1081 13025 1133
rect 13077 1081 13094 1133
rect 13146 1081 13163 1133
rect 13215 1081 13216 1133
rect 12886 1075 13216 1081
rect 12153 1026 12205 1038
rect 12153 968 12205 974
rect 14823 997 14875 1003
rect 10737 888 10743 940
rect 10795 888 10807 940
rect 10859 888 10865 940
rect 14823 931 14875 945
rect 986 738 992 790
rect 1044 738 1061 790
rect 1113 738 1130 790
rect 1182 738 1199 790
rect 1251 738 1268 790
rect 1320 738 1337 790
rect 1389 738 1405 790
rect 1457 738 1473 790
rect 1525 738 1531 790
rect 986 696 1531 738
rect 986 644 992 696
rect 1044 644 1061 696
rect 1113 644 1130 696
rect 1182 644 1199 696
rect 1251 644 1268 696
rect 1320 644 1337 696
rect 1389 644 1405 696
rect 1457 644 1473 696
rect 1525 644 1531 696
rect 986 643 1531 644
rect 12255 591 12264 647
rect 12320 591 12344 647
rect 12400 592 12423 647
rect 12255 540 12363 591
rect 12415 540 12423 592
tri 14812 563 14823 574 se
rect 14823 563 14875 879
rect 12255 528 12423 540
rect 12255 504 12363 528
tri 12255 476 12283 504 ne
rect 12283 476 12363 504
rect 12415 476 12423 528
rect 12786 514 12812 563
tri 14789 540 14812 563 se
rect 14812 540 14875 563
tri 12283 466 12293 476 ne
rect 12293 466 12423 476
tri 12745 405 12773 433 se
rect 12773 411 12825 505
rect 13257 485 13306 500
rect 12773 405 12819 411
tri 12819 405 12825 411 nw
tri -155 379 -129 405 se
rect -129 386 -74 405
rect -129 379 -123 386
tri -389 341 -351 379 se
rect -351 341 -315 379
tri -315 341 -277 379 nw
tri -193 341 -155 379 se
rect -155 341 -123 379
rect -389 340 -316 341
tri -316 340 -315 341 nw
tri -194 340 -193 341 se
rect -193 340 -123 341
rect -389 50 -333 340
tri -333 323 -316 340 nw
tri -197 337 -194 340 se
rect -194 337 -123 340
tri -123 337 -74 386 nw
rect 12334 379 12793 405
tri 12793 379 12819 405 nw
rect 12334 362 12767 379
rect -197 323 -137 337
tri -137 323 -123 337 nw
rect -389 -30 -333 -6
rect -389 -95 -333 -86
rect -197 -95 -145 323
tri -145 315 -137 323 nw
rect 12390 353 12767 362
tri 12767 353 12793 379 nw
rect 12390 341 12420 353
tri 12420 341 12432 353 nw
rect 12390 340 12419 341
tri 12419 340 12420 341 nw
rect 12390 323 12402 340
tri 12402 323 12419 340 nw
tri 13238 323 13255 340 se
rect 13255 323 13307 485
rect 13425 445 13474 498
rect 14747 488 14753 540
rect 14805 488 14817 540
rect 14869 488 14875 540
rect 13617 397 13652 442
rect 13789 394 13823 443
rect 14263 399 14307 448
tri 12390 311 12402 323 nw
tri 13226 311 13238 323 se
rect 13238 318 13307 323
rect 13238 311 13296 318
tri 13222 307 13226 311 se
rect 13226 307 13296 311
tri 13296 307 13307 318 nw
rect 12334 282 12390 306
rect 12428 255 12434 307
rect 12486 255 12498 307
rect 12550 255 13244 307
tri 13244 255 13296 307 nw
rect 12334 217 12390 226
tri -145 -95 -124 -74 sw
rect -197 -96 -124 -95
tri -124 -96 -123 -95 sw
tri -197 -170 -123 -96 ne
tri -123 -155 -64 -96 sw
rect -123 -170 -64 -155
tri -64 -170 -49 -155 sw
tri -123 -213 -80 -170 ne
rect -80 -207 -49 -170
tri -49 -207 -12 -170 sw
rect -80 -213 -12 -207
tri -80 -229 -64 -213 ne
tri -138 -1219 -64 -1145 se
rect -64 -1167 -12 -213
tri 11400 -315 11502 -213 sw
rect 11348 -371 11357 -315
rect 11413 -371 11437 -315
rect 11493 -371 11502 -315
tri 11400 -473 11502 -371 nw
tri -64 -1219 -12 -1167 nw
tri -197 -1278 -138 -1219 se
rect -138 -1278 -123 -1219
tri -123 -1278 -64 -1219 nw
rect -197 -1529 -145 -1278
tri -145 -1300 -123 -1278 nw
tri -145 -1529 -99 -1483 sw
tri -200 -1532 -197 -1529 se
rect -197 -1532 -99 -1529
tri -99 -1532 -96 -1529 sw
rect -200 -1588 -191 -1532
rect -135 -1588 -111 -1532
rect -55 -1588 -46 -1532
<< via2 >>
rect -374 631 -318 687
rect -374 551 -318 607
rect 3154 3979 3156 3987
rect 3156 3979 3208 3987
rect 3208 3979 3210 3987
rect 3250 3979 3272 3987
rect 3272 3979 3284 3987
rect 3284 3979 3306 3987
rect 3346 3979 3348 3987
rect 3348 3979 3400 3987
rect 3400 3979 3402 3987
rect 3442 3979 3464 3987
rect 3464 3979 3476 3987
rect 3476 3979 3498 3987
rect 3538 3979 3540 3987
rect 3540 3979 3592 3987
rect 3592 3979 3594 3987
rect 3154 3931 3210 3979
rect 3250 3931 3306 3979
rect 3346 3931 3402 3979
rect 3442 3931 3498 3979
rect 3538 3931 3594 3979
rect 3154 3850 3210 3906
rect 3250 3850 3306 3906
rect 3346 3850 3402 3906
rect 3442 3850 3498 3906
rect 3538 3850 3594 3906
rect 3154 3769 3210 3825
rect 3250 3769 3306 3825
rect 3346 3769 3402 3825
rect 3442 3769 3498 3825
rect 3538 3769 3594 3825
rect 3154 3688 3210 3744
rect 3250 3688 3306 3744
rect 3346 3688 3402 3744
rect 3442 3688 3498 3744
rect 3538 3688 3594 3744
rect 3154 3607 3210 3663
rect 3250 3607 3306 3663
rect 3346 3607 3402 3663
rect 3442 3607 3498 3663
rect 3538 3607 3594 3663
rect 3154 3526 3210 3582
rect 3250 3526 3306 3582
rect 3346 3526 3402 3582
rect 3442 3526 3498 3582
rect 3538 3526 3594 3582
rect 3154 3445 3210 3501
rect 3250 3445 3306 3501
rect 3346 3445 3402 3501
rect 3442 3445 3498 3501
rect 3538 3445 3594 3501
rect 3154 3364 3210 3420
rect 3250 3364 3306 3420
rect 3346 3364 3402 3420
rect 3442 3364 3498 3420
rect 3538 3364 3594 3420
rect 3154 3283 3210 3339
rect 3250 3283 3306 3339
rect 3346 3283 3402 3339
rect 3442 3283 3498 3339
rect 3538 3283 3594 3339
rect 3154 3202 3210 3258
rect 3250 3202 3306 3258
rect 3346 3202 3402 3258
rect 3442 3202 3498 3258
rect 3538 3202 3594 3258
rect 3154 3121 3210 3177
rect 3250 3121 3306 3177
rect 3346 3121 3402 3177
rect 3442 3121 3498 3177
rect 3538 3121 3594 3177
rect 3154 3057 3210 3096
rect 3250 3057 3306 3096
rect 3346 3057 3402 3096
rect 3442 3057 3498 3096
rect 3538 3057 3594 3096
rect 3154 3040 3156 3057
rect 3156 3040 3208 3057
rect 3208 3040 3210 3057
rect 3250 3040 3272 3057
rect 3272 3040 3284 3057
rect 3284 3040 3306 3057
rect 3346 3040 3348 3057
rect 3348 3040 3400 3057
rect 3400 3040 3402 3057
rect 3442 3040 3464 3057
rect 3464 3040 3476 3057
rect 3476 3040 3498 3057
rect 3538 3040 3540 3057
rect 3540 3040 3592 3057
rect 3592 3040 3594 3057
rect 3154 3005 3156 3015
rect 3156 3005 3208 3015
rect 3208 3005 3210 3015
rect 3250 3005 3272 3015
rect 3272 3005 3284 3015
rect 3284 3005 3306 3015
rect 3346 3005 3348 3015
rect 3348 3005 3400 3015
rect 3400 3005 3402 3015
rect 3442 3005 3464 3015
rect 3464 3005 3476 3015
rect 3476 3005 3498 3015
rect 3538 3005 3540 3015
rect 3540 3005 3592 3015
rect 3592 3005 3594 3015
rect 3154 2981 3210 3005
rect 3250 2981 3306 3005
rect 3346 2981 3402 3005
rect 3442 2981 3498 3005
rect 3538 2981 3594 3005
rect 3154 2959 3156 2981
rect 3156 2959 3208 2981
rect 3208 2959 3210 2981
rect 3250 2959 3272 2981
rect 3272 2959 3284 2981
rect 3284 2959 3306 2981
rect 3346 2959 3348 2981
rect 3348 2959 3400 2981
rect 3400 2959 3402 2981
rect 3442 2959 3464 2981
rect 3464 2959 3476 2981
rect 3476 2959 3498 2981
rect 3538 2959 3540 2981
rect 3540 2959 3592 2981
rect 3592 2959 3594 2981
rect 3154 2929 3156 2934
rect 3156 2929 3208 2934
rect 3208 2929 3210 2934
rect 3250 2929 3272 2934
rect 3272 2929 3284 2934
rect 3284 2929 3306 2934
rect 3346 2929 3348 2934
rect 3348 2929 3400 2934
rect 3400 2929 3402 2934
rect 3442 2929 3464 2934
rect 3464 2929 3476 2934
rect 3476 2929 3498 2934
rect 3538 2929 3540 2934
rect 3540 2929 3592 2934
rect 3592 2929 3594 2934
rect 3154 2878 3210 2929
rect 3250 2878 3306 2929
rect 3346 2878 3402 2929
rect 3442 2878 3498 2929
rect 3538 2878 3594 2929
rect 3154 2797 3210 2853
rect 3250 2797 3306 2853
rect 3346 2797 3402 2853
rect 3442 2797 3498 2853
rect 3538 2797 3594 2853
rect 3154 2716 3210 2772
rect 3250 2716 3306 2772
rect 3346 2716 3402 2772
rect 3442 2716 3498 2772
rect 3538 2716 3594 2772
rect 3154 2635 3210 2691
rect 3250 2635 3306 2691
rect 3346 2635 3402 2691
rect 3442 2635 3498 2691
rect 3538 2635 3594 2691
rect 3154 2554 3210 2610
rect 3250 2554 3306 2610
rect 3346 2554 3402 2610
rect 3442 2554 3498 2610
rect 3538 2554 3594 2610
rect 3154 2473 3210 2529
rect 3250 2473 3306 2529
rect 3346 2473 3402 2529
rect 3442 2473 3498 2529
rect 3538 2473 3594 2529
rect 3154 2442 3210 2447
rect 3250 2442 3306 2447
rect 3346 2442 3402 2447
rect 3442 2442 3498 2447
rect 3538 2442 3594 2447
rect 3154 2391 3156 2442
rect 3156 2391 3208 2442
rect 3208 2391 3210 2442
rect 3250 2391 3272 2442
rect 3272 2391 3284 2442
rect 3284 2391 3306 2442
rect 3346 2391 3348 2442
rect 3348 2391 3400 2442
rect 3400 2391 3402 2442
rect 3442 2391 3464 2442
rect 3464 2391 3476 2442
rect 3476 2391 3498 2442
rect 3538 2391 3540 2442
rect 3540 2391 3592 2442
rect 3592 2391 3594 2442
rect 3154 2364 3210 2365
rect 3250 2364 3306 2365
rect 3346 2364 3402 2365
rect 3442 2364 3498 2365
rect 3538 2364 3594 2365
rect 3154 2312 3156 2364
rect 3156 2312 3208 2364
rect 3208 2312 3210 2364
rect 3250 2312 3272 2364
rect 3272 2312 3284 2364
rect 3284 2312 3306 2364
rect 3346 2312 3348 2364
rect 3348 2312 3400 2364
rect 3400 2312 3402 2364
rect 3442 2312 3464 2364
rect 3464 2312 3476 2364
rect 3476 2312 3498 2364
rect 3538 2312 3540 2364
rect 3540 2312 3592 2364
rect 3592 2312 3594 2364
rect 3154 2309 3210 2312
rect 3250 2309 3306 2312
rect 3346 2309 3402 2312
rect 3442 2309 3498 2312
rect 3538 2309 3594 2312
rect 3154 2227 3210 2283
rect 3250 2227 3306 2283
rect 3346 2227 3402 2283
rect 3442 2227 3498 2283
rect 3538 2227 3594 2283
rect 3154 2145 3210 2201
rect 3250 2145 3306 2201
rect 3346 2145 3402 2201
rect 3442 2145 3498 2201
rect 3538 2145 3594 2201
rect 3154 2063 3210 2119
rect 3250 2063 3306 2119
rect 3346 2063 3402 2119
rect 3442 2063 3498 2119
rect 3538 2063 3594 2119
rect 3154 2029 3210 2037
rect 3250 2029 3306 2037
rect 3346 2029 3402 2037
rect 3442 2029 3498 2037
rect 3538 2029 3594 2037
rect 3154 1981 3156 2029
rect 3156 1981 3208 2029
rect 3208 1981 3210 2029
rect 3250 1981 3272 2029
rect 3272 1981 3284 2029
rect 3284 1981 3306 2029
rect 3346 1981 3348 2029
rect 3348 1981 3400 2029
rect 3400 1981 3402 2029
rect 3442 1981 3464 2029
rect 3464 1981 3476 2029
rect 3476 1981 3498 2029
rect 3538 1981 3540 2029
rect 3540 1981 3592 2029
rect 3592 1981 3594 2029
rect 3154 1903 3156 1955
rect 3156 1903 3208 1955
rect 3208 1903 3210 1955
rect 3250 1903 3272 1955
rect 3272 1903 3284 1955
rect 3284 1903 3306 1955
rect 3346 1903 3348 1955
rect 3348 1903 3400 1955
rect 3400 1903 3402 1955
rect 3442 1903 3464 1955
rect 3464 1903 3476 1955
rect 3476 1903 3498 1955
rect 3538 1903 3540 1955
rect 3540 1903 3592 1955
rect 3592 1903 3594 1955
rect 3154 1899 3210 1903
rect 3250 1899 3306 1903
rect 3346 1899 3402 1903
rect 3442 1899 3498 1903
rect 3538 1899 3594 1903
rect 3154 1829 3156 1873
rect 3156 1829 3208 1873
rect 3208 1829 3210 1873
rect 3250 1829 3272 1873
rect 3272 1829 3284 1873
rect 3284 1829 3306 1873
rect 3346 1829 3348 1873
rect 3348 1829 3400 1873
rect 3400 1829 3402 1873
rect 3442 1829 3464 1873
rect 3464 1829 3476 1873
rect 3476 1829 3498 1873
rect 3538 1829 3540 1873
rect 3540 1829 3592 1873
rect 3592 1829 3594 1873
rect 3154 1817 3210 1829
rect 3250 1817 3306 1829
rect 3346 1817 3402 1829
rect 3442 1817 3498 1829
rect 3538 1817 3594 1829
rect 3154 1735 3210 1791
rect 3250 1735 3306 1791
rect 3346 1735 3402 1791
rect 3442 1735 3498 1791
rect 3538 1735 3594 1791
rect 3154 1653 3210 1709
rect 3250 1653 3306 1709
rect 3346 1653 3402 1709
rect 3442 1653 3498 1709
rect 3538 1653 3594 1709
rect 12264 591 12320 647
rect 12344 592 12400 647
rect 12344 591 12363 592
rect 12363 591 12400 592
rect -389 -6 -333 50
rect -389 -86 -333 -30
rect 12334 306 12390 362
rect 12334 226 12390 282
rect 11357 -371 11413 -315
rect 11437 -371 11493 -315
rect -191 -1588 -135 -1532
rect -111 -1588 -55 -1532
<< metal3 >>
rect 3146 3987 3602 3992
rect 3146 3931 3154 3987
rect 3210 3931 3250 3987
rect 3306 3931 3346 3987
rect 3402 3931 3442 3987
rect 3498 3931 3538 3987
rect 3594 3931 3602 3987
rect 3146 3906 3602 3931
rect 3146 3850 3154 3906
rect 3210 3850 3250 3906
rect 3306 3850 3346 3906
rect 3402 3850 3442 3906
rect 3498 3850 3538 3906
rect 3594 3850 3602 3906
rect 3146 3825 3602 3850
rect 3146 3769 3154 3825
rect 3210 3769 3250 3825
rect 3306 3769 3346 3825
rect 3402 3769 3442 3825
rect 3498 3769 3538 3825
rect 3594 3769 3602 3825
rect 3146 3744 3602 3769
rect 3146 3688 3154 3744
rect 3210 3688 3250 3744
rect 3306 3688 3346 3744
rect 3402 3688 3442 3744
rect 3498 3688 3538 3744
rect 3594 3688 3602 3744
rect 3146 3663 3602 3688
rect 3146 3607 3154 3663
rect 3210 3607 3250 3663
rect 3306 3607 3346 3663
rect 3402 3607 3442 3663
rect 3498 3607 3538 3663
rect 3594 3607 3602 3663
rect 3146 3582 3602 3607
rect 3146 3526 3154 3582
rect 3210 3526 3250 3582
rect 3306 3526 3346 3582
rect 3402 3526 3442 3582
rect 3498 3526 3538 3582
rect 3594 3526 3602 3582
rect 3146 3501 3602 3526
rect 3146 3445 3154 3501
rect 3210 3445 3250 3501
rect 3306 3445 3346 3501
rect 3402 3445 3442 3501
rect 3498 3445 3538 3501
rect 3594 3445 3602 3501
rect 3146 3420 3602 3445
rect 3146 3364 3154 3420
rect 3210 3364 3250 3420
rect 3306 3364 3346 3420
rect 3402 3364 3442 3420
rect 3498 3364 3538 3420
rect 3594 3364 3602 3420
rect 3146 3339 3602 3364
rect 3146 3283 3154 3339
rect 3210 3283 3250 3339
rect 3306 3283 3346 3339
rect 3402 3283 3442 3339
rect 3498 3283 3538 3339
rect 3594 3283 3602 3339
rect 3146 3258 3602 3283
rect 3146 3202 3154 3258
rect 3210 3202 3250 3258
rect 3306 3202 3346 3258
rect 3402 3202 3442 3258
rect 3498 3202 3538 3258
rect 3594 3202 3602 3258
rect 3146 3177 3602 3202
rect 3146 3121 3154 3177
rect 3210 3121 3250 3177
rect 3306 3121 3346 3177
rect 3402 3121 3442 3177
rect 3498 3121 3538 3177
rect 3594 3121 3602 3177
rect 3146 3096 3602 3121
rect 3146 3040 3154 3096
rect 3210 3040 3250 3096
rect 3306 3040 3346 3096
rect 3402 3040 3442 3096
rect 3498 3040 3538 3096
rect 3594 3040 3602 3096
rect 3146 3015 3602 3040
rect 3146 2959 3154 3015
rect 3210 2959 3250 3015
rect 3306 2959 3346 3015
rect 3402 2959 3442 3015
rect 3498 2959 3538 3015
rect 3594 2959 3602 3015
rect 3146 2934 3602 2959
rect 3146 2554 3154 2934
rect 3210 2895 3250 2934
rect 3306 2895 3346 2934
rect 3402 2895 3442 2934
rect 3498 2895 3538 2934
rect 3218 2831 3248 2895
rect 3312 2831 3342 2895
rect 3406 2831 3436 2895
rect 3500 2831 3530 2895
rect 3210 2809 3250 2831
rect 3306 2809 3346 2831
rect 3402 2809 3442 2831
rect 3498 2809 3538 2831
rect 3218 2745 3248 2809
rect 3312 2745 3342 2809
rect 3406 2745 3436 2809
rect 3500 2745 3530 2809
rect 3210 2723 3250 2745
rect 3306 2723 3346 2745
rect 3402 2723 3442 2745
rect 3498 2723 3538 2745
rect 3218 2659 3248 2723
rect 3312 2659 3342 2723
rect 3406 2659 3436 2723
rect 3500 2659 3530 2723
rect 3210 2637 3250 2659
rect 3306 2637 3346 2659
rect 3402 2637 3442 2659
rect 3498 2637 3538 2659
rect 3218 2573 3248 2637
rect 3312 2573 3342 2637
rect 3406 2573 3436 2637
rect 3500 2573 3530 2637
rect 3210 2554 3250 2573
rect 3306 2554 3346 2573
rect 3402 2554 3442 2573
rect 3498 2554 3538 2573
rect 3594 2554 3602 2934
rect 3146 2551 3602 2554
rect 3146 2473 3154 2551
rect 3218 2487 3248 2551
rect 3312 2487 3342 2551
rect 3406 2487 3436 2551
rect 3500 2487 3530 2551
rect 3210 2473 3250 2487
rect 3306 2473 3346 2487
rect 3402 2473 3442 2487
rect 3498 2473 3538 2487
rect 3594 2473 3602 2551
rect 3146 2465 3602 2473
rect 3146 2391 3154 2465
rect 3218 2401 3248 2465
rect 3312 2401 3342 2465
rect 3406 2401 3436 2465
rect 3500 2401 3530 2465
rect 3210 2391 3250 2401
rect 3306 2391 3346 2401
rect 3402 2391 3442 2401
rect 3498 2391 3538 2401
rect 3594 2391 3602 2465
rect 3146 2379 3602 2391
rect 3146 2309 3154 2379
rect 3218 2315 3248 2379
rect 3312 2315 3342 2379
rect 3406 2315 3436 2379
rect 3500 2315 3530 2379
rect 3210 2309 3250 2315
rect 3306 2309 3346 2315
rect 3402 2309 3442 2315
rect 3498 2309 3538 2315
rect 3594 2309 3602 2379
rect 3146 2292 3602 2309
rect 3146 2227 3154 2292
rect 3218 2228 3248 2292
rect 3312 2228 3342 2292
rect 3406 2228 3436 2292
rect 3500 2228 3530 2292
rect 3210 2227 3250 2228
rect 3306 2227 3346 2228
rect 3402 2227 3442 2228
rect 3498 2227 3538 2228
rect 3594 2227 3602 2292
rect 3146 2205 3602 2227
rect 3146 2141 3154 2205
rect 3218 2141 3248 2205
rect 3312 2141 3342 2205
rect 3406 2141 3436 2205
rect 3500 2141 3530 2205
rect 3594 2141 3602 2205
rect 3146 2119 3602 2141
rect 3146 2054 3154 2119
rect 3210 2118 3250 2119
rect 3306 2118 3346 2119
rect 3402 2118 3442 2119
rect 3498 2118 3538 2119
rect 3218 2054 3248 2118
rect 3312 2054 3342 2118
rect 3406 2054 3436 2118
rect 3500 2054 3530 2118
rect 3594 2054 3602 2119
rect 3146 2037 3602 2054
rect 3146 1967 3154 2037
rect 3210 2031 3250 2037
rect 3306 2031 3346 2037
rect 3402 2031 3442 2037
rect 3498 2031 3538 2037
rect 3218 1967 3248 2031
rect 3312 1967 3342 2031
rect 3406 1967 3436 2031
rect 3500 1967 3530 2031
rect 3594 1967 3602 2037
rect 3146 1955 3602 1967
rect 3146 1899 3154 1955
rect 3210 1899 3250 1955
rect 3306 1899 3346 1955
rect 3402 1899 3442 1955
rect 3498 1899 3538 1955
rect 3594 1899 3602 1955
rect 3146 1873 3602 1899
rect 3146 1817 3154 1873
rect 3210 1817 3250 1873
rect 3306 1817 3346 1873
rect 3402 1817 3442 1873
rect 3498 1817 3538 1873
rect 3594 1817 3602 1873
rect 3146 1791 3602 1817
rect 3146 1735 3154 1791
rect 3210 1735 3250 1791
rect 3306 1735 3346 1791
rect 3402 1735 3442 1791
rect 3498 1735 3538 1791
rect 3594 1735 3602 1791
rect 3146 1709 3602 1735
rect 3146 1653 3154 1709
rect 3210 1653 3250 1709
rect 3306 1653 3346 1709
rect 3402 1653 3442 1709
rect 3498 1653 3538 1709
rect 3594 1653 3602 1709
rect 3146 1648 3602 1653
rect -413 687 -257 692
rect -413 650 -374 687
rect -318 650 -257 687
rect -413 586 -407 650
rect -343 607 -327 631
rect -263 586 -257 650
rect 12249 650 12405 652
rect 12249 586 12255 650
rect 12319 647 12335 650
rect 12399 647 12405 650
rect 12320 591 12335 647
rect 12400 591 12405 647
rect 12319 586 12335 591
rect 12399 586 12405 591
rect -413 551 -374 586
rect -318 551 -257 586
rect -413 545 -257 551
rect 12329 362 12395 367
rect 12329 306 12334 362
rect 12390 306 12395 362
rect 12329 282 12395 306
rect 12329 226 12334 282
rect 12390 226 12395 282
rect -394 50 -328 55
rect -394 -6 -389 50
rect -333 -6 -328 50
rect -394 -30 -328 -6
rect -394 -86 -389 -30
rect -333 -86 -328 -30
tri -412 -273 -394 -255 se
rect -394 -273 -328 -86
tri -448 -309 -412 -273 se
rect -412 -309 -328 -273
tri -328 -309 -292 -273 sw
rect -448 -373 -442 -309
rect -378 -373 -362 -309
rect -298 -373 -292 -309
rect 11348 -373 11357 -309
rect 11421 -373 11437 -309
rect 11501 -373 11516 -309
rect 11348 -376 11516 -373
tri 12240 -1527 12329 -1438 se
rect 12329 -1527 12395 226
rect -204 -1528 -47 -1527
rect -204 -1592 -198 -1528
rect -134 -1592 -118 -1528
rect -54 -1592 -47 -1528
tri 12239 -1528 12240 -1527 se
rect 12240 -1528 12395 -1527
rect 12239 -1592 12245 -1528
rect 12309 -1592 12325 -1528
rect 12389 -1592 12395 -1528
rect -204 -1593 -47 -1592
<< via3 >>
rect 3154 2878 3210 2895
rect 3210 2878 3218 2895
rect 3154 2853 3218 2878
rect 3154 2831 3210 2853
rect 3210 2831 3218 2853
rect 3248 2878 3250 2895
rect 3250 2878 3306 2895
rect 3306 2878 3312 2895
rect 3248 2853 3312 2878
rect 3248 2831 3250 2853
rect 3250 2831 3306 2853
rect 3306 2831 3312 2853
rect 3342 2878 3346 2895
rect 3346 2878 3402 2895
rect 3402 2878 3406 2895
rect 3342 2853 3406 2878
rect 3342 2831 3346 2853
rect 3346 2831 3402 2853
rect 3402 2831 3406 2853
rect 3436 2878 3442 2895
rect 3442 2878 3498 2895
rect 3498 2878 3500 2895
rect 3436 2853 3500 2878
rect 3436 2831 3442 2853
rect 3442 2831 3498 2853
rect 3498 2831 3500 2853
rect 3530 2878 3538 2895
rect 3538 2878 3594 2895
rect 3530 2853 3594 2878
rect 3530 2831 3538 2853
rect 3538 2831 3594 2853
rect 3154 2797 3210 2809
rect 3210 2797 3218 2809
rect 3154 2772 3218 2797
rect 3154 2745 3210 2772
rect 3210 2745 3218 2772
rect 3248 2797 3250 2809
rect 3250 2797 3306 2809
rect 3306 2797 3312 2809
rect 3248 2772 3312 2797
rect 3248 2745 3250 2772
rect 3250 2745 3306 2772
rect 3306 2745 3312 2772
rect 3342 2797 3346 2809
rect 3346 2797 3402 2809
rect 3402 2797 3406 2809
rect 3342 2772 3406 2797
rect 3342 2745 3346 2772
rect 3346 2745 3402 2772
rect 3402 2745 3406 2772
rect 3436 2797 3442 2809
rect 3442 2797 3498 2809
rect 3498 2797 3500 2809
rect 3436 2772 3500 2797
rect 3436 2745 3442 2772
rect 3442 2745 3498 2772
rect 3498 2745 3500 2772
rect 3530 2797 3538 2809
rect 3538 2797 3594 2809
rect 3530 2772 3594 2797
rect 3530 2745 3538 2772
rect 3538 2745 3594 2772
rect 3154 2716 3210 2723
rect 3210 2716 3218 2723
rect 3154 2691 3218 2716
rect 3154 2659 3210 2691
rect 3210 2659 3218 2691
rect 3248 2716 3250 2723
rect 3250 2716 3306 2723
rect 3306 2716 3312 2723
rect 3248 2691 3312 2716
rect 3248 2659 3250 2691
rect 3250 2659 3306 2691
rect 3306 2659 3312 2691
rect 3342 2716 3346 2723
rect 3346 2716 3402 2723
rect 3402 2716 3406 2723
rect 3342 2691 3406 2716
rect 3342 2659 3346 2691
rect 3346 2659 3402 2691
rect 3402 2659 3406 2691
rect 3436 2716 3442 2723
rect 3442 2716 3498 2723
rect 3498 2716 3500 2723
rect 3436 2691 3500 2716
rect 3436 2659 3442 2691
rect 3442 2659 3498 2691
rect 3498 2659 3500 2691
rect 3530 2716 3538 2723
rect 3538 2716 3594 2723
rect 3530 2691 3594 2716
rect 3530 2659 3538 2691
rect 3538 2659 3594 2691
rect 3154 2635 3210 2637
rect 3210 2635 3218 2637
rect 3154 2610 3218 2635
rect 3154 2573 3210 2610
rect 3210 2573 3218 2610
rect 3248 2635 3250 2637
rect 3250 2635 3306 2637
rect 3306 2635 3312 2637
rect 3248 2610 3312 2635
rect 3248 2573 3250 2610
rect 3250 2573 3306 2610
rect 3306 2573 3312 2610
rect 3342 2635 3346 2637
rect 3346 2635 3402 2637
rect 3402 2635 3406 2637
rect 3342 2610 3406 2635
rect 3342 2573 3346 2610
rect 3346 2573 3402 2610
rect 3402 2573 3406 2610
rect 3436 2635 3442 2637
rect 3442 2635 3498 2637
rect 3498 2635 3500 2637
rect 3436 2610 3500 2635
rect 3436 2573 3442 2610
rect 3442 2573 3498 2610
rect 3498 2573 3500 2610
rect 3530 2635 3538 2637
rect 3538 2635 3594 2637
rect 3530 2610 3594 2635
rect 3530 2573 3538 2610
rect 3538 2573 3594 2610
rect 3154 2529 3218 2551
rect 3154 2487 3210 2529
rect 3210 2487 3218 2529
rect 3248 2529 3312 2551
rect 3248 2487 3250 2529
rect 3250 2487 3306 2529
rect 3306 2487 3312 2529
rect 3342 2529 3406 2551
rect 3342 2487 3346 2529
rect 3346 2487 3402 2529
rect 3402 2487 3406 2529
rect 3436 2529 3500 2551
rect 3436 2487 3442 2529
rect 3442 2487 3498 2529
rect 3498 2487 3500 2529
rect 3530 2529 3594 2551
rect 3530 2487 3538 2529
rect 3538 2487 3594 2529
rect 3154 2447 3218 2465
rect 3154 2401 3210 2447
rect 3210 2401 3218 2447
rect 3248 2447 3312 2465
rect 3248 2401 3250 2447
rect 3250 2401 3306 2447
rect 3306 2401 3312 2447
rect 3342 2447 3406 2465
rect 3342 2401 3346 2447
rect 3346 2401 3402 2447
rect 3402 2401 3406 2447
rect 3436 2447 3500 2465
rect 3436 2401 3442 2447
rect 3442 2401 3498 2447
rect 3498 2401 3500 2447
rect 3530 2447 3594 2465
rect 3530 2401 3538 2447
rect 3538 2401 3594 2447
rect 3154 2365 3218 2379
rect 3154 2315 3210 2365
rect 3210 2315 3218 2365
rect 3248 2365 3312 2379
rect 3248 2315 3250 2365
rect 3250 2315 3306 2365
rect 3306 2315 3312 2365
rect 3342 2365 3406 2379
rect 3342 2315 3346 2365
rect 3346 2315 3402 2365
rect 3402 2315 3406 2365
rect 3436 2365 3500 2379
rect 3436 2315 3442 2365
rect 3442 2315 3498 2365
rect 3498 2315 3500 2365
rect 3530 2365 3594 2379
rect 3530 2315 3538 2365
rect 3538 2315 3594 2365
rect 3154 2283 3218 2292
rect 3154 2228 3210 2283
rect 3210 2228 3218 2283
rect 3248 2283 3312 2292
rect 3248 2228 3250 2283
rect 3250 2228 3306 2283
rect 3306 2228 3312 2283
rect 3342 2283 3406 2292
rect 3342 2228 3346 2283
rect 3346 2228 3402 2283
rect 3402 2228 3406 2283
rect 3436 2283 3500 2292
rect 3436 2228 3442 2283
rect 3442 2228 3498 2283
rect 3498 2228 3500 2283
rect 3530 2283 3594 2292
rect 3530 2228 3538 2283
rect 3538 2228 3594 2283
rect 3154 2201 3218 2205
rect 3154 2145 3210 2201
rect 3210 2145 3218 2201
rect 3154 2141 3218 2145
rect 3248 2201 3312 2205
rect 3248 2145 3250 2201
rect 3250 2145 3306 2201
rect 3306 2145 3312 2201
rect 3248 2141 3312 2145
rect 3342 2201 3406 2205
rect 3342 2145 3346 2201
rect 3346 2145 3402 2201
rect 3402 2145 3406 2201
rect 3342 2141 3406 2145
rect 3436 2201 3500 2205
rect 3436 2145 3442 2201
rect 3442 2145 3498 2201
rect 3498 2145 3500 2201
rect 3436 2141 3500 2145
rect 3530 2201 3594 2205
rect 3530 2145 3538 2201
rect 3538 2145 3594 2201
rect 3530 2141 3594 2145
rect 3154 2063 3210 2118
rect 3210 2063 3218 2118
rect 3154 2054 3218 2063
rect 3248 2063 3250 2118
rect 3250 2063 3306 2118
rect 3306 2063 3312 2118
rect 3248 2054 3312 2063
rect 3342 2063 3346 2118
rect 3346 2063 3402 2118
rect 3402 2063 3406 2118
rect 3342 2054 3406 2063
rect 3436 2063 3442 2118
rect 3442 2063 3498 2118
rect 3498 2063 3500 2118
rect 3436 2054 3500 2063
rect 3530 2063 3538 2118
rect 3538 2063 3594 2118
rect 3530 2054 3594 2063
rect 3154 1981 3210 2031
rect 3210 1981 3218 2031
rect 3154 1967 3218 1981
rect 3248 1981 3250 2031
rect 3250 1981 3306 2031
rect 3306 1981 3312 2031
rect 3248 1967 3312 1981
rect 3342 1981 3346 2031
rect 3346 1981 3402 2031
rect 3402 1981 3406 2031
rect 3342 1967 3406 1981
rect 3436 1981 3442 2031
rect 3442 1981 3498 2031
rect 3498 1981 3500 2031
rect 3436 1967 3500 1981
rect 3530 1981 3538 2031
rect 3538 1981 3594 2031
rect 3530 1967 3594 1981
rect -407 631 -374 650
rect -374 631 -343 650
rect -327 631 -318 650
rect -318 631 -263 650
rect -407 607 -343 631
rect -327 607 -263 631
rect -407 586 -374 607
rect -374 586 -343 607
rect -327 586 -318 607
rect -318 586 -263 607
rect 12255 647 12319 650
rect 12335 647 12399 650
rect 12255 591 12264 647
rect 12264 591 12319 647
rect 12335 591 12344 647
rect 12344 591 12399 647
rect 12255 586 12319 591
rect 12335 586 12399 591
rect -442 -373 -378 -309
rect -362 -373 -298 -309
rect 11357 -315 11421 -309
rect 11357 -371 11413 -315
rect 11413 -371 11421 -315
rect 11357 -373 11421 -371
rect 11437 -315 11501 -309
rect 11437 -371 11493 -315
rect 11493 -371 11501 -315
rect 11437 -373 11501 -371
rect -198 -1532 -134 -1528
rect -198 -1588 -191 -1532
rect -191 -1588 -135 -1532
rect -135 -1588 -134 -1532
rect -198 -1592 -134 -1588
rect -118 -1532 -54 -1528
rect -118 -1588 -111 -1532
rect -111 -1588 -55 -1532
rect -55 -1588 -54 -1532
rect -118 -1592 -54 -1588
rect 12245 -1592 12309 -1528
rect 12325 -1592 12389 -1528
<< metal4 >>
rect 3150 2895 3598 2896
rect 3150 2831 3154 2895
rect 3218 2831 3248 2895
rect 3312 2831 3342 2895
rect 3406 2831 3436 2895
rect 3500 2831 3530 2895
rect 3594 2831 3598 2895
rect 3150 2809 3598 2831
rect 3150 2745 3154 2809
rect 3218 2745 3248 2809
rect 3312 2745 3342 2809
rect 3406 2745 3436 2809
rect 3500 2745 3530 2809
rect 3594 2745 3598 2809
rect 3150 2723 3598 2745
rect 3150 2659 3154 2723
rect 3218 2659 3248 2723
rect 3312 2659 3342 2723
rect 3406 2659 3436 2723
rect 3500 2659 3530 2723
rect 3594 2659 3598 2723
rect 3150 2637 3598 2659
rect 3150 2573 3154 2637
rect 3218 2573 3248 2637
rect 3312 2573 3342 2637
rect 3406 2573 3436 2637
rect 3500 2573 3530 2637
rect 3594 2573 3598 2637
rect 3150 2551 3598 2573
rect 3150 2487 3154 2551
rect 3218 2487 3248 2551
rect 3312 2487 3342 2551
rect 3406 2487 3436 2551
rect 3500 2487 3530 2551
rect 3594 2487 3598 2551
rect 3150 2465 3598 2487
rect 3150 2401 3154 2465
rect 3218 2401 3248 2465
rect 3312 2401 3342 2465
rect 3406 2401 3436 2465
rect 3500 2401 3530 2465
rect 3594 2401 3598 2465
rect 3150 2379 3598 2401
rect 3150 2315 3154 2379
rect 3218 2315 3248 2379
rect 3312 2315 3342 2379
rect 3406 2315 3436 2379
rect 3500 2315 3530 2379
rect 3594 2315 3598 2379
rect 3150 2292 3598 2315
rect 3150 2228 3154 2292
rect 3218 2228 3248 2292
rect 3312 2228 3342 2292
rect 3406 2228 3436 2292
rect 3500 2228 3530 2292
rect 3594 2228 3598 2292
rect 3150 2205 3598 2228
rect 3150 2141 3154 2205
rect 3218 2141 3248 2205
rect 3312 2141 3342 2205
rect 3406 2141 3436 2205
rect 3500 2141 3530 2205
rect 3594 2141 3598 2205
rect 3150 2118 3598 2141
rect 3150 2054 3154 2118
rect 3218 2054 3248 2118
rect 3312 2054 3342 2118
rect 3406 2054 3436 2118
rect 3500 2054 3530 2118
rect 3594 2054 3598 2118
rect 3150 2031 3598 2054
rect 3150 1967 3154 2031
rect 3218 1967 3248 2031
rect 3312 1967 3342 2031
rect 3406 1967 3436 2031
rect 3500 1967 3530 2031
rect 3594 1967 3598 2031
rect 3150 1966 3598 1967
rect -408 650 12400 651
rect -408 586 -407 650
rect -343 586 -327 650
rect -263 586 12255 650
rect 12319 586 12335 650
rect 12399 586 12400 650
rect -408 585 12400 586
rect -443 -309 11502 -308
rect -443 -373 -442 -309
rect -378 -373 -362 -309
rect -298 -373 11357 -309
rect 11421 -373 11437 -309
rect 11501 -373 11502 -309
rect -443 -374 11502 -373
rect -199 -1528 12394 -1527
rect -199 -1592 -198 -1528
rect -134 -1592 -118 -1528
rect -54 -1592 12245 -1528
rect 12309 -1592 12325 -1528
rect 12389 -1592 12394 -1528
rect -199 -1593 12394 -1592
use sky130_fd_io__com_opath_datoev2  sky130_fd_io__com_opath_datoev2_0
timestamp 1648127584
transform 1 0 467 0 -1 6943
box -349 -1098 12658 2562
use sky130_fd_io__gpiov2_obpredrvr  sky130_fd_io__gpiov2_obpredrvr_0
timestamp 1648127584
transform 1 0 288 0 -1 5207
box -958 -720 12780 4968
use sky130_fd_io__gpiov2_octl  sky130_fd_io__gpiov2_octl_0
timestamp 1648127584
transform 1 0 8821 0 -1 7867
box -9346 1177 6467 7642
<< labels >>
flabel metal1 s 14854 6410 14989 6527 3 FreeSans 520 180 0 0 VPWR
port 1 nsew
flabel metal1 s 12123 2928 12165 3058 7 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 9029 3979 9071 4181 7 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 470 3979 512 4181 3 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 1264 2928 1306 3058 3 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 1264 2312 1306 2442 3 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 12634 1302 12676 1504 7 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 12639 644 12676 790 7 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 12634 3453 12676 3655 7 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 1264 3453 1306 3655 3 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 288 644 325 790 3 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 288 1302 330 1504 3 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 12158 1828 12200 2030 7 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 12258 2312 12300 2442 7 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 12140 2928 12182 3058 7 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 491 4080 491 4080 3 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 1285 2993 1285 2993 3 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 1285 2377 1285 2377 3 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 951 1828 993 2030 3 FreeSans 300 0 0 0 VGND_IO
port 2 nsew
flabel metal1 s 12655 1403 12655 1403 7 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 12657 717 12657 717 7 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 12655 3554 12655 3554 7 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 1285 3554 1285 3554 3 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 306 717 306 717 3 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 309 1403 309 1403 3 FreeSans 300 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 5854 6502 5921 6850 3 FreeSans 520 0 0 0 VPWR_KA
port 4 nsew
flabel metal1 s 524 4938 564 5068 3 FreeSans 300 180 0 0 VGND
port 5 nsew
flabel metal1 s 288 5857 328 6059 3 FreeSans 300 180 0 0 VGND
port 5 nsew
flabel metal1 s 288 4708 328 4910 3 FreeSans 300 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 12991 4708 13031 4910 3 FreeSans 300 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 5900 6502 5967 6850 3 FreeSans 520 0 0 0 VPWR_KA
port 4 nsew
flabel metal1 s 544 5003 544 5003 3 FreeSans 300 180 0 0 VGND
port 5 nsew
flabel metal1 s 12900 4938 12940 5068 3 FreeSans 300 180 0 0 VGND
port 5 nsew
flabel metal1 s 308 5958 308 5958 3 FreeSans 300 180 0 0 VGND
port 5 nsew
flabel metal1 s 13102 5787 13142 5989 3 FreeSans 300 180 0 0 VGND
port 5 nsew
flabel metal1 s 308 4809 308 4809 3 FreeSans 300 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 13011 4809 13011 4809 3 FreeSans 300 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 13170 5809 13337 5965 3 FreeSans 520 180 0 0 VGND
port 5 nsew
flabel metal1 s 14840 4258 15007 4414 3 FreeSans 520 0 0 0 VGND
port 5 nsew
flabel metal1 s 14840 2226 15007 2382 3 FreeSans 520 0 0 0 VGND
port 5 nsew
flabel metal1 s 14840 260 15007 416 3 FreeSans 520 0 0 0 VGND
port 5 nsew
flabel metal1 s 13251 4812 13562 4987 3 FreeSans 520 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 14697 3248 15008 3480 3 FreeSans 520 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 14697 1137 15008 1369 3 FreeSans 520 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 14923 4336 14923 4336 3 FreeSans 520 0 0 0 VGND
port 5 nsew
flabel metal1 s 14923 2304 14923 2304 3 FreeSans 520 0 0 0 VGND
port 5 nsew
flabel metal1 s 14923 338 14923 338 3 FreeSans 520 0 0 0 VGND
port 5 nsew
flabel metal1 s 13406 4899 13406 4899 3 FreeSans 520 180 0 0 VCC_IO
port 3 nsew
flabel metal1 s 14852 3364 14852 3364 3 FreeSans 520 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 14852 1253 14852 1253 3 FreeSans 520 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 15042 5345 15116 5380 3 FreeSans 520 180 0 0 SLOW
port 6 nsew
flabel metal1 s 14478 5304 14522 5348 3 FreeSans 520 180 0 0 HLD_I_H_N
port 7 nsew
flabel metal1 s 15079 5362 15079 5362 3 FreeSans 520 180 0 0 SLOW
port 6 nsew
flabel metal1 s 14501 5326 14501 5326 3 FreeSans 520 180 0 0 HLD_I_H_N
port 7 nsew
flabel metal1 s 5095 6957 5128 6995 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 8 nsew
flabel metal1 s 5111 6976 5111 6976 3 FreeSans 520 0 0 0 HLD_I_OVR_H
port 8 nsew
flabel metal1 s 15079 5362 15079 5362 3 FreeSans 520 180 0 0 SLOW
port 6 nsew
flabel metal1 s 14824 6126 14868 6164 3 FreeSans 520 180 0 0 OD_H
port 9 nsew
flabel metal1 s 14501 5326 14501 5326 3 FreeSans 520 180 0 0 HLD_I_H_N
port 7 nsew
flabel metal1 s 13425 5630 13492 5674 3 FreeSans 520 180 0 0 SLOW_H_N
port 10 nsew
flabel metal1 s 8283 5096 8333 5148 3 FreeSans 300 180 0 0 DRVHI_H
port 11 nsew
flabel metal1 s 8308 5122 8308 5122 3 FreeSans 300 180 0 0 DRVHI_H
port 11 nsew
flabel metal1 s 6190 1228 6231 1274 3 FreeSans 300 0 0 0 PU_H_N[3]
port 12 nsew
flabel metal1 s 6054 1228 6094 1274 7 FreeSans 300 0 0 0 PU_H_N[2]
port 13 nsew
flabel metal1 s 10362 1072 10402 1118 3 FreeSans 300 0 0 0 PU_H_N[1]
port 14 nsew
flabel metal1 s 7956 1148 7996 1194 3 FreeSans 300 0 0 0 PU_H_N[0]
port 15 nsew
flabel metal1 s 9390 1030 9436 1076 3 FreeSans 300 0 0 0 PD_H[1]
port 16 nsew
flabel metal1 s 8148 1030 8194 1076 3 FreeSans 300 0 0 0 PD_H[0]
port 17 nsew
flabel metal1 s 11863 2475 11928 2502 3 FreeSans 520 0 0 0 PD_H[4]
port 18 nsew
flabel metal1 s 8242 4238 8242 4238 0 FreeSans 440 0 0 0 DRVLO_H_N
port 19 nsew
flabel metal2 s 13617 397 13652 442 3 FreeSans 520 90 0 0 DM_H_N[2]
port 20 nsew
flabel metal2 s 14263 399 14307 448 3 FreeSans 520 90 0 0 DM_H_N[0]
port 21 nsew
flabel metal2 s 12786 514 12812 563 3 FreeSans 520 90 0 0 DM_H[2]
port 22 nsew
flabel metal2 s 13425 445 13474 498 3 FreeSans 520 90 0 0 DM_H[1]
port 23 nsew
flabel metal2 s 13257 437 13306 500 3 FreeSans 520 90 0 0 DM_H[0]
port 24 nsew
flabel metal2 s 13634 419 13634 419 3 FreeSans 520 90 0 0 DM_H_N[2]
port 20 nsew
flabel metal2 s 14285 423 14285 423 3 FreeSans 520 90 0 0 DM_H_N[0]
port 21 nsew
flabel metal2 s 13449 471 13449 471 3 FreeSans 520 90 0 0 DM_H[1]
port 23 nsew
flabel metal2 s 3827 6885 3879 6924 3 FreeSans 520 0 0 0 OUT
port 25 nsew
flabel metal2 s 3354 6878 3400 6924 7 FreeSans 300 0 0 0 OE_N
port 26 nsew
flabel metal2 s 3848 6898 3848 6898 3 FreeSans 520 0 0 0 OUT
port 25 nsew
flabel metal2 s 3377 6901 3377 6901 7 FreeSans 300 0 0 0 OE_N
port 26 nsew
flabel metal2 s -367 5535 -318 5598 3 FreeSans 520 90 0 0 DM_H[0]
port 24 nsew
flabel metal2 s 13634 419 13634 419 3 FreeSans 520 90 0 0 DM_H_N[2]
port 20 nsew
flabel metal2 s 13789 394 13823 443 3 FreeSans 520 90 0 0 DM_H_N[1]
port 27 nsew
flabel metal2 s 14285 423 14285 423 3 FreeSans 520 90 0 0 DM_H_N[0]
port 21 nsew
flabel metal2 s 13449 471 13449 471 3 FreeSans 520 90 0 0 DM_H[1]
port 23 nsew
flabel metal2 s 11401 2065 11449 2117 3 FreeSans 300 0 0 0 PD_H[3]
port 28 nsew
flabel metal2 s 1 5402 27 5451 3 FreeSans 520 90 0 0 DM_H[2]
port 22 nsew
flabel metal2 s -193 5390 -144 5443 3 FreeSans 520 90 0 0 DM_H[1]
port 23 nsew
flabel metal2 s 10919 2470 10967 2522 3 FreeSans 300 0 0 0 PD_H[2]
port 29 nsew
<< properties >>
string GDS_END 7685534
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7611198
<< end >>
