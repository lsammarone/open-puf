magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< obsli1 >>
rect 228 1186 266 1220
rect 300 1186 338 1220
rect 372 1186 410 1220
rect 444 1186 482 1220
rect 516 1186 554 1220
rect 588 1186 626 1220
rect 660 1186 698 1220
rect 732 1186 736 1220
rect 38 1033 72 1071
rect 38 961 72 999
rect 38 889 72 927
rect 38 817 72 855
rect 38 745 72 783
rect 38 673 72 711
rect 38 601 72 639
rect 38 529 72 567
rect 38 457 72 495
rect 38 385 72 423
rect 38 313 72 351
rect 38 241 72 279
rect 38 135 72 207
rect 149 111 183 1129
rect 233 111 339 1129
rect 387 111 493 1129
rect 541 111 647 1129
rect 697 111 731 1129
rect 811 135 845 1105
rect 228 20 266 54
rect 300 20 338 54
rect 372 20 410 54
rect 444 20 482 54
rect 516 20 554 54
rect 588 20 626 54
rect 660 20 698 54
rect 732 20 736 54
<< obsli1c >>
rect 194 1186 228 1220
rect 266 1186 300 1220
rect 338 1186 372 1220
rect 410 1186 444 1220
rect 482 1186 516 1220
rect 554 1186 588 1220
rect 626 1186 660 1220
rect 698 1186 732 1220
rect 38 1071 72 1105
rect 38 999 72 1033
rect 38 927 72 961
rect 38 855 72 889
rect 38 783 72 817
rect 38 711 72 745
rect 38 639 72 673
rect 38 567 72 601
rect 38 495 72 529
rect 38 423 72 457
rect 38 351 72 385
rect 38 279 72 313
rect 38 207 72 241
rect 194 20 228 54
rect 266 20 300 54
rect 338 20 372 54
rect 410 20 444 54
rect 482 20 516 54
rect 554 20 588 54
rect 626 20 660 54
rect 698 20 732 54
<< metal1 >>
rect 182 1220 744 1232
rect 182 1186 194 1220
rect 228 1186 266 1220
rect 300 1186 338 1220
rect 372 1186 410 1220
rect 444 1186 482 1220
rect 516 1186 554 1220
rect 588 1186 626 1220
rect 660 1186 698 1220
rect 732 1186 744 1220
rect 182 1174 744 1186
rect 26 1105 84 1117
rect 26 1071 38 1105
rect 72 1071 84 1105
rect 26 1033 84 1071
rect 26 999 38 1033
rect 72 999 84 1033
rect 26 961 84 999
rect 26 927 38 961
rect 72 927 84 961
rect 26 889 84 927
rect 26 855 38 889
rect 72 855 84 889
rect 26 817 84 855
rect 26 783 38 817
rect 72 783 84 817
rect 26 745 84 783
rect 26 711 38 745
rect 72 711 84 745
rect 26 673 84 711
rect 26 639 38 673
rect 72 639 84 673
rect 26 601 84 639
rect 26 567 38 601
rect 72 567 84 601
rect 26 529 84 567
rect 26 495 38 529
rect 72 495 84 529
rect 26 457 84 495
rect 26 423 38 457
rect 72 423 84 457
rect 26 385 84 423
rect 26 351 38 385
rect 72 351 84 385
rect 26 313 84 351
rect 26 279 38 313
rect 72 279 84 313
rect 26 241 84 279
rect 26 207 38 241
rect 72 207 84 241
rect 26 123 84 207
rect 182 54 744 66
rect 182 20 194 54
rect 228 20 266 54
rect 300 20 338 54
rect 372 20 410 54
rect 444 20 482 54
rect 516 20 554 54
rect 588 20 626 54
rect 660 20 698 54
rect 732 20 744 54
rect 182 8 744 20
<< obsm1 >>
rect 140 1117 192 1128
rect 382 1117 498 1129
rect 688 1117 740 1129
rect 140 123 195 1117
rect 223 123 349 1117
rect 377 123 503 1117
rect 531 123 657 1117
rect 685 123 743 1117
rect 799 123 857 1117
rect 140 112 192 123
rect 382 112 498 123
rect 688 112 740 123
<< metal2 >>
rect 0 872 884 1129
rect 0 396 884 844
rect 0 112 884 368
<< labels >>
rlabel metal2 s 0 396 884 844 6 DRAIN
port 1 nsew
rlabel metal1 s 182 1174 744 1232 6 GATE
port 2 nsew
rlabel metal1 s 182 8 744 66 6 GATE
port 2 nsew
rlabel metal2 s 0 872 884 1129 6 SOURCE
port 3 nsew
rlabel metal2 s 0 112 884 368 6 SOURCE
port 3 nsew
rlabel metal1 s 26 123 84 1117 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 4 884 1236
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7186134
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7156630
<< end >>
