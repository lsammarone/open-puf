.subckt NBR128 VDD VSS OUT
+ C[127] C[126] C[125] C[124] C[123] C[122] C[121] C[120] C[119] C[118] C[117] C[116] C[115] C[114] C[113] C[112] C[111] C[110] C[109] C[108] C[107] C[106] C[105] C[104] C[103] C[102] C[101] C[100] C[99] C[98] C[97] C[96] C[95] C[94] C[93] C[92] C[91] C[90] C[89] C[88] C[87] C[86] C[85] C[84] C[83] C[82] C[81] C[80] C[79] C[78] C[77] C[76] C[75] C[74] C[73] C[72] C[71] C[70] C[69] C[68] C[67] C[66] C[65] C[64] C[63] C[62] C[61] C[60] C[59] C[58] C[57] C[56] C[55] C[54] C[53] C[52] C[51] C[50] C[49] C[48] C[47] C[46] C[45] C[44] C[43] C[42] C[41] C[40] C[39] C[38] C[37] C[36] C[35] C[34] C[33] C[32] C[31] C[30] C[29] C[28] C[27] C[26] C[25] C[24] C[23] C[22] C[21] C[20] C[19] C[18] C[17] C[16] C[15] C[14] C[13] C[12] C[11] C[10] C[9] C[8] C[7] C[6] C[5] C[4] C[3] C[2] C[1] C[0] RESET
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin
*+ C[127],C[126],C[125],C[124],C[123],C[122],C[121],C[120],C[119],C[118],C[117],C[116],C[115],C[114],C[113],C[112],C[111],C[110],C[109],C[108],C[107],C[106],C[105],C[104],C[103],C[102],C[101],C[100],C[99],C[98],C[97],C[96],C[95],C[94],C[93],C[92],C[91],C[90],C[89],C[88],C[87],C[86],C[85],C[84],C[83],C[82],C[81],C[80],C[79],C[78],C[77],C[76],C[75],C[74],C[73],C[72],C[71],C[70],C[69],C[68],C[67],C[66],C[65],C[64],C[63],C[62],C[61],C[60],C[59],C[58],C[57],C[56],C[55],C[54],C[53],C[52],C[51],C[50],C[49],C[48],C[47],C[46],C[45],C[44],C[43],C[42],C[41],C[40],C[39],C[38],C[37],C[36],C[35],C[34],C[33],C[32],C[31],C[30],C[29],C[28],C[27],C[26],C[25],C[24],C[23],C[22],C[21],C[20],C[19],C[18],C[17],C[16],C[15],C[14],C[13],C[12],C[11],C[10],C[9],C[8],C[7],C[6],C[5],C[4],C[3],C[2],C[1],C[0]
*.ipin RESET
x47 net1 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x48 net1 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x4 net1 VSS VSS VDD VDD r1 sky130_fd_sc_hd__inv_16
x5 net1 VSS VSS VDD VDD r2 sky130_fd_sc_hd__inv_16
x6 net1 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x7 net1 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x8 net1 VSS VSS VDD VDD r3 sky130_fd_sc_hd__inv_16
x10 net1 VSS VSS VDD VDD r4 sky130_fd_sc_hd__inv_16
x11 net2 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_16
x12 net2 VSS VSS VDD VDD net1 sky130_fd_sc_hd__inv_16
x13 net3 VSS VSS VDD VDD r6 sky130_fd_sc_hd__inv_16
x14 net3 VSS VSS VDD VDD r5 sky130_fd_sc_hd__inv_16
x15 net3 VSS VSS VDD VDD r5 sky130_fd_sc_hd__inv_16
x16 net3 VSS VSS VDD VDD r6 sky130_fd_sc_hd__inv_16
x17 net3 VSS VSS VDD VDD r8 sky130_fd_sc_hd__inv_16
x18 net3 VSS VSS VDD VDD r7 sky130_fd_sc_hd__inv_16
x19 net3 VSS VSS VDD VDD r7 sky130_fd_sc_hd__inv_16
x20 net3 VSS VSS VDD VDD r8 sky130_fd_sc_hd__inv_16
x21 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_16
x22 net2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__inv_16
x23 net6 VSS VSS VDD VDD net2 sky130_fd_sc_hd__inv_16
x3[7] r1 VDD VSS out[8] out[7] net8[7] C[7] out2[7] out2[8] singlestage_nbr
x3[6] r1 VDD VSS out[7] out[6] net8[6] C[6] out2[6] out2[7] singlestage_nbr
x3[5] r1 VDD VSS out[6] out[5] net8[5] C[5] out2[5] out2[6] singlestage_nbr
x3[4] r1 VDD VSS out[5] out[4] net8[4] C[4] out2[4] out2[5] singlestage_nbr
x3[3] r1 VDD VSS out[4] out[3] net8[3] C[3] out2[3] out2[4] singlestage_nbr
x3[2] r1 VDD VSS out[3] out[2] net8[2] C[2] out2[2] out2[3] singlestage_nbr
x3[1] r1 VDD VSS out[2] out[1] net8[1] C[1] out2[1] out2[2] singlestage_nbr
x3[0] r1 VDD VSS out[1] out[0] net8[0] C[0] out2[0] out2[1] singlestage_nbr
x1[15] r2 VDD VSS out[16] out[15] net9[7] C[15] out2[15] out2[16] singlestage_nbr
x1[14] r2 VDD VSS out[15] out[14] net9[6] C[14] out2[14] out2[15] singlestage_nbr
x1[13] r2 VDD VSS out[14] out[13] net9[5] C[13] out2[13] out2[14] singlestage_nbr
x1[12] r2 VDD VSS out[13] out[12] net9[4] C[12] out2[12] out2[13] singlestage_nbr
x1[11] r2 VDD VSS out[12] out[11] net9[3] C[11] out2[11] out2[12] singlestage_nbr
x1[10] r2 VDD VSS out[11] out[10] net9[2] C[10] out2[10] out2[11] singlestage_nbr
x1[9] r2 VDD VSS out[10] out[9] net9[1] C[9] out2[9] out2[10] singlestage_nbr
x1[8] r2 VDD VSS out[9] out[8] net9[0] C[8] out2[8] out2[9] singlestage_nbr
x2[23] r5 VDD VSS out[24] out[23] net10[7] C[23] out2[23] out2[24] singlestage_nbr
x2[22] r5 VDD VSS out[23] out[22] net10[6] C[22] out2[22] out2[23] singlestage_nbr
x2[21] r5 VDD VSS out[22] out[21] net10[5] C[21] out2[21] out2[22] singlestage_nbr
x2[20] r5 VDD VSS out[21] out[20] net10[4] C[20] out2[20] out2[21] singlestage_nbr
x2[19] r5 VDD VSS out[20] out[19] net10[3] C[19] out2[19] out2[20] singlestage_nbr
x2[18] r5 VDD VSS out[19] out[18] net10[2] C[18] out2[18] out2[19] singlestage_nbr
x2[17] r5 VDD VSS out[18] out[17] net10[1] C[17] out2[17] out2[18] singlestage_nbr
x2[16] r5 VDD VSS out[17] out[16] net10[0] C[16] out2[16] out2[17] singlestage_nbr
x4[31] r6 VDD VSS out[32] out[31] net11[7] C[31] out2[31] out2[32] singlestage_nbr
x4[30] r6 VDD VSS out[31] out[30] net11[6] C[30] out2[30] out2[31] singlestage_nbr
x4[29] r6 VDD VSS out[30] out[29] net11[5] C[29] out2[29] out2[30] singlestage_nbr
x4[28] r6 VDD VSS out[29] out[28] net11[4] C[28] out2[28] out2[29] singlestage_nbr
x4[27] r6 VDD VSS out[28] out[27] net11[3] C[27] out2[27] out2[28] singlestage_nbr
x4[26] r6 VDD VSS out[27] out[26] net11[2] C[26] out2[26] out2[27] singlestage_nbr
x4[25] r6 VDD VSS out[26] out[25] net11[1] C[25] out2[25] out2[26] singlestage_nbr
x4[24] r6 VDD VSS out[25] out[24] net11[0] C[24] out2[24] out2[25] singlestage_nbr
x5[62] r13 VDD VSS out[63] out[62] net15[7] C[62] out2[62] out2[63] singlestage_nbr
x5[61] r13 VDD VSS out[62] out[61] net15[6] C[61] out2[61] out2[62] singlestage_nbr
x5[60] r13 VDD VSS out[61] out[60] net15[5] C[60] out2[60] out2[61] singlestage_nbr
x5[59] r13 VDD VSS out[60] out[59] net15[4] C[59] out2[59] out2[60] singlestage_nbr
x5[58] r13 VDD VSS out[59] out[58] net15[3] C[58] out2[58] out2[59] singlestage_nbr
x5[57] r13 VDD VSS out[58] out[57] net15[2] C[57] out2[57] out2[58] singlestage_nbr
x5[56] r13 VDD VSS out[57] out[56] net15[1] C[56] out2[56] out2[57] singlestage_nbr
x5[55] r13 VDD VSS out[56] out[55] net15[0] C[55] out2[55] out2[56] singlestage_nbr
x6[54] r14 VDD VSS out[55] out[54] net14[7] C[54] out2[54] out2[55] singlestage_nbr
x6[53] r14 VDD VSS out[54] out[53] net14[6] C[53] out2[53] out2[54] singlestage_nbr
x6[52] r14 VDD VSS out[53] out[52] net14[5] C[52] out2[52] out2[53] singlestage_nbr
x6[51] r14 VDD VSS out[52] out[51] net14[4] C[51] out2[51] out2[52] singlestage_nbr
x6[50] r14 VDD VSS out[51] out[50] net14[3] C[50] out2[50] out2[51] singlestage_nbr
x6[49] r14 VDD VSS out[50] out[49] net14[2] C[49] out2[49] out2[50] singlestage_nbr
x6[48] r14 VDD VSS out[49] out[48] net14[1] C[48] out2[48] out2[49] singlestage_nbr
x6[47] r14 VDD VSS out[48] out[47] net14[0] C[47] out2[47] out2[48] singlestage_nbr
x7[46] r9 VDD VSS out[47] out[46] net13[7] C[46] out2[46] out2[47] singlestage_nbr
x7[45] r9 VDD VSS out[46] out[45] net13[6] C[45] out2[45] out2[46] singlestage_nbr
x7[44] r9 VDD VSS out[45] out[44] net13[5] C[44] out2[44] out2[45] singlestage_nbr
x7[43] r9 VDD VSS out[44] out[43] net13[4] C[43] out2[43] out2[44] singlestage_nbr
x7[42] r9 VDD VSS out[43] out[42] net13[3] C[42] out2[42] out2[43] singlestage_nbr
x7[41] r9 VDD VSS out[42] out[41] net13[2] C[41] out2[41] out2[42] singlestage_nbr
x7[40] r9 VDD VSS out[41] out[40] net13[1] C[40] out2[40] out2[41] singlestage_nbr
x7[39] r9 VDD VSS out[40] out[39] net13[0] C[39] out2[39] out2[40] singlestage_nbr
x8[38] r10 VDD VSS out[39] out[38] net12[6] C[38] out2[38] out2[39] singlestage_nbr
x8[37] r10 VDD VSS out[38] out[37] net12[5] C[37] out2[37] out2[38] singlestage_nbr
x8[36] r10 VDD VSS out[37] out[36] net12[4] C[36] out2[36] out2[37] singlestage_nbr
x8[35] r10 VDD VSS out[36] out[35] net12[3] C[35] out2[35] out2[36] singlestage_nbr
x8[34] r10 VDD VSS out[35] out[34] net12[2] C[34] out2[34] out2[35] singlestage_nbr
x8[33] r10 VDD VSS out[34] out[33] net12[1] C[33] out2[33] out2[34] singlestage_nbr
x8[32] r10 VDD VSS out[33] out[32] net12[0] C[32] out2[32] out2[33] singlestage_nbr
x1 net6 VSS VSS VDD VDD net2 sky130_fd_sc_hd__inv_16
x2 net4 VSS VSS VDD VDD r10 sky130_fd_sc_hd__inv_16
x3 net4 VSS VSS VDD VDD r9 sky130_fd_sc_hd__inv_16
x9 net4 VSS VSS VDD VDD r9 sky130_fd_sc_hd__inv_16
x24 net4 VSS VSS VDD VDD r10 sky130_fd_sc_hd__inv_16
x25 net4 VSS VSS VDD VDD r12 sky130_fd_sc_hd__inv_16
x26 net4 VSS VSS VDD VDD r11 sky130_fd_sc_hd__inv_16
x27 net4 VSS VSS VDD VDD r11 sky130_fd_sc_hd__inv_16
x28 net4 VSS VSS VDD VDD r12 sky130_fd_sc_hd__inv_16
x29 net2 VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_16
x30 net2 VSS VSS VDD VDD net4 sky130_fd_sc_hd__inv_16
x31 net5 VSS VSS VDD VDD r14 sky130_fd_sc_hd__inv_16
x32 net5 VSS VSS VDD VDD r13 sky130_fd_sc_hd__inv_16
x33 net5 VSS VSS VDD VDD r13 sky130_fd_sc_hd__inv_16
x34 net5 VSS VSS VDD VDD r14 sky130_fd_sc_hd__inv_16
x35 net5 VSS VSS VDD VDD r16 sky130_fd_sc_hd__inv_16
x36 net5 VSS VSS VDD VDD r15 sky130_fd_sc_hd__inv_16
x37 net5 VSS VSS VDD VDD r15 sky130_fd_sc_hd__inv_16
x38 net5 VSS VSS VDD VDD r16 sky130_fd_sc_hd__inv_16
x39 net2 VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_16
x40 net2 VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_16
x6[70] r16 VDD VSS out[71] out[70] net16[7] C[70] out2[70] out2[71] singlestage_nbr
x6[69] r16 VDD VSS out[70] out[69] net16[6] C[69] out2[69] out2[70] singlestage_nbr
x6[68] r16 VDD VSS out[69] out[68] net16[5] C[68] out2[68] out2[69] singlestage_nbr
x6[67] r16 VDD VSS out[68] out[67] net16[4] C[67] out2[67] out2[68] singlestage_nbr
x6[66] r16 VDD VSS out[67] out[66] net16[3] C[66] out2[66] out2[67] singlestage_nbr
x6[65] r16 VDD VSS out[66] out[65] net16[2] C[65] out2[65] out2[66] singlestage_nbr
x6[64] r16 VDD VSS out[65] out[64] net16[1] C[64] out2[64] out2[65] singlestage_nbr
x6[63] r16 VDD VSS out[64] out[63] net16[0] C[63] out2[63] out2[64] singlestage_nbr
x7[78] r15 VDD VSS out[79] out[78] net17[7] C[78] out2[78] out2[79] singlestage_nbr
x7[77] r15 VDD VSS out[78] out[77] net17[6] C[77] out2[77] out2[78] singlestage_nbr
x7[76] r15 VDD VSS out[77] out[76] net17[5] C[76] out2[76] out2[77] singlestage_nbr
x7[75] r15 VDD VSS out[76] out[75] net17[4] C[75] out2[75] out2[76] singlestage_nbr
x7[74] r15 VDD VSS out[75] out[74] net17[3] C[74] out2[74] out2[75] singlestage_nbr
x7[73] r15 VDD VSS out[74] out[73] net17[2] C[73] out2[73] out2[74] singlestage_nbr
x7[72] r15 VDD VSS out[73] out[72] net17[1] C[72] out2[72] out2[73] singlestage_nbr
x7[71] r15 VDD VSS out[72] out[71] net17[0] C[71] out2[71] out2[72] singlestage_nbr
x8[86] r12 VDD VSS out[87] out[86] net18[7] C[86] out2[86] out2[87] singlestage_nbr
x8[85] r12 VDD VSS out[86] out[85] net18[6] C[85] out2[85] out2[86] singlestage_nbr
x8[84] r12 VDD VSS out[85] out[84] net18[5] C[84] out2[84] out2[85] singlestage_nbr
x8[83] r12 VDD VSS out[84] out[83] net18[4] C[83] out2[83] out2[84] singlestage_nbr
x8[82] r12 VDD VSS out[83] out[82] net18[3] C[82] out2[82] out2[83] singlestage_nbr
x8[81] r12 VDD VSS out[82] out[81] net18[2] C[81] out2[81] out2[82] singlestage_nbr
x8[80] r12 VDD VSS out[81] out[80] net18[1] C[80] out2[80] out2[81] singlestage_nbr
x8[79] r12 VDD VSS out[80] out[79] net18[0] C[79] out2[79] out2[80] singlestage_nbr
x9[94] r11 VDD VSS out[95] out[94] net22[7] C[94] out2[94] out2[95] singlestage_nbr
x9[93] r11 VDD VSS out[94] out[93] net22[6] C[93] out2[93] out2[94] singlestage_nbr
x9[92] r11 VDD VSS out[93] out[92] net22[5] C[92] out2[92] out2[93] singlestage_nbr
x9[91] r11 VDD VSS out[92] out[91] net22[4] C[91] out2[91] out2[92] singlestage_nbr
x9[90] r11 VDD VSS out[91] out[90] net22[3] C[90] out2[90] out2[91] singlestage_nbr
x9[89] r11 VDD VSS out[90] out[89] net22[2] C[89] out2[89] out2[90] singlestage_nbr
x9[88] r11 VDD VSS out[89] out[88] net22[1] C[88] out2[88] out2[89] singlestage_nbr
x9[87] r11 VDD VSS out[88] out[87] net22[0] C[87] out2[87] out2[88] singlestage_nbr
x1[127] r3 VDD VSS out[0] out[127] OUT C[127] out2[127] out2[0] singlestage_nbr
x1[126] r3 VDD VSS out[127] out[126] buf_out[7] C[126] out2[126] out2[127] singlestage_nbr
x1[125] r3 VDD VSS out[126] out[125] buf_out[6] C[125] out2[125] out2[126] singlestage_nbr
x1[124] r3 VDD VSS out[125] out[124] buf_out[5] C[124] out2[124] out2[125] singlestage_nbr
x1[123] r3 VDD VSS out[124] out[123] buf_out[4] C[123] out2[123] out2[124] singlestage_nbr
x1[122] r3 VDD VSS out[123] out[122] buf_out[3] C[122] out2[122] out2[123] singlestage_nbr
x1[121] r3 VDD VSS out[122] out[121] buf_out[2] C[121] out2[121] out2[122] singlestage_nbr
x1[120] r3 VDD VSS out[121] out[120] buf_out[1] C[120] out2[120] out2[121] singlestage_nbr
x1[119] r3 VDD VSS out[120] out[119] buf_out[0] C[119] out2[119] out2[120] singlestage_nbr
x2[118] r4 VDD VSS out[119] out[118] net21[7] C[118] out2[118] out2[119] singlestage_nbr
x2[117] r4 VDD VSS out[118] out[117] net21[6] C[117] out2[117] out2[118] singlestage_nbr
x2[116] r4 VDD VSS out[117] out[116] net21[5] C[116] out2[116] out2[117] singlestage_nbr
x2[115] r4 VDD VSS out[116] out[115] net21[4] C[115] out2[115] out2[116] singlestage_nbr
x2[114] r4 VDD VSS out[115] out[114] net21[3] C[114] out2[114] out2[115] singlestage_nbr
x2[113] r4 VDD VSS out[114] out[113] net21[2] C[113] out2[113] out2[114] singlestage_nbr
x2[112] r4 VDD VSS out[113] out[112] net21[1] C[112] out2[112] out2[113] singlestage_nbr
x2[111] r4 VDD VSS out[112] out[111] net21[0] C[111] out2[111] out2[112] singlestage_nbr
x3[110] r8 VDD VSS out[111] out[110] net20[7] C[110] out2[110] out2[111] singlestage_nbr
x3[109] r8 VDD VSS out[110] out[109] net20[6] C[109] out2[109] out2[110] singlestage_nbr
x3[108] r8 VDD VSS out[109] out[108] net20[5] C[108] out2[108] out2[109] singlestage_nbr
x3[107] r8 VDD VSS out[108] out[107] net20[4] C[107] out2[107] out2[108] singlestage_nbr
x3[106] r8 VDD VSS out[107] out[106] net20[3] C[106] out2[106] out2[107] singlestage_nbr
x3[105] r8 VDD VSS out[106] out[105] net20[2] C[105] out2[105] out2[106] singlestage_nbr
x3[104] r8 VDD VSS out[105] out[104] net20[1] C[104] out2[104] out2[105] singlestage_nbr
x3[103] r8 VDD VSS out[104] out[103] net20[0] C[103] out2[103] out2[104] singlestage_nbr
x4[102] r7 VDD VSS out[103] out[102] net19[7] C[102] out2[102] out2[103] singlestage_nbr
x4[101] r7 VDD VSS out[102] out[101] net19[6] C[101] out2[101] out2[102] singlestage_nbr
x4[100] r7 VDD VSS out[101] out[100] net19[5] C[100] out2[100] out2[101] singlestage_nbr
x4[99] r7 VDD VSS out[100] out[99] net19[4] C[99] out2[99] out2[100] singlestage_nbr
x4[98] r7 VDD VSS out[99] out[98] net19[3] C[98] out2[98] out2[99] singlestage_nbr
x4[97] r7 VDD VSS out[98] out[97] net19[2] C[97] out2[97] out2[98] singlestage_nbr
x4[96] r7 VDD VSS out[97] out[96] net19[1] C[96] out2[96] out2[97] singlestage_nbr
x4[95] r7 VDD VSS out[96] out[95] net19[0] C[95] out2[95] out2[96] singlestage_nbr
x41 RESET VSS VSS VDD VDD net7 sky130_fd_sc_hd__buf_2
x42 net7 VSS VSS VDD VDD net6 sky130_fd_sc_hd__inv_8
.ends

* expanding   symbol:  singlestage_nbr.sym # of pins=9
* sym_path: /home/users/lsammaro/open-puf/design/singlestage_nbr.sym
* sch_path: /home/users/lsammaro/open-puf/design/singlestage_nbr.sch
.subckt singlestage_nbr  RESET VDD VSS OUT1 IN1 buf_out C IN2 OUT2
*.ipin IN1
*.ipin C
*.ipin RESET
*.iopin VSS
*.iopin VDD
*.opin OUT2
*.opin buf_out
*.opin OUT1
*.ipin IN2
x1 RESET IN1 VSS VSS VDD VDD net1 sky130_fd_sc_hd__nor2_1
x2 RESET IN2 VSS VSS VDD VDD net2 sky130_fd_sc_hd__nor2_1
x5 Cb VSS VSS VDD VDD Cbb sky130_fd_sc_hd__inv_1
x6 C VSS VSS VDD VDD Cb sky130_fd_sc_hd__inv_1
x7 OUT2 VSS VSS VDD VDD net3 sky130_fd_sc_hd__buf_1
x3 Cbb VSS net1 VDD OUT2 Cb net2 mux2-1
x4 Cbb VSS net2 VDD OUT1 Cb net1 mux2-1
x8 OUT1 VSS VSS VDD VDD buf_out sky130_fd_sc_hd__buf_1
.ends


* expanding   symbol:  mux2-1.sym # of pins=7
* sym_path: /home/users/lsammaro/open-puf/design/mux2-1.sym
* sch_path: /home/users/lsammaro/open-puf/design/mux2-1.sch
.subckt mux2-1  S VSS IN1 VDD OUT Sbar IN2
*.ipin IN1
*.ipin IN2
*.ipin Sbar
*.ipin S
*.opin OUT
*.iopin VSS
*.iopin VDD
XM2 IN1 S OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 IN2 Sbar OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 IN1 Sbar OUT VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 IN2 S OUT VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends

** flattened .save nodes

