magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< pwell >>
rect 10 10 634 146
<< nmoslvt >>
rect 92 36 122 120
rect 178 36 208 120
rect 264 36 294 120
rect 350 36 380 120
rect 436 36 466 120
rect 522 36 552 120
<< ndiff >>
rect 36 101 92 120
rect 36 67 47 101
rect 81 67 92 101
rect 36 36 92 67
rect 122 101 178 120
rect 122 67 133 101
rect 167 67 178 101
rect 122 36 178 67
rect 208 101 264 120
rect 208 67 219 101
rect 253 67 264 101
rect 208 36 264 67
rect 294 101 350 120
rect 294 67 305 101
rect 339 67 350 101
rect 294 36 350 67
rect 380 101 436 120
rect 380 67 391 101
rect 425 67 436 101
rect 380 36 436 67
rect 466 101 522 120
rect 466 67 477 101
rect 511 67 522 101
rect 466 36 522 67
rect 552 101 608 120
rect 552 67 563 101
rect 597 67 608 101
rect 552 36 608 67
<< ndiffc >>
rect 47 67 81 101
rect 133 67 167 101
rect 219 67 253 101
rect 305 67 339 101
rect 391 67 425 101
rect 477 67 511 101
rect 563 67 597 101
<< poly >>
rect 92 201 552 217
rect 92 167 135 201
rect 169 167 203 201
rect 237 167 271 201
rect 305 167 339 201
rect 373 167 407 201
rect 441 167 475 201
rect 509 167 552 201
rect 92 146 552 167
rect 92 120 122 146
rect 178 120 208 146
rect 264 120 294 146
rect 350 120 380 146
rect 436 120 466 146
rect 522 120 552 146
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
rect 436 10 466 36
rect 522 10 552 36
<< polycont >>
rect 135 167 169 201
rect 203 167 237 201
rect 271 167 305 201
rect 339 167 373 201
rect 407 167 441 201
rect 475 167 509 201
<< locali >>
rect 119 201 525 217
rect 119 167 125 201
rect 169 167 197 201
rect 237 167 269 201
rect 305 167 339 201
rect 375 167 407 201
rect 447 167 475 201
rect 519 167 525 201
rect 119 151 525 167
rect 47 101 81 117
rect 47 51 81 67
rect 133 101 167 117
rect 133 51 167 67
rect 219 101 253 117
rect 219 51 253 67
rect 305 101 339 117
rect 305 51 339 67
rect 391 101 425 117
rect 391 51 425 67
rect 477 101 511 117
rect 477 51 511 67
rect 563 101 597 117
rect 563 51 597 67
<< viali >>
rect 125 167 135 201
rect 135 167 159 201
rect 197 167 203 201
rect 203 167 231 201
rect 269 167 271 201
rect 271 167 303 201
rect 341 167 373 201
rect 373 167 375 201
rect 413 167 441 201
rect 441 167 447 201
rect 485 167 509 201
rect 509 167 519 201
rect 47 67 81 101
rect 133 67 167 101
rect 219 67 253 101
rect 305 67 339 101
rect 391 67 425 101
rect 477 67 511 101
rect 563 67 597 101
<< metal1 >>
rect 113 201 531 213
rect 113 167 125 201
rect 159 167 197 201
rect 231 167 269 201
rect 303 167 341 201
rect 375 167 413 201
rect 447 167 485 201
rect 519 167 531 201
rect 113 155 531 167
rect 41 101 87 117
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 124 108 176 117
rect 124 49 176 56
rect 213 101 259 117
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 296 108 348 117
rect 296 49 348 56
rect 385 101 431 117
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 468 108 520 117
rect 468 49 520 56
rect 557 101 603 117
rect 557 67 563 101
rect 597 67 603 101
rect 557 -29 603 67
rect 41 -89 603 -29
<< via1 >>
rect 124 101 176 108
rect 124 67 133 101
rect 133 67 167 101
rect 167 67 176 101
rect 124 56 176 67
rect 296 101 348 108
rect 296 67 305 101
rect 305 67 339 101
rect 339 67 348 101
rect 296 56 348 67
rect 468 101 520 108
rect 468 67 477 101
rect 477 67 511 101
rect 511 67 520 101
rect 468 56 520 67
<< metal2 >>
rect 122 108 178 115
rect 122 106 124 108
rect 176 106 178 108
rect 122 41 178 50
rect 294 108 350 115
rect 294 106 296 108
rect 348 106 350 108
rect 294 41 350 50
rect 466 108 522 115
rect 466 106 468 108
rect 520 106 522 108
rect 466 41 522 50
<< via2 >>
rect 122 56 124 106
rect 124 56 176 106
rect 176 56 178 106
rect 122 50 178 56
rect 294 56 296 106
rect 296 56 348 106
rect 348 56 350 106
rect 294 50 350 56
rect 466 56 468 106
rect 468 56 520 106
rect 520 56 522 106
rect 466 50 522 56
<< metal3 >>
rect 117 106 527 111
rect 117 50 122 106
rect 178 50 294 106
rect 350 50 466 106
rect 522 50 527 106
rect 117 45 527 50
<< labels >>
flabel metal3 s 117 45 527 111 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 41 -89 603 -29 0 FreeSans 400 0 0 0 SOURCE
port 2 nsew
flabel metal1 s 113 155 531 213 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel pwell s 77 128 90 142 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 5904622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5897008
string path 1.600 2.925 1.600 -2.225 
<< end >>
