magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 13 43 764 283
rect -26 -43 794 43
<< locali >>
rect 121 435 313 498
rect 673 435 743 751
rect 121 162 187 329
rect 223 162 451 329
rect 682 99 743 435
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 112 735 302 741
rect 112 701 118 735
rect 152 701 190 735
rect 224 701 262 735
rect 296 701 302 735
rect 26 399 76 609
rect 112 534 302 701
rect 440 735 630 751
rect 440 701 446 735
rect 480 701 518 735
rect 552 701 590 735
rect 624 701 630 735
rect 354 399 404 609
rect 440 435 630 701
rect 26 365 648 399
rect 26 165 85 365
rect 582 333 648 365
rect 487 113 648 265
rect 487 79 497 113
rect 531 79 603 113
rect 637 79 648 113
rect 487 73 648 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 118 701 152 735
rect 190 701 224 735
rect 262 701 296 735
rect 446 701 480 735
rect 518 701 552 735
rect 590 701 624 735
rect 497 79 531 113
rect 603 79 637 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 118 735
rect 152 701 190 735
rect 224 701 262 735
rect 296 701 446 735
rect 480 701 518 735
rect 552 701 590 735
rect 624 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 497 113
rect 531 79 603 113
rect 637 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel locali s 121 162 187 329 6 A
port 1 nsew signal input
rlabel locali s 121 435 313 498 6 B
port 2 nsew signal input
rlabel locali s 223 162 451 329 6 C
port 3 nsew signal input
rlabel metal1 s 0 51 768 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 768 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 794 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 13 43 764 283 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 768 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 834 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 768 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 682 99 743 435 6 X
port 8 nsew signal output
rlabel locali s 673 435 743 751 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 768 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 813630
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 803460
<< end >>
