magic
tech sky130A
magscale 1 2
timestamp 1654292831
<< nwell >>
rect 27786 -2335 28723 -2334
rect 27706 -2656 28723 -2335
rect 30250 -2656 30618 -2335
<< nsubdiff >>
rect 30374 -2466 30508 -2449
rect 30374 -2500 30402 -2466
rect 30436 -2500 30508 -2466
rect 30374 -2519 30508 -2500
<< nsubdiffcont >>
rect 30402 -2500 30436 -2466
<< locali >>
rect 30363 -2457 30522 -2425
rect 30171 -2466 30522 -2457
rect 30171 -2500 30402 -2466
rect 30436 -2500 30522 -2466
rect 30171 -2514 30522 -2500
rect 30363 -2533 30522 -2514
<< viali >>
rect 27597 -2580 27631 -2546
rect 29040 -2563 29074 -2529
rect 29208 -2563 29242 -2529
rect 29376 -2563 29410 -2529
rect 29544 -2563 29578 -2529
rect 29712 -2563 29746 -2529
rect 29880 -2563 29914 -2529
rect 30048 -2563 30082 -2529
rect 30788 -2564 30822 -2530
rect 30956 -2564 30990 -2530
rect 31124 -2564 31158 -2530
rect 31292 -2564 31326 -2530
rect 31460 -2564 31494 -2530
rect 31628 -2564 31662 -2530
rect 31796 -2564 31830 -2530
rect 28049 -2700 28083 -2666
rect 28135 -2700 28169 -2666
rect 28609 -2702 28643 -2668
rect 28800 -2698 28834 -2664
rect 28919 -2698 28953 -2664
rect 29038 -2698 29072 -2664
rect 29157 -2698 29191 -2664
rect 29276 -2698 29310 -2664
rect 29395 -2698 29429 -2664
rect 29514 -2698 29548 -2664
rect 30724 -2696 30758 -2662
rect 30843 -2696 30877 -2662
rect 30962 -2696 30996 -2662
rect 31081 -2696 31115 -2662
rect 31200 -2696 31234 -2662
rect 31319 -2696 31353 -2662
rect 31438 -2696 31472 -2662
<< metal1 >>
rect 86 1593 444 1613
rect 86 1592 386 1593
rect 86 1540 110 1592
rect 162 1541 386 1592
rect 438 1541 444 1593
rect 162 1540 444 1541
rect 86 1516 444 1540
rect 60809 851 61053 929
rect 27668 -2421 28740 -2325
rect 30212 -2421 30678 -2325
rect 27578 -2546 27642 -2505
rect 27578 -2580 27597 -2546
rect 27631 -2580 27642 -2546
rect -317 -2720 27469 -2646
rect 27578 -2647 27642 -2580
rect 29028 -2529 31845 -2504
rect 29028 -2563 29040 -2529
rect 29074 -2563 29208 -2529
rect 29242 -2563 29376 -2529
rect 29410 -2563 29544 -2529
rect 29578 -2563 29712 -2529
rect 29746 -2563 29880 -2529
rect 29914 -2563 30048 -2529
rect 30082 -2530 31845 -2529
rect 30082 -2538 30788 -2530
rect 30082 -2563 30260 -2538
rect 29028 -2590 30260 -2563
rect 30312 -2590 30363 -2538
rect 30415 -2590 30466 -2538
rect 30518 -2590 30569 -2538
rect 30621 -2564 30788 -2538
rect 30822 -2564 30956 -2530
rect 30990 -2564 31124 -2530
rect 31158 -2564 31292 -2530
rect 31326 -2564 31460 -2530
rect 31494 -2564 31628 -2530
rect 31662 -2564 31796 -2530
rect 31830 -2564 31845 -2530
rect 30621 -2590 31845 -2564
rect 29028 -2612 31845 -2590
rect 27578 -2666 28256 -2647
rect 27578 -2700 28049 -2666
rect 28083 -2700 28135 -2666
rect 28169 -2700 28256 -2666
rect 27578 -2711 28256 -2700
rect 28587 -2662 31768 -2653
rect 28587 -2664 30724 -2662
rect 28587 -2668 28800 -2664
rect 28587 -2702 28609 -2668
rect 28643 -2698 28800 -2668
rect 28834 -2698 28919 -2664
rect 28953 -2698 29038 -2664
rect 29072 -2698 29157 -2664
rect 29191 -2698 29276 -2664
rect 29310 -2698 29395 -2664
rect 29429 -2698 29514 -2664
rect 29548 -2696 30724 -2664
rect 30758 -2696 30843 -2662
rect 30877 -2696 30962 -2662
rect 30996 -2696 31081 -2662
rect 31115 -2696 31200 -2662
rect 31234 -2696 31319 -2662
rect 31353 -2696 31438 -2662
rect 31472 -2696 31768 -2662
rect 29548 -2698 31768 -2696
rect 28643 -2702 31768 -2698
rect 28587 -2710 31768 -2702
rect 27668 -2965 28773 -2869
rect 30212 -2965 30678 -2869
rect -167 -6186 614 -6171
rect -167 -6194 555 -6186
rect -167 -6246 -150 -6194
rect -98 -6238 555 -6194
rect 607 -6238 614 -6186
rect -98 -6246 614 -6238
rect -167 -6264 614 -6246
<< via1 >>
rect 30296 3154 30348 3206
rect 30413 3154 30465 3206
rect 30530 3154 30582 3206
rect 110 1540 162 1592
rect 386 1541 438 1593
rect 31363 -2407 31415 -2355
rect 31493 -2407 31545 -2355
rect 31623 -2407 31675 -2355
rect 30260 -2590 30312 -2538
rect 30363 -2590 30415 -2538
rect 30466 -2590 30518 -2538
rect 30569 -2590 30621 -2538
rect 31353 -2937 31405 -2885
rect 31466 -2937 31518 -2885
rect 31579 -2937 31631 -2885
rect 31692 -2937 31744 -2885
rect 31805 -2937 31857 -2885
rect 31353 -4826 31405 -4774
rect 31466 -4826 31518 -4774
rect 31579 -4826 31631 -4774
rect 31692 -4826 31744 -4774
rect 31805 -4826 31857 -4774
rect 31353 -4931 31405 -4879
rect 31466 -4931 31518 -4879
rect 31579 -4931 31631 -4879
rect 31692 -4931 31744 -4879
rect 31805 -4931 31857 -4879
rect -150 -6246 -98 -6194
rect 555 -6238 607 -6186
rect 30285 -9075 30337 -9023
rect 30368 -9075 30420 -9023
rect 30451 -9075 30503 -9023
rect 30534 -9075 30586 -9023
<< metal2 >>
rect 1839 6719 1883 7341
rect 3727 6719 3771 7341
rect 5615 6719 5659 7341
rect 7503 6719 7547 7341
rect 9391 6719 9435 7341
rect 11279 6719 11323 7341
rect 13167 6719 13211 7341
rect 15055 6719 15099 7341
rect 16943 6719 16987 7341
rect 18831 6719 18875 7341
rect 20719 6719 20763 7341
rect 22607 6719 22651 7341
rect 24495 6719 24539 7341
rect 26383 6719 26427 7341
rect 28271 6719 28315 7341
rect 30159 6719 30203 7341
rect 32047 6719 32091 7341
rect 33935 6719 33979 7341
rect 35823 6719 35867 7341
rect 37711 6719 37755 7341
rect 39599 6719 39643 7341
rect 41487 6719 41531 7341
rect 43375 6719 43419 7341
rect 45263 6719 45307 7341
rect 47151 6719 47195 7341
rect 49039 6719 49083 7341
rect 50927 6719 50971 7341
rect 52815 6719 52859 7341
rect 54703 6719 54747 7341
rect 56591 6719 56635 7341
rect 58479 6719 58523 7341
rect 60367 6719 60411 7341
rect 60942 6037 60978 6070
rect -159 6001 555 6037
rect 60231 6001 60978 6037
rect -159 -6171 -123 6001
rect 30232 3261 30628 3290
rect 30232 3205 30263 3261
rect 30319 3206 30372 3261
rect 30428 3206 30481 3261
rect 30537 3206 30628 3261
rect 30348 3205 30372 3206
rect 30465 3205 30481 3206
rect 30232 3159 30296 3205
rect 30348 3159 30413 3205
rect 30465 3159 30530 3205
rect 30232 3103 30263 3159
rect 30348 3154 30372 3159
rect 30465 3154 30481 3159
rect 30582 3154 30628 3206
rect 30319 3103 30372 3154
rect 30428 3103 30481 3154
rect 30537 3103 30628 3154
rect 30232 3082 30628 3103
rect 75 1592 173 1619
rect 75 1540 110 1592
rect 162 1540 173 1592
rect 75 1500 173 1540
rect 373 1593 477 1616
rect 373 1541 386 1593
rect 438 1581 477 1593
rect 60942 1581 60978 6001
rect 438 1545 649 1581
rect 60325 1545 60978 1581
rect 438 1541 477 1545
rect 373 1516 477 1541
rect -160 -6194 -49 -6171
rect -160 -6246 -150 -6194
rect -98 -6246 -49 -6194
rect -160 -6286 -49 -6246
rect 107 -10650 143 1500
rect 469 241 513 863
rect 2357 241 2401 863
rect 4245 241 4289 863
rect 6133 241 6177 863
rect 8021 241 8065 863
rect 9909 241 9953 863
rect 11797 241 11841 863
rect 13685 241 13729 863
rect 15573 241 15617 863
rect 17461 241 17505 863
rect 19349 241 19393 863
rect 21237 241 21281 863
rect 23125 241 23169 863
rect 25013 241 25057 863
rect 26901 241 26945 863
rect 28789 241 28833 863
rect 30677 241 30721 863
rect 32565 241 32609 863
rect 34453 241 34497 863
rect 36341 241 36385 863
rect 38229 241 38273 863
rect 40117 241 40161 863
rect 42005 241 42049 863
rect 43893 241 43937 863
rect 45781 241 45825 863
rect 47669 241 47713 863
rect 49557 241 49601 863
rect 51445 241 51489 863
rect 53333 241 53377 863
rect 55221 241 55265 863
rect 57109 241 57153 863
rect 58997 241 59041 863
rect 30233 -1921 30630 -1882
rect 30233 -1977 30256 -1921
rect 30312 -1977 30360 -1921
rect 30416 -1977 30464 -1921
rect 30520 -1977 30568 -1921
rect 30624 -1977 30630 -1921
rect 30233 -2020 30630 -1977
rect 30233 -2076 30256 -2020
rect 30312 -2076 30360 -2020
rect 30416 -2076 30464 -2020
rect 30520 -2076 30568 -2020
rect 30624 -2076 30630 -2020
rect 30233 -2538 30630 -2076
rect 31324 -2351 31725 -2326
rect 31324 -2407 31363 -2351
rect 31419 -2407 31492 -2351
rect 31548 -2407 31621 -2351
rect 31677 -2407 31725 -2351
rect 31324 -2420 31725 -2407
rect 30233 -2590 30260 -2538
rect 30312 -2590 30363 -2538
rect 30415 -2590 30466 -2538
rect 30518 -2590 30569 -2538
rect 30621 -2590 30630 -2538
rect 30233 -3250 30630 -2590
rect 30233 -3306 30269 -3250
rect 30325 -3306 30357 -3250
rect 30413 -3306 30445 -3250
rect 30501 -3306 30533 -3250
rect 30589 -3306 30630 -3250
rect 30233 -3345 30630 -3306
rect 30233 -3401 30269 -3345
rect 30325 -3401 30357 -3345
rect 30413 -3401 30445 -3345
rect 30501 -3401 30533 -3345
rect 30589 -3401 30630 -3345
rect 30233 -3432 30630 -3401
rect 31298 -2885 31965 -2868
rect 31298 -2937 31353 -2885
rect 31405 -2937 31466 -2885
rect 31518 -2937 31579 -2885
rect 31631 -2937 31692 -2885
rect 31744 -2937 31805 -2885
rect 31857 -2937 31965 -2885
rect 31298 -4774 31965 -2937
rect 31298 -4826 31353 -4774
rect 31405 -4826 31466 -4774
rect 31518 -4826 31579 -4774
rect 31631 -4826 31692 -4774
rect 31744 -4826 31805 -4774
rect 31857 -4826 31965 -4774
rect 31298 -4879 31965 -4826
rect 698 -5512 742 -4890
rect 2586 -5512 2630 -4890
rect 4474 -5512 4518 -4890
rect 6362 -5512 6406 -4890
rect 8250 -5512 8294 -4890
rect 10138 -5512 10182 -4890
rect 12026 -5512 12070 -4890
rect 13914 -5512 13958 -4890
rect 15802 -5512 15846 -4890
rect 17690 -5512 17734 -4890
rect 19578 -5512 19622 -4890
rect 21466 -5512 21510 -4890
rect 23354 -5512 23398 -4890
rect 25242 -5512 25286 -4890
rect 27130 -5512 27174 -4890
rect 29018 -5512 29062 -4890
rect 30906 -5512 30950 -4890
rect 31298 -4931 31353 -4879
rect 31405 -4931 31466 -4879
rect 31518 -4931 31579 -4879
rect 31631 -4931 31692 -4879
rect 31744 -4931 31805 -4879
rect 31857 -4931 31965 -4879
rect 31298 -4979 31965 -4931
rect 32794 -5512 32838 -4890
rect 34682 -5512 34726 -4890
rect 36570 -5512 36614 -4890
rect 38458 -5512 38502 -4890
rect 40346 -5512 40390 -4890
rect 42234 -5512 42278 -4890
rect 44122 -5512 44166 -4890
rect 46010 -5512 46054 -4890
rect 47898 -5512 47942 -4890
rect 49786 -5512 49830 -4890
rect 51674 -5512 51718 -4890
rect 53562 -5512 53606 -4890
rect 55450 -5512 55494 -4890
rect 57338 -5512 57382 -4890
rect 59226 -5512 59270 -4890
rect 548 -6186 618 -6165
rect 548 -6238 555 -6186
rect 607 -6194 618 -6186
rect 607 -6230 878 -6194
rect 60554 -6230 61279 -6194
rect 607 -6238 618 -6230
rect 548 -6269 618 -6238
rect 30233 -8974 30630 -8941
rect 30233 -9030 30274 -8974
rect 30330 -9023 30366 -8974
rect 30422 -9023 30458 -8974
rect 30514 -9023 30550 -8974
rect 30337 -9030 30366 -9023
rect 30422 -9030 30451 -9023
rect 30514 -9030 30534 -9023
rect 30606 -9030 30630 -8974
rect 30233 -9065 30285 -9030
rect 30337 -9065 30368 -9030
rect 30420 -9065 30451 -9030
rect 30503 -9065 30534 -9030
rect 30586 -9065 30630 -9030
rect 30233 -9121 30274 -9065
rect 30337 -9075 30366 -9065
rect 30422 -9075 30451 -9065
rect 30514 -9075 30534 -9065
rect 30330 -9121 30366 -9075
rect 30422 -9121 30458 -9075
rect 30514 -9121 30550 -9075
rect 30606 -9121 30630 -9065
rect 30233 -9147 30630 -9121
rect 61243 -10650 61279 -6230
rect 107 -10686 784 -10650
rect 60460 -10686 61279 -10650
rect 61243 -10697 61279 -10686
rect 2068 -11990 2112 -11368
rect 3956 -11990 4000 -11368
rect 5844 -11990 5888 -11368
rect 7732 -11990 7776 -11368
rect 9620 -11990 9664 -11368
rect 11508 -11990 11552 -11368
rect 13396 -11990 13440 -11368
rect 15284 -11990 15328 -11368
rect 17172 -11990 17216 -11368
rect 19060 -11990 19104 -11368
rect 20948 -11990 20992 -11368
rect 22836 -11990 22880 -11368
rect 24724 -11990 24768 -11368
rect 26612 -11990 26656 -11368
rect 28500 -11990 28544 -11368
rect 30388 -11990 30432 -11368
rect 32276 -11990 32320 -11368
rect 34164 -11990 34208 -11368
rect 36052 -11990 36096 -11368
rect 37940 -11990 37984 -11368
rect 39828 -11990 39872 -11368
rect 41716 -11990 41760 -11368
rect 43604 -11990 43648 -11368
rect 45492 -11990 45536 -11368
rect 47380 -11990 47424 -11368
rect 49268 -11990 49312 -11368
rect 51156 -11990 51200 -11368
rect 53044 -11990 53088 -11368
rect 54932 -11990 54976 -11368
rect 56820 -11990 56864 -11368
rect 58708 -11990 58752 -11368
rect 60596 -11990 60640 -11368
<< via2 >>
rect 30263 3206 30319 3261
rect 30372 3206 30428 3261
rect 30481 3206 30537 3261
rect 30263 3205 30296 3206
rect 30296 3205 30319 3206
rect 30372 3205 30413 3206
rect 30413 3205 30428 3206
rect 30481 3205 30530 3206
rect 30530 3205 30537 3206
rect 30263 3154 30296 3159
rect 30296 3154 30319 3159
rect 30372 3154 30413 3159
rect 30413 3154 30428 3159
rect 30481 3154 30530 3159
rect 30530 3154 30537 3159
rect 30263 3103 30319 3154
rect 30372 3103 30428 3154
rect 30481 3103 30537 3154
rect 30256 -1977 30312 -1921
rect 30360 -1977 30416 -1921
rect 30464 -1977 30520 -1921
rect 30568 -1977 30624 -1921
rect 30256 -2076 30312 -2020
rect 30360 -2076 30416 -2020
rect 30464 -2076 30520 -2020
rect 30568 -2076 30624 -2020
rect 31363 -2355 31419 -2351
rect 31363 -2407 31415 -2355
rect 31415 -2407 31419 -2355
rect 31492 -2355 31548 -2351
rect 31492 -2407 31493 -2355
rect 31493 -2407 31545 -2355
rect 31545 -2407 31548 -2355
rect 31621 -2355 31677 -2351
rect 31621 -2407 31623 -2355
rect 31623 -2407 31675 -2355
rect 31675 -2407 31677 -2355
rect 30269 -3306 30325 -3250
rect 30357 -3306 30413 -3250
rect 30445 -3306 30501 -3250
rect 30533 -3306 30589 -3250
rect 30269 -3401 30325 -3345
rect 30357 -3401 30413 -3345
rect 30445 -3401 30501 -3345
rect 30533 -3401 30589 -3345
rect 30274 -9023 30330 -8974
rect 30366 -9023 30422 -8974
rect 30458 -9023 30514 -8974
rect 30550 -9023 30606 -8974
rect 30274 -9030 30285 -9023
rect 30285 -9030 30330 -9023
rect 30366 -9030 30368 -9023
rect 30368 -9030 30420 -9023
rect 30420 -9030 30422 -9023
rect 30458 -9030 30503 -9023
rect 30503 -9030 30514 -9023
rect 30550 -9030 30586 -9023
rect 30586 -9030 30606 -9023
rect 30274 -9075 30285 -9065
rect 30285 -9075 30330 -9065
rect 30366 -9075 30368 -9065
rect 30368 -9075 30420 -9065
rect 30420 -9075 30422 -9065
rect 30458 -9075 30503 -9065
rect 30503 -9075 30514 -9065
rect 30550 -9075 30586 -9065
rect 30586 -9075 30606 -9065
rect 30274 -9121 30330 -9075
rect 30366 -9121 30422 -9075
rect 30458 -9121 30514 -9075
rect 30550 -9121 30606 -9075
<< metal3 >>
rect 30232 3261 30627 3290
rect 30232 3205 30263 3261
rect 30319 3238 30372 3261
rect 30428 3205 30481 3261
rect 30537 3205 30627 3261
rect 30232 3159 30306 3205
rect 30402 3159 30627 3205
rect 30232 3103 30263 3159
rect 30319 3103 30372 3130
rect 30428 3103 30481 3159
rect 30537 3103 30627 3159
rect 30232 3082 30627 3103
rect 30232 -1921 30629 -1879
rect 30232 -1977 30256 -1921
rect 30312 -1946 30360 -1921
rect 30416 -1977 30464 -1921
rect 30520 -1946 30568 -1921
rect 30624 -1977 30629 -1921
rect 30232 -2020 30297 -1977
rect 30393 -2020 30479 -1977
rect 30575 -2020 30629 -1977
rect 30232 -2076 30256 -2020
rect 30312 -2076 30360 -2054
rect 30416 -2076 30464 -2020
rect 30520 -2076 30568 -2054
rect 30624 -2076 30629 -2020
rect 30232 -2103 30629 -2076
rect 31324 -2337 31725 -2326
rect 31324 -2351 31445 -2337
rect 31619 -2351 31725 -2337
rect 31324 -2407 31363 -2351
rect 31419 -2401 31445 -2351
rect 31619 -2401 31621 -2351
rect 31419 -2407 31492 -2401
rect 31548 -2407 31621 -2401
rect 31677 -2407 31725 -2351
rect 31324 -2420 31725 -2407
rect 30233 -3250 30630 -3192
rect 30233 -3306 30269 -3250
rect 30325 -3269 30357 -3250
rect 30413 -3306 30445 -3250
rect 30501 -3269 30533 -3250
rect 30589 -3306 30630 -3250
rect 30233 -3345 30289 -3306
rect 30385 -3345 30479 -3306
rect 30575 -3345 30630 -3306
rect 30233 -3401 30269 -3345
rect 30325 -3401 30357 -3377
rect 30413 -3401 30445 -3345
rect 30501 -3401 30533 -3377
rect 30589 -3401 30630 -3345
rect 30233 -3432 30630 -3401
rect 30233 -8974 30630 -8941
rect 30233 -9030 30274 -8974
rect 30330 -8998 30366 -8974
rect 30422 -9030 30458 -8974
rect 30514 -8997 30550 -8974
rect 30606 -9030 30630 -8974
rect 30233 -9065 30301 -9030
rect 30397 -9065 30475 -9030
rect 30571 -9065 30630 -9030
rect 30233 -9121 30274 -9065
rect 30330 -9121 30366 -9106
rect 30422 -9121 30458 -9065
rect 30514 -9121 30550 -9105
rect 30606 -9121 30630 -9065
rect 30233 -9147 30630 -9121
<< via3 >>
rect 30306 3205 30319 3238
rect 30319 3205 30372 3238
rect 30372 3205 30402 3238
rect 30306 3159 30402 3205
rect 30306 3130 30319 3159
rect 30319 3130 30372 3159
rect 30372 3130 30402 3159
rect 31369 2236 31493 2402
rect 31568 2236 31692 2402
rect 30297 -1977 30312 -1946
rect 30312 -1977 30360 -1946
rect 30360 -1977 30393 -1946
rect 30479 -1977 30520 -1946
rect 30520 -1977 30568 -1946
rect 30568 -1977 30575 -1946
rect 30297 -2020 30393 -1977
rect 30479 -2020 30575 -1977
rect 30297 -2054 30312 -2020
rect 30312 -2054 30360 -2020
rect 30360 -2054 30393 -2020
rect 30479 -2054 30520 -2020
rect 30520 -2054 30568 -2020
rect 30568 -2054 30575 -2020
rect 31445 -2351 31619 -2337
rect 31445 -2401 31492 -2351
rect 31492 -2401 31548 -2351
rect 31548 -2401 31619 -2351
rect 30289 -3306 30325 -3269
rect 30325 -3306 30357 -3269
rect 30357 -3306 30385 -3269
rect 30479 -3306 30501 -3269
rect 30501 -3306 30533 -3269
rect 30533 -3306 30575 -3269
rect 30289 -3345 30385 -3306
rect 30479 -3345 30575 -3306
rect 30289 -3377 30325 -3345
rect 30325 -3377 30357 -3345
rect 30357 -3377 30385 -3345
rect 30479 -3377 30501 -3345
rect 30501 -3377 30533 -3345
rect 30533 -3377 30575 -3345
rect 3205 -4914 3374 -4777
rect 1911 -7041 2080 -6904
rect 30301 -9030 30330 -8998
rect 30330 -9030 30366 -8998
rect 30366 -9030 30397 -8998
rect 30475 -9030 30514 -8997
rect 30514 -9030 30550 -8997
rect 30550 -9030 30571 -8997
rect 30301 -9065 30397 -9030
rect 30475 -9065 30571 -9030
rect 30301 -9106 30330 -9065
rect 30330 -9106 30366 -9065
rect 30366 -9106 30397 -9065
rect 30475 -9105 30514 -9065
rect 30514 -9105 30550 -9065
rect 30550 -9105 30571 -9065
rect 1920 -9981 2089 -9844
rect 3218 -12106 3387 -11969
<< metal4 >>
rect 1683 -6904 2301 5164
rect 1683 -7041 1911 -6904
rect 2080 -7041 2301 -6904
rect 1683 -9844 2301 -7041
rect 1683 -9981 1920 -9844
rect 2089 -9981 2301 -9844
rect 1683 -10071 2301 -9981
rect 2916 -4777 3700 7281
rect 30232 3238 30629 3350
rect 30232 3130 30306 3238
rect 30402 3130 30629 3238
rect 30232 -1442 30629 3130
rect 30231 -1803 30629 -1442
rect 30232 -1946 30629 -1803
rect 30232 -2054 30297 -1946
rect 30393 -2054 30479 -1946
rect 30575 -2054 30629 -1946
rect 30232 -2103 30629 -2054
rect 31317 2402 31721 2521
rect 31317 2236 31369 2402
rect 31493 2236 31568 2402
rect 31692 2236 31721 2402
rect 31317 -2017 31721 2236
rect 31317 -2148 31725 -2017
rect 31324 -2337 31725 -2148
rect 31324 -2401 31445 -2337
rect 31619 -2401 31725 -2337
rect 31324 -2420 31725 -2401
rect 2916 -4914 3205 -4777
rect 3374 -4914 3700 -4777
rect 2916 -11969 3700 -4914
rect 30234 -3269 30630 -3193
rect 30234 -3377 30289 -3269
rect 30385 -3377 30479 -3269
rect 30575 -3377 30630 -3269
rect 30234 -8997 30630 -3377
rect 30234 -8998 30475 -8997
rect 30234 -9106 30301 -8998
rect 30397 -9105 30475 -8998
rect 30571 -9105 30630 -8997
rect 30397 -9106 30630 -9105
rect 30234 -9209 30630 -9106
rect 2916 -12106 3218 -11969
rect 3387 -12106 3700 -11969
rect 2916 -12294 3700 -12106
use BR128half  BR128half_0
timestamp 1654224521
transform 1 0 449 0 1 71
box -430 -58 60604 7443
use BR128half  BR128half_1
timestamp 1654224521
transform -1 0 60660 0 1 -12160
box -430 -58 60604 7443
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 27372 0 1 -2917
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1650294714
transform 1 0 27850 0 1 -2918
box -38 -48 866 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654066915
transform 1 0 28740 0 1 -2917
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654066915
transform 1 0 30656 0 1 -2917
box -38 -48 1510 592
<< labels >>
flabel metal1 60809 851 61053 929 1 FreeSans 800 0 0 0 OUT
port 3 n
flabel metal2 60367 6719 60411 7341 1 FreeSans 800 0 0 0 C[0]
port 131 n
flabel metal2 58479 6719 58523 7341 1 FreeSans 800 0 0 0 C[1]
port 130 n
flabel metal2 56591 6719 56635 7341 1 FreeSans 800 0 0 0 C[2]
port 129 n
flabel metal2 54703 6719 54747 7341 1 FreeSans 800 0 0 0 C[3]
port 128 n
flabel metal2 52815 6719 52859 7341 1 FreeSans 800 0 0 0 C[4]
port 127 n
flabel metal2 50927 6719 50971 7341 1 FreeSans 800 0 0 0 C[5]
port 126 n
flabel metal2 49039 6719 49083 7341 1 FreeSans 800 0 0 0 C[6]
port 125 n
flabel metal2 47151 6719 47195 7341 1 FreeSans 800 0 0 0 C[7]
port 124 n
flabel metal2 45263 6719 45307 7341 1 FreeSans 800 0 0 0 C[8]
port 123 n
flabel metal2 43375 6719 43419 7341 1 FreeSans 800 0 0 0 C[9]
port 122 n
flabel metal2 41487 6719 41531 7341 1 FreeSans 800 0 0 0 C[10]
port 121 n
flabel metal2 39599 6719 39643 7341 1 FreeSans 800 0 0 0 C[11]
port 120 n
flabel metal2 37711 6719 37755 7341 1 FreeSans 800 0 0 0 C[12]
port 119 n
flabel metal2 35823 6719 35867 7341 1 FreeSans 800 0 0 0 C[13]
port 118 n
flabel metal2 33935 6719 33979 7341 1 FreeSans 800 0 0 0 C[14]
port 117 n
flabel metal2 32047 6719 32091 7341 1 FreeSans 800 0 0 0 C[15]
port 116 n
flabel metal2 30159 6719 30203 7341 1 FreeSans 800 0 0 0 C[16]
port 115 n
flabel metal2 28271 6719 28315 7341 1 FreeSans 800 0 0 0 C[17]
port 114 n
flabel metal2 26383 6719 26427 7341 1 FreeSans 800 0 0 0 C[18]
port 113 n
flabel metal2 24495 6719 24539 7341 1 FreeSans 800 0 0 0 C[19]
port 112 n
flabel metal2 22607 6719 22651 7341 1 FreeSans 800 0 0 0 C[20]
port 111 n
flabel metal2 20719 6719 20763 7341 1 FreeSans 800 0 0 0 C[21]
port 110 n
flabel metal2 18831 6719 18875 7341 1 FreeSans 800 0 0 0 C[22]
port 109 n
flabel metal2 16943 6719 16987 7341 1 FreeSans 800 0 0 0 C[23]
port 108 n
flabel metal2 15055 6719 15099 7341 1 FreeSans 800 0 0 0 C[24]
port 107 n
flabel metal2 13167 6719 13211 7341 1 FreeSans 800 0 0 0 C[25]
port 106 n
flabel metal2 11279 6719 11323 7341 1 FreeSans 800 0 0 0 C[26]
port 105 n
flabel metal2 9391 6719 9435 7341 1 FreeSans 800 0 0 0 C[27]
port 104 n
flabel metal2 7503 6719 7547 7341 1 FreeSans 800 0 0 0 C[28]
port 103 n
flabel metal2 5615 6719 5659 7341 1 FreeSans 800 0 0 0 C[29]
port 102 n
flabel metal2 3727 6719 3771 7341 1 FreeSans 800 0 0 0 C[30]
port 101 n
flabel metal2 1839 6719 1883 7341 1 FreeSans 800 0 0 0 C[31]
port 100 n
flabel metal2 698 -5512 742 -4890 1 FreeSans 800 0 0 0 C[32]
port 99 n
flabel metal2 2586 -5512 2630 -4890 1 FreeSans 800 0 0 0 C[33]
port 98 n
flabel metal2 4474 -5512 4518 -4890 1 FreeSans 800 0 0 0 C[34]
port 97 n
flabel metal2 6362 -5512 6406 -4890 1 FreeSans 800 0 0 0 C[35]
port 96 n
flabel metal2 8250 -5512 8294 -4890 1 FreeSans 800 0 0 0 C[36]
port 95 n
flabel metal2 10138 -5512 10182 -4890 1 FreeSans 800 0 0 0 C[37]
port 94 n
flabel metal2 12026 -5512 12070 -4890 1 FreeSans 800 0 0 0 C[38]
port 93 n
flabel metal2 13914 -5512 13958 -4890 1 FreeSans 800 0 0 0 C[39]
port 92 n
flabel metal2 15802 -5512 15846 -4890 1 FreeSans 800 0 0 0 C[40]
port 91 n
flabel metal2 17690 -5512 17734 -4890 1 FreeSans 800 0 0 0 C[41]
port 90 n
flabel metal2 19578 -5512 19622 -4890 1 FreeSans 800 0 0 0 C[42]
port 89 n
flabel metal2 21466 -5512 21510 -4890 1 FreeSans 800 0 0 0 C[43]
port 88 n
flabel metal2 23354 -5512 23398 -4890 1 FreeSans 800 0 0 0 C[44]
port 87 n
flabel metal2 25242 -5512 25286 -4890 1 FreeSans 800 0 0 0 C[45]
port 86 n
flabel metal2 27130 -5512 27174 -4890 1 FreeSans 800 0 0 0 C[46]
port 85 n
flabel metal2 29018 -5512 29062 -4890 1 FreeSans 800 0 0 0 C[47]
port 84 n
flabel metal2 30906 -5512 30950 -4890 1 FreeSans 800 0 0 0 C[48]
port 83 n
flabel metal2 32794 -5512 32838 -4890 1 FreeSans 800 0 0 0 C[49]
port 82 n
flabel metal2 34682 -5512 34726 -4890 1 FreeSans 800 0 0 0 C[50]
port 81 n
flabel metal2 36570 -5512 36614 -4890 1 FreeSans 800 0 0 0 C[51]
port 80 n
flabel metal2 38458 -5512 38502 -4890 1 FreeSans 800 0 0 0 C[52]
port 79 n
flabel metal2 40346 -5512 40390 -4890 1 FreeSans 800 0 0 0 C[53]
port 78 n
flabel metal2 42234 -5512 42278 -4890 1 FreeSans 800 0 0 0 C[54]
port 77 n
flabel metal2 44122 -5512 44166 -4890 1 FreeSans 800 0 0 0 C[55]
port 76 n
flabel metal2 46010 -5512 46054 -4890 1 FreeSans 800 0 0 0 C[56]
port 75 n
flabel metal2 47898 -5512 47942 -4890 1 FreeSans 800 0 0 0 C[57]
port 74 n
flabel metal2 49786 -5512 49830 -4890 1 FreeSans 800 0 0 0 C[58]
port 73 n
flabel metal2 51674 -5512 51718 -4890 1 FreeSans 800 0 0 0 C[59]
port 72 n
flabel metal2 53562 -5512 53606 -4890 1 FreeSans 800 0 0 0 C[60]
port 71 n
flabel metal2 55450 -5512 55494 -4890 1 FreeSans 800 0 0 0 C[61]
port 70 n
flabel metal2 57338 -5512 57382 -4890 1 FreeSans 800 0 0 0 C[62]
port 69 n
flabel metal2 59226 -5512 59270 -4890 1 FreeSans 800 0 0 0 C[63]
port 68 n
flabel metal2 60596 -11990 60640 -11368 1 FreeSans 800 0 0 0 C[64]
port 67 n
flabel metal2 58708 -11990 58752 -11368 1 FreeSans 800 0 0 0 C[65]
port 66 n
flabel metal2 56820 -11990 56864 -11368 1 FreeSans 800 0 0 0 C[66]
port 65 n
flabel metal2 54932 -11990 54976 -11368 1 FreeSans 800 0 0 0 C[67]
port 64 n
flabel metal2 53044 -11990 53088 -11368 1 FreeSans 800 0 0 0 C[68]
port 63 n
flabel metal2 51156 -11990 51200 -11368 1 FreeSans 800 0 0 0 C[69]
port 62 n
flabel metal2 49268 -11990 49312 -11368 1 FreeSans 800 0 0 0 C[70]
port 61 n
flabel metal2 47380 -11990 47424 -11368 1 FreeSans 800 0 0 0 C[71]
port 60 n
flabel metal2 45492 -11990 45536 -11368 1 FreeSans 800 0 0 0 C[72]
port 59 n
flabel metal2 43604 -11990 43648 -11368 1 FreeSans 800 0 0 0 C[73]
port 58 n
flabel metal2 41716 -11990 41760 -11368 1 FreeSans 800 0 0 0 C[74]
port 57 n
flabel metal2 39828 -11990 39872 -11368 1 FreeSans 800 0 0 0 C[75]
port 56 n
flabel metal2 37940 -11990 37984 -11368 1 FreeSans 800 0 0 0 C[76]
port 55 n
flabel metal2 36052 -11990 36096 -11368 1 FreeSans 800 0 0 0 C[77]
port 54 n
flabel metal2 34164 -11990 34208 -11368 1 FreeSans 800 0 0 0 C[78]
port 53 n
flabel metal2 32276 -11990 32320 -11368 1 FreeSans 800 0 0 0 C[79]
port 52 n
flabel metal2 30388 -11990 30432 -11368 1 FreeSans 800 0 0 0 C[80]
port 51 n
flabel metal2 28500 -11990 28544 -11368 1 FreeSans 800 0 0 0 C[81]
port 50 n
flabel metal2 26612 -11990 26656 -11368 1 FreeSans 800 0 0 0 C[82]
port 49 n
flabel metal2 24724 -11990 24768 -11368 1 FreeSans 800 0 0 0 C[83]
port 48 n
flabel metal2 22836 -11990 22880 -11368 1 FreeSans 800 0 0 0 C[84]
port 47 n
flabel metal2 20948 -11990 20992 -11368 1 FreeSans 800 0 0 0 C[85]
port 46 n
flabel metal2 19060 -11990 19104 -11368 1 FreeSans 800 0 0 0 C[86]
port 45 n
flabel metal2 17172 -11990 17216 -11368 1 FreeSans 800 0 0 0 C[87]
port 44 n
flabel metal2 15284 -11990 15328 -11368 1 FreeSans 800 0 0 0 C[88]
port 43 n
flabel metal2 13396 -11990 13440 -11368 1 FreeSans 800 0 0 0 C[89]
port 42 n
flabel metal2 11508 -11990 11552 -11368 1 FreeSans 800 0 0 0 C[90]
port 41 n
flabel metal2 9620 -11990 9664 -11368 1 FreeSans 800 0 0 0 C[91]
port 40 n
flabel metal2 7732 -11990 7776 -11368 1 FreeSans 800 0 0 0 C[92]
port 39 n
flabel metal2 5844 -11990 5888 -11368 1 FreeSans 800 0 0 0 C[93]
port 38 n
flabel metal2 3956 -11990 4000 -11368 1 FreeSans 800 0 0 0 C[94]
port 37 n
flabel metal2 2068 -11990 2112 -11368 1 FreeSans 800 0 0 0 C[95]
port 36 n
flabel metal2 469 241 513 863 1 FreeSans 800 0 0 0 C[96]
port 35 n
flabel metal2 2357 241 2401 863 1 FreeSans 800 0 0 0 C[97]
port 34 n
flabel metal2 4245 241 4289 863 1 FreeSans 800 0 0 0 C[98]
port 33 n
flabel metal2 6133 241 6177 863 1 FreeSans 800 0 0 0 C[99]
port 32 n
flabel metal2 8021 241 8065 863 1 FreeSans 800 0 0 0 C[100]
port 31 n
flabel metal2 9909 241 9953 863 1 FreeSans 800 0 0 0 C[101]
port 30 n
flabel metal2 11797 241 11841 863 1 FreeSans 800 0 0 0 C[102]
port 29 n
flabel metal2 13685 241 13729 863 1 FreeSans 800 0 0 0 C[103]
port 28 n
flabel metal2 15573 241 15617 863 1 FreeSans 800 0 0 0 C[104]
port 27 n
flabel metal2 17461 241 17505 863 1 FreeSans 800 0 0 0 C[105]
port 26 n
flabel metal2 19349 241 19393 863 1 FreeSans 800 0 0 0 C[106]
port 25 n
flabel metal2 21237 241 21281 863 1 FreeSans 800 0 0 0 C[107]
port 24 n
flabel metal2 23125 241 23169 863 1 FreeSans 800 0 0 0 C[108]
port 23 n
flabel metal2 25013 241 25057 863 1 FreeSans 800 0 0 0 C[109]
port 22 n
flabel metal2 26901 241 26945 863 1 FreeSans 800 0 0 0 C[110]
port 21 n
flabel metal2 28789 241 28833 863 1 FreeSans 800 0 0 0 C[111]
port 20 n
flabel metal2 30677 241 30721 863 1 FreeSans 800 0 0 0 C[112]
port 19 n
flabel metal2 32565 241 32609 863 1 FreeSans 800 0 0 0 C[113]
port 18 n
flabel metal2 34453 241 34497 863 1 FreeSans 800 0 0 0 C[114]
port 17 n
flabel metal2 36341 241 36385 863 1 FreeSans 800 0 0 0 C[115]
port 16 n
flabel metal2 38229 241 38273 863 1 FreeSans 800 0 0 0 C[116]
port 15 n
flabel metal2 40117 241 40161 863 1 FreeSans 800 0 0 0 C[117]
port 14 n
flabel metal2 42005 241 42049 863 1 FreeSans 800 0 0 0 C[118]
port 13 n
flabel metal2 43893 241 43937 863 1 FreeSans 800 0 0 0 C[119]
port 12 n
flabel metal2 45781 241 45825 863 1 FreeSans 800 0 0 0 C[120]
port 11 n
flabel metal2 47669 241 47713 863 1 FreeSans 800 0 0 0 C[121]
port 10 n
flabel metal2 49557 241 49601 863 1 FreeSans 800 0 0 0 C[122]
port 9 n
flabel metal2 51445 241 51489 863 1 FreeSans 800 0 0 0 C[123]
port 8 n
flabel metal2 53333 241 53377 863 1 FreeSans 800 0 0 0 C[124]
port 7 n
flabel metal2 55221 241 55265 863 1 FreeSans 800 0 0 0 C[125]
port 6 n
flabel metal2 57109 241 57153 863 1 FreeSans 800 0 0 0 C[126]
port 5 n
flabel metal2 58997 241 59041 863 1 FreeSans 800 0 0 0 C[127]
port 4 n
flabel metal4 1683 -6904 2301 5164 1 FreeSans 1600 0 0 0 VDD
port 1 n
flabel metal4 2916 -4777 3700 7281 1 FreeSans 1600 0 0 0 VSS
port 2 n
flabel metal1 -317 -2720 -187 -2646 1 FreeSans 800 0 0 0 RESET
port 132 n
<< end >>
