* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pnp_05v5_W3p40L3p40__bf_slope = 0.0
.param sky130_fd_pr__pnp_05v5_W3p40L3p40__is_slope = 0.0
.param sky130_fd_pr__pnp_05v5_W3p40L3p40__xti_slope = 0.0
*  statistics {
*   mismatch {
*     vary  sky130_fd_pr__pnp_05v5_W3p40L3p40__bf_slope dist=gauss std=0.05537
*     vary  sky130_fd_pr__pnp_05v5_W3p40L3p40__is_slope dist=gauss std=0.01662
*     vary  sky130_fd_pr__pnp_05v5_W3p40L3p40__xti_slope dist=gauss std=0.06
*   }
* }
.subckt  sky130_fd_pr__pnp_05v5_W3p40L3p40 Collector Base Emitter
+ 
.param  mult = 1.0
+ sky130_fd_pr__pnp_05v5_W3p40L3p40__bf_mm = {(16.603*dkbfpp5x*sky130_fd_pr__pnp_05v5_W3p40L3p40__bf_slope*0.45/sqrt(mult))}
+ sky130_fd_pr__pnp_05v5_W3p40L3p40__is_mm = {(7.1190e-018*1.00*dkispp5x*sky130_fd_pr__pnp_05v5_W3p40L3p40__is_slope*0.13/sqrt(mult))}
+ sky130_fd_pr__pnp_05v5_W3p40L3p40__xti_mm = {(5*sky130_fd_pr__pnp_05v5_W3p40L3p40__xti_slope/sqrt(mult))}
qsky130_fd_pr__pnp_05v5_W3p40L3p40 Collector Base Emitter Collector sky130_fd_pr__pnp_05v5_W3p40L3p40__model
.model sky130_fd_pr__pnp_05v5_W3p40L3p40__model pnp level = 1.0
* General Parameters
+ tref = 30 subs = 1.0
* Capacitance Parameters
+ cjc = '9.155e-17*5.17*5.17*sky130_fd_pr__model__parasitic__diode_ps2nw__ajunction_mult+5.822e-16*4*5.17*sky130_fd_pr__model__parasitic__diode_ps2nw__pjunction_mult' cje = '7.4079e-16*3.4*3.4*sky130_fd_pr__pfet_01v8__ajunction_mult+9.88e-17*4*3.4*sky130_fd_pr__pfet_01v8__pjunction_mult' cjs = 0.0
+ fc = 0.5 mjc = 0.24 mje = 0.3 mjs = 0.24
+ vjc = 0.54 vje = 0.74 vjs = 0.54 xcjc = 1.0
+ ptf = 0 tf = 6.15385e-010 tr = 5e-008 vtf = 1.0e-12
+ xtf = 0.0
* Noise Parameters
+ af = 1.30180 kf = 4.9435066e-11
* DC Parameters
+ is = '7.1190e-018*dkispp5x+sky130_fd_pr__pnp_05v5_W3p40L3p40__is_mm' rb = 73.32 re = 5.3848 irb = 0.0002
+ rc = 100.0 rbm = 25.19 bf = '16.603*dkbfpp5x+sky130_fd_pr__pnp_05v5_W3p40L3p40__bf_mm' nf = '1.000*dknfpp5x'
+ vaf = 111.6 ikf = 0.00038589 ise = '1.0310e-015*dkisepp5x' ne = 1.64
+ ns = 1 br = 0.2675 iss = 0 nr = 1.0
+ var = 4.3 ikr = 0.0043 nkf = 0.426 isc = 1.9855e-15
+ nc = 1.000
* Temperature Parameters
+ xtb = 1.692 xti = '5.0+sky130_fd_pr__pnp_05v5_W3p40L3p40__xti_mm' eg = 1.125 tnf1 = 5.972e-6
+ tikf1 = -0.002456 tnf2 = -3.0e-8
.ends sky130_fd_pr__pnp_05v5_W3p40L3p40
